magic
tech sky130A
timestamp 1640891559
<< nwell >>
rect -680 4800 4720 5480
rect -680 2880 4720 3560
rect -680 960 4720 1640
<< pmoslvt >>
rect -480 5200 -280 5300
rect -480 4980 -280 5080
rect 0 5200 200 5300
rect 320 5200 520 5300
rect 640 5200 840 5300
rect 960 5200 1160 5300
rect 0 4980 200 5080
rect 320 4980 520 5080
rect 640 4980 840 5080
rect 960 4980 1160 5080
rect 1440 5200 1640 5300
rect 1760 5200 1960 5300
rect 2080 5200 2280 5300
rect 2400 5200 2600 5300
rect 1440 4980 1640 5080
rect 1760 4980 1960 5080
rect 2080 4980 2280 5080
rect 2400 4980 2600 5080
rect 2880 5200 3080 5300
rect 3200 5200 3400 5300
rect 3520 5200 3720 5300
rect 3840 5200 4040 5300
rect 2880 4980 3080 5080
rect 3200 4980 3400 5080
rect 3520 4980 3720 5080
rect 3840 4980 4040 5080
rect 4320 5200 4520 5300
rect 4320 4980 4520 5080
rect -480 3280 -280 3380
rect -480 3060 -280 3160
rect 0 3280 200 3380
rect 320 3280 520 3380
rect 640 3280 840 3380
rect 960 3280 1160 3380
rect 0 3060 200 3160
rect 320 3060 520 3160
rect 640 3060 840 3160
rect 960 3060 1160 3160
rect 1440 3280 1640 3380
rect 1760 3280 1960 3380
rect 2080 3280 2280 3380
rect 2400 3280 2600 3380
rect 1440 3060 1640 3160
rect 1760 3060 1960 3160
rect 2080 3060 2280 3160
rect 2400 3060 2600 3160
rect 2880 3280 3080 3380
rect 3200 3280 3400 3380
rect 3520 3280 3720 3380
rect 3840 3280 4040 3380
rect 2880 3060 3080 3160
rect 3200 3060 3400 3160
rect 3520 3060 3720 3160
rect 3840 3060 4040 3160
rect 4320 3280 4520 3380
rect 4320 3060 4520 3160
rect -480 1360 -280 1460
rect -480 1140 -280 1240
rect 0 1360 200 1460
rect 320 1360 520 1460
rect 640 1360 840 1460
rect 960 1360 1160 1460
rect 0 1140 200 1240
rect 320 1140 520 1240
rect 640 1140 840 1240
rect 960 1140 1160 1240
rect 1440 1360 1640 1460
rect 1760 1360 1960 1460
rect 2080 1360 2280 1460
rect 2400 1360 2600 1460
rect 1440 1140 1640 1240
rect 1760 1140 1960 1240
rect 2080 1140 2280 1240
rect 2400 1140 2600 1240
rect 2880 1360 3080 1460
rect 3200 1360 3400 1460
rect 3520 1360 3720 1460
rect 3840 1360 4040 1460
rect 2880 1140 3080 1240
rect 3200 1140 3400 1240
rect 3520 1140 3720 1240
rect 3840 1140 4040 1240
rect 4320 1360 4520 1460
rect 4320 1140 4520 1240
<< nmoslvt >>
rect -480 3840 -280 3940
rect 0 3840 200 3940
rect 320 3840 520 3940
rect 640 3840 840 3940
rect 960 3840 1160 3940
rect 1440 3840 1640 3940
rect 1760 3840 1960 3940
rect 2080 3840 2280 3940
rect 2400 3840 2600 3940
rect 2880 3840 3080 3940
rect 3200 3840 3400 3940
rect 3520 3840 3720 3940
rect 3840 3840 4040 3940
rect 4320 3840 4520 3940
rect -480 1920 -280 2020
rect 0 1920 200 2020
rect 320 1920 520 2020
rect 640 1920 840 2020
rect 960 1920 1160 2020
rect 1440 1920 1640 2020
rect 1760 1920 1960 2020
rect 2080 1920 2280 2020
rect 2400 1920 2600 2020
rect 2880 1920 3080 2020
rect 3200 1920 3400 2020
rect 3520 1920 3720 2020
rect 3840 1920 4040 2020
rect 4320 1920 4520 2020
rect -480 0 -280 100
rect 0 0 200 100
rect 320 0 520 100
rect 640 0 840 100
rect 960 0 1160 100
rect 1440 0 1640 100
rect 1760 0 1960 100
rect 2080 0 2280 100
rect 2400 0 2600 100
rect 2880 0 3080 100
rect 3200 0 3400 100
rect 3520 0 3720 100
rect 3840 0 4040 100
rect 4320 0 4520 100
<< ndiff >>
rect -560 3930 -480 3940
rect -560 3850 -555 3930
rect -525 3850 -480 3930
rect -560 3840 -480 3850
rect -280 3930 -200 3940
rect -280 3850 -235 3930
rect -205 3850 -200 3930
rect -280 3840 -200 3850
rect -80 3930 0 3940
rect -80 3850 -75 3930
rect -45 3850 0 3930
rect -80 3840 0 3850
rect 200 3930 320 3940
rect 200 3850 245 3930
rect 275 3850 320 3930
rect 200 3840 320 3850
rect 520 3930 640 3940
rect 520 3850 565 3930
rect 595 3850 640 3930
rect 520 3840 640 3850
rect 840 3930 960 3940
rect 840 3850 885 3930
rect 915 3850 960 3930
rect 840 3840 960 3850
rect 1160 3930 1240 3940
rect 1160 3850 1205 3930
rect 1235 3850 1240 3930
rect 1160 3840 1240 3850
rect 1360 3930 1440 3940
rect 1360 3850 1365 3930
rect 1395 3850 1440 3930
rect 1360 3840 1440 3850
rect 1640 3930 1760 3940
rect 1640 3850 1685 3930
rect 1715 3850 1760 3930
rect 1640 3840 1760 3850
rect 1960 3930 2080 3940
rect 1960 3850 2005 3930
rect 2035 3850 2080 3930
rect 1960 3840 2080 3850
rect 2280 3930 2400 3940
rect 2280 3850 2325 3930
rect 2355 3850 2400 3930
rect 2280 3840 2400 3850
rect 2600 3930 2680 3940
rect 2600 3850 2645 3930
rect 2675 3850 2680 3930
rect 2600 3840 2680 3850
rect 2800 3930 2880 3940
rect 2800 3850 2805 3930
rect 2835 3850 2880 3930
rect 2800 3840 2880 3850
rect 3080 3930 3200 3940
rect 3080 3850 3125 3930
rect 3155 3850 3200 3930
rect 3080 3840 3200 3850
rect 3400 3930 3520 3940
rect 3400 3850 3445 3930
rect 3475 3850 3520 3930
rect 3400 3840 3520 3850
rect 3720 3930 3840 3940
rect 3720 3850 3765 3930
rect 3795 3850 3840 3930
rect 3720 3840 3840 3850
rect 4040 3930 4120 3940
rect 4040 3850 4085 3930
rect 4115 3850 4120 3930
rect 4040 3840 4120 3850
rect 4240 3930 4320 3940
rect 4240 3850 4245 3930
rect 4275 3850 4320 3930
rect 4240 3840 4320 3850
rect 4520 3930 4600 3940
rect 4520 3850 4565 3930
rect 4595 3850 4600 3930
rect 4520 3840 4600 3850
rect -560 2010 -480 2020
rect -560 1930 -555 2010
rect -525 1930 -480 2010
rect -560 1920 -480 1930
rect -280 2010 -200 2020
rect -280 1930 -235 2010
rect -205 1930 -200 2010
rect -280 1920 -200 1930
rect -80 2010 0 2020
rect -80 1930 -75 2010
rect -45 1930 0 2010
rect -80 1920 0 1930
rect 200 2010 320 2020
rect 200 1930 245 2010
rect 275 1930 320 2010
rect 200 1920 320 1930
rect 520 2010 640 2020
rect 520 1930 565 2010
rect 595 1930 640 2010
rect 520 1920 640 1930
rect 840 2010 960 2020
rect 840 1930 885 2010
rect 915 1930 960 2010
rect 840 1920 960 1930
rect 1160 2010 1240 2020
rect 1160 1930 1205 2010
rect 1235 1930 1240 2010
rect 1160 1920 1240 1930
rect 1360 2010 1440 2020
rect 1360 1930 1365 2010
rect 1395 1930 1440 2010
rect 1360 1920 1440 1930
rect 1640 2010 1760 2020
rect 1640 1930 1685 2010
rect 1715 1930 1760 2010
rect 1640 1920 1760 1930
rect 1960 2010 2080 2020
rect 1960 1930 2005 2010
rect 2035 1930 2080 2010
rect 1960 1920 2080 1930
rect 2280 2010 2400 2020
rect 2280 1930 2325 2010
rect 2355 1930 2400 2010
rect 2280 1920 2400 1930
rect 2600 2010 2680 2020
rect 2600 1930 2645 2010
rect 2675 1930 2680 2010
rect 2600 1920 2680 1930
rect 2800 2010 2880 2020
rect 2800 1930 2805 2010
rect 2835 1930 2880 2010
rect 2800 1920 2880 1930
rect 3080 2010 3200 2020
rect 3080 1930 3125 2010
rect 3155 1930 3200 2010
rect 3080 1920 3200 1930
rect 3400 2010 3520 2020
rect 3400 1930 3445 2010
rect 3475 1930 3520 2010
rect 3400 1920 3520 1930
rect 3720 2010 3840 2020
rect 3720 1930 3765 2010
rect 3795 1930 3840 2010
rect 3720 1920 3840 1930
rect 4040 2010 4120 2020
rect 4040 1930 4085 2010
rect 4115 1930 4120 2010
rect 4040 1920 4120 1930
rect 4240 2010 4320 2020
rect 4240 1930 4245 2010
rect 4275 1930 4320 2010
rect 4240 1920 4320 1930
rect 4520 2010 4600 2020
rect 4520 1930 4565 2010
rect 4595 1930 4600 2010
rect 4520 1920 4600 1930
rect -560 90 -480 100
rect -560 10 -555 90
rect -525 10 -480 90
rect -560 0 -480 10
rect -280 90 -200 100
rect -280 10 -235 90
rect -205 10 -200 90
rect -280 0 -200 10
rect -80 90 0 100
rect -80 10 -75 90
rect -45 10 0 90
rect -80 0 0 10
rect 200 90 320 100
rect 200 10 245 90
rect 275 10 320 90
rect 200 0 320 10
rect 520 90 640 100
rect 520 10 565 90
rect 595 10 640 90
rect 520 0 640 10
rect 840 90 960 100
rect 840 10 885 90
rect 915 10 960 90
rect 840 0 960 10
rect 1160 90 1240 100
rect 1160 10 1205 90
rect 1235 10 1240 90
rect 1160 0 1240 10
rect 1360 90 1440 100
rect 1360 10 1365 90
rect 1395 10 1440 90
rect 1360 0 1440 10
rect 1640 90 1760 100
rect 1640 10 1685 90
rect 1715 10 1760 90
rect 1640 0 1760 10
rect 1960 90 2080 100
rect 1960 10 2005 90
rect 2035 10 2080 90
rect 1960 0 2080 10
rect 2280 90 2400 100
rect 2280 10 2325 90
rect 2355 10 2400 90
rect 2280 0 2400 10
rect 2600 90 2680 100
rect 2600 10 2645 90
rect 2675 10 2680 90
rect 2600 0 2680 10
rect 2800 90 2880 100
rect 2800 10 2805 90
rect 2835 10 2880 90
rect 2800 0 2880 10
rect 3080 90 3200 100
rect 3080 10 3125 90
rect 3155 10 3200 90
rect 3080 0 3200 10
rect 3400 90 3520 100
rect 3400 10 3445 90
rect 3475 10 3520 90
rect 3400 0 3520 10
rect 3720 90 3840 100
rect 3720 10 3765 90
rect 3795 10 3840 90
rect 3720 0 3840 10
rect 4040 90 4120 100
rect 4040 10 4085 90
rect 4115 10 4120 90
rect 4040 0 4120 10
rect 4240 90 4320 100
rect 4240 10 4245 90
rect 4275 10 4320 90
rect 4240 0 4320 10
rect 4520 90 4600 100
rect 4520 10 4565 90
rect 4595 10 4600 90
rect 4520 0 4600 10
<< pdiff >>
rect -560 5290 -480 5300
rect -560 5210 -555 5290
rect -525 5210 -480 5290
rect -560 5200 -480 5210
rect -280 5290 -200 5300
rect -280 5210 -235 5290
rect -205 5210 -200 5290
rect -280 5200 -200 5210
rect -560 5070 -480 5080
rect -560 4990 -555 5070
rect -525 4990 -480 5070
rect -560 4980 -480 4990
rect -280 5070 -200 5080
rect -280 4990 -235 5070
rect -205 4990 -200 5070
rect -280 4980 -200 4990
rect -80 5290 0 5300
rect -80 5210 -75 5290
rect -45 5210 0 5290
rect -80 5200 0 5210
rect 200 5290 320 5300
rect 200 5210 245 5290
rect 275 5210 320 5290
rect 200 5200 320 5210
rect 520 5290 640 5300
rect 520 5210 565 5290
rect 595 5210 640 5290
rect 520 5200 640 5210
rect 840 5290 960 5300
rect 840 5210 885 5290
rect 915 5210 960 5290
rect 840 5200 960 5210
rect 1160 5290 1240 5300
rect 1160 5210 1205 5290
rect 1235 5210 1240 5290
rect 1160 5200 1240 5210
rect -80 5070 0 5080
rect -80 4990 -75 5070
rect -45 4990 0 5070
rect -80 4980 0 4990
rect 200 5070 320 5080
rect 200 4990 245 5070
rect 275 4990 320 5070
rect 200 4980 320 4990
rect 520 5070 640 5080
rect 520 4990 565 5070
rect 595 4990 640 5070
rect 520 4980 640 4990
rect 840 5070 960 5080
rect 840 4990 885 5070
rect 915 4990 960 5070
rect 840 4980 960 4990
rect 1160 5070 1240 5080
rect 1160 4990 1205 5070
rect 1235 4990 1240 5070
rect 1160 4980 1240 4990
rect 1360 5290 1440 5300
rect 1360 5210 1365 5290
rect 1395 5210 1440 5290
rect 1360 5200 1440 5210
rect 1640 5290 1760 5300
rect 1640 5210 1685 5290
rect 1715 5210 1760 5290
rect 1640 5200 1760 5210
rect 1960 5290 2080 5300
rect 1960 5210 2005 5290
rect 2035 5210 2080 5290
rect 1960 5200 2080 5210
rect 2280 5290 2400 5300
rect 2280 5210 2325 5290
rect 2355 5210 2400 5290
rect 2280 5200 2400 5210
rect 2600 5290 2680 5300
rect 2600 5210 2645 5290
rect 2675 5210 2680 5290
rect 2600 5200 2680 5210
rect 1360 5070 1440 5080
rect 1360 4990 1365 5070
rect 1395 4990 1440 5070
rect 1360 4980 1440 4990
rect 1640 5070 1760 5080
rect 1640 4990 1685 5070
rect 1715 4990 1760 5070
rect 1640 4980 1760 4990
rect 1960 5070 2080 5080
rect 1960 4990 2005 5070
rect 2035 4990 2080 5070
rect 1960 4980 2080 4990
rect 2280 5070 2400 5080
rect 2280 4990 2325 5070
rect 2355 4990 2400 5070
rect 2280 4980 2400 4990
rect 2600 5070 2680 5080
rect 2600 4990 2645 5070
rect 2675 4990 2680 5070
rect 2600 4980 2680 4990
rect 2800 5290 2880 5300
rect 2800 5210 2805 5290
rect 2835 5210 2880 5290
rect 2800 5200 2880 5210
rect 3080 5290 3200 5300
rect 3080 5210 3125 5290
rect 3155 5210 3200 5290
rect 3080 5200 3200 5210
rect 3400 5290 3520 5300
rect 3400 5210 3445 5290
rect 3475 5210 3520 5290
rect 3400 5200 3520 5210
rect 3720 5290 3840 5300
rect 3720 5210 3765 5290
rect 3795 5210 3840 5290
rect 3720 5200 3840 5210
rect 4040 5290 4120 5300
rect 4040 5210 4085 5290
rect 4115 5210 4120 5290
rect 4040 5200 4120 5210
rect 2800 5070 2880 5080
rect 2800 4990 2805 5070
rect 2835 4990 2880 5070
rect 2800 4980 2880 4990
rect 3080 5070 3200 5080
rect 3080 4990 3125 5070
rect 3155 4990 3200 5070
rect 3080 4980 3200 4990
rect 3400 5070 3520 5080
rect 3400 4990 3445 5070
rect 3475 4990 3520 5070
rect 3400 4980 3520 4990
rect 3720 5070 3840 5080
rect 3720 4990 3765 5070
rect 3795 4990 3840 5070
rect 3720 4980 3840 4990
rect 4040 5070 4120 5080
rect 4040 4990 4085 5070
rect 4115 4990 4120 5070
rect 4040 4980 4120 4990
rect 4240 5290 4320 5300
rect 4240 5210 4245 5290
rect 4275 5210 4320 5290
rect 4240 5200 4320 5210
rect 4520 5290 4600 5300
rect 4520 5210 4565 5290
rect 4595 5210 4600 5290
rect 4520 5200 4600 5210
rect 4240 5070 4320 5080
rect 4240 4990 4245 5070
rect 4275 4990 4320 5070
rect 4240 4980 4320 4990
rect 4520 5070 4600 5080
rect 4520 4990 4565 5070
rect 4595 4990 4600 5070
rect 4520 4980 4600 4990
rect -560 3370 -480 3380
rect -560 3290 -555 3370
rect -525 3290 -480 3370
rect -560 3280 -480 3290
rect -280 3370 -200 3380
rect -280 3290 -235 3370
rect -205 3290 -200 3370
rect -280 3280 -200 3290
rect -560 3150 -480 3160
rect -560 3070 -555 3150
rect -525 3070 -480 3150
rect -560 3060 -480 3070
rect -280 3150 -200 3160
rect -280 3070 -235 3150
rect -205 3070 -200 3150
rect -280 3060 -200 3070
rect -80 3370 0 3380
rect -80 3290 -75 3370
rect -45 3290 0 3370
rect -80 3280 0 3290
rect 200 3370 320 3380
rect 200 3290 245 3370
rect 275 3290 320 3370
rect 200 3280 320 3290
rect 520 3370 640 3380
rect 520 3290 565 3370
rect 595 3290 640 3370
rect 520 3280 640 3290
rect 840 3370 960 3380
rect 840 3290 885 3370
rect 915 3290 960 3370
rect 840 3280 960 3290
rect 1160 3370 1240 3380
rect 1160 3290 1205 3370
rect 1235 3290 1240 3370
rect 1160 3280 1240 3290
rect -80 3150 0 3160
rect -80 3070 -75 3150
rect -45 3070 0 3150
rect -80 3060 0 3070
rect 200 3150 320 3160
rect 200 3070 245 3150
rect 275 3070 320 3150
rect 200 3060 320 3070
rect 520 3150 640 3160
rect 520 3070 565 3150
rect 595 3070 640 3150
rect 520 3060 640 3070
rect 840 3150 960 3160
rect 840 3070 885 3150
rect 915 3070 960 3150
rect 840 3060 960 3070
rect 1160 3150 1240 3160
rect 1160 3070 1205 3150
rect 1235 3070 1240 3150
rect 1160 3060 1240 3070
rect 1360 3370 1440 3380
rect 1360 3290 1365 3370
rect 1395 3290 1440 3370
rect 1360 3280 1440 3290
rect 1640 3370 1760 3380
rect 1640 3290 1685 3370
rect 1715 3290 1760 3370
rect 1640 3280 1760 3290
rect 1960 3370 2080 3380
rect 1960 3290 2005 3370
rect 2035 3290 2080 3370
rect 1960 3280 2080 3290
rect 2280 3370 2400 3380
rect 2280 3290 2325 3370
rect 2355 3290 2400 3370
rect 2280 3280 2400 3290
rect 2600 3370 2680 3380
rect 2600 3290 2645 3370
rect 2675 3290 2680 3370
rect 2600 3280 2680 3290
rect 1360 3150 1440 3160
rect 1360 3070 1365 3150
rect 1395 3070 1440 3150
rect 1360 3060 1440 3070
rect 1640 3150 1760 3160
rect 1640 3070 1685 3150
rect 1715 3070 1760 3150
rect 1640 3060 1760 3070
rect 1960 3150 2080 3160
rect 1960 3070 2005 3150
rect 2035 3070 2080 3150
rect 1960 3060 2080 3070
rect 2280 3150 2400 3160
rect 2280 3070 2325 3150
rect 2355 3070 2400 3150
rect 2280 3060 2400 3070
rect 2600 3150 2680 3160
rect 2600 3070 2645 3150
rect 2675 3070 2680 3150
rect 2600 3060 2680 3070
rect 2800 3370 2880 3380
rect 2800 3290 2805 3370
rect 2835 3290 2880 3370
rect 2800 3280 2880 3290
rect 3080 3370 3200 3380
rect 3080 3290 3125 3370
rect 3155 3290 3200 3370
rect 3080 3280 3200 3290
rect 3400 3370 3520 3380
rect 3400 3290 3445 3370
rect 3475 3290 3520 3370
rect 3400 3280 3520 3290
rect 3720 3370 3840 3380
rect 3720 3290 3765 3370
rect 3795 3290 3840 3370
rect 3720 3280 3840 3290
rect 4040 3370 4120 3380
rect 4040 3290 4085 3370
rect 4115 3290 4120 3370
rect 4040 3280 4120 3290
rect 2800 3150 2880 3160
rect 2800 3070 2805 3150
rect 2835 3070 2880 3150
rect 2800 3060 2880 3070
rect 3080 3150 3200 3160
rect 3080 3070 3125 3150
rect 3155 3070 3200 3150
rect 3080 3060 3200 3070
rect 3400 3150 3520 3160
rect 3400 3070 3445 3150
rect 3475 3070 3520 3150
rect 3400 3060 3520 3070
rect 3720 3150 3840 3160
rect 3720 3070 3765 3150
rect 3795 3070 3840 3150
rect 3720 3060 3840 3070
rect 4040 3150 4120 3160
rect 4040 3070 4085 3150
rect 4115 3070 4120 3150
rect 4040 3060 4120 3070
rect 4240 3370 4320 3380
rect 4240 3290 4245 3370
rect 4275 3290 4320 3370
rect 4240 3280 4320 3290
rect 4520 3370 4600 3380
rect 4520 3290 4565 3370
rect 4595 3290 4600 3370
rect 4520 3280 4600 3290
rect 4240 3150 4320 3160
rect 4240 3070 4245 3150
rect 4275 3070 4320 3150
rect 4240 3060 4320 3070
rect 4520 3150 4600 3160
rect 4520 3070 4565 3150
rect 4595 3070 4600 3150
rect 4520 3060 4600 3070
rect -560 1450 -480 1460
rect -560 1370 -555 1450
rect -525 1370 -480 1450
rect -560 1360 -480 1370
rect -280 1450 -200 1460
rect -280 1370 -235 1450
rect -205 1370 -200 1450
rect -280 1360 -200 1370
rect -560 1230 -480 1240
rect -560 1150 -555 1230
rect -525 1150 -480 1230
rect -560 1140 -480 1150
rect -280 1230 -200 1240
rect -280 1150 -235 1230
rect -205 1150 -200 1230
rect -280 1140 -200 1150
rect -80 1450 0 1460
rect -80 1370 -75 1450
rect -45 1370 0 1450
rect -80 1360 0 1370
rect 200 1450 320 1460
rect 200 1370 245 1450
rect 275 1370 320 1450
rect 200 1360 320 1370
rect 520 1450 640 1460
rect 520 1370 565 1450
rect 595 1370 640 1450
rect 520 1360 640 1370
rect 840 1450 960 1460
rect 840 1370 885 1450
rect 915 1370 960 1450
rect 840 1360 960 1370
rect 1160 1450 1240 1460
rect 1160 1370 1205 1450
rect 1235 1370 1240 1450
rect 1160 1360 1240 1370
rect -80 1230 0 1240
rect -80 1150 -75 1230
rect -45 1150 0 1230
rect -80 1140 0 1150
rect 200 1230 320 1240
rect 200 1150 245 1230
rect 275 1150 320 1230
rect 200 1140 320 1150
rect 520 1230 640 1240
rect 520 1150 565 1230
rect 595 1150 640 1230
rect 520 1140 640 1150
rect 840 1230 960 1240
rect 840 1150 885 1230
rect 915 1150 960 1230
rect 840 1140 960 1150
rect 1160 1230 1240 1240
rect 1160 1150 1205 1230
rect 1235 1150 1240 1230
rect 1160 1140 1240 1150
rect 1360 1450 1440 1460
rect 1360 1370 1365 1450
rect 1395 1370 1440 1450
rect 1360 1360 1440 1370
rect 1640 1450 1760 1460
rect 1640 1370 1685 1450
rect 1715 1370 1760 1450
rect 1640 1360 1760 1370
rect 1960 1450 2080 1460
rect 1960 1370 2005 1450
rect 2035 1370 2080 1450
rect 1960 1360 2080 1370
rect 2280 1450 2400 1460
rect 2280 1370 2325 1450
rect 2355 1370 2400 1450
rect 2280 1360 2400 1370
rect 2600 1450 2680 1460
rect 2600 1370 2645 1450
rect 2675 1370 2680 1450
rect 2600 1360 2680 1370
rect 1360 1230 1440 1240
rect 1360 1150 1365 1230
rect 1395 1150 1440 1230
rect 1360 1140 1440 1150
rect 1640 1230 1760 1240
rect 1640 1150 1685 1230
rect 1715 1150 1760 1230
rect 1640 1140 1760 1150
rect 1960 1230 2080 1240
rect 1960 1150 2005 1230
rect 2035 1150 2080 1230
rect 1960 1140 2080 1150
rect 2280 1230 2400 1240
rect 2280 1150 2325 1230
rect 2355 1150 2400 1230
rect 2280 1140 2400 1150
rect 2600 1230 2680 1240
rect 2600 1150 2645 1230
rect 2675 1150 2680 1230
rect 2600 1140 2680 1150
rect 2800 1450 2880 1460
rect 2800 1370 2805 1450
rect 2835 1370 2880 1450
rect 2800 1360 2880 1370
rect 3080 1450 3200 1460
rect 3080 1370 3125 1450
rect 3155 1370 3200 1450
rect 3080 1360 3200 1370
rect 3400 1450 3520 1460
rect 3400 1370 3445 1450
rect 3475 1370 3520 1450
rect 3400 1360 3520 1370
rect 3720 1450 3840 1460
rect 3720 1370 3765 1450
rect 3795 1370 3840 1450
rect 3720 1360 3840 1370
rect 4040 1450 4120 1460
rect 4040 1370 4085 1450
rect 4115 1370 4120 1450
rect 4040 1360 4120 1370
rect 2800 1230 2880 1240
rect 2800 1150 2805 1230
rect 2835 1150 2880 1230
rect 2800 1140 2880 1150
rect 3080 1230 3200 1240
rect 3080 1150 3125 1230
rect 3155 1150 3200 1230
rect 3080 1140 3200 1150
rect 3400 1230 3520 1240
rect 3400 1150 3445 1230
rect 3475 1150 3520 1230
rect 3400 1140 3520 1150
rect 3720 1230 3840 1240
rect 3720 1150 3765 1230
rect 3795 1150 3840 1230
rect 3720 1140 3840 1150
rect 4040 1230 4120 1240
rect 4040 1150 4085 1230
rect 4115 1150 4120 1230
rect 4040 1140 4120 1150
rect 4240 1450 4320 1460
rect 4240 1370 4245 1450
rect 4275 1370 4320 1450
rect 4240 1360 4320 1370
rect 4520 1450 4600 1460
rect 4520 1370 4565 1450
rect 4595 1370 4600 1450
rect 4520 1360 4600 1370
rect 4240 1230 4320 1240
rect 4240 1150 4245 1230
rect 4275 1150 4320 1230
rect 4240 1140 4320 1150
rect 4520 1230 4600 1240
rect 4520 1150 4565 1230
rect 4595 1150 4600 1230
rect 4520 1140 4600 1150
<< ndiffc >>
rect -555 3850 -525 3930
rect -235 3850 -205 3930
rect -75 3850 -45 3930
rect 245 3850 275 3930
rect 565 3850 595 3930
rect 885 3850 915 3930
rect 1205 3850 1235 3930
rect 1365 3850 1395 3930
rect 1685 3850 1715 3930
rect 2005 3850 2035 3930
rect 2325 3850 2355 3930
rect 2645 3850 2675 3930
rect 2805 3850 2835 3930
rect 3125 3850 3155 3930
rect 3445 3850 3475 3930
rect 3765 3850 3795 3930
rect 4085 3850 4115 3930
rect 4245 3850 4275 3930
rect 4565 3850 4595 3930
rect -555 1930 -525 2010
rect -235 1930 -205 2010
rect -75 1930 -45 2010
rect 245 1930 275 2010
rect 565 1930 595 2010
rect 885 1930 915 2010
rect 1205 1930 1235 2010
rect 1365 1930 1395 2010
rect 1685 1930 1715 2010
rect 2005 1930 2035 2010
rect 2325 1930 2355 2010
rect 2645 1930 2675 2010
rect 2805 1930 2835 2010
rect 3125 1930 3155 2010
rect 3445 1930 3475 2010
rect 3765 1930 3795 2010
rect 4085 1930 4115 2010
rect 4245 1930 4275 2010
rect 4565 1930 4595 2010
rect -555 10 -525 90
rect -235 10 -205 90
rect -75 10 -45 90
rect 245 10 275 90
rect 565 10 595 90
rect 885 10 915 90
rect 1205 10 1235 90
rect 1365 10 1395 90
rect 1685 10 1715 90
rect 2005 10 2035 90
rect 2325 10 2355 90
rect 2645 10 2675 90
rect 2805 10 2835 90
rect 3125 10 3155 90
rect 3445 10 3475 90
rect 3765 10 3795 90
rect 4085 10 4115 90
rect 4245 10 4275 90
rect 4565 10 4595 90
<< pdiffc >>
rect -555 5210 -525 5290
rect -235 5210 -205 5290
rect -555 4990 -525 5070
rect -235 4990 -205 5070
rect -75 5210 -45 5290
rect 245 5210 275 5290
rect 565 5210 595 5290
rect 885 5210 915 5290
rect 1205 5210 1235 5290
rect -75 4990 -45 5070
rect 245 4990 275 5070
rect 565 4990 595 5070
rect 885 4990 915 5070
rect 1205 4990 1235 5070
rect 1365 5210 1395 5290
rect 1685 5210 1715 5290
rect 2005 5210 2035 5290
rect 2325 5210 2355 5290
rect 2645 5210 2675 5290
rect 1365 4990 1395 5070
rect 1685 4990 1715 5070
rect 2005 4990 2035 5070
rect 2325 4990 2355 5070
rect 2645 4990 2675 5070
rect 2805 5210 2835 5290
rect 3125 5210 3155 5290
rect 3445 5210 3475 5290
rect 3765 5210 3795 5290
rect 4085 5210 4115 5290
rect 2805 4990 2835 5070
rect 3125 4990 3155 5070
rect 3445 4990 3475 5070
rect 3765 4990 3795 5070
rect 4085 4990 4115 5070
rect 4245 5210 4275 5290
rect 4565 5210 4595 5290
rect 4245 4990 4275 5070
rect 4565 4990 4595 5070
rect -555 3290 -525 3370
rect -235 3290 -205 3370
rect -555 3070 -525 3150
rect -235 3070 -205 3150
rect -75 3290 -45 3370
rect 245 3290 275 3370
rect 565 3290 595 3370
rect 885 3290 915 3370
rect 1205 3290 1235 3370
rect -75 3070 -45 3150
rect 245 3070 275 3150
rect 565 3070 595 3150
rect 885 3070 915 3150
rect 1205 3070 1235 3150
rect 1365 3290 1395 3370
rect 1685 3290 1715 3370
rect 2005 3290 2035 3370
rect 2325 3290 2355 3370
rect 2645 3290 2675 3370
rect 1365 3070 1395 3150
rect 1685 3070 1715 3150
rect 2005 3070 2035 3150
rect 2325 3070 2355 3150
rect 2645 3070 2675 3150
rect 2805 3290 2835 3370
rect 3125 3290 3155 3370
rect 3445 3290 3475 3370
rect 3765 3290 3795 3370
rect 4085 3290 4115 3370
rect 2805 3070 2835 3150
rect 3125 3070 3155 3150
rect 3445 3070 3475 3150
rect 3765 3070 3795 3150
rect 4085 3070 4115 3150
rect 4245 3290 4275 3370
rect 4565 3290 4595 3370
rect 4245 3070 4275 3150
rect 4565 3070 4595 3150
rect -555 1370 -525 1450
rect -235 1370 -205 1450
rect -555 1150 -525 1230
rect -235 1150 -205 1230
rect -75 1370 -45 1450
rect 245 1370 275 1450
rect 565 1370 595 1450
rect 885 1370 915 1450
rect 1205 1370 1235 1450
rect -75 1150 -45 1230
rect 245 1150 275 1230
rect 565 1150 595 1230
rect 885 1150 915 1230
rect 1205 1150 1235 1230
rect 1365 1370 1395 1450
rect 1685 1370 1715 1450
rect 2005 1370 2035 1450
rect 2325 1370 2355 1450
rect 2645 1370 2675 1450
rect 1365 1150 1395 1230
rect 1685 1150 1715 1230
rect 2005 1150 2035 1230
rect 2325 1150 2355 1230
rect 2645 1150 2675 1230
rect 2805 1370 2835 1450
rect 3125 1370 3155 1450
rect 3445 1370 3475 1450
rect 3765 1370 3795 1450
rect 4085 1370 4115 1450
rect 2805 1150 2835 1230
rect 3125 1150 3155 1230
rect 3445 1150 3475 1230
rect 3765 1150 3795 1230
rect 4085 1150 4115 1230
rect 4245 1370 4275 1450
rect 4565 1370 4595 1450
rect 4245 1150 4275 1230
rect 4565 1150 4595 1230
<< psubdiff >>
rect -800 5560 -680 5600
rect 4760 5560 4840 5600
rect -800 4680 -680 4720
rect 4760 4680 4840 4720
rect -800 4040 -560 4080
rect -200 4040 -80 4080
rect 1240 4040 1360 4080
rect 2680 4040 2800 4080
rect 4120 4040 4240 4080
rect 4600 4040 4840 4080
rect -800 3720 -560 3760
rect -200 3720 -80 3760
rect 1240 3720 1360 3760
rect 2680 3720 2800 3760
rect 4120 3720 4240 3760
rect 4600 3720 4840 3760
rect -800 3680 -760 3720
rect 4800 3680 4840 3720
rect -800 3640 -680 3680
rect 4760 3640 4840 3680
rect -800 2760 -680 2800
rect 4760 2760 4840 2800
rect -800 2120 -560 2160
rect -200 2120 -80 2160
rect 1240 2120 1360 2160
rect 2680 2120 2800 2160
rect 4120 2120 4240 2160
rect 4600 2120 4840 2160
rect -800 1800 -560 1840
rect -200 1800 -80 1840
rect 1240 1800 1360 1840
rect 2680 1800 2800 1840
rect 4120 1800 4240 1840
rect 4600 1800 4840 1840
rect -800 1760 -760 1800
rect 4800 1760 4840 1800
rect -800 1720 -680 1760
rect 4760 1720 4840 1760
rect -800 840 -680 880
rect 4760 840 4840 880
rect -800 200 -560 240
rect -200 200 -80 240
rect 1240 200 1360 240
rect 2680 200 2800 240
rect 4120 200 4240 240
rect 4600 200 4840 240
rect -800 -120 -560 -80
rect -200 -120 -80 -80
rect 1240 -120 1360 -80
rect 2680 -120 2800 -80
rect 4120 -120 4240 -80
rect 4600 -120 4840 -80
<< nsubdiff >>
rect -640 5400 -560 5440
rect -200 5400 -80 5440
rect 1240 5400 1360 5440
rect 2680 5400 2800 5440
rect 4120 5400 4240 5440
rect 4600 5400 4680 5440
rect -640 4840 -560 4880
rect -200 4840 -80 4880
rect 1240 4840 1360 4880
rect 2680 4840 2800 4880
rect 4120 4840 4240 4880
rect 4600 4840 4680 4880
rect -640 3480 -560 3520
rect -200 3480 -80 3520
rect 1240 3480 1360 3520
rect 2680 3480 2800 3520
rect 4120 3480 4240 3520
rect 4600 3480 4680 3520
rect -640 2920 -560 2960
rect -200 2920 -80 2960
rect 1240 2920 1360 2960
rect 2680 2920 2800 2960
rect 4120 2920 4240 2960
rect 4600 2920 4680 2960
rect -640 1560 -560 1600
rect -200 1560 -80 1600
rect 1240 1560 1360 1600
rect 2680 1560 2800 1600
rect 4120 1560 4240 1600
rect 4600 1560 4680 1600
rect -640 1000 -560 1040
rect -200 1000 -80 1040
rect 1240 1000 1360 1040
rect 2680 1000 2800 1040
rect 4120 1000 4240 1040
rect 4600 1000 4680 1040
<< psubdiffcont >>
rect -680 5560 4760 5600
rect -800 4720 -760 5560
rect 4800 4720 4840 5560
rect -680 4680 4760 4720
rect -800 4080 -760 4680
rect 4800 4080 4840 4680
rect -560 4040 -200 4080
rect -80 4040 1240 4080
rect 1360 4040 2680 4080
rect 2800 4040 4120 4080
rect 4240 4040 4600 4080
rect -800 3760 -760 4040
rect -640 3760 -600 4040
rect -160 3760 -120 4040
rect 1280 3760 1320 4040
rect 2720 3760 2760 4040
rect 4160 3760 4200 4040
rect 4640 3760 4680 4040
rect 4800 3760 4840 4040
rect -560 3720 -200 3760
rect -80 3720 1240 3760
rect 1360 3720 2680 3760
rect 2800 3720 4120 3760
rect 4240 3720 4600 3760
rect -680 3640 4760 3680
rect -800 2800 -760 3640
rect 4800 2800 4840 3640
rect -680 2760 4760 2800
rect -800 2160 -760 2760
rect 4800 2160 4840 2760
rect -560 2120 -200 2160
rect -80 2120 1240 2160
rect 1360 2120 2680 2160
rect 2800 2120 4120 2160
rect 4240 2120 4600 2160
rect -800 1840 -760 2120
rect -640 1840 -600 2120
rect -160 1840 -120 2120
rect 1280 1840 1320 2120
rect 2720 1840 2760 2120
rect 4160 1840 4200 2120
rect 4640 1840 4680 2120
rect 4800 1840 4840 2120
rect -560 1800 -200 1840
rect -80 1800 1240 1840
rect 1360 1800 2680 1840
rect 2800 1800 4120 1840
rect 4240 1800 4600 1840
rect -680 1720 4760 1760
rect -800 880 -760 1720
rect 4800 880 4840 1720
rect -680 840 4760 880
rect -800 240 -760 840
rect 4800 240 4840 840
rect -560 200 -200 240
rect -80 200 1240 240
rect 1360 200 2680 240
rect 2800 200 4120 240
rect 4240 200 4600 240
rect -800 -80 -760 200
rect -640 -80 -600 200
rect -160 -80 -120 200
rect 1280 -80 1320 200
rect 2720 -80 2760 200
rect 4160 -80 4200 200
rect 4640 -80 4680 200
rect 4800 -80 4840 200
rect -560 -120 -200 -80
rect -80 -120 1240 -80
rect 1360 -120 2680 -80
rect 2800 -120 4120 -80
rect 4240 -120 4600 -80
<< nsubdiffcont >>
rect -560 5400 -200 5440
rect -80 5400 1240 5440
rect 1360 5400 2680 5440
rect 2800 5400 4120 5440
rect 4240 5400 4600 5440
rect -640 4880 -600 5400
rect -160 4880 -120 5400
rect 1280 4880 1320 5400
rect 2720 4880 2760 5400
rect 4160 4880 4200 5400
rect 4640 4880 4680 5400
rect -560 4840 -200 4880
rect -80 4840 1240 4880
rect 1360 4840 2680 4880
rect 2800 4840 4120 4880
rect 4240 4840 4600 4880
rect -560 3480 -200 3520
rect -80 3480 1240 3520
rect 1360 3480 2680 3520
rect 2800 3480 4120 3520
rect 4240 3480 4600 3520
rect -640 2960 -600 3480
rect -160 2960 -120 3480
rect 1280 2960 1320 3480
rect 2720 2960 2760 3480
rect 4160 2960 4200 3480
rect 4640 2960 4680 3480
rect -560 2920 -200 2960
rect -80 2920 1240 2960
rect 1360 2920 2680 2960
rect 2800 2920 4120 2960
rect 4240 2920 4600 2960
rect -560 1560 -200 1600
rect -80 1560 1240 1600
rect 1360 1560 2680 1600
rect 2800 1560 4120 1600
rect 4240 1560 4600 1600
rect -640 1040 -600 1560
rect -160 1040 -120 1560
rect 1280 1040 1320 1560
rect 2720 1040 2760 1560
rect 4160 1040 4200 1560
rect 4640 1040 4680 1560
rect -560 1000 -200 1040
rect -80 1000 1240 1040
rect 1360 1000 2680 1040
rect 2800 1000 4120 1040
rect 4240 1000 4600 1040
<< poly >>
rect -480 5355 -280 5360
rect -480 5325 -470 5355
rect -290 5325 -280 5355
rect -480 5300 -280 5325
rect -480 5180 -280 5200
rect -480 5080 -280 5100
rect -480 4955 -280 4980
rect -480 4925 -470 4955
rect -290 4925 -280 4955
rect -480 4920 -280 4925
rect 0 5355 200 5360
rect 0 5325 10 5355
rect 190 5325 200 5355
rect 0 5300 200 5325
rect 320 5355 520 5360
rect 320 5325 330 5355
rect 510 5325 520 5355
rect 320 5300 520 5325
rect 640 5355 840 5360
rect 640 5325 650 5355
rect 830 5325 840 5355
rect 640 5300 840 5325
rect 960 5355 1160 5360
rect 960 5325 970 5355
rect 1150 5325 1160 5355
rect 960 5300 1160 5325
rect 0 5180 200 5200
rect 320 5180 520 5200
rect 640 5180 840 5200
rect 960 5180 1160 5200
rect 0 5080 200 5100
rect 320 5080 520 5100
rect 640 5080 840 5100
rect 960 5080 1160 5100
rect 0 4955 200 4980
rect 0 4925 10 4955
rect 190 4925 200 4955
rect 0 4920 200 4925
rect 320 4955 520 4980
rect 320 4925 330 4955
rect 510 4925 520 4955
rect 320 4920 520 4925
rect 640 4955 840 4980
rect 640 4925 650 4955
rect 830 4925 840 4955
rect 640 4920 840 4925
rect 960 4955 1160 4980
rect 960 4925 970 4955
rect 1150 4925 1160 4955
rect 960 4920 1160 4925
rect 1440 5355 1640 5360
rect 1440 5325 1450 5355
rect 1630 5325 1640 5355
rect 1440 5300 1640 5325
rect 1760 5355 1960 5360
rect 1760 5325 1770 5355
rect 1950 5325 1960 5355
rect 1760 5300 1960 5325
rect 2080 5355 2280 5360
rect 2080 5325 2090 5355
rect 2270 5325 2280 5355
rect 2080 5300 2280 5325
rect 2400 5355 2600 5360
rect 2400 5325 2410 5355
rect 2590 5325 2600 5355
rect 2400 5300 2600 5325
rect 1440 5180 1640 5200
rect 1760 5180 1960 5200
rect 2080 5180 2280 5200
rect 2400 5180 2600 5200
rect 1440 5080 1640 5100
rect 1760 5080 1960 5100
rect 2080 5080 2280 5100
rect 2400 5080 2600 5100
rect 1440 4955 1640 4980
rect 1440 4925 1450 4955
rect 1630 4925 1640 4955
rect 1440 4920 1640 4925
rect 1760 4955 1960 4980
rect 1760 4925 1770 4955
rect 1950 4925 1960 4955
rect 1760 4920 1960 4925
rect 2080 4955 2280 4980
rect 2080 4925 2090 4955
rect 2270 4925 2280 4955
rect 2080 4920 2280 4925
rect 2400 4955 2600 4980
rect 2400 4925 2410 4955
rect 2590 4925 2600 4955
rect 2400 4920 2600 4925
rect 2880 5355 3080 5360
rect 2880 5325 2890 5355
rect 3070 5325 3080 5355
rect 2880 5300 3080 5325
rect 3200 5355 3400 5360
rect 3200 5325 3210 5355
rect 3390 5325 3400 5355
rect 3200 5300 3400 5325
rect 3520 5355 3720 5360
rect 3520 5325 3530 5355
rect 3710 5325 3720 5355
rect 3520 5300 3720 5325
rect 3840 5355 4040 5360
rect 3840 5325 3850 5355
rect 4030 5325 4040 5355
rect 3840 5300 4040 5325
rect 2880 5180 3080 5200
rect 3200 5180 3400 5200
rect 3520 5180 3720 5200
rect 3840 5180 4040 5200
rect 2880 5080 3080 5100
rect 3200 5080 3400 5100
rect 3520 5080 3720 5100
rect 3840 5080 4040 5100
rect 2880 4955 3080 4980
rect 2880 4925 2890 4955
rect 3070 4925 3080 4955
rect 2880 4920 3080 4925
rect 3200 4955 3400 4980
rect 3200 4925 3210 4955
rect 3390 4925 3400 4955
rect 3200 4920 3400 4925
rect 3520 4955 3720 4980
rect 3520 4925 3530 4955
rect 3710 4925 3720 4955
rect 3520 4920 3720 4925
rect 3840 4955 4040 4980
rect 3840 4925 3850 4955
rect 4030 4925 4040 4955
rect 3840 4920 4040 4925
rect 4320 5355 4520 5360
rect 4320 5325 4330 5355
rect 4510 5325 4520 5355
rect 4320 5300 4520 5325
rect 4320 5180 4520 5200
rect 4320 5080 4520 5100
rect 4320 4955 4520 4980
rect 4320 4925 4330 4955
rect 4510 4925 4520 4955
rect 4320 4920 4520 4925
rect -480 3995 -280 4000
rect -480 3965 -470 3995
rect -290 3965 -280 3995
rect -480 3940 -280 3965
rect -480 3820 -280 3840
rect 0 3995 200 4000
rect 0 3965 10 3995
rect 190 3965 200 3995
rect 0 3940 200 3965
rect 320 3995 520 4000
rect 320 3965 330 3995
rect 510 3965 520 3995
rect 320 3940 520 3965
rect 640 3995 840 4000
rect 640 3965 650 3995
rect 830 3965 840 3995
rect 640 3940 840 3965
rect 960 3995 1160 4000
rect 960 3965 970 3995
rect 1150 3965 1160 3995
rect 960 3940 1160 3965
rect 0 3820 200 3840
rect 320 3820 520 3840
rect 640 3820 840 3840
rect 960 3820 1160 3840
rect 1440 3995 1640 4000
rect 1440 3965 1450 3995
rect 1630 3965 1640 3995
rect 1440 3940 1640 3965
rect 1760 3995 1960 4000
rect 1760 3965 1770 3995
rect 1950 3965 1960 3995
rect 1760 3940 1960 3965
rect 2080 3995 2280 4000
rect 2080 3965 2090 3995
rect 2270 3965 2280 3995
rect 2080 3940 2280 3965
rect 2400 3995 2600 4000
rect 2400 3965 2410 3995
rect 2590 3965 2600 3995
rect 2400 3940 2600 3965
rect 1440 3820 1640 3840
rect 1760 3820 1960 3840
rect 2080 3820 2280 3840
rect 2400 3820 2600 3840
rect 2880 3995 3080 4000
rect 2880 3965 2890 3995
rect 3070 3965 3080 3995
rect 2880 3940 3080 3965
rect 3200 3995 3400 4000
rect 3200 3965 3210 3995
rect 3390 3965 3400 3995
rect 3200 3940 3400 3965
rect 3520 3995 3720 4000
rect 3520 3965 3530 3995
rect 3710 3965 3720 3995
rect 3520 3940 3720 3965
rect 3840 3995 4040 4000
rect 3840 3965 3850 3995
rect 4030 3965 4040 3995
rect 3840 3940 4040 3965
rect 2880 3820 3080 3840
rect 3200 3820 3400 3840
rect 3520 3820 3720 3840
rect 3840 3820 4040 3840
rect 4320 3995 4520 4000
rect 4320 3965 4330 3995
rect 4510 3965 4520 3995
rect 4320 3940 4520 3965
rect 4320 3820 4520 3840
rect -480 3435 -280 3440
rect -480 3405 -470 3435
rect -290 3405 -280 3435
rect -480 3380 -280 3405
rect -480 3260 -280 3280
rect -480 3160 -280 3180
rect -480 3035 -280 3060
rect -480 3005 -470 3035
rect -290 3005 -280 3035
rect -480 3000 -280 3005
rect 0 3435 200 3440
rect 0 3405 10 3435
rect 190 3405 200 3435
rect 0 3380 200 3405
rect 320 3435 520 3440
rect 320 3405 330 3435
rect 510 3405 520 3435
rect 320 3380 520 3405
rect 640 3435 840 3440
rect 640 3405 650 3435
rect 830 3405 840 3435
rect 640 3380 840 3405
rect 960 3435 1160 3440
rect 960 3405 970 3435
rect 1150 3405 1160 3435
rect 960 3380 1160 3405
rect 0 3260 200 3280
rect 320 3260 520 3280
rect 640 3260 840 3280
rect 960 3260 1160 3280
rect 0 3160 200 3180
rect 320 3160 520 3180
rect 640 3160 840 3180
rect 960 3160 1160 3180
rect 0 3035 200 3060
rect 0 3005 10 3035
rect 190 3005 200 3035
rect 0 3000 200 3005
rect 320 3035 520 3060
rect 320 3005 330 3035
rect 510 3005 520 3035
rect 320 3000 520 3005
rect 640 3035 840 3060
rect 640 3005 650 3035
rect 830 3005 840 3035
rect 640 3000 840 3005
rect 960 3035 1160 3060
rect 960 3005 970 3035
rect 1150 3005 1160 3035
rect 960 3000 1160 3005
rect 1440 3435 1640 3440
rect 1440 3405 1450 3435
rect 1630 3405 1640 3435
rect 1440 3380 1640 3405
rect 1760 3435 1960 3440
rect 1760 3405 1770 3435
rect 1950 3405 1960 3435
rect 1760 3380 1960 3405
rect 2080 3435 2280 3440
rect 2080 3405 2090 3435
rect 2270 3405 2280 3435
rect 2080 3380 2280 3405
rect 2400 3435 2600 3440
rect 2400 3405 2410 3435
rect 2590 3405 2600 3435
rect 2400 3380 2600 3405
rect 1440 3260 1640 3280
rect 1760 3260 1960 3280
rect 2080 3260 2280 3280
rect 2400 3260 2600 3280
rect 1440 3160 1640 3180
rect 1760 3160 1960 3180
rect 2080 3160 2280 3180
rect 2400 3160 2600 3180
rect 1440 3035 1640 3060
rect 1440 3005 1450 3035
rect 1630 3005 1640 3035
rect 1440 3000 1640 3005
rect 1760 3035 1960 3060
rect 1760 3005 1770 3035
rect 1950 3005 1960 3035
rect 1760 3000 1960 3005
rect 2080 3035 2280 3060
rect 2080 3005 2090 3035
rect 2270 3005 2280 3035
rect 2080 3000 2280 3005
rect 2400 3035 2600 3060
rect 2400 3005 2410 3035
rect 2590 3005 2600 3035
rect 2400 3000 2600 3005
rect 2880 3435 3080 3440
rect 2880 3405 2890 3435
rect 3070 3405 3080 3435
rect 2880 3380 3080 3405
rect 3200 3435 3400 3440
rect 3200 3405 3210 3435
rect 3390 3405 3400 3435
rect 3200 3380 3400 3405
rect 3520 3435 3720 3440
rect 3520 3405 3530 3435
rect 3710 3405 3720 3435
rect 3520 3380 3720 3405
rect 3840 3435 4040 3440
rect 3840 3405 3850 3435
rect 4030 3405 4040 3435
rect 3840 3380 4040 3405
rect 2880 3260 3080 3280
rect 3200 3260 3400 3280
rect 3520 3260 3720 3280
rect 3840 3260 4040 3280
rect 2880 3160 3080 3180
rect 3200 3160 3400 3180
rect 3520 3160 3720 3180
rect 3840 3160 4040 3180
rect 2880 3035 3080 3060
rect 2880 3005 2890 3035
rect 3070 3005 3080 3035
rect 2880 3000 3080 3005
rect 3200 3035 3400 3060
rect 3200 3005 3210 3035
rect 3390 3005 3400 3035
rect 3200 3000 3400 3005
rect 3520 3035 3720 3060
rect 3520 3005 3530 3035
rect 3710 3005 3720 3035
rect 3520 3000 3720 3005
rect 3840 3035 4040 3060
rect 3840 3005 3850 3035
rect 4030 3005 4040 3035
rect 3840 3000 4040 3005
rect 4320 3435 4520 3440
rect 4320 3405 4330 3435
rect 4510 3405 4520 3435
rect 4320 3380 4520 3405
rect 4320 3260 4520 3280
rect 4320 3160 4520 3180
rect 4320 3035 4520 3060
rect 4320 3005 4330 3035
rect 4510 3005 4520 3035
rect 4320 3000 4520 3005
rect -480 2075 -280 2080
rect -480 2045 -470 2075
rect -290 2045 -280 2075
rect -480 2020 -280 2045
rect -480 1900 -280 1920
rect 0 2075 200 2080
rect 0 2045 10 2075
rect 190 2045 200 2075
rect 0 2020 200 2045
rect 320 2075 520 2080
rect 320 2045 330 2075
rect 510 2045 520 2075
rect 320 2020 520 2045
rect 640 2075 840 2080
rect 640 2045 650 2075
rect 830 2045 840 2075
rect 640 2020 840 2045
rect 960 2075 1160 2080
rect 960 2045 970 2075
rect 1150 2045 1160 2075
rect 960 2020 1160 2045
rect 0 1900 200 1920
rect 320 1900 520 1920
rect 640 1900 840 1920
rect 960 1900 1160 1920
rect 1440 2075 1640 2080
rect 1440 2045 1450 2075
rect 1630 2045 1640 2075
rect 1440 2020 1640 2045
rect 1760 2075 1960 2080
rect 1760 2045 1770 2075
rect 1950 2045 1960 2075
rect 1760 2020 1960 2045
rect 2080 2075 2280 2080
rect 2080 2045 2090 2075
rect 2270 2045 2280 2075
rect 2080 2020 2280 2045
rect 2400 2075 2600 2080
rect 2400 2045 2410 2075
rect 2590 2045 2600 2075
rect 2400 2020 2600 2045
rect 1440 1900 1640 1920
rect 1760 1900 1960 1920
rect 2080 1900 2280 1920
rect 2400 1900 2600 1920
rect 2880 2075 3080 2080
rect 2880 2045 2890 2075
rect 3070 2045 3080 2075
rect 2880 2020 3080 2045
rect 3200 2075 3400 2080
rect 3200 2045 3210 2075
rect 3390 2045 3400 2075
rect 3200 2020 3400 2045
rect 3520 2075 3720 2080
rect 3520 2045 3530 2075
rect 3710 2045 3720 2075
rect 3520 2020 3720 2045
rect 3840 2075 4040 2080
rect 3840 2045 3850 2075
rect 4030 2045 4040 2075
rect 3840 2020 4040 2045
rect 2880 1900 3080 1920
rect 3200 1900 3400 1920
rect 3520 1900 3720 1920
rect 3840 1900 4040 1920
rect 4320 2075 4520 2080
rect 4320 2045 4330 2075
rect 4510 2045 4520 2075
rect 4320 2020 4520 2045
rect 4320 1900 4520 1920
rect -480 1515 -280 1520
rect -480 1485 -470 1515
rect -290 1485 -280 1515
rect -480 1460 -280 1485
rect -480 1340 -280 1360
rect -480 1240 -280 1260
rect -480 1115 -280 1140
rect -480 1085 -470 1115
rect -290 1085 -280 1115
rect -480 1080 -280 1085
rect 0 1515 200 1520
rect 0 1485 10 1515
rect 190 1485 200 1515
rect 0 1460 200 1485
rect 320 1515 520 1520
rect 320 1485 330 1515
rect 510 1485 520 1515
rect 320 1460 520 1485
rect 640 1515 840 1520
rect 640 1485 650 1515
rect 830 1485 840 1515
rect 640 1460 840 1485
rect 960 1515 1160 1520
rect 960 1485 970 1515
rect 1150 1485 1160 1515
rect 960 1460 1160 1485
rect 0 1340 200 1360
rect 320 1340 520 1360
rect 640 1340 840 1360
rect 960 1340 1160 1360
rect 0 1240 200 1260
rect 320 1240 520 1260
rect 640 1240 840 1260
rect 960 1240 1160 1260
rect 0 1115 200 1140
rect 0 1085 10 1115
rect 190 1085 200 1115
rect 0 1080 200 1085
rect 320 1115 520 1140
rect 320 1085 330 1115
rect 510 1085 520 1115
rect 320 1080 520 1085
rect 640 1115 840 1140
rect 640 1085 650 1115
rect 830 1085 840 1115
rect 640 1080 840 1085
rect 960 1115 1160 1140
rect 960 1085 970 1115
rect 1150 1085 1160 1115
rect 960 1080 1160 1085
rect 1440 1515 1640 1520
rect 1440 1485 1450 1515
rect 1630 1485 1640 1515
rect 1440 1460 1640 1485
rect 1760 1515 1960 1520
rect 1760 1485 1770 1515
rect 1950 1485 1960 1515
rect 1760 1460 1960 1485
rect 2080 1515 2280 1520
rect 2080 1485 2090 1515
rect 2270 1485 2280 1515
rect 2080 1460 2280 1485
rect 2400 1515 2600 1520
rect 2400 1485 2410 1515
rect 2590 1485 2600 1515
rect 2400 1460 2600 1485
rect 1440 1340 1640 1360
rect 1760 1340 1960 1360
rect 2080 1340 2280 1360
rect 2400 1340 2600 1360
rect 1440 1240 1640 1260
rect 1760 1240 1960 1260
rect 2080 1240 2280 1260
rect 2400 1240 2600 1260
rect 1440 1115 1640 1140
rect 1440 1085 1450 1115
rect 1630 1085 1640 1115
rect 1440 1080 1640 1085
rect 1760 1115 1960 1140
rect 1760 1085 1770 1115
rect 1950 1085 1960 1115
rect 1760 1080 1960 1085
rect 2080 1115 2280 1140
rect 2080 1085 2090 1115
rect 2270 1085 2280 1115
rect 2080 1080 2280 1085
rect 2400 1115 2600 1140
rect 2400 1085 2410 1115
rect 2590 1085 2600 1115
rect 2400 1080 2600 1085
rect 2880 1515 3080 1520
rect 2880 1485 2890 1515
rect 3070 1485 3080 1515
rect 2880 1460 3080 1485
rect 3200 1515 3400 1520
rect 3200 1485 3210 1515
rect 3390 1485 3400 1515
rect 3200 1460 3400 1485
rect 3520 1515 3720 1520
rect 3520 1485 3530 1515
rect 3710 1485 3720 1515
rect 3520 1460 3720 1485
rect 3840 1515 4040 1520
rect 3840 1485 3850 1515
rect 4030 1485 4040 1515
rect 3840 1460 4040 1485
rect 2880 1340 3080 1360
rect 3200 1340 3400 1360
rect 3520 1340 3720 1360
rect 3840 1340 4040 1360
rect 2880 1240 3080 1260
rect 3200 1240 3400 1260
rect 3520 1240 3720 1260
rect 3840 1240 4040 1260
rect 2880 1115 3080 1140
rect 2880 1085 2890 1115
rect 3070 1085 3080 1115
rect 2880 1080 3080 1085
rect 3200 1115 3400 1140
rect 3200 1085 3210 1115
rect 3390 1085 3400 1115
rect 3200 1080 3400 1085
rect 3520 1115 3720 1140
rect 3520 1085 3530 1115
rect 3710 1085 3720 1115
rect 3520 1080 3720 1085
rect 3840 1115 4040 1140
rect 3840 1085 3850 1115
rect 4030 1085 4040 1115
rect 3840 1080 4040 1085
rect 4320 1515 4520 1520
rect 4320 1485 4330 1515
rect 4510 1485 4520 1515
rect 4320 1460 4520 1485
rect 4320 1340 4520 1360
rect 4320 1240 4520 1260
rect 4320 1115 4520 1140
rect 4320 1085 4330 1115
rect 4510 1085 4520 1115
rect 4320 1080 4520 1085
rect -480 155 -280 160
rect -480 125 -470 155
rect -290 125 -280 155
rect -480 100 -280 125
rect -480 -20 -280 0
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 100 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 100 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 100 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 100 1160 125
rect 0 -20 200 0
rect 320 -20 520 0
rect 640 -20 840 0
rect 960 -20 1160 0
rect 1440 155 1640 160
rect 1440 125 1450 155
rect 1630 125 1640 155
rect 1440 100 1640 125
rect 1760 155 1960 160
rect 1760 125 1770 155
rect 1950 125 1960 155
rect 1760 100 1960 125
rect 2080 155 2280 160
rect 2080 125 2090 155
rect 2270 125 2280 155
rect 2080 100 2280 125
rect 2400 155 2600 160
rect 2400 125 2410 155
rect 2590 125 2600 155
rect 2400 100 2600 125
rect 1440 -20 1640 0
rect 1760 -20 1960 0
rect 2080 -20 2280 0
rect 2400 -20 2600 0
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 100 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 100 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 100 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 100 4040 125
rect 2880 -20 3080 0
rect 3200 -20 3400 0
rect 3520 -20 3720 0
rect 3840 -20 4040 0
rect 4320 155 4520 160
rect 4320 125 4330 155
rect 4510 125 4520 155
rect 4320 100 4520 125
rect 4320 -20 4520 0
<< polycont >>
rect -470 5325 -290 5355
rect -470 4925 -290 4955
rect 10 5325 190 5355
rect 330 5325 510 5355
rect 650 5325 830 5355
rect 970 5325 1150 5355
rect 10 4925 190 4955
rect 330 4925 510 4955
rect 650 4925 830 4955
rect 970 4925 1150 4955
rect 1450 5325 1630 5355
rect 1770 5325 1950 5355
rect 2090 5325 2270 5355
rect 2410 5325 2590 5355
rect 1450 4925 1630 4955
rect 1770 4925 1950 4955
rect 2090 4925 2270 4955
rect 2410 4925 2590 4955
rect 2890 5325 3070 5355
rect 3210 5325 3390 5355
rect 3530 5325 3710 5355
rect 3850 5325 4030 5355
rect 2890 4925 3070 4955
rect 3210 4925 3390 4955
rect 3530 4925 3710 4955
rect 3850 4925 4030 4955
rect 4330 5325 4510 5355
rect 4330 4925 4510 4955
rect -470 3965 -290 3995
rect 10 3965 190 3995
rect 330 3965 510 3995
rect 650 3965 830 3995
rect 970 3965 1150 3995
rect 1450 3965 1630 3995
rect 1770 3965 1950 3995
rect 2090 3965 2270 3995
rect 2410 3965 2590 3995
rect 2890 3965 3070 3995
rect 3210 3965 3390 3995
rect 3530 3965 3710 3995
rect 3850 3965 4030 3995
rect 4330 3965 4510 3995
rect -470 3405 -290 3435
rect -470 3005 -290 3035
rect 10 3405 190 3435
rect 330 3405 510 3435
rect 650 3405 830 3435
rect 970 3405 1150 3435
rect 10 3005 190 3035
rect 330 3005 510 3035
rect 650 3005 830 3035
rect 970 3005 1150 3035
rect 1450 3405 1630 3435
rect 1770 3405 1950 3435
rect 2090 3405 2270 3435
rect 2410 3405 2590 3435
rect 1450 3005 1630 3035
rect 1770 3005 1950 3035
rect 2090 3005 2270 3035
rect 2410 3005 2590 3035
rect 2890 3405 3070 3435
rect 3210 3405 3390 3435
rect 3530 3405 3710 3435
rect 3850 3405 4030 3435
rect 2890 3005 3070 3035
rect 3210 3005 3390 3035
rect 3530 3005 3710 3035
rect 3850 3005 4030 3035
rect 4330 3405 4510 3435
rect 4330 3005 4510 3035
rect -470 2045 -290 2075
rect 10 2045 190 2075
rect 330 2045 510 2075
rect 650 2045 830 2075
rect 970 2045 1150 2075
rect 1450 2045 1630 2075
rect 1770 2045 1950 2075
rect 2090 2045 2270 2075
rect 2410 2045 2590 2075
rect 2890 2045 3070 2075
rect 3210 2045 3390 2075
rect 3530 2045 3710 2075
rect 3850 2045 4030 2075
rect 4330 2045 4510 2075
rect -470 1485 -290 1515
rect -470 1085 -290 1115
rect 10 1485 190 1515
rect 330 1485 510 1515
rect 650 1485 830 1515
rect 970 1485 1150 1515
rect 10 1085 190 1115
rect 330 1085 510 1115
rect 650 1085 830 1115
rect 970 1085 1150 1115
rect 1450 1485 1630 1515
rect 1770 1485 1950 1515
rect 2090 1485 2270 1515
rect 2410 1485 2590 1515
rect 1450 1085 1630 1115
rect 1770 1085 1950 1115
rect 2090 1085 2270 1115
rect 2410 1085 2590 1115
rect 2890 1485 3070 1515
rect 3210 1485 3390 1515
rect 3530 1485 3710 1515
rect 3850 1485 4030 1515
rect 2890 1085 3070 1115
rect 3210 1085 3390 1115
rect 3530 1085 3710 1115
rect 3850 1085 4030 1115
rect 4330 1485 4510 1515
rect 4330 1085 4510 1115
rect -470 125 -290 155
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect 1450 125 1630 155
rect 1770 125 1950 155
rect 2090 125 2270 155
rect 2410 125 2590 155
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3850 125 4030 155
rect 4330 125 4510 155
<< locali >>
rect -800 5560 -680 5600
rect 4760 5560 4840 5600
rect -640 5400 -560 5440
rect -200 5400 -80 5440
rect 1240 5400 1360 5440
rect 2680 5400 2800 5440
rect 4120 5400 4240 5440
rect 4600 5400 4680 5440
rect -560 5290 -520 5400
rect -480 5355 -200 5360
rect -480 5325 -470 5355
rect -290 5325 -200 5355
rect -480 5320 -200 5325
rect -560 5210 -555 5290
rect -525 5210 -520 5290
rect -560 5070 -520 5210
rect -560 4990 -555 5070
rect -525 4990 -520 5070
rect -560 4880 -520 4990
rect -240 5290 -200 5320
rect -240 5210 -235 5290
rect -205 5210 -200 5290
rect -240 5070 -200 5210
rect -240 4990 -235 5070
rect -205 4990 -200 5070
rect -240 4960 -200 4990
rect -480 4955 -200 4960
rect -480 4925 -470 4955
rect -290 4925 -200 4955
rect -480 4920 -200 4925
rect 0 5355 200 5360
rect 0 5325 10 5355
rect 190 5325 200 5355
rect 0 5320 200 5325
rect 320 5355 520 5360
rect 320 5325 330 5355
rect 510 5325 520 5355
rect 320 5320 520 5325
rect 640 5355 840 5360
rect 640 5325 650 5355
rect 830 5325 840 5355
rect 640 5320 840 5325
rect 960 5355 1160 5360
rect 960 5325 970 5355
rect 1150 5325 1160 5355
rect 960 5320 1160 5325
rect -80 5290 -40 5300
rect -80 5210 -75 5290
rect -45 5210 -40 5290
rect -80 5200 -40 5210
rect 240 5290 280 5300
rect 240 5210 245 5290
rect 275 5210 280 5290
rect 240 5200 280 5210
rect 560 5290 600 5300
rect 560 5210 565 5290
rect 595 5210 600 5290
rect 560 5200 600 5210
rect 880 5290 920 5300
rect 880 5210 885 5290
rect 915 5210 920 5290
rect 880 5200 920 5210
rect 1200 5290 1240 5300
rect 1200 5210 1205 5290
rect 1235 5210 1240 5290
rect 1200 5200 1240 5210
rect -80 5070 -40 5080
rect -80 4990 -75 5070
rect -45 4990 -40 5070
rect -80 4980 -40 4990
rect 240 5070 280 5080
rect 240 4990 245 5070
rect 275 4990 280 5070
rect 240 4980 280 4990
rect 560 5070 600 5080
rect 560 4990 565 5070
rect 595 4990 600 5070
rect 560 4980 600 4990
rect 880 5070 920 5080
rect 880 4990 885 5070
rect 915 4990 920 5070
rect 880 4980 920 4990
rect 1200 5070 1240 5080
rect 1200 4990 1205 5070
rect 1235 4990 1240 5070
rect 1200 4980 1240 4990
rect 0 4955 200 4960
rect 0 4925 10 4955
rect 190 4925 200 4955
rect 0 4920 200 4925
rect 320 4955 520 4960
rect 320 4925 330 4955
rect 510 4925 520 4955
rect 320 4920 520 4925
rect 640 4955 840 4960
rect 640 4925 650 4955
rect 830 4925 840 4955
rect 640 4920 840 4925
rect 960 4955 1160 4960
rect 960 4925 970 4955
rect 1150 4925 1160 4955
rect 960 4920 1160 4925
rect 1440 5355 1640 5360
rect 1440 5325 1450 5355
rect 1630 5325 1640 5355
rect 1440 5320 1640 5325
rect 1760 5355 1960 5360
rect 1760 5325 1770 5355
rect 1950 5325 1960 5355
rect 1760 5320 1960 5325
rect 2080 5355 2280 5360
rect 2080 5325 2090 5355
rect 2270 5325 2280 5355
rect 2080 5320 2280 5325
rect 2400 5355 2600 5360
rect 2400 5325 2410 5355
rect 2590 5325 2600 5355
rect 2400 5320 2600 5325
rect 1360 5290 1400 5300
rect 1360 5210 1365 5290
rect 1395 5210 1400 5290
rect 1360 5200 1400 5210
rect 1680 5290 1720 5300
rect 1680 5210 1685 5290
rect 1715 5210 1720 5290
rect 1680 5200 1720 5210
rect 2000 5290 2040 5300
rect 2000 5210 2005 5290
rect 2035 5210 2040 5290
rect 2000 5200 2040 5210
rect 2320 5290 2360 5300
rect 2320 5210 2325 5290
rect 2355 5210 2360 5290
rect 2320 5200 2360 5210
rect 2640 5290 2680 5300
rect 2640 5210 2645 5290
rect 2675 5210 2680 5290
rect 2640 5200 2680 5210
rect 1360 5070 1400 5080
rect 1360 4990 1365 5070
rect 1395 4990 1400 5070
rect 1360 4980 1400 4990
rect 1680 5070 1720 5080
rect 1680 4990 1685 5070
rect 1715 4990 1720 5070
rect 1680 4980 1720 4990
rect 2000 5070 2040 5080
rect 2000 4990 2005 5070
rect 2035 4990 2040 5070
rect 2000 4980 2040 4990
rect 2320 5070 2360 5080
rect 2320 4990 2325 5070
rect 2355 4990 2360 5070
rect 2320 4980 2360 4990
rect 2640 5070 2680 5080
rect 2640 4990 2645 5070
rect 2675 4990 2680 5070
rect 2640 4980 2680 4990
rect 1440 4955 1640 4960
rect 1440 4925 1450 4955
rect 1630 4925 1640 4955
rect 1440 4920 1640 4925
rect 1760 4955 1960 4960
rect 1760 4925 1770 4955
rect 1950 4925 1960 4955
rect 1760 4920 1960 4925
rect 2080 4955 2280 4960
rect 2080 4925 2090 4955
rect 2270 4925 2280 4955
rect 2080 4920 2280 4925
rect 2400 4955 2600 4960
rect 2400 4925 2410 4955
rect 2590 4925 2600 4955
rect 2400 4920 2600 4925
rect 2880 5355 3080 5360
rect 2880 5325 2890 5355
rect 3070 5325 3080 5355
rect 2880 5320 3080 5325
rect 3200 5355 3400 5360
rect 3200 5325 3210 5355
rect 3390 5325 3400 5355
rect 3200 5320 3400 5325
rect 3520 5355 3720 5360
rect 3520 5325 3530 5355
rect 3710 5325 3720 5355
rect 3520 5320 3720 5325
rect 3840 5355 4040 5360
rect 3840 5325 3850 5355
rect 4030 5325 4040 5355
rect 3840 5320 4040 5325
rect 2800 5290 2840 5300
rect 2800 5210 2805 5290
rect 2835 5210 2840 5290
rect 2800 5200 2840 5210
rect 3120 5290 3160 5300
rect 3120 5210 3125 5290
rect 3155 5210 3160 5290
rect 3120 5200 3160 5210
rect 3440 5290 3480 5300
rect 3440 5210 3445 5290
rect 3475 5210 3480 5290
rect 3440 5200 3480 5210
rect 3760 5290 3800 5300
rect 3760 5210 3765 5290
rect 3795 5210 3800 5290
rect 3760 5200 3800 5210
rect 4080 5290 4120 5300
rect 4080 5210 4085 5290
rect 4115 5210 4120 5290
rect 4080 5200 4120 5210
rect 2800 5070 2840 5080
rect 2800 4990 2805 5070
rect 2835 4990 2840 5070
rect 2800 4980 2840 4990
rect 3120 5070 3160 5080
rect 3120 4990 3125 5070
rect 3155 4990 3160 5070
rect 3120 4980 3160 4990
rect 3440 5070 3480 5080
rect 3440 4990 3445 5070
rect 3475 4990 3480 5070
rect 3440 4980 3480 4990
rect 3760 5070 3800 5080
rect 3760 4990 3765 5070
rect 3795 4990 3800 5070
rect 3760 4980 3800 4990
rect 4080 5070 4120 5080
rect 4080 4990 4085 5070
rect 4115 4990 4120 5070
rect 4080 4980 4120 4990
rect 2880 4955 3080 4960
rect 2880 4925 2890 4955
rect 3070 4925 3080 4955
rect 2880 4920 3080 4925
rect 3200 4955 3400 4960
rect 3200 4925 3210 4955
rect 3390 4925 3400 4955
rect 3200 4920 3400 4925
rect 3520 4955 3720 4960
rect 3520 4925 3530 4955
rect 3710 4925 3720 4955
rect 3520 4920 3720 4925
rect 3840 4955 4040 4960
rect 3840 4925 3850 4955
rect 4030 4925 4040 4955
rect 3840 4920 4040 4925
rect 4240 5355 4520 5360
rect 4240 5325 4330 5355
rect 4510 5325 4520 5355
rect 4240 5320 4520 5325
rect 4240 5290 4280 5320
rect 4240 5210 4245 5290
rect 4275 5210 4280 5290
rect 4240 5070 4280 5210
rect 4240 4990 4245 5070
rect 4275 4990 4280 5070
rect 4240 4960 4280 4990
rect 4560 5290 4600 5400
rect 4560 5210 4565 5290
rect 4595 5210 4600 5290
rect 4560 5070 4600 5210
rect 4560 4990 4565 5070
rect 4595 4990 4600 5070
rect 4240 4955 4520 4960
rect 4240 4925 4330 4955
rect 4510 4925 4520 4955
rect 4240 4920 4520 4925
rect 4560 4880 4600 4990
rect -640 4840 -560 4880
rect -200 4840 -80 4880
rect 1240 4840 1360 4880
rect 2680 4840 2800 4880
rect 4120 4840 4240 4880
rect 4600 4840 4680 4880
rect -800 4680 -680 4720
rect 4760 4680 4840 4720
rect -800 4040 -560 4080
rect -200 4040 -80 4080
rect 1240 4040 1360 4080
rect 2680 4040 2800 4080
rect 4120 4040 4240 4080
rect 4600 4040 4840 4080
rect -560 3930 -520 4040
rect -480 3995 -200 4000
rect -480 3965 -470 3995
rect -290 3965 -200 3995
rect -480 3960 -200 3965
rect -560 3850 -555 3930
rect -525 3850 -520 3930
rect -560 3760 -520 3850
rect -240 3930 -200 3960
rect -240 3850 -235 3930
rect -205 3850 -200 3930
rect -240 3840 -200 3850
rect 0 3995 200 4000
rect 0 3965 10 3995
rect 190 3965 200 3995
rect 0 3960 200 3965
rect 320 3995 520 4000
rect 320 3965 330 3995
rect 510 3965 520 3995
rect 320 3960 520 3965
rect 640 3995 840 4000
rect 640 3965 650 3995
rect 830 3965 840 3995
rect 640 3960 840 3965
rect 960 3995 1160 4000
rect 960 3965 970 3995
rect 1150 3965 1160 3995
rect 960 3960 1160 3965
rect -80 3930 -40 3940
rect -80 3850 -75 3930
rect -45 3850 -40 3930
rect -80 3840 -40 3850
rect 240 3930 280 3940
rect 240 3850 245 3930
rect 275 3850 280 3930
rect 240 3840 280 3850
rect 560 3930 600 3940
rect 560 3850 565 3930
rect 595 3850 600 3930
rect 560 3840 600 3850
rect 880 3930 920 3940
rect 880 3850 885 3930
rect 915 3850 920 3930
rect 880 3840 920 3850
rect 1200 3930 1240 3940
rect 1200 3850 1205 3930
rect 1235 3850 1240 3930
rect 1200 3840 1240 3850
rect 1440 3995 1640 4000
rect 1440 3965 1450 3995
rect 1630 3965 1640 3995
rect 1440 3960 1640 3965
rect 1760 3995 1960 4000
rect 1760 3965 1770 3995
rect 1950 3965 1960 3995
rect 1760 3960 1960 3965
rect 2080 3995 2280 4000
rect 2080 3965 2090 3995
rect 2270 3965 2280 3995
rect 2080 3960 2280 3965
rect 2400 3995 2600 4000
rect 2400 3965 2410 3995
rect 2590 3965 2600 3995
rect 2400 3960 2600 3965
rect 1360 3930 1400 3940
rect 1360 3850 1365 3930
rect 1395 3850 1400 3930
rect 1360 3840 1400 3850
rect 1680 3930 1720 3940
rect 1680 3850 1685 3930
rect 1715 3850 1720 3930
rect 1680 3840 1720 3850
rect 2000 3930 2040 3940
rect 2000 3850 2005 3930
rect 2035 3850 2040 3930
rect 2000 3840 2040 3850
rect 2320 3930 2360 3940
rect 2320 3850 2325 3930
rect 2355 3850 2360 3930
rect 2320 3840 2360 3850
rect 2640 3930 2680 3940
rect 2640 3850 2645 3930
rect 2675 3850 2680 3930
rect 2640 3840 2680 3850
rect 2880 3995 3080 4000
rect 2880 3965 2890 3995
rect 3070 3965 3080 3995
rect 2880 3960 3080 3965
rect 3200 3995 3400 4000
rect 3200 3965 3210 3995
rect 3390 3965 3400 3995
rect 3200 3960 3400 3965
rect 3520 3995 3720 4000
rect 3520 3965 3530 3995
rect 3710 3965 3720 3995
rect 3520 3960 3720 3965
rect 3840 3995 4040 4000
rect 3840 3965 3850 3995
rect 4030 3965 4040 3995
rect 3840 3960 4040 3965
rect 2800 3930 2840 3940
rect 2800 3850 2805 3930
rect 2835 3850 2840 3930
rect 2800 3840 2840 3850
rect 3120 3930 3160 3940
rect 3120 3850 3125 3930
rect 3155 3850 3160 3930
rect 3120 3840 3160 3850
rect 3440 3930 3480 3940
rect 3440 3850 3445 3930
rect 3475 3850 3480 3930
rect 3440 3840 3480 3850
rect 3760 3930 3800 3940
rect 3760 3850 3765 3930
rect 3795 3850 3800 3930
rect 3760 3840 3800 3850
rect 4080 3930 4120 3940
rect 4080 3850 4085 3930
rect 4115 3850 4120 3930
rect 4080 3840 4120 3850
rect 4240 3995 4520 4000
rect 4240 3965 4330 3995
rect 4510 3965 4520 3995
rect 4240 3960 4520 3965
rect 4240 3930 4280 3960
rect 4240 3850 4245 3930
rect 4275 3850 4280 3930
rect 4240 3840 4280 3850
rect 4560 3930 4600 4040
rect 4560 3850 4565 3930
rect 4595 3850 4600 3930
rect 4560 3760 4600 3850
rect -800 3720 -560 3760
rect -200 3720 -80 3760
rect 1240 3720 1360 3760
rect 2680 3720 2800 3760
rect 4120 3720 4240 3760
rect 4600 3720 4840 3760
rect -800 3680 -760 3720
rect 4800 3680 4840 3720
rect -800 3640 -680 3680
rect 4760 3640 4840 3680
rect -640 3480 -560 3520
rect -200 3480 -80 3520
rect 1240 3480 1360 3520
rect 2680 3480 2800 3520
rect 4120 3480 4240 3520
rect 4600 3480 4680 3520
rect -560 3370 -520 3480
rect -480 3435 -200 3440
rect -480 3405 -470 3435
rect -290 3405 -200 3435
rect -480 3400 -200 3405
rect -560 3290 -555 3370
rect -525 3290 -520 3370
rect -560 3150 -520 3290
rect -560 3070 -555 3150
rect -525 3070 -520 3150
rect -560 2960 -520 3070
rect -240 3370 -200 3400
rect -240 3290 -235 3370
rect -205 3290 -200 3370
rect -240 3150 -200 3290
rect -240 3070 -235 3150
rect -205 3070 -200 3150
rect -240 3040 -200 3070
rect -480 3035 -200 3040
rect -480 3005 -470 3035
rect -290 3005 -200 3035
rect -480 3000 -200 3005
rect 0 3435 200 3440
rect 0 3405 10 3435
rect 190 3405 200 3435
rect 0 3400 200 3405
rect 320 3435 520 3440
rect 320 3405 330 3435
rect 510 3405 520 3435
rect 320 3400 520 3405
rect 640 3435 840 3440
rect 640 3405 650 3435
rect 830 3405 840 3435
rect 640 3400 840 3405
rect 960 3435 1160 3440
rect 960 3405 970 3435
rect 1150 3405 1160 3435
rect 960 3400 1160 3405
rect -80 3370 -40 3380
rect -80 3290 -75 3370
rect -45 3290 -40 3370
rect -80 3280 -40 3290
rect 240 3370 280 3380
rect 240 3290 245 3370
rect 275 3290 280 3370
rect 240 3280 280 3290
rect 560 3370 600 3380
rect 560 3290 565 3370
rect 595 3290 600 3370
rect 560 3280 600 3290
rect 880 3370 920 3380
rect 880 3290 885 3370
rect 915 3290 920 3370
rect 880 3280 920 3290
rect 1200 3370 1240 3380
rect 1200 3290 1205 3370
rect 1235 3290 1240 3370
rect 1200 3280 1240 3290
rect -80 3150 -40 3160
rect -80 3070 -75 3150
rect -45 3070 -40 3150
rect -80 3060 -40 3070
rect 240 3150 280 3160
rect 240 3070 245 3150
rect 275 3070 280 3150
rect 240 3060 280 3070
rect 560 3150 600 3160
rect 560 3070 565 3150
rect 595 3070 600 3150
rect 560 3060 600 3070
rect 880 3150 920 3160
rect 880 3070 885 3150
rect 915 3070 920 3150
rect 880 3060 920 3070
rect 1200 3150 1240 3160
rect 1200 3070 1205 3150
rect 1235 3070 1240 3150
rect 1200 3060 1240 3070
rect 0 3035 200 3040
rect 0 3005 10 3035
rect 190 3005 200 3035
rect 0 3000 200 3005
rect 320 3035 520 3040
rect 320 3005 330 3035
rect 510 3005 520 3035
rect 320 3000 520 3005
rect 640 3035 840 3040
rect 640 3005 650 3035
rect 830 3005 840 3035
rect 640 3000 840 3005
rect 960 3035 1160 3040
rect 960 3005 970 3035
rect 1150 3005 1160 3035
rect 960 3000 1160 3005
rect 1440 3435 1640 3440
rect 1440 3405 1450 3435
rect 1630 3405 1640 3435
rect 1440 3400 1640 3405
rect 1760 3435 1960 3440
rect 1760 3405 1770 3435
rect 1950 3405 1960 3435
rect 1760 3400 1960 3405
rect 2080 3435 2280 3440
rect 2080 3405 2090 3435
rect 2270 3405 2280 3435
rect 2080 3400 2280 3405
rect 2400 3435 2600 3440
rect 2400 3405 2410 3435
rect 2590 3405 2600 3435
rect 2400 3400 2600 3405
rect 1360 3370 1400 3380
rect 1360 3290 1365 3370
rect 1395 3290 1400 3370
rect 1360 3280 1400 3290
rect 1680 3370 1720 3380
rect 1680 3290 1685 3370
rect 1715 3290 1720 3370
rect 1680 3280 1720 3290
rect 2000 3370 2040 3380
rect 2000 3290 2005 3370
rect 2035 3290 2040 3370
rect 2000 3280 2040 3290
rect 2320 3370 2360 3380
rect 2320 3290 2325 3370
rect 2355 3290 2360 3370
rect 2320 3280 2360 3290
rect 2640 3370 2680 3380
rect 2640 3290 2645 3370
rect 2675 3290 2680 3370
rect 2640 3280 2680 3290
rect 1360 3150 1400 3160
rect 1360 3070 1365 3150
rect 1395 3070 1400 3150
rect 1360 3060 1400 3070
rect 1680 3150 1720 3160
rect 1680 3070 1685 3150
rect 1715 3070 1720 3150
rect 1680 3060 1720 3070
rect 2000 3150 2040 3160
rect 2000 3070 2005 3150
rect 2035 3070 2040 3150
rect 2000 3060 2040 3070
rect 2320 3150 2360 3160
rect 2320 3070 2325 3150
rect 2355 3070 2360 3150
rect 2320 3060 2360 3070
rect 2640 3150 2680 3160
rect 2640 3070 2645 3150
rect 2675 3070 2680 3150
rect 2640 3060 2680 3070
rect 1440 3035 1640 3040
rect 1440 3005 1450 3035
rect 1630 3005 1640 3035
rect 1440 3000 1640 3005
rect 1760 3035 1960 3040
rect 1760 3005 1770 3035
rect 1950 3005 1960 3035
rect 1760 3000 1960 3005
rect 2080 3035 2280 3040
rect 2080 3005 2090 3035
rect 2270 3005 2280 3035
rect 2080 3000 2280 3005
rect 2400 3035 2600 3040
rect 2400 3005 2410 3035
rect 2590 3005 2600 3035
rect 2400 3000 2600 3005
rect 2880 3435 4120 3440
rect 2880 3405 2890 3435
rect 3070 3405 3210 3435
rect 3390 3405 3530 3435
rect 3710 3405 3850 3435
rect 4030 3405 4120 3435
rect 2880 3400 4120 3405
rect 2800 3370 2840 3380
rect 2800 3290 2805 3370
rect 2835 3290 2840 3370
rect 2800 3280 2840 3290
rect 3120 3370 3160 3380
rect 3120 3290 3125 3370
rect 3155 3290 3160 3370
rect 3120 3280 3160 3290
rect 3440 3370 3480 3380
rect 3440 3290 3445 3370
rect 3475 3290 3480 3370
rect 3440 3280 3480 3290
rect 3760 3370 3800 3380
rect 3760 3290 3765 3370
rect 3795 3290 3800 3370
rect 3760 3280 3800 3290
rect 4080 3370 4120 3400
rect 4080 3290 4085 3370
rect 4115 3290 4120 3370
rect 4080 3280 4120 3290
rect 2800 3150 2840 3160
rect 2800 3070 2805 3150
rect 2835 3070 2840 3150
rect 2800 3060 2840 3070
rect 3120 3150 3160 3160
rect 3120 3070 3125 3150
rect 3155 3070 3160 3150
rect 3120 3060 3160 3070
rect 3440 3150 3480 3160
rect 3440 3070 3445 3150
rect 3475 3070 3480 3150
rect 3440 3060 3480 3070
rect 3760 3150 3800 3160
rect 3760 3070 3765 3150
rect 3795 3070 3800 3150
rect 3760 3060 3800 3070
rect 4080 3150 4120 3160
rect 4080 3070 4085 3150
rect 4115 3070 4120 3150
rect 4080 3060 4120 3070
rect 2880 3035 3080 3040
rect 2880 3005 2890 3035
rect 3070 3005 3080 3035
rect 2880 3000 3080 3005
rect 3200 3035 3400 3040
rect 3200 3005 3210 3035
rect 3390 3005 3400 3035
rect 3200 3000 3400 3005
rect 3520 3035 3720 3040
rect 3520 3005 3530 3035
rect 3710 3005 3720 3035
rect 3520 3000 3720 3005
rect 3840 3035 4040 3040
rect 3840 3005 3850 3035
rect 4030 3005 4040 3035
rect 3840 3000 4040 3005
rect 4240 3435 4520 3440
rect 4240 3405 4330 3435
rect 4510 3405 4520 3435
rect 4240 3400 4520 3405
rect 4240 3370 4280 3400
rect 4240 3290 4245 3370
rect 4275 3290 4280 3370
rect 4240 3150 4280 3290
rect 4240 3070 4245 3150
rect 4275 3070 4280 3150
rect 4240 3040 4280 3070
rect 4560 3370 4600 3480
rect 4560 3290 4565 3370
rect 4595 3290 4600 3370
rect 4560 3150 4600 3290
rect 4560 3070 4565 3150
rect 4595 3070 4600 3150
rect 4240 3035 4520 3040
rect 4240 3005 4330 3035
rect 4510 3005 4520 3035
rect 4240 3000 4520 3005
rect 4560 2960 4600 3070
rect -640 2920 -560 2960
rect -200 2920 -80 2960
rect 1240 2920 1360 2960
rect 2680 2920 2800 2960
rect 4120 2920 4240 2960
rect 4600 2920 4680 2960
rect -800 2760 -680 2800
rect 4760 2760 4840 2800
rect -800 2120 -560 2160
rect -200 2120 -80 2160
rect 1240 2120 1360 2160
rect 2680 2120 2800 2160
rect 4120 2120 4240 2160
rect 4600 2120 4840 2160
rect -560 2010 -520 2120
rect -480 2075 -200 2080
rect -480 2045 -470 2075
rect -290 2045 -200 2075
rect -480 2040 -200 2045
rect -560 1930 -555 2010
rect -525 1930 -520 2010
rect -560 1840 -520 1930
rect -240 2010 -200 2040
rect -240 1930 -235 2010
rect -205 1930 -200 2010
rect -240 1920 -200 1930
rect 0 2075 200 2080
rect 0 2045 10 2075
rect 190 2045 200 2075
rect 0 2040 200 2045
rect 320 2075 520 2080
rect 320 2045 330 2075
rect 510 2045 520 2075
rect 320 2040 520 2045
rect 640 2075 840 2080
rect 640 2045 650 2075
rect 830 2045 840 2075
rect 640 2040 840 2045
rect 960 2075 1160 2080
rect 960 2045 970 2075
rect 1150 2045 1160 2075
rect 960 2040 1160 2045
rect -80 2010 -40 2020
rect -80 1930 -75 2010
rect -45 1930 -40 2010
rect -80 1920 -40 1930
rect 240 2010 280 2020
rect 240 1930 245 2010
rect 275 1930 280 2010
rect 240 1920 280 1930
rect 560 2010 600 2020
rect 560 1930 565 2010
rect 595 1930 600 2010
rect 560 1920 600 1930
rect 880 2010 920 2020
rect 880 1930 885 2010
rect 915 1930 920 2010
rect 880 1920 920 1930
rect 1200 2010 1240 2020
rect 1200 1930 1205 2010
rect 1235 1930 1240 2010
rect 1200 1920 1240 1930
rect 1440 2075 1640 2080
rect 1440 2045 1450 2075
rect 1630 2045 1640 2075
rect 1440 2040 1640 2045
rect 1760 2075 1960 2080
rect 1760 2045 1770 2075
rect 1950 2045 1960 2075
rect 1760 2040 1960 2045
rect 2080 2075 2280 2080
rect 2080 2045 2090 2075
rect 2270 2045 2280 2075
rect 2080 2040 2280 2045
rect 2400 2075 2600 2080
rect 2400 2045 2410 2075
rect 2590 2045 2600 2075
rect 2400 2040 2600 2045
rect 1360 2010 1400 2020
rect 1360 1930 1365 2010
rect 1395 1930 1400 2010
rect 1360 1920 1400 1930
rect 1680 2010 1720 2020
rect 1680 1930 1685 2010
rect 1715 1930 1720 2010
rect 1680 1920 1720 1930
rect 2000 2010 2040 2020
rect 2000 1930 2005 2010
rect 2035 1930 2040 2010
rect 2000 1920 2040 1930
rect 2320 2010 2360 2020
rect 2320 1930 2325 2010
rect 2355 1930 2360 2010
rect 2320 1920 2360 1930
rect 2640 2010 2680 2020
rect 2640 1930 2645 2010
rect 2675 1930 2680 2010
rect 2640 1920 2680 1930
rect 2880 2075 3080 2080
rect 2880 2045 2890 2075
rect 3070 2045 3080 2075
rect 2880 2040 3080 2045
rect 3200 2075 3400 2080
rect 3200 2045 3210 2075
rect 3390 2045 3400 2075
rect 3200 2040 3400 2045
rect 3520 2075 3720 2080
rect 3520 2045 3530 2075
rect 3710 2045 3720 2075
rect 3520 2040 3720 2045
rect 3840 2075 4040 2080
rect 3840 2045 3850 2075
rect 4030 2045 4040 2075
rect 3840 2040 4040 2045
rect 2800 2010 2840 2020
rect 2800 1930 2805 2010
rect 2835 1930 2840 2010
rect 2800 1920 2840 1930
rect 3120 2010 3160 2020
rect 3120 1930 3125 2010
rect 3155 1930 3160 2010
rect 3120 1920 3160 1930
rect 3440 2010 3480 2020
rect 3440 1930 3445 2010
rect 3475 1930 3480 2010
rect 3440 1920 3480 1930
rect 3760 2010 3800 2020
rect 3760 1930 3765 2010
rect 3795 1930 3800 2010
rect 3760 1920 3800 1930
rect 4080 2010 4120 2020
rect 4080 1930 4085 2010
rect 4115 1930 4120 2010
rect 4080 1920 4120 1930
rect 4240 2075 4520 2080
rect 4240 2045 4330 2075
rect 4510 2045 4520 2075
rect 4240 2040 4520 2045
rect 4240 2010 4280 2040
rect 4240 1930 4245 2010
rect 4275 1930 4280 2010
rect 4240 1920 4280 1930
rect 4560 2010 4600 2120
rect 4560 1930 4565 2010
rect 4595 1930 4600 2010
rect 4560 1840 4600 1930
rect -800 1800 -560 1840
rect -200 1800 -80 1840
rect 1240 1800 1360 1840
rect 2680 1800 2800 1840
rect 4120 1800 4240 1840
rect 4600 1800 4840 1840
rect -800 1760 -760 1800
rect 4800 1760 4840 1800
rect -800 1720 -680 1760
rect 4760 1720 4840 1760
rect -640 1560 -560 1600
rect -200 1560 -80 1600
rect 1240 1560 1360 1600
rect 2680 1560 2800 1600
rect 4120 1560 4240 1600
rect 4600 1560 4680 1600
rect -560 1450 -520 1560
rect -480 1515 -200 1520
rect -480 1485 -470 1515
rect -290 1485 -200 1515
rect -480 1480 -200 1485
rect -560 1370 -555 1450
rect -525 1370 -520 1450
rect -560 1230 -520 1370
rect -560 1150 -555 1230
rect -525 1150 -520 1230
rect -560 1040 -520 1150
rect -240 1450 -200 1480
rect -240 1370 -235 1450
rect -205 1370 -200 1450
rect -240 1230 -200 1370
rect -240 1150 -235 1230
rect -205 1150 -200 1230
rect -240 1120 -200 1150
rect -480 1115 -200 1120
rect -480 1085 -470 1115
rect -290 1085 -200 1115
rect -480 1080 -200 1085
rect 0 1515 200 1520
rect 0 1485 10 1515
rect 190 1485 200 1515
rect 0 1480 200 1485
rect 320 1515 520 1520
rect 320 1485 330 1515
rect 510 1485 520 1515
rect 320 1480 520 1485
rect 640 1515 840 1520
rect 640 1485 650 1515
rect 830 1485 840 1515
rect 640 1480 840 1485
rect 960 1515 1160 1520
rect 960 1485 970 1515
rect 1150 1485 1160 1515
rect 960 1480 1160 1485
rect -80 1450 -40 1460
rect -80 1370 -75 1450
rect -45 1370 -40 1450
rect -80 1360 -40 1370
rect 240 1450 280 1460
rect 240 1370 245 1450
rect 275 1370 280 1450
rect 240 1360 280 1370
rect 560 1450 600 1460
rect 560 1370 565 1450
rect 595 1370 600 1450
rect 560 1360 600 1370
rect 880 1450 920 1460
rect 880 1370 885 1450
rect 915 1370 920 1450
rect 880 1360 920 1370
rect 1200 1450 1240 1460
rect 1200 1370 1205 1450
rect 1235 1370 1240 1450
rect 1200 1360 1240 1370
rect -80 1230 -40 1240
rect -80 1150 -75 1230
rect -45 1150 -40 1230
rect -80 1140 -40 1150
rect 240 1230 280 1240
rect 240 1150 245 1230
rect 275 1150 280 1230
rect 240 1140 280 1150
rect 560 1230 600 1240
rect 560 1150 565 1230
rect 595 1150 600 1230
rect 560 1140 600 1150
rect 880 1230 920 1240
rect 880 1150 885 1230
rect 915 1150 920 1230
rect 880 1140 920 1150
rect 1200 1230 1240 1240
rect 1200 1150 1205 1230
rect 1235 1150 1240 1230
rect 1200 1140 1240 1150
rect 0 1115 200 1120
rect 0 1085 10 1115
rect 190 1085 200 1115
rect 0 1080 200 1085
rect 320 1115 520 1120
rect 320 1085 330 1115
rect 510 1085 520 1115
rect 320 1080 520 1085
rect 640 1115 840 1120
rect 640 1085 650 1115
rect 830 1085 840 1115
rect 640 1080 840 1085
rect 960 1115 1160 1120
rect 960 1085 970 1115
rect 1150 1085 1160 1115
rect 960 1080 1160 1085
rect 1440 1515 1640 1520
rect 1440 1485 1450 1515
rect 1630 1485 1640 1515
rect 1440 1480 1640 1485
rect 1760 1515 1960 1520
rect 1760 1485 1770 1515
rect 1950 1485 1960 1515
rect 1760 1480 1960 1485
rect 2080 1515 2280 1520
rect 2080 1485 2090 1515
rect 2270 1485 2280 1515
rect 2080 1480 2280 1485
rect 2400 1515 2600 1520
rect 2400 1485 2410 1515
rect 2590 1485 2600 1515
rect 2400 1480 2600 1485
rect 1360 1450 1400 1460
rect 1360 1370 1365 1450
rect 1395 1370 1400 1450
rect 1360 1360 1400 1370
rect 1680 1450 1720 1460
rect 1680 1370 1685 1450
rect 1715 1370 1720 1450
rect 1680 1360 1720 1370
rect 2000 1450 2040 1460
rect 2000 1370 2005 1450
rect 2035 1370 2040 1450
rect 2000 1360 2040 1370
rect 2320 1450 2360 1460
rect 2320 1370 2325 1450
rect 2355 1370 2360 1450
rect 2320 1360 2360 1370
rect 2640 1450 2680 1460
rect 2640 1370 2645 1450
rect 2675 1370 2680 1450
rect 2640 1360 2680 1370
rect 1360 1230 1400 1240
rect 1360 1150 1365 1230
rect 1395 1150 1400 1230
rect 1360 1140 1400 1150
rect 1680 1230 1720 1240
rect 1680 1150 1685 1230
rect 1715 1150 1720 1230
rect 1680 1140 1720 1150
rect 2000 1230 2040 1240
rect 2000 1150 2005 1230
rect 2035 1150 2040 1230
rect 2000 1140 2040 1150
rect 2320 1230 2360 1240
rect 2320 1150 2325 1230
rect 2355 1150 2360 1230
rect 2320 1140 2360 1150
rect 2640 1230 2680 1240
rect 2640 1150 2645 1230
rect 2675 1150 2680 1230
rect 2640 1140 2680 1150
rect 1440 1115 1640 1120
rect 1440 1085 1450 1115
rect 1630 1085 1640 1115
rect 1440 1080 1640 1085
rect 1760 1115 1960 1120
rect 1760 1085 1770 1115
rect 1950 1085 1960 1115
rect 1760 1080 1960 1085
rect 2080 1115 2280 1120
rect 2080 1085 2090 1115
rect 2270 1085 2280 1115
rect 2080 1080 2280 1085
rect 2400 1115 2600 1120
rect 2400 1085 2410 1115
rect 2590 1085 2600 1115
rect 2400 1080 2600 1085
rect 2880 1515 3080 1520
rect 2880 1485 2890 1515
rect 3070 1485 3080 1515
rect 2880 1480 3080 1485
rect 3200 1515 3400 1520
rect 3200 1485 3210 1515
rect 3390 1485 3400 1515
rect 3200 1480 3400 1485
rect 3520 1515 3720 1520
rect 3520 1485 3530 1515
rect 3710 1485 3720 1515
rect 3520 1480 3720 1485
rect 3840 1515 4040 1520
rect 3840 1485 3850 1515
rect 4030 1485 4040 1515
rect 3840 1480 4040 1485
rect 2800 1450 2840 1460
rect 2800 1370 2805 1450
rect 2835 1370 2840 1450
rect 2800 1360 2840 1370
rect 3120 1450 3160 1460
rect 3120 1370 3125 1450
rect 3155 1370 3160 1450
rect 3120 1360 3160 1370
rect 3440 1450 3480 1460
rect 3440 1370 3445 1450
rect 3475 1370 3480 1450
rect 3440 1360 3480 1370
rect 3760 1450 3800 1460
rect 3760 1370 3765 1450
rect 3795 1370 3800 1450
rect 3760 1360 3800 1370
rect 4080 1450 4120 1460
rect 4080 1370 4085 1450
rect 4115 1370 4120 1450
rect 4080 1360 4120 1370
rect 2800 1230 2840 1240
rect 2800 1150 2805 1230
rect 2835 1150 2840 1230
rect 2800 1140 2840 1150
rect 3120 1230 3160 1240
rect 3120 1150 3125 1230
rect 3155 1150 3160 1230
rect 3120 1140 3160 1150
rect 3440 1230 3480 1240
rect 3440 1150 3445 1230
rect 3475 1150 3480 1230
rect 3440 1140 3480 1150
rect 3760 1230 3800 1240
rect 3760 1150 3765 1230
rect 3795 1150 3800 1230
rect 3760 1140 3800 1150
rect 4080 1230 4120 1240
rect 4080 1150 4085 1230
rect 4115 1150 4120 1230
rect 4080 1140 4120 1150
rect 2880 1115 3080 1120
rect 2880 1085 2890 1115
rect 3070 1085 3080 1115
rect 2880 1080 3080 1085
rect 3200 1115 3400 1120
rect 3200 1085 3210 1115
rect 3390 1085 3400 1115
rect 3200 1080 3400 1085
rect 3520 1115 3720 1120
rect 3520 1085 3530 1115
rect 3710 1085 3720 1115
rect 3520 1080 3720 1085
rect 3840 1115 4040 1120
rect 3840 1085 3850 1115
rect 4030 1085 4040 1115
rect 3840 1080 4040 1085
rect 4240 1515 4520 1520
rect 4240 1485 4330 1515
rect 4510 1485 4520 1515
rect 4240 1480 4520 1485
rect 4240 1450 4280 1480
rect 4240 1370 4245 1450
rect 4275 1370 4280 1450
rect 4240 1230 4280 1370
rect 4240 1150 4245 1230
rect 4275 1150 4280 1230
rect 4240 1120 4280 1150
rect 4560 1450 4600 1560
rect 4560 1370 4565 1450
rect 4595 1370 4600 1450
rect 4560 1230 4600 1370
rect 4560 1150 4565 1230
rect 4595 1150 4600 1230
rect 4240 1115 4520 1120
rect 4240 1085 4330 1115
rect 4510 1085 4520 1115
rect 4240 1080 4520 1085
rect 4560 1040 4600 1150
rect -640 1000 -560 1040
rect -200 1000 -80 1040
rect 1240 1000 1360 1040
rect 2680 1000 2800 1040
rect 4120 1000 4240 1040
rect 4600 1000 4680 1040
rect -800 840 -680 880
rect 4760 840 4840 880
rect -800 200 -560 240
rect -200 200 -80 240
rect 1240 200 1360 240
rect 2680 200 2800 240
rect 4120 200 4240 240
rect 4600 200 4840 240
rect -560 90 -520 200
rect -480 155 -200 160
rect -480 125 -470 155
rect -290 125 -200 155
rect -480 120 -200 125
rect -560 10 -555 90
rect -525 10 -520 90
rect -560 -80 -520 10
rect -240 90 -200 120
rect -240 10 -235 90
rect -205 10 -200 90
rect -240 0 -200 10
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 120 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 120 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 120 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 120 1160 125
rect -80 90 -40 100
rect -80 10 -75 90
rect -45 10 -40 90
rect -80 0 -40 10
rect 240 90 280 100
rect 240 10 245 90
rect 275 10 280 90
rect 240 0 280 10
rect 560 90 600 100
rect 560 10 565 90
rect 595 10 600 90
rect 560 0 600 10
rect 880 90 920 100
rect 880 10 885 90
rect 915 10 920 90
rect 880 0 920 10
rect 1200 90 1240 100
rect 1200 10 1205 90
rect 1235 10 1240 90
rect 1200 0 1240 10
rect 1440 155 1640 160
rect 1440 125 1450 155
rect 1630 125 1640 155
rect 1440 120 1640 125
rect 1760 155 1960 160
rect 1760 125 1770 155
rect 1950 125 1960 155
rect 1760 120 1960 125
rect 2080 155 2280 160
rect 2080 125 2090 155
rect 2270 125 2280 155
rect 2080 120 2280 125
rect 2400 155 2600 160
rect 2400 125 2410 155
rect 2590 125 2600 155
rect 2400 120 2600 125
rect 1360 90 1400 100
rect 1360 10 1365 90
rect 1395 10 1400 90
rect 1360 0 1400 10
rect 1680 90 1720 100
rect 1680 10 1685 90
rect 1715 10 1720 90
rect 1680 0 1720 10
rect 2000 90 2040 100
rect 2000 10 2005 90
rect 2035 10 2040 90
rect 2000 0 2040 10
rect 2320 90 2360 100
rect 2320 10 2325 90
rect 2355 10 2360 90
rect 2320 0 2360 10
rect 2640 90 2680 100
rect 2640 10 2645 90
rect 2675 10 2680 90
rect 2640 0 2680 10
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 120 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 120 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 120 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 120 4040 125
rect 2800 90 2840 100
rect 2800 10 2805 90
rect 2835 10 2840 90
rect 2800 0 2840 10
rect 3120 90 3160 100
rect 3120 10 3125 90
rect 3155 10 3160 90
rect 3120 0 3160 10
rect 3440 90 3480 100
rect 3440 10 3445 90
rect 3475 10 3480 90
rect 3440 0 3480 10
rect 3760 90 3800 100
rect 3760 10 3765 90
rect 3795 10 3800 90
rect 3760 0 3800 10
rect 4080 90 4120 100
rect 4080 10 4085 90
rect 4115 10 4120 90
rect 4080 0 4120 10
rect 4240 155 4520 160
rect 4240 125 4330 155
rect 4510 125 4520 155
rect 4240 120 4520 125
rect 4240 90 4280 120
rect 4240 10 4245 90
rect 4275 10 4280 90
rect 4240 0 4280 10
rect 4560 90 4600 200
rect 4560 10 4565 90
rect 4595 10 4600 90
rect 4560 -80 4600 10
rect -800 -120 -560 -80
rect -200 -120 -80 -80
rect 1240 -120 1360 -80
rect 2680 -120 2800 -80
rect 4120 -120 4240 -80
rect 4600 -120 4840 -80
<< viali >>
rect -470 5325 -290 5355
rect -555 5210 -525 5290
rect -555 4990 -525 5070
rect -235 5210 -205 5290
rect -235 4990 -205 5070
rect -470 4925 -290 4955
rect 10 5325 190 5355
rect 330 5325 510 5355
rect 650 5325 830 5355
rect 970 5325 1150 5355
rect -75 5210 -45 5290
rect 245 5210 275 5290
rect 565 5210 595 5290
rect 885 5210 915 5290
rect 1205 5210 1235 5290
rect -75 4990 -45 5070
rect 245 4990 275 5070
rect 565 4990 595 5070
rect 885 4990 915 5070
rect 1205 4990 1235 5070
rect 10 4925 190 4955
rect 330 4925 510 4955
rect 650 4925 830 4955
rect 970 4925 1150 4955
rect 1450 5325 1630 5355
rect 1770 5325 1950 5355
rect 2090 5325 2270 5355
rect 2410 5325 2590 5355
rect 1365 5210 1395 5290
rect 1685 5210 1715 5290
rect 2005 5210 2035 5290
rect 2325 5210 2355 5290
rect 2645 5210 2675 5290
rect 1365 4990 1395 5070
rect 1685 4990 1715 5070
rect 2005 4990 2035 5070
rect 2325 4990 2355 5070
rect 2645 4990 2675 5070
rect 1450 4925 1630 4955
rect 1770 4925 1950 4955
rect 2090 4925 2270 4955
rect 2410 4925 2590 4955
rect 2890 5325 3070 5355
rect 3210 5325 3390 5355
rect 3530 5325 3710 5355
rect 3850 5325 4030 5355
rect 2805 5210 2835 5290
rect 3125 5210 3155 5290
rect 3445 5210 3475 5290
rect 3765 5210 3795 5290
rect 4085 5210 4115 5290
rect 2805 4990 2835 5070
rect 3125 4990 3155 5070
rect 3445 4990 3475 5070
rect 3765 4990 3795 5070
rect 4085 4990 4115 5070
rect 2890 4925 3070 4955
rect 3210 4925 3390 4955
rect 3530 4925 3710 4955
rect 3850 4925 4030 4955
rect 4330 5325 4510 5355
rect 4245 5210 4275 5290
rect 4245 4990 4275 5070
rect 4565 5210 4595 5290
rect 4565 4990 4595 5070
rect 4330 4925 4510 4955
rect -470 3965 -290 3995
rect -555 3850 -525 3930
rect -235 3850 -205 3930
rect 10 3965 190 3995
rect 330 3965 510 3995
rect 650 3965 830 3995
rect 970 3965 1150 3995
rect -75 3850 -45 3930
rect 245 3850 275 3930
rect 565 3850 595 3930
rect 885 3850 915 3930
rect 1205 3850 1235 3930
rect 1450 3965 1630 3995
rect 1770 3965 1950 3995
rect 2090 3965 2270 3995
rect 2410 3965 2590 3995
rect 1365 3850 1395 3930
rect 1685 3850 1715 3930
rect 2005 3850 2035 3930
rect 2325 3850 2355 3930
rect 2645 3850 2675 3930
rect 2890 3965 3070 3995
rect 3210 3965 3390 3995
rect 3530 3965 3710 3995
rect 3850 3965 4030 3995
rect 2805 3850 2835 3930
rect 3125 3850 3155 3930
rect 3445 3850 3475 3930
rect 3765 3850 3795 3930
rect 4085 3850 4115 3930
rect 4330 3965 4510 3995
rect 4245 3850 4275 3930
rect 4565 3850 4595 3930
rect -470 3405 -290 3435
rect -555 3290 -525 3370
rect -555 3070 -525 3150
rect -235 3290 -205 3370
rect -235 3070 -205 3150
rect -470 3005 -290 3035
rect 10 3405 190 3435
rect 330 3405 510 3435
rect 650 3405 830 3435
rect 970 3405 1150 3435
rect -75 3290 -45 3370
rect 245 3290 275 3370
rect 565 3290 595 3370
rect 885 3290 915 3370
rect 1205 3290 1235 3370
rect -75 3070 -45 3150
rect 245 3070 275 3150
rect 565 3070 595 3150
rect 885 3070 915 3150
rect 1205 3070 1235 3150
rect 10 3005 190 3035
rect 330 3005 510 3035
rect 650 3005 830 3035
rect 970 3005 1150 3035
rect 1450 3405 1630 3435
rect 1770 3405 1950 3435
rect 2090 3405 2270 3435
rect 2410 3405 2590 3435
rect 1365 3290 1395 3370
rect 1685 3290 1715 3370
rect 2005 3290 2035 3370
rect 2325 3290 2355 3370
rect 2645 3290 2675 3370
rect 1365 3070 1395 3150
rect 1685 3070 1715 3150
rect 2005 3070 2035 3150
rect 2325 3070 2355 3150
rect 2645 3070 2675 3150
rect 1450 3005 1630 3035
rect 1770 3005 1950 3035
rect 2090 3005 2270 3035
rect 2410 3005 2590 3035
rect 2890 3405 3070 3435
rect 3210 3405 3390 3435
rect 3530 3405 3710 3435
rect 3850 3405 4030 3435
rect 2805 3290 2835 3370
rect 3125 3290 3155 3370
rect 3445 3290 3475 3370
rect 3765 3290 3795 3370
rect 4085 3290 4115 3370
rect 2805 3070 2835 3150
rect 3125 3070 3155 3150
rect 3445 3070 3475 3150
rect 3765 3070 3795 3150
rect 4085 3070 4115 3150
rect 2890 3005 3070 3035
rect 3210 3005 3390 3035
rect 3530 3005 3710 3035
rect 3850 3005 4030 3035
rect 4330 3405 4510 3435
rect 4245 3290 4275 3370
rect 4245 3070 4275 3150
rect 4565 3290 4595 3370
rect 4565 3070 4595 3150
rect 4330 3005 4510 3035
rect -470 2045 -290 2075
rect -555 1930 -525 2010
rect -235 1930 -205 2010
rect 10 2045 190 2075
rect 330 2045 510 2075
rect 650 2045 830 2075
rect 970 2045 1150 2075
rect -75 1930 -45 2010
rect 245 1930 275 2010
rect 565 1930 595 2010
rect 885 1930 915 2010
rect 1205 1930 1235 2010
rect 1450 2045 1630 2075
rect 1770 2045 1950 2075
rect 2090 2045 2270 2075
rect 2410 2045 2590 2075
rect 1365 1930 1395 2010
rect 1685 1930 1715 2010
rect 2005 1930 2035 2010
rect 2325 1930 2355 2010
rect 2645 1930 2675 2010
rect 2890 2045 3070 2075
rect 3210 2045 3390 2075
rect 3530 2045 3710 2075
rect 3850 2045 4030 2075
rect 2805 1930 2835 2010
rect 3125 1930 3155 2010
rect 3445 1930 3475 2010
rect 3765 1930 3795 2010
rect 4085 1930 4115 2010
rect 4330 2045 4510 2075
rect 4245 1930 4275 2010
rect 4565 1930 4595 2010
rect -470 1485 -290 1515
rect -555 1370 -525 1450
rect -555 1150 -525 1230
rect -235 1370 -205 1450
rect -235 1150 -205 1230
rect -470 1085 -290 1115
rect 10 1485 190 1515
rect 330 1485 510 1515
rect 650 1485 830 1515
rect 970 1485 1150 1515
rect -75 1370 -45 1450
rect 245 1370 275 1450
rect 565 1370 595 1450
rect 885 1370 915 1450
rect 1205 1370 1235 1450
rect -75 1150 -45 1230
rect 245 1150 275 1230
rect 565 1150 595 1230
rect 885 1150 915 1230
rect 1205 1150 1235 1230
rect 10 1085 190 1115
rect 330 1085 510 1115
rect 650 1085 830 1115
rect 970 1085 1150 1115
rect 1450 1485 1630 1515
rect 1770 1485 1950 1515
rect 2090 1485 2270 1515
rect 2410 1485 2590 1515
rect 1365 1370 1395 1450
rect 1685 1370 1715 1450
rect 2005 1370 2035 1450
rect 2325 1370 2355 1450
rect 2645 1370 2675 1450
rect 1365 1150 1395 1230
rect 1685 1150 1715 1230
rect 2005 1150 2035 1230
rect 2325 1150 2355 1230
rect 2645 1150 2675 1230
rect 1450 1085 1630 1115
rect 1770 1085 1950 1115
rect 2090 1085 2270 1115
rect 2410 1085 2590 1115
rect 2890 1485 3070 1515
rect 3210 1485 3390 1515
rect 3530 1485 3710 1515
rect 3850 1485 4030 1515
rect 2805 1370 2835 1450
rect 3125 1370 3155 1450
rect 3445 1370 3475 1450
rect 3765 1370 3795 1450
rect 4085 1370 4115 1450
rect 2805 1150 2835 1230
rect 3125 1150 3155 1230
rect 3445 1150 3475 1230
rect 3765 1150 3795 1230
rect 4085 1150 4115 1230
rect 2890 1085 3070 1115
rect 3210 1085 3390 1115
rect 3530 1085 3710 1115
rect 3850 1085 4030 1115
rect 4330 1485 4510 1515
rect 4245 1370 4275 1450
rect 4245 1150 4275 1230
rect 4565 1370 4595 1450
rect 4565 1150 4595 1230
rect 4330 1085 4510 1115
rect -470 125 -290 155
rect -555 10 -525 90
rect -235 10 -205 90
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect -75 10 -45 90
rect 245 10 275 90
rect 565 10 595 90
rect 885 10 915 90
rect 1205 10 1235 90
rect 1450 125 1630 155
rect 1770 125 1950 155
rect 2090 125 2270 155
rect 2410 125 2590 155
rect 1365 10 1395 90
rect 1685 10 1715 90
rect 2005 10 2035 90
rect 2325 10 2355 90
rect 2645 10 2675 90
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3850 125 4030 155
rect 2805 10 2835 90
rect 3125 10 3155 90
rect 3445 10 3475 90
rect 3765 10 3795 90
rect 4085 10 4115 90
rect 4330 125 4510 155
rect 4245 10 4275 90
rect 4565 10 4595 90
<< metal1 >>
rect -480 5355 -280 5360
rect -480 5325 -470 5355
rect -290 5325 -280 5355
rect -480 5320 -280 5325
rect 0 5355 200 5360
rect 0 5325 10 5355
rect 190 5325 200 5355
rect 0 5320 200 5325
rect 320 5355 520 5360
rect 320 5325 330 5355
rect 510 5325 520 5355
rect 320 5320 520 5325
rect 640 5355 840 5360
rect 640 5325 650 5355
rect 830 5325 840 5355
rect 640 5320 840 5325
rect 960 5355 1160 5360
rect 960 5325 970 5355
rect 1150 5325 1160 5355
rect 960 5320 1160 5325
rect 1440 5355 1640 5360
rect 1440 5325 1450 5355
rect 1630 5325 1640 5355
rect 1440 5320 1640 5325
rect 1760 5355 1960 5360
rect 1760 5325 1770 5355
rect 1950 5325 1960 5355
rect 1760 5320 1960 5325
rect 2080 5355 2280 5360
rect 2080 5325 2090 5355
rect 2270 5325 2280 5355
rect 2080 5320 2280 5325
rect 2400 5355 2600 5360
rect 2400 5325 2410 5355
rect 2590 5325 2600 5355
rect 2400 5320 2600 5325
rect 2880 5355 3080 5360
rect 2880 5325 2890 5355
rect 3070 5325 3080 5355
rect 2880 5320 3080 5325
rect 3200 5355 3400 5360
rect 3200 5325 3210 5355
rect 3390 5325 3400 5355
rect 3200 5320 3400 5325
rect 3520 5355 3720 5360
rect 3520 5325 3530 5355
rect 3710 5325 3720 5355
rect 3520 5320 3720 5325
rect 3840 5355 4040 5360
rect 3840 5325 3850 5355
rect 4030 5325 4040 5355
rect 3840 5320 4040 5325
rect 4320 5355 4520 5360
rect 4320 5325 4330 5355
rect 4510 5325 4520 5355
rect 4320 5320 4520 5325
rect -560 5290 -520 5300
rect -560 5210 -555 5290
rect -525 5210 -520 5290
rect -560 5195 -520 5210
rect -560 5165 -555 5195
rect -525 5165 -520 5195
rect -560 5115 -520 5165
rect -560 5085 -555 5115
rect -525 5085 -520 5115
rect -560 5070 -520 5085
rect -560 4990 -555 5070
rect -525 4990 -520 5070
rect -560 4980 -520 4990
rect -240 5290 -200 5300
rect -240 5210 -235 5290
rect -205 5210 -200 5290
rect -240 5070 -200 5210
rect -240 4990 -235 5070
rect -205 4990 -200 5070
rect -240 4980 -200 4990
rect -80 5290 -40 5300
rect -80 5210 -75 5290
rect -45 5210 -40 5290
rect -80 5070 -40 5210
rect 240 5290 280 5300
rect 240 5210 245 5290
rect 275 5210 280 5290
rect 240 5200 280 5210
rect 560 5290 600 5300
rect 560 5210 565 5290
rect 595 5210 600 5290
rect 560 5195 600 5210
rect 880 5290 920 5300
rect 880 5210 885 5290
rect 915 5210 920 5290
rect 880 5200 920 5210
rect 1200 5290 1240 5300
rect 1200 5210 1205 5290
rect 1235 5210 1240 5290
rect 560 5165 565 5195
rect 595 5165 600 5195
rect 560 5160 600 5165
rect -80 4990 -75 5070
rect -45 4990 -40 5070
rect -80 4980 -40 4990
rect 240 5070 280 5080
rect 240 4990 245 5070
rect 275 4990 280 5070
rect 240 4980 280 4990
rect 560 5070 600 5080
rect 560 4990 565 5070
rect 595 4990 600 5070
rect -480 4955 -280 4960
rect -480 4925 -470 4955
rect -290 4925 -280 4955
rect -480 4920 -280 4925
rect 0 4955 200 4960
rect 0 4925 10 4955
rect 190 4925 200 4955
rect 0 4920 200 4925
rect 320 4955 520 4960
rect 320 4925 330 4955
rect 510 4925 520 4955
rect 320 4920 520 4925
rect 80 4795 120 4800
rect 80 4765 85 4795
rect 115 4765 120 4795
rect -80 4155 -40 4160
rect -80 4125 -75 4155
rect -45 4125 -40 4155
rect -800 4075 -760 4080
rect -800 4045 -795 4075
rect -765 4045 -760 4075
rect -800 3915 -760 4045
rect -480 3995 -280 4000
rect -480 3965 -470 3995
rect -290 3965 -280 3995
rect -480 3960 -280 3965
rect -800 3885 -795 3915
rect -765 3885 -760 3915
rect -800 3835 -760 3885
rect -800 3805 -795 3835
rect -765 3805 -760 3835
rect -800 3755 -760 3805
rect -560 3930 -520 3940
rect -560 3850 -555 3930
rect -525 3850 -520 3930
rect -560 3835 -520 3850
rect -240 3930 -200 3940
rect -240 3850 -235 3930
rect -205 3850 -200 3930
rect -240 3840 -200 3850
rect -160 3915 -120 4000
rect -160 3885 -155 3915
rect -125 3885 -120 3915
rect -560 3805 -555 3835
rect -525 3805 -520 3835
rect -560 3800 -520 3805
rect -160 3835 -120 3885
rect -80 3930 -40 4125
rect 80 4000 120 4765
rect 400 4795 440 4800
rect 400 4765 405 4795
rect 435 4765 440 4795
rect 240 4555 280 4560
rect 240 4525 245 4555
rect 275 4525 280 4555
rect 0 3995 200 4000
rect 0 3965 10 3995
rect 190 3965 200 3995
rect 0 3960 200 3965
rect -80 3850 -75 3930
rect -45 3850 -40 3930
rect -80 3840 -40 3850
rect 240 3930 280 4525
rect 400 4000 440 4765
rect 560 4315 600 4990
rect 880 5070 920 5080
rect 880 4990 885 5070
rect 915 4990 920 5070
rect 880 4980 920 4990
rect 1200 5070 1240 5210
rect 1200 4990 1205 5070
rect 1235 4990 1240 5070
rect 1200 4980 1240 4990
rect 1360 5290 1400 5300
rect 1360 5210 1365 5290
rect 1395 5210 1400 5290
rect 1360 5195 1400 5210
rect 1360 5165 1365 5195
rect 1395 5165 1400 5195
rect 1360 5115 1400 5165
rect 1360 5085 1365 5115
rect 1395 5085 1400 5115
rect 1360 5070 1400 5085
rect 1360 4990 1365 5070
rect 1395 4990 1400 5070
rect 1360 4980 1400 4990
rect 1520 4960 1560 5320
rect 1680 5290 1720 5300
rect 1680 5210 1685 5290
rect 1715 5210 1720 5290
rect 1680 5200 1720 5210
rect 1680 5070 1720 5080
rect 1680 4990 1685 5070
rect 1715 4990 1720 5070
rect 1680 4980 1720 4990
rect 1840 4960 1880 5320
rect 2000 5290 2040 5300
rect 2000 5210 2005 5290
rect 2035 5210 2040 5290
rect 2000 5200 2040 5210
rect 2000 5070 2040 5080
rect 2000 4990 2005 5070
rect 2035 4990 2040 5070
rect 2000 4980 2040 4990
rect 2160 4960 2200 5320
rect 2320 5290 2360 5300
rect 2320 5210 2325 5290
rect 2355 5210 2360 5290
rect 2320 5200 2360 5210
rect 2320 5070 2360 5080
rect 2320 4990 2325 5070
rect 2355 4990 2360 5070
rect 2320 4980 2360 4990
rect 2480 4960 2520 5320
rect 2640 5290 2680 5300
rect 2640 5210 2645 5290
rect 2675 5210 2680 5290
rect 2640 5195 2680 5210
rect 2640 5165 2645 5195
rect 2675 5165 2680 5195
rect 2640 5115 2680 5165
rect 2640 5085 2645 5115
rect 2675 5085 2680 5115
rect 2640 5070 2680 5085
rect 2640 4990 2645 5070
rect 2675 4990 2680 5070
rect 2640 4980 2680 4990
rect 2800 5290 2840 5300
rect 2800 5210 2805 5290
rect 2835 5210 2840 5290
rect 2800 5195 2840 5210
rect 2800 5165 2805 5195
rect 2835 5165 2840 5195
rect 2800 5115 2840 5165
rect 2800 5085 2805 5115
rect 2835 5085 2840 5115
rect 2800 5070 2840 5085
rect 2800 4990 2805 5070
rect 2835 4990 2840 5070
rect 2800 4980 2840 4990
rect 2960 4960 3000 5320
rect 3120 5290 3160 5300
rect 3120 5210 3125 5290
rect 3155 5210 3160 5290
rect 3120 5200 3160 5210
rect 3120 5070 3160 5080
rect 3120 4990 3125 5070
rect 3155 4990 3160 5070
rect 3120 4980 3160 4990
rect 3280 4960 3320 5320
rect 3440 5290 3480 5300
rect 3440 5210 3445 5290
rect 3475 5210 3480 5290
rect 3440 5200 3480 5210
rect 3440 5070 3480 5080
rect 3440 4990 3445 5070
rect 3475 4990 3480 5070
rect 3440 4980 3480 4990
rect 3600 4960 3640 5320
rect 3760 5290 3800 5300
rect 3760 5210 3765 5290
rect 3795 5210 3800 5290
rect 3760 5200 3800 5210
rect 3760 5070 3800 5080
rect 3760 4990 3765 5070
rect 3795 4990 3800 5070
rect 3760 4980 3800 4990
rect 3920 4960 3960 5320
rect 4080 5290 4120 5300
rect 4080 5210 4085 5290
rect 4115 5210 4120 5290
rect 4080 5195 4120 5210
rect 4080 5165 4085 5195
rect 4115 5165 4120 5195
rect 4080 5115 4120 5165
rect 4080 5085 4085 5115
rect 4115 5085 4120 5115
rect 4080 5070 4120 5085
rect 4080 4990 4085 5070
rect 4115 4990 4120 5070
rect 4080 4980 4120 4990
rect 4240 5290 4280 5300
rect 4240 5210 4245 5290
rect 4275 5210 4280 5290
rect 4240 5070 4280 5210
rect 4240 4990 4245 5070
rect 4275 4990 4280 5070
rect 4240 4980 4280 4990
rect 4560 5290 4600 5300
rect 4560 5210 4565 5290
rect 4595 5210 4600 5290
rect 4560 5195 4600 5210
rect 4560 5165 4565 5195
rect 4595 5165 4600 5195
rect 4560 5115 4600 5165
rect 4560 5085 4565 5115
rect 4595 5085 4600 5115
rect 4560 5070 4600 5085
rect 4560 4990 4565 5070
rect 4595 4990 4600 5070
rect 4560 4980 4600 4990
rect 640 4955 840 4960
rect 640 4925 650 4955
rect 830 4925 840 4955
rect 640 4920 840 4925
rect 960 4955 1160 4960
rect 960 4925 970 4955
rect 1150 4925 1160 4955
rect 960 4920 1160 4925
rect 1440 4955 1640 4960
rect 1440 4925 1450 4955
rect 1630 4925 1640 4955
rect 1440 4920 1640 4925
rect 1760 4955 1960 4960
rect 1760 4925 1770 4955
rect 1950 4925 1960 4955
rect 1760 4920 1960 4925
rect 2080 4955 2280 4960
rect 2080 4925 2090 4955
rect 2270 4925 2280 4955
rect 2080 4920 2280 4925
rect 2400 4955 2600 4960
rect 2400 4925 2410 4955
rect 2590 4925 2600 4955
rect 2400 4920 2600 4925
rect 2880 4955 3080 4960
rect 2880 4925 2890 4955
rect 3070 4925 3080 4955
rect 2880 4920 3080 4925
rect 3200 4955 3400 4960
rect 3200 4925 3210 4955
rect 3390 4925 3400 4955
rect 3200 4920 3400 4925
rect 3520 4955 3720 4960
rect 3520 4925 3530 4955
rect 3710 4925 3720 4955
rect 3520 4920 3720 4925
rect 3840 4955 4040 4960
rect 3840 4925 3850 4955
rect 4030 4925 4040 4955
rect 3840 4920 4040 4925
rect 4320 4955 4520 4960
rect 4320 4925 4330 4955
rect 4510 4925 4520 4955
rect 4320 4920 4520 4925
rect 560 4285 565 4315
rect 595 4285 600 4315
rect 560 4280 600 4285
rect 720 4795 760 4800
rect 720 4765 725 4795
rect 755 4765 760 4795
rect 560 4155 600 4160
rect 560 4125 565 4155
rect 595 4125 600 4155
rect 320 3995 520 4000
rect 320 3965 330 3995
rect 510 3965 520 3995
rect 320 3960 520 3965
rect 560 3960 600 4125
rect 720 4000 760 4765
rect 1040 4795 1080 4800
rect 1040 4765 1045 4795
rect 1075 4765 1080 4795
rect 880 4555 920 4560
rect 880 4525 885 4555
rect 915 4525 920 4555
rect 640 3995 840 4000
rect 640 3965 650 3995
rect 830 3965 840 3995
rect 640 3960 840 3965
rect 240 3850 245 3930
rect 275 3850 280 3930
rect 240 3840 280 3850
rect 560 3930 600 3940
rect 560 3850 565 3930
rect 595 3850 600 3930
rect 560 3840 600 3850
rect 880 3930 920 4525
rect 1040 4000 1080 4765
rect 1520 4795 1560 4920
rect 1520 4765 1525 4795
rect 1555 4765 1560 4795
rect 1200 4155 1240 4160
rect 1200 4125 1205 4155
rect 1235 4125 1240 4155
rect 960 3995 1160 4000
rect 960 3965 970 3995
rect 1150 3965 1160 3995
rect 960 3960 1160 3965
rect 880 3850 885 3930
rect 915 3850 920 3930
rect 880 3840 920 3850
rect 1200 3930 1240 4125
rect 1360 4155 1400 4160
rect 1360 4125 1365 4155
rect 1395 4125 1400 4155
rect 1200 3850 1205 3930
rect 1235 3850 1240 3930
rect 1200 3840 1240 3850
rect 1280 3915 1320 4000
rect 1280 3885 1285 3915
rect 1315 3885 1320 3915
rect -160 3805 -155 3835
rect -125 3805 -120 3835
rect -800 3725 -795 3755
rect -765 3725 -760 3755
rect -800 3720 -760 3725
rect -160 3755 -120 3805
rect -160 3725 -155 3755
rect -125 3725 -120 3755
rect -160 3720 -120 3725
rect 1280 3835 1320 3885
rect 1280 3805 1285 3835
rect 1315 3805 1320 3835
rect 1280 3755 1320 3805
rect 1360 3930 1400 4125
rect 1520 4000 1560 4765
rect 1840 4795 1880 4920
rect 1840 4765 1845 4795
rect 1875 4765 1880 4795
rect 1680 4555 1720 4560
rect 1680 4525 1685 4555
rect 1715 4525 1720 4555
rect 1440 3995 1640 4000
rect 1440 3965 1450 3995
rect 1630 3965 1640 3995
rect 1440 3960 1640 3965
rect 1360 3850 1365 3930
rect 1395 3850 1400 3930
rect 1360 3800 1400 3850
rect 1680 3930 1720 4525
rect 1840 4000 1880 4765
rect 2160 4795 2200 4920
rect 2160 4765 2165 4795
rect 2195 4765 2200 4795
rect 2000 4155 2040 4160
rect 2000 4125 2005 4155
rect 2035 4125 2040 4155
rect 1760 3995 1960 4000
rect 1760 3965 1770 3995
rect 1950 3965 1960 3995
rect 1760 3960 1960 3965
rect 1680 3850 1685 3930
rect 1715 3850 1720 3930
rect 1680 3840 1720 3850
rect 2000 3930 2040 4125
rect 2160 4000 2200 4765
rect 2480 4795 2520 4920
rect 2480 4765 2485 4795
rect 2515 4765 2520 4795
rect 2320 4555 2360 4560
rect 2320 4525 2325 4555
rect 2355 4525 2360 4555
rect 2080 3995 2280 4000
rect 2080 3965 2090 3995
rect 2270 3965 2280 3995
rect 2080 3960 2280 3965
rect 2000 3850 2005 3930
rect 2035 3850 2040 3930
rect 2000 3840 2040 3850
rect 2320 3930 2360 4525
rect 2480 4000 2520 4765
rect 2960 4795 3000 4920
rect 2960 4765 2965 4795
rect 2995 4765 3000 4795
rect 2960 4760 3000 4765
rect 3280 4795 3320 4920
rect 3280 4765 3285 4795
rect 3315 4765 3320 4795
rect 3280 4760 3320 4765
rect 3600 4795 3640 4920
rect 3600 4765 3605 4795
rect 3635 4765 3640 4795
rect 3600 4760 3640 4765
rect 3920 4795 3960 4920
rect 3920 4765 3925 4795
rect 3955 4765 3960 4795
rect 3920 4760 3960 4765
rect 4080 4795 4120 4800
rect 4080 4765 4085 4795
rect 4115 4765 4120 4795
rect 2640 4155 2680 4160
rect 2640 4125 2645 4155
rect 2675 4125 2680 4155
rect 2400 3995 2600 4000
rect 2400 3965 2410 3995
rect 2590 3965 2600 3995
rect 2400 3960 2600 3965
rect 2320 3850 2325 3930
rect 2355 3850 2360 3930
rect 2320 3840 2360 3850
rect 2640 3930 2680 4125
rect 2960 4155 3000 4160
rect 2960 4125 2965 4155
rect 2995 4125 3000 4155
rect 2960 4000 3000 4125
rect 3280 4155 3320 4160
rect 3280 4125 3285 4155
rect 3315 4125 3320 4155
rect 3280 4000 3320 4125
rect 3600 4155 3640 4160
rect 3600 4125 3605 4155
rect 3635 4125 3640 4155
rect 3600 4000 3640 4125
rect 3920 4155 3960 4160
rect 3920 4125 3925 4155
rect 3955 4125 3960 4155
rect 3920 4000 3960 4125
rect 2640 3850 2645 3930
rect 2675 3850 2680 3930
rect 2640 3840 2680 3850
rect 2720 3915 2760 4000
rect 2880 3995 3080 4000
rect 2880 3965 2890 3995
rect 3070 3965 3080 3995
rect 2880 3960 3080 3965
rect 3200 3995 3400 4000
rect 3200 3965 3210 3995
rect 3390 3965 3400 3995
rect 3200 3960 3400 3965
rect 2720 3885 2725 3915
rect 2755 3885 2760 3915
rect 2720 3835 2760 3885
rect 2720 3805 2725 3835
rect 2755 3805 2760 3835
rect 1280 3725 1285 3755
rect 1315 3725 1320 3755
rect 1280 3720 1320 3725
rect 2720 3755 2760 3805
rect 2800 3930 2840 3940
rect 2800 3850 2805 3930
rect 2835 3850 2840 3930
rect 2800 3835 2840 3850
rect 3120 3930 3160 3940
rect 3120 3850 3125 3930
rect 3155 3850 3160 3930
rect 3120 3840 3160 3850
rect 3440 3930 3480 4000
rect 3520 3995 3720 4000
rect 3520 3965 3530 3995
rect 3710 3965 3720 3995
rect 3520 3960 3720 3965
rect 3840 3995 4040 4000
rect 3840 3965 3850 3995
rect 4030 3965 4040 3995
rect 3840 3960 4040 3965
rect 3440 3850 3445 3930
rect 3475 3850 3480 3930
rect 3440 3840 3480 3850
rect 3760 3930 3800 3940
rect 3760 3850 3765 3930
rect 3795 3850 3800 3930
rect 3760 3840 3800 3850
rect 4080 3930 4120 4765
rect 4080 3850 4085 3930
rect 4115 3850 4120 3930
rect 4080 3840 4120 3850
rect 4160 3915 4200 4000
rect 4320 3995 4520 4000
rect 4320 3965 4330 3995
rect 4510 3965 4520 3995
rect 4320 3960 4520 3965
rect 4160 3885 4165 3915
rect 4195 3885 4200 3915
rect 2800 3805 2805 3835
rect 2835 3805 2840 3835
rect 2800 3800 2840 3805
rect 4160 3835 4200 3885
rect 4240 3930 4280 3940
rect 4240 3850 4245 3930
rect 4275 3850 4280 3930
rect 4240 3840 4280 3850
rect 4560 3930 4600 3940
rect 4560 3850 4565 3930
rect 4595 3850 4600 3930
rect 4160 3805 4165 3835
rect 4195 3805 4200 3835
rect 2720 3725 2725 3755
rect 2755 3725 2760 3755
rect 2720 3720 2760 3725
rect 4160 3755 4200 3805
rect 4560 3835 4600 3850
rect 4560 3805 4565 3835
rect 4595 3805 4600 3835
rect 4560 3800 4600 3805
rect 4640 3915 4680 4000
rect 4640 3885 4645 3915
rect 4675 3885 4680 3915
rect 4640 3835 4680 3885
rect 4640 3805 4645 3835
rect 4675 3805 4680 3835
rect 4160 3725 4165 3755
rect 4195 3725 4200 3755
rect 4160 3720 4200 3725
rect 4640 3755 4680 3805
rect 4640 3725 4645 3755
rect 4675 3725 4680 3755
rect 4640 3720 4680 3725
rect -800 3675 -760 3680
rect -800 3645 -795 3675
rect -765 3645 -760 3675
rect -800 3640 -760 3645
rect -480 3435 -280 3440
rect -480 3405 -470 3435
rect -290 3405 -280 3435
rect -480 3400 -280 3405
rect 0 3435 200 3440
rect 0 3405 10 3435
rect 190 3405 200 3435
rect 0 3400 200 3405
rect 320 3435 520 3440
rect 320 3405 330 3435
rect 510 3405 520 3435
rect 320 3400 520 3405
rect 640 3435 840 3440
rect 640 3405 650 3435
rect 830 3405 840 3435
rect 640 3400 840 3405
rect 960 3435 1160 3440
rect 960 3405 970 3435
rect 1150 3405 1160 3435
rect 960 3400 1160 3405
rect 1440 3435 1640 3440
rect 1440 3405 1450 3435
rect 1630 3405 1640 3435
rect 1440 3400 1640 3405
rect 1760 3435 1960 3440
rect 1760 3405 1770 3435
rect 1950 3405 1960 3435
rect 1760 3400 1960 3405
rect 2080 3435 2280 3440
rect 2080 3405 2090 3435
rect 2270 3405 2280 3435
rect 2080 3400 2280 3405
rect 2400 3435 2600 3440
rect 2400 3405 2410 3435
rect 2590 3405 2600 3435
rect 2400 3400 2600 3405
rect 2880 3435 3080 3440
rect 2880 3405 2890 3435
rect 3070 3405 3080 3435
rect 2880 3400 3080 3405
rect 3200 3435 3400 3440
rect 3200 3405 3210 3435
rect 3390 3405 3400 3435
rect 3200 3400 3400 3405
rect 3520 3435 3720 3440
rect 3520 3405 3530 3435
rect 3710 3405 3720 3435
rect 3520 3400 3720 3405
rect 3840 3435 4040 3440
rect 3840 3405 3850 3435
rect 4030 3405 4040 3435
rect 3840 3400 4040 3405
rect 4320 3435 4520 3440
rect 4320 3405 4330 3435
rect 4510 3405 4520 3435
rect 4320 3400 4520 3405
rect -560 3370 -520 3380
rect -560 3290 -555 3370
rect -525 3290 -520 3370
rect -560 3275 -520 3290
rect -560 3245 -555 3275
rect -525 3245 -520 3275
rect -560 3195 -520 3245
rect -560 3165 -555 3195
rect -525 3165 -520 3195
rect -560 3150 -520 3165
rect -560 3070 -555 3150
rect -525 3070 -520 3150
rect -560 3060 -520 3070
rect -240 3370 -200 3380
rect -240 3290 -235 3370
rect -205 3290 -200 3370
rect -240 3150 -200 3290
rect -240 3070 -235 3150
rect -205 3070 -200 3150
rect -240 3060 -200 3070
rect -80 3370 -40 3380
rect -80 3290 -75 3370
rect -45 3290 -40 3370
rect -80 3150 -40 3290
rect 240 3370 280 3380
rect 240 3290 245 3370
rect 275 3290 280 3370
rect 240 3280 280 3290
rect 560 3370 600 3380
rect 560 3290 565 3370
rect 595 3290 600 3370
rect 560 3275 600 3290
rect 880 3370 920 3380
rect 880 3290 885 3370
rect 915 3290 920 3370
rect 880 3280 920 3290
rect 1200 3370 1240 3380
rect 1200 3290 1205 3370
rect 1235 3290 1240 3370
rect 560 3245 565 3275
rect 595 3245 600 3275
rect 560 3240 600 3245
rect -80 3070 -75 3150
rect -45 3070 -40 3150
rect -80 3060 -40 3070
rect 240 3150 280 3160
rect 240 3070 245 3150
rect 275 3070 280 3150
rect 240 3060 280 3070
rect 560 3150 600 3160
rect 560 3070 565 3150
rect 595 3070 600 3150
rect -480 3035 -280 3040
rect -480 3005 -470 3035
rect -290 3005 -280 3035
rect -480 3000 -280 3005
rect 0 3035 200 3040
rect 0 3005 10 3035
rect 190 3005 200 3035
rect 0 3000 200 3005
rect 320 3035 520 3040
rect 320 3005 330 3035
rect 510 3005 520 3035
rect 320 3000 520 3005
rect 560 2635 600 3070
rect 880 3150 920 3160
rect 880 3070 885 3150
rect 915 3070 920 3150
rect 880 3060 920 3070
rect 1200 3150 1240 3290
rect 1200 3070 1205 3150
rect 1235 3070 1240 3150
rect 1200 3060 1240 3070
rect 1360 3370 1400 3380
rect 1360 3290 1365 3370
rect 1395 3290 1400 3370
rect 1360 3150 1400 3290
rect 1680 3370 1720 3380
rect 1680 3290 1685 3370
rect 1715 3290 1720 3370
rect 1680 3280 1720 3290
rect 2000 3370 2040 3380
rect 2000 3290 2005 3370
rect 2035 3290 2040 3370
rect 2000 3275 2040 3290
rect 2320 3370 2360 3380
rect 2320 3290 2325 3370
rect 2355 3290 2360 3370
rect 2320 3280 2360 3290
rect 2640 3370 2680 3380
rect 2640 3290 2645 3370
rect 2675 3290 2680 3370
rect 2000 3245 2005 3275
rect 2035 3245 2040 3275
rect 2000 3240 2040 3245
rect 1360 3070 1365 3150
rect 1395 3070 1400 3150
rect 1360 3060 1400 3070
rect 1680 3150 1720 3160
rect 1680 3070 1685 3150
rect 1715 3070 1720 3150
rect 1680 3060 1720 3070
rect 2000 3150 2040 3160
rect 2000 3070 2005 3150
rect 2035 3070 2040 3150
rect 640 3035 840 3040
rect 640 3005 650 3035
rect 830 3005 840 3035
rect 640 3000 840 3005
rect 960 3035 1160 3040
rect 960 3005 970 3035
rect 1150 3005 1160 3035
rect 960 3000 1160 3005
rect 1440 3035 1640 3040
rect 1440 3005 1450 3035
rect 1630 3005 1640 3035
rect 1440 3000 1640 3005
rect 1760 3035 1960 3040
rect 1760 3005 1770 3035
rect 1950 3005 1960 3035
rect 1760 3000 1960 3005
rect 2000 2875 2040 3070
rect 2320 3150 2360 3160
rect 2320 3070 2325 3150
rect 2355 3070 2360 3150
rect 2320 3060 2360 3070
rect 2640 3150 2680 3290
rect 2640 3070 2645 3150
rect 2675 3070 2680 3150
rect 2640 3060 2680 3070
rect 2800 3370 2840 3380
rect 2800 3290 2805 3370
rect 2835 3290 2840 3370
rect 2800 3275 2840 3290
rect 3120 3370 3160 3380
rect 3120 3290 3125 3370
rect 3155 3290 3160 3370
rect 3120 3280 3160 3290
rect 3440 3370 3480 3380
rect 3440 3290 3445 3370
rect 3475 3290 3480 3370
rect 3440 3280 3480 3290
rect 3760 3370 3800 3380
rect 3760 3290 3765 3370
rect 3795 3290 3800 3370
rect 3760 3280 3800 3290
rect 4080 3370 4120 3380
rect 4080 3290 4085 3370
rect 4115 3290 4120 3370
rect 2800 3245 2805 3275
rect 2835 3245 2840 3275
rect 2800 3195 2840 3245
rect 2800 3165 2805 3195
rect 2835 3165 2840 3195
rect 2800 3150 2840 3165
rect 2800 3070 2805 3150
rect 2835 3070 2840 3150
rect 2800 3060 2840 3070
rect 3120 3150 3160 3160
rect 3120 3070 3125 3150
rect 3155 3070 3160 3150
rect 3120 3060 3160 3070
rect 3440 3150 3480 3160
rect 3440 3070 3445 3150
rect 3475 3070 3480 3150
rect 3440 3060 3480 3070
rect 3760 3150 3800 3160
rect 3760 3070 3765 3150
rect 3795 3070 3800 3150
rect 3760 3060 3800 3070
rect 4080 3150 4120 3290
rect 4080 3070 4085 3150
rect 4115 3070 4120 3150
rect 2080 3035 2280 3040
rect 2080 3005 2090 3035
rect 2270 3005 2280 3035
rect 2080 3000 2280 3005
rect 2400 3035 2600 3040
rect 2400 3005 2410 3035
rect 2590 3005 2600 3035
rect 2400 3000 2600 3005
rect 2880 3035 3080 3040
rect 2880 3005 2890 3035
rect 3070 3005 3080 3035
rect 2880 3000 3080 3005
rect 3200 3035 3400 3040
rect 3200 3005 3210 3035
rect 3390 3005 3400 3035
rect 3200 3000 3400 3005
rect 3440 3035 3480 3040
rect 3440 3005 3445 3035
rect 3475 3005 3480 3035
rect 2000 2845 2005 2875
rect 2035 2845 2040 2875
rect 2000 2840 2040 2845
rect 2640 2875 2680 2880
rect 2640 2845 2645 2875
rect 2675 2845 2680 2875
rect 560 2605 565 2635
rect 595 2605 600 2635
rect 560 2600 600 2605
rect 1200 2635 1240 2640
rect 1200 2605 1205 2635
rect 1235 2605 1240 2635
rect -160 2475 -120 2480
rect -160 2445 -155 2475
rect -125 2445 -120 2475
rect -160 2315 -120 2445
rect -160 2285 -155 2315
rect -125 2285 -120 2315
rect -160 2155 -120 2285
rect -160 2125 -155 2155
rect -125 2125 -120 2155
rect -480 2075 -280 2080
rect -480 2045 -470 2075
rect -290 2045 -280 2075
rect -480 2040 -280 2045
rect -560 2010 -520 2020
rect -560 1930 -555 2010
rect -525 1930 -520 2010
rect -560 1915 -520 1930
rect -240 2010 -200 2020
rect -240 1930 -235 2010
rect -205 1930 -200 2010
rect -240 1920 -200 1930
rect -160 1995 -120 2125
rect 80 2395 120 2400
rect 80 2365 85 2395
rect 115 2365 120 2395
rect 80 2080 120 2365
rect 400 2395 440 2400
rect 400 2365 405 2395
rect 435 2365 440 2395
rect 400 2080 440 2365
rect 720 2395 760 2400
rect 720 2365 725 2395
rect 755 2365 760 2395
rect 720 2080 760 2365
rect 1040 2395 1080 2400
rect 1040 2365 1045 2395
rect 1075 2365 1080 2395
rect 1040 2080 1080 2365
rect 0 2075 200 2080
rect 0 2045 10 2075
rect 190 2045 200 2075
rect 0 2040 200 2045
rect 320 2075 520 2080
rect 320 2045 330 2075
rect 510 2045 520 2075
rect 320 2040 520 2045
rect 640 2075 840 2080
rect 640 2045 650 2075
rect 830 2045 840 2075
rect 640 2040 840 2045
rect 960 2075 1160 2080
rect 960 2045 970 2075
rect 1150 2045 1160 2075
rect 960 2040 1160 2045
rect -160 1965 -155 1995
rect -125 1965 -120 1995
rect -560 1885 -555 1915
rect -525 1885 -520 1915
rect -560 1880 -520 1885
rect -160 1915 -120 1965
rect -160 1885 -155 1915
rect -125 1885 -120 1915
rect -160 1835 -120 1885
rect -80 2010 -40 2020
rect -80 1930 -75 2010
rect -45 1930 -40 2010
rect -80 1915 -40 1930
rect 240 2010 280 2020
rect 240 1930 245 2010
rect 275 1930 280 2010
rect 240 1920 280 1930
rect 560 2010 600 2020
rect 560 1930 565 2010
rect 595 1930 600 2010
rect 560 1920 600 1930
rect 880 2010 920 2020
rect 880 1930 885 2010
rect 915 1930 920 2010
rect 880 1920 920 1930
rect 1200 2010 1240 2605
rect 1200 1930 1205 2010
rect 1235 1930 1240 2010
rect 1200 1920 1240 1930
rect 1280 2475 1320 2480
rect 1280 2445 1285 2475
rect 1315 2445 1320 2475
rect 1280 2315 1320 2445
rect 1280 2285 1285 2315
rect 1315 2285 1320 2315
rect 1280 2155 1320 2285
rect 1280 2125 1285 2155
rect 1315 2125 1320 2155
rect 1280 1995 1320 2125
rect 1520 2235 1560 2240
rect 1520 2205 1525 2235
rect 1555 2205 1560 2235
rect 1520 2080 1560 2205
rect 1840 2235 1880 2240
rect 1840 2205 1845 2235
rect 1875 2205 1880 2235
rect 1840 2080 1880 2205
rect 2160 2235 2200 2240
rect 2160 2205 2165 2235
rect 2195 2205 2200 2235
rect 2160 2080 2200 2205
rect 2480 2235 2520 2240
rect 2480 2205 2485 2235
rect 2515 2205 2520 2235
rect 2480 2080 2520 2205
rect 1440 2075 1640 2080
rect 1440 2045 1450 2075
rect 1630 2045 1640 2075
rect 1440 2040 1640 2045
rect 1760 2075 1960 2080
rect 1760 2045 1770 2075
rect 1950 2045 1960 2075
rect 1760 2040 1960 2045
rect 2080 2075 2280 2080
rect 2080 2045 2090 2075
rect 2270 2045 2280 2075
rect 2080 2040 2280 2045
rect 2400 2075 2600 2080
rect 2400 2045 2410 2075
rect 2590 2045 2600 2075
rect 2400 2040 2600 2045
rect 1280 1965 1285 1995
rect 1315 1965 1320 1995
rect -80 1885 -75 1915
rect -45 1885 -40 1915
rect -80 1880 -40 1885
rect 1280 1915 1320 1965
rect 1280 1885 1285 1915
rect 1315 1885 1320 1915
rect -160 1805 -155 1835
rect -125 1805 -120 1835
rect -160 1800 -120 1805
rect 1280 1835 1320 1885
rect 1360 2010 1400 2020
rect 1360 1930 1365 2010
rect 1395 1930 1400 2010
rect 1360 1915 1400 1930
rect 1680 2010 1720 2020
rect 1680 1930 1685 2010
rect 1715 1930 1720 2010
rect 1680 1920 1720 1930
rect 2000 2010 2040 2020
rect 2000 1930 2005 2010
rect 2035 1930 2040 2010
rect 2000 1920 2040 1930
rect 2320 2010 2360 2020
rect 2320 1930 2325 2010
rect 2355 1930 2360 2010
rect 2320 1920 2360 1930
rect 2640 2010 2680 2845
rect 2640 1930 2645 2010
rect 2675 1930 2680 2010
rect 2640 1920 2680 1930
rect 2720 2475 2760 2480
rect 2720 2445 2725 2475
rect 2755 2445 2760 2475
rect 2720 2315 2760 2445
rect 2720 2285 2725 2315
rect 2755 2285 2760 2315
rect 2720 2155 2760 2285
rect 2720 2125 2725 2155
rect 2755 2125 2760 2155
rect 2720 1995 2760 2125
rect 2960 2235 3000 2240
rect 2960 2205 2965 2235
rect 2995 2205 3000 2235
rect 2960 2080 3000 2205
rect 3280 2235 3320 2240
rect 3280 2205 3285 2235
rect 3315 2205 3320 2235
rect 3280 2080 3320 2205
rect 2880 2075 3080 2080
rect 2880 2045 2890 2075
rect 3070 2045 3080 2075
rect 2880 2040 3080 2045
rect 3200 2075 3400 2080
rect 3200 2045 3210 2075
rect 3390 2045 3400 2075
rect 3200 2040 3400 2045
rect 2720 1965 2725 1995
rect 2755 1965 2760 1995
rect 1360 1885 1365 1915
rect 1395 1885 1400 1915
rect 1360 1880 1400 1885
rect 2720 1915 2760 1965
rect 2720 1885 2725 1915
rect 2755 1885 2760 1915
rect 1280 1805 1285 1835
rect 1315 1805 1320 1835
rect 1280 1800 1320 1805
rect 2720 1835 2760 1885
rect 2800 2010 2840 2020
rect 2800 1930 2805 2010
rect 2835 1930 2840 2010
rect 2800 1915 2840 1930
rect 3120 2010 3160 2020
rect 3120 1930 3125 2010
rect 3155 1930 3160 2010
rect 3120 1920 3160 1930
rect 3440 2010 3480 3005
rect 3520 3035 3720 3040
rect 3520 3005 3530 3035
rect 3710 3005 3720 3035
rect 3520 3000 3720 3005
rect 3840 3035 4040 3040
rect 3840 3005 3850 3035
rect 4030 3005 4040 3035
rect 3840 3000 4040 3005
rect 4080 3035 4120 3070
rect 4240 3370 4280 3380
rect 4240 3290 4245 3370
rect 4275 3290 4280 3370
rect 4240 3150 4280 3290
rect 4240 3070 4245 3150
rect 4275 3070 4280 3150
rect 4240 3060 4280 3070
rect 4560 3370 4600 3380
rect 4560 3290 4565 3370
rect 4595 3290 4600 3370
rect 4560 3275 4600 3290
rect 4560 3245 4565 3275
rect 4595 3245 4600 3275
rect 4560 3195 4600 3245
rect 4560 3165 4565 3195
rect 4595 3165 4600 3195
rect 4560 3150 4600 3165
rect 4560 3070 4565 3150
rect 4595 3070 4600 3150
rect 4560 3060 4600 3070
rect 4080 3005 4085 3035
rect 4115 3005 4120 3035
rect 4080 3000 4120 3005
rect 4320 3035 4520 3040
rect 4320 3005 4330 3035
rect 4510 3005 4520 3035
rect 4320 3000 4520 3005
rect 4160 2475 4200 2480
rect 4160 2445 4165 2475
rect 4195 2445 4200 2475
rect 4160 2315 4200 2445
rect 4160 2285 4165 2315
rect 4195 2285 4200 2315
rect 3600 2235 3640 2240
rect 3600 2205 3605 2235
rect 3635 2205 3640 2235
rect 3600 2080 3640 2205
rect 3920 2235 3960 2240
rect 3920 2205 3925 2235
rect 3955 2205 3960 2235
rect 3920 2080 3960 2205
rect 4160 2155 4200 2285
rect 4160 2125 4165 2155
rect 4195 2125 4200 2155
rect 3520 2075 3720 2080
rect 3520 2045 3530 2075
rect 3710 2045 3720 2075
rect 3520 2040 3720 2045
rect 3840 2075 4040 2080
rect 3840 2045 3850 2075
rect 4030 2045 4040 2075
rect 3840 2040 4040 2045
rect 3440 1930 3445 2010
rect 3475 1930 3480 2010
rect 3440 1920 3480 1930
rect 3760 2010 3800 2020
rect 3760 1930 3765 2010
rect 3795 1930 3800 2010
rect 3760 1920 3800 1930
rect 4080 2010 4120 2020
rect 4080 1930 4085 2010
rect 4115 1930 4120 2010
rect 2800 1885 2805 1915
rect 2835 1885 2840 1915
rect 2800 1880 2840 1885
rect 4080 1915 4120 1930
rect 4080 1885 4085 1915
rect 4115 1885 4120 1915
rect 4080 1880 4120 1885
rect 4160 1995 4200 2125
rect 4640 2475 4680 2480
rect 4640 2445 4645 2475
rect 4675 2445 4680 2475
rect 4640 2315 4680 2445
rect 4640 2285 4645 2315
rect 4675 2285 4680 2315
rect 4640 2155 4680 2285
rect 4640 2125 4645 2155
rect 4675 2125 4680 2155
rect 4320 2075 4520 2080
rect 4320 2045 4330 2075
rect 4510 2045 4520 2075
rect 4320 2040 4520 2045
rect 4160 1965 4165 1995
rect 4195 1965 4200 1995
rect 4160 1915 4200 1965
rect 4240 2010 4280 2020
rect 4240 1930 4245 2010
rect 4275 1930 4280 2010
rect 4240 1920 4280 1930
rect 4560 2010 4600 2020
rect 4560 1930 4565 2010
rect 4595 1930 4600 2010
rect 4160 1885 4165 1915
rect 4195 1885 4200 1915
rect 2720 1805 2725 1835
rect 2755 1805 2760 1835
rect 2720 1800 2760 1805
rect 4160 1835 4200 1885
rect 4560 1915 4600 1930
rect 4560 1885 4565 1915
rect 4595 1885 4600 1915
rect 4560 1880 4600 1885
rect 4640 1995 4680 2125
rect 4640 1965 4645 1995
rect 4675 1965 4680 1995
rect 4640 1915 4680 1965
rect 4640 1885 4645 1915
rect 4675 1885 4680 1915
rect 4160 1805 4165 1835
rect 4195 1805 4200 1835
rect 4160 1800 4200 1805
rect 4640 1835 4680 1885
rect 4640 1805 4645 1835
rect 4675 1805 4680 1835
rect 4640 1800 4680 1805
rect -480 1515 -280 1520
rect -480 1485 -470 1515
rect -290 1485 -280 1515
rect -480 1480 -280 1485
rect 0 1515 200 1520
rect 0 1485 10 1515
rect 190 1485 200 1515
rect 0 1480 200 1485
rect 320 1515 520 1520
rect 320 1485 330 1515
rect 510 1485 520 1515
rect 320 1480 520 1485
rect 640 1515 840 1520
rect 640 1485 650 1515
rect 830 1485 840 1515
rect 640 1480 840 1485
rect 960 1515 1160 1520
rect 960 1485 970 1515
rect 1150 1485 1160 1515
rect 960 1480 1160 1485
rect 1440 1515 1640 1520
rect 1440 1485 1450 1515
rect 1630 1485 1640 1515
rect 1440 1480 1640 1485
rect 1760 1515 1960 1520
rect 1760 1485 1770 1515
rect 1950 1485 1960 1515
rect 1760 1480 1960 1485
rect 2080 1515 2280 1520
rect 2080 1485 2090 1515
rect 2270 1485 2280 1515
rect 2080 1480 2280 1485
rect 2400 1515 2600 1520
rect 2400 1485 2410 1515
rect 2590 1485 2600 1515
rect 2400 1480 2600 1485
rect 2880 1515 3080 1520
rect 2880 1485 2890 1515
rect 3070 1485 3080 1515
rect 2880 1480 3080 1485
rect 3200 1515 3400 1520
rect 3200 1485 3210 1515
rect 3390 1485 3400 1515
rect 3200 1480 3400 1485
rect 3520 1515 3720 1520
rect 3520 1485 3530 1515
rect 3710 1485 3720 1515
rect 3520 1480 3720 1485
rect 3840 1515 4040 1520
rect 3840 1485 3850 1515
rect 4030 1485 4040 1515
rect 3840 1480 4040 1485
rect 4320 1515 4520 1520
rect 4320 1485 4330 1515
rect 4510 1485 4520 1515
rect 4320 1480 4520 1485
rect -560 1450 -520 1460
rect -560 1370 -555 1450
rect -525 1370 -520 1450
rect -560 1355 -520 1370
rect -560 1325 -555 1355
rect -525 1325 -520 1355
rect -560 1275 -520 1325
rect -560 1245 -555 1275
rect -525 1245 -520 1275
rect -560 1230 -520 1245
rect -560 1150 -555 1230
rect -525 1150 -520 1230
rect -560 1140 -520 1150
rect -240 1450 -200 1460
rect -240 1370 -235 1450
rect -205 1370 -200 1450
rect -240 1230 -200 1370
rect -240 1150 -235 1230
rect -205 1150 -200 1230
rect -240 1140 -200 1150
rect -80 1450 -40 1460
rect -80 1370 -75 1450
rect -45 1370 -40 1450
rect -80 1230 -40 1370
rect 240 1450 280 1460
rect 240 1370 245 1450
rect 275 1370 280 1450
rect 240 1355 280 1370
rect 240 1325 245 1355
rect 275 1325 280 1355
rect 240 1320 280 1325
rect 560 1450 600 1460
rect 560 1370 565 1450
rect 595 1370 600 1450
rect -80 1150 -75 1230
rect -45 1150 -40 1230
rect -80 1140 -40 1150
rect 240 1230 280 1240
rect 240 1150 245 1230
rect 275 1150 280 1230
rect -480 1115 -280 1120
rect -480 1085 -470 1115
rect -290 1085 -280 1115
rect -480 1080 -280 1085
rect 0 1115 200 1120
rect 0 1085 10 1115
rect 190 1085 200 1115
rect 0 1080 200 1085
rect -160 875 -120 880
rect -160 845 -155 875
rect -125 845 -120 875
rect -160 715 -120 845
rect -160 685 -155 715
rect -125 685 -120 715
rect -160 555 -120 685
rect -160 525 -155 555
rect -125 525 -120 555
rect -160 395 -120 525
rect -160 365 -155 395
rect -125 365 -120 395
rect -160 235 -120 365
rect -160 205 -155 235
rect -125 205 -120 235
rect -480 155 -280 160
rect -480 125 -470 155
rect -290 125 -280 155
rect -480 120 -280 125
rect -560 90 -520 100
rect -560 10 -555 90
rect -525 10 -520 90
rect -560 -5 -520 10
rect -240 90 -200 100
rect -240 10 -235 90
rect -205 10 -200 90
rect -240 0 -200 10
rect -160 75 -120 205
rect 80 795 120 800
rect 80 765 85 795
rect 115 765 120 795
rect 80 160 120 765
rect 240 795 280 1150
rect 560 1230 600 1370
rect 880 1450 920 1460
rect 880 1370 885 1450
rect 915 1370 920 1450
rect 880 1355 920 1370
rect 880 1325 885 1355
rect 915 1325 920 1355
rect 880 1320 920 1325
rect 1200 1450 1240 1460
rect 1200 1370 1205 1450
rect 1235 1370 1240 1450
rect 560 1150 565 1230
rect 595 1150 600 1230
rect 560 1140 600 1150
rect 880 1230 920 1240
rect 880 1150 885 1230
rect 915 1150 920 1230
rect 320 1115 520 1120
rect 320 1085 330 1115
rect 510 1085 520 1115
rect 320 1080 520 1085
rect 640 1115 840 1120
rect 640 1085 650 1115
rect 830 1085 840 1115
rect 640 1080 840 1085
rect 240 765 245 795
rect 275 765 280 795
rect 240 760 280 765
rect 400 795 440 800
rect 400 765 405 795
rect 435 765 440 795
rect 400 160 440 765
rect 720 795 760 800
rect 720 765 725 795
rect 755 765 760 795
rect 560 475 600 480
rect 560 445 565 475
rect 595 445 600 475
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 120 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 120 520 125
rect -160 45 -155 75
rect -125 45 -120 75
rect -560 -35 -555 -5
rect -525 -35 -520 -5
rect -560 -40 -520 -35
rect -160 -5 -120 45
rect -160 -35 -155 -5
rect -125 -35 -120 -5
rect -160 -85 -120 -35
rect -80 90 -40 100
rect -80 10 -75 90
rect -45 10 -40 90
rect -80 -5 -40 10
rect 240 90 280 100
rect 240 10 245 90
rect 275 10 280 90
rect 240 0 280 10
rect 560 90 600 445
rect 720 160 760 765
rect 880 795 920 1150
rect 1200 1230 1240 1370
rect 1200 1150 1205 1230
rect 1235 1150 1240 1230
rect 1200 1140 1240 1150
rect 1360 1450 1400 1460
rect 1360 1370 1365 1450
rect 1395 1370 1400 1450
rect 1360 1230 1400 1370
rect 1680 1450 1720 1460
rect 1680 1370 1685 1450
rect 1715 1370 1720 1450
rect 1680 1360 1720 1370
rect 2000 1450 2040 1460
rect 2000 1370 2005 1450
rect 2035 1370 2040 1450
rect 2000 1355 2040 1370
rect 2320 1450 2360 1460
rect 2320 1370 2325 1450
rect 2355 1370 2360 1450
rect 2320 1360 2360 1370
rect 2640 1450 2680 1460
rect 2640 1370 2645 1450
rect 2675 1370 2680 1450
rect 2000 1325 2005 1355
rect 2035 1325 2040 1355
rect 2000 1320 2040 1325
rect 1360 1150 1365 1230
rect 1395 1150 1400 1230
rect 1360 1140 1400 1150
rect 1680 1230 1720 1240
rect 1680 1150 1685 1230
rect 1715 1150 1720 1230
rect 1680 1140 1720 1150
rect 2000 1230 2040 1240
rect 2000 1150 2005 1230
rect 2035 1150 2040 1230
rect 960 1115 1160 1120
rect 960 1085 970 1115
rect 1150 1085 1160 1115
rect 960 1080 1160 1085
rect 1440 1115 1640 1120
rect 1440 1085 1450 1115
rect 1630 1085 1640 1115
rect 1440 1080 1640 1085
rect 1760 1115 1960 1120
rect 1760 1085 1770 1115
rect 1950 1085 1960 1115
rect 1760 1080 1960 1085
rect 1280 875 1320 880
rect 1280 845 1285 875
rect 1315 845 1320 875
rect 880 765 885 795
rect 915 765 920 795
rect 880 760 920 765
rect 1040 795 1080 800
rect 1040 765 1045 795
rect 1075 765 1080 795
rect 1040 160 1080 765
rect 1200 795 1240 800
rect 1200 765 1205 795
rect 1235 765 1240 795
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 120 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 120 1160 125
rect 560 10 565 90
rect 595 10 600 90
rect 560 0 600 10
rect 880 90 920 100
rect 880 10 885 90
rect 915 10 920 90
rect 880 0 920 10
rect 1200 90 1240 765
rect 1200 10 1205 90
rect 1235 10 1240 90
rect 1200 0 1240 10
rect 1280 715 1320 845
rect 1280 685 1285 715
rect 1315 685 1320 715
rect 1280 555 1320 685
rect 1280 525 1285 555
rect 1315 525 1320 555
rect 1280 395 1320 525
rect 1280 365 1285 395
rect 1315 365 1320 395
rect 1280 235 1320 365
rect 1280 205 1285 235
rect 1315 205 1320 235
rect 1280 75 1320 205
rect 1520 795 1560 800
rect 1520 765 1525 795
rect 1555 765 1560 795
rect 1520 160 1560 765
rect 1840 795 1880 800
rect 1840 765 1845 795
rect 1875 765 1880 795
rect 1840 160 1880 765
rect 2000 635 2040 1150
rect 2320 1230 2360 1240
rect 2320 1150 2325 1230
rect 2355 1150 2360 1230
rect 2320 1140 2360 1150
rect 2640 1230 2680 1370
rect 2640 1150 2645 1230
rect 2675 1150 2680 1230
rect 2640 1140 2680 1150
rect 2800 1450 2840 1460
rect 2800 1370 2805 1450
rect 2835 1370 2840 1450
rect 2800 1230 2840 1370
rect 3120 1450 3160 1460
rect 3120 1370 3125 1450
rect 3155 1370 3160 1450
rect 3120 1360 3160 1370
rect 3440 1450 3480 1460
rect 3440 1370 3445 1450
rect 3475 1370 3480 1450
rect 3440 1355 3480 1370
rect 3760 1450 3800 1460
rect 3760 1370 3765 1450
rect 3795 1370 3800 1450
rect 3760 1360 3800 1370
rect 4080 1450 4120 1460
rect 4080 1370 4085 1450
rect 4115 1370 4120 1450
rect 3440 1325 3445 1355
rect 3475 1325 3480 1355
rect 3440 1320 3480 1325
rect 2800 1150 2805 1230
rect 2835 1150 2840 1230
rect 2800 1140 2840 1150
rect 3120 1230 3160 1240
rect 3120 1150 3125 1230
rect 3155 1150 3160 1230
rect 3120 1140 3160 1150
rect 3440 1230 3480 1240
rect 3440 1150 3445 1230
rect 3475 1150 3480 1230
rect 2080 1115 2280 1120
rect 2080 1085 2090 1115
rect 2270 1085 2280 1115
rect 2080 1080 2280 1085
rect 2400 1115 2600 1120
rect 2400 1085 2410 1115
rect 2590 1085 2600 1115
rect 2400 1080 2600 1085
rect 2880 1115 3080 1120
rect 2880 1085 2890 1115
rect 3070 1085 3080 1115
rect 2880 1080 3080 1085
rect 3200 1115 3400 1120
rect 3200 1085 3210 1115
rect 3390 1085 3400 1115
rect 3200 1080 3400 1085
rect 2720 875 2760 880
rect 2720 845 2725 875
rect 2755 845 2760 875
rect 2720 715 2760 845
rect 2720 685 2725 715
rect 2755 685 2760 715
rect 2000 605 2005 635
rect 2035 605 2040 635
rect 2000 600 2040 605
rect 2160 635 2200 640
rect 2160 605 2165 635
rect 2195 605 2200 635
rect 2000 475 2040 480
rect 2000 445 2005 475
rect 2035 445 2040 475
rect 1440 155 1640 160
rect 1440 125 1450 155
rect 1630 125 1640 155
rect 1440 120 1640 125
rect 1760 155 1960 160
rect 1760 125 1770 155
rect 1950 125 1960 155
rect 1760 120 1960 125
rect 1280 45 1285 75
rect 1315 45 1320 75
rect -80 -35 -75 -5
rect -45 -35 -40 -5
rect -80 -40 -40 -35
rect 1280 -5 1320 45
rect 1280 -35 1285 -5
rect 1315 -35 1320 -5
rect -160 -115 -155 -85
rect -125 -115 -120 -85
rect -160 -120 -120 -115
rect 1280 -85 1320 -35
rect 1360 90 1400 100
rect 1360 10 1365 90
rect 1395 10 1400 90
rect 1360 -5 1400 10
rect 1680 90 1720 100
rect 1680 10 1685 90
rect 1715 10 1720 90
rect 1680 0 1720 10
rect 2000 90 2040 445
rect 2160 160 2200 605
rect 2480 635 2520 640
rect 2480 605 2485 635
rect 2515 605 2520 635
rect 2480 160 2520 605
rect 2640 635 2680 640
rect 2640 605 2645 635
rect 2675 605 2680 635
rect 2080 155 2280 160
rect 2080 125 2090 155
rect 2270 125 2280 155
rect 2080 120 2280 125
rect 2400 155 2600 160
rect 2400 125 2410 155
rect 2590 125 2600 155
rect 2400 120 2600 125
rect 2000 10 2005 90
rect 2035 10 2040 90
rect 2000 0 2040 10
rect 2320 90 2360 100
rect 2320 10 2325 90
rect 2355 10 2360 90
rect 2320 0 2360 10
rect 2640 90 2680 605
rect 2640 10 2645 90
rect 2675 10 2680 90
rect 2640 0 2680 10
rect 2720 555 2760 685
rect 2720 525 2725 555
rect 2755 525 2760 555
rect 2720 395 2760 525
rect 2720 365 2725 395
rect 2755 365 2760 395
rect 2720 235 2760 365
rect 2720 205 2725 235
rect 2755 205 2760 235
rect 2720 75 2760 205
rect 2960 315 3000 320
rect 2960 285 2965 315
rect 2995 285 3000 315
rect 2960 160 3000 285
rect 3280 315 3320 320
rect 3280 285 3285 315
rect 3315 285 3320 315
rect 3280 160 3320 285
rect 3440 315 3480 1150
rect 3760 1230 3800 1240
rect 3760 1150 3765 1230
rect 3795 1150 3800 1230
rect 3760 1140 3800 1150
rect 4080 1230 4120 1370
rect 4080 1150 4085 1230
rect 4115 1150 4120 1230
rect 4080 1140 4120 1150
rect 4240 1450 4280 1460
rect 4240 1370 4245 1450
rect 4275 1370 4280 1450
rect 4240 1230 4280 1370
rect 4240 1150 4245 1230
rect 4275 1150 4280 1230
rect 4240 1140 4280 1150
rect 4560 1450 4600 1460
rect 4560 1370 4565 1450
rect 4595 1370 4600 1450
rect 4560 1355 4600 1370
rect 4560 1325 4565 1355
rect 4595 1325 4600 1355
rect 4560 1275 4600 1325
rect 4560 1245 4565 1275
rect 4595 1245 4600 1275
rect 4560 1230 4600 1245
rect 4560 1150 4565 1230
rect 4595 1150 4600 1230
rect 4560 1140 4600 1150
rect 3520 1115 3720 1120
rect 3520 1085 3530 1115
rect 3710 1085 3720 1115
rect 3520 1080 3720 1085
rect 3840 1115 4040 1120
rect 3840 1085 3850 1115
rect 4030 1085 4040 1115
rect 3840 1080 4040 1085
rect 4320 1115 4520 1120
rect 4320 1085 4330 1115
rect 4510 1085 4520 1115
rect 4320 1080 4520 1085
rect 4160 875 4200 880
rect 4160 845 4165 875
rect 4195 845 4200 875
rect 4160 715 4200 845
rect 4160 685 4165 715
rect 4195 685 4200 715
rect 4160 555 4200 685
rect 4160 525 4165 555
rect 4195 525 4200 555
rect 4160 395 4200 525
rect 4160 365 4165 395
rect 4195 365 4200 395
rect 3440 285 3445 315
rect 3475 285 3480 315
rect 3440 280 3480 285
rect 3600 315 3640 320
rect 3600 285 3605 315
rect 3635 285 3640 315
rect 3600 160 3640 285
rect 3920 315 3960 320
rect 3920 285 3925 315
rect 3955 285 3960 315
rect 3920 160 3960 285
rect 4080 315 4120 320
rect 4080 285 4085 315
rect 4115 285 4120 315
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 120 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 120 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 120 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 120 4040 125
rect 2720 45 2725 75
rect 2755 45 2760 75
rect 1360 -35 1365 -5
rect 1395 -35 1400 -5
rect 1360 -40 1400 -35
rect 2720 -5 2760 45
rect 2720 -35 2725 -5
rect 2755 -35 2760 -5
rect 1280 -115 1285 -85
rect 1315 -115 1320 -85
rect 1280 -120 1320 -115
rect 2720 -85 2760 -35
rect 2800 90 2840 100
rect 2800 10 2805 90
rect 2835 10 2840 90
rect 2800 -5 2840 10
rect 3120 90 3160 100
rect 3120 10 3125 90
rect 3155 10 3160 90
rect 3120 0 3160 10
rect 3440 90 3480 100
rect 3440 10 3445 90
rect 3475 10 3480 90
rect 3440 0 3480 10
rect 3760 90 3800 100
rect 3760 10 3765 90
rect 3795 10 3800 90
rect 3760 0 3800 10
rect 4080 90 4120 285
rect 4080 10 4085 90
rect 4115 10 4120 90
rect 4080 0 4120 10
rect 4160 235 4200 365
rect 4160 205 4165 235
rect 4195 205 4200 235
rect 4160 75 4200 205
rect 4640 875 4680 880
rect 4640 845 4645 875
rect 4675 845 4680 875
rect 4640 715 4680 845
rect 4640 685 4645 715
rect 4675 685 4680 715
rect 4640 555 4680 685
rect 4640 525 4645 555
rect 4675 525 4680 555
rect 4640 395 4680 525
rect 4640 365 4645 395
rect 4675 365 4680 395
rect 4640 235 4680 365
rect 4640 205 4645 235
rect 4675 205 4680 235
rect 4320 155 4520 160
rect 4320 125 4330 155
rect 4510 125 4520 155
rect 4320 120 4520 125
rect 4160 45 4165 75
rect 4195 45 4200 75
rect 2800 -35 2805 -5
rect 2835 -35 2840 -5
rect 2800 -40 2840 -35
rect 4160 -5 4200 45
rect 4240 90 4280 100
rect 4240 10 4245 90
rect 4275 10 4280 90
rect 4240 0 4280 10
rect 4560 90 4600 100
rect 4560 10 4565 90
rect 4595 10 4600 90
rect 4160 -35 4165 -5
rect 4195 -35 4200 -5
rect 2720 -115 2725 -85
rect 2755 -115 2760 -85
rect 2720 -120 2760 -115
rect 4160 -85 4200 -35
rect 4560 -5 4600 10
rect 4560 -35 4565 -5
rect 4595 -35 4600 -5
rect 4560 -40 4600 -35
rect 4640 75 4680 205
rect 4640 45 4645 75
rect 4675 45 4680 75
rect 4640 -5 4680 45
rect 4640 -35 4645 -5
rect 4675 -35 4680 -5
rect 4160 -115 4165 -85
rect 4195 -115 4200 -85
rect 4160 -120 4200 -115
rect 4640 -85 4680 -35
rect 4640 -115 4645 -85
rect 4675 -115 4680 -85
rect 4640 -120 4680 -115
<< via1 >>
rect 10 5325 190 5355
rect 330 5325 510 5355
rect 650 5325 830 5355
rect 970 5325 1150 5355
rect -555 5165 -525 5195
rect -555 5085 -525 5115
rect 565 5245 595 5275
rect 565 5165 595 5195
rect 10 4925 190 4955
rect 330 4925 510 4955
rect 85 4765 115 4795
rect -75 4125 -45 4155
rect -795 4045 -765 4075
rect -795 3885 -765 3915
rect -795 3805 -765 3835
rect -555 3885 -525 3915
rect -155 3885 -125 3915
rect -555 3805 -525 3835
rect 405 4765 435 4795
rect 245 4525 275 4555
rect 1365 5165 1395 5195
rect 1365 5085 1395 5115
rect 2005 5245 2035 5275
rect 2645 5165 2675 5195
rect 2645 5085 2675 5115
rect 2805 5245 2835 5275
rect 2805 5165 2835 5195
rect 2805 5085 2835 5115
rect 2805 5005 2835 5035
rect 4085 5165 4115 5195
rect 4085 5085 4115 5115
rect 4565 5165 4595 5195
rect 4565 5085 4595 5115
rect 650 4925 830 4955
rect 970 4925 1150 4955
rect 565 4285 595 4315
rect 725 4765 755 4795
rect 565 4125 595 4155
rect 1045 4765 1075 4795
rect 885 4525 915 4555
rect 1525 4765 1555 4795
rect 1205 4125 1235 4155
rect 1365 4125 1395 4155
rect 1285 3885 1315 3915
rect -155 3805 -125 3835
rect -795 3725 -765 3755
rect -155 3725 -125 3755
rect 1285 3805 1315 3835
rect 1845 4765 1875 4795
rect 1685 4525 1715 4555
rect 2165 4765 2195 4795
rect 2005 4125 2035 4155
rect 2485 4765 2515 4795
rect 2325 4525 2355 4555
rect 2965 4765 2995 4795
rect 3285 4765 3315 4795
rect 3605 4765 3635 4795
rect 3925 4765 3955 4795
rect 4085 4765 4115 4795
rect 2645 4125 2675 4155
rect 2965 4125 2995 4155
rect 3285 4125 3315 4155
rect 3605 4125 3635 4155
rect 3925 4125 3955 4155
rect 2725 3885 2755 3915
rect 2725 3805 2755 3835
rect 1285 3725 1315 3755
rect 2805 3885 2835 3915
rect 4165 3885 4195 3915
rect 2805 3805 2835 3835
rect 4565 3885 4595 3915
rect 4165 3805 4195 3835
rect 2725 3725 2755 3755
rect 4565 3805 4595 3835
rect 4645 3885 4675 3915
rect 4645 3805 4675 3835
rect 4165 3725 4195 3755
rect 4645 3725 4675 3755
rect -795 3645 -765 3675
rect 10 3405 190 3435
rect 330 3405 510 3435
rect 650 3405 830 3435
rect 970 3405 1150 3435
rect 1450 3405 1630 3435
rect 1770 3405 1950 3435
rect 2090 3405 2270 3435
rect 2410 3405 2590 3435
rect -555 3245 -525 3275
rect -555 3165 -525 3195
rect 565 3325 595 3355
rect 565 3245 595 3275
rect 10 3005 190 3035
rect 330 3005 510 3035
rect 2005 3325 2035 3355
rect 2005 3245 2035 3275
rect 650 3005 830 3035
rect 970 3005 1150 3035
rect 1450 3005 1630 3035
rect 1770 3005 1950 3035
rect 2805 3325 2835 3355
rect 2805 3245 2835 3275
rect 2805 3165 2835 3195
rect 2805 3085 2835 3115
rect 2090 3005 2270 3035
rect 2410 3005 2590 3035
rect 2890 3005 3070 3035
rect 3210 3005 3390 3035
rect 3445 3005 3475 3035
rect 2005 2845 2035 2875
rect 2645 2845 2675 2875
rect 565 2605 595 2635
rect 1205 2605 1235 2635
rect -155 2445 -125 2475
rect -155 2285 -125 2315
rect -155 2125 -125 2155
rect -555 1965 -525 1995
rect 85 2365 115 2395
rect 405 2365 435 2395
rect 725 2365 755 2395
rect 1045 2365 1075 2395
rect -155 1965 -125 1995
rect -555 1885 -525 1915
rect -155 1885 -125 1915
rect -75 1965 -45 1995
rect 1285 2445 1315 2475
rect 1285 2285 1315 2315
rect 1285 2125 1315 2155
rect 1525 2205 1555 2235
rect 1845 2205 1875 2235
rect 2165 2205 2195 2235
rect 2485 2205 2515 2235
rect 1285 1965 1315 1995
rect -75 1885 -45 1915
rect 1285 1885 1315 1915
rect -155 1805 -125 1835
rect 1365 1965 1395 1995
rect 2725 2445 2755 2475
rect 2725 2285 2755 2315
rect 2725 2125 2755 2155
rect 2965 2205 2995 2235
rect 3285 2205 3315 2235
rect 2725 1965 2755 1995
rect 1365 1885 1395 1915
rect 2725 1885 2755 1915
rect 1285 1805 1315 1835
rect 2805 1965 2835 1995
rect 3530 3005 3710 3035
rect 3850 3005 4030 3035
rect 4565 3245 4595 3275
rect 4565 3165 4595 3195
rect 4085 3005 4115 3035
rect 4165 2445 4195 2475
rect 4165 2285 4195 2315
rect 3605 2205 3635 2235
rect 3925 2205 3955 2235
rect 4165 2125 4195 2155
rect 4085 1965 4115 1995
rect 2805 1885 2835 1915
rect 4085 1885 4115 1915
rect 4645 2445 4675 2475
rect 4645 2285 4675 2315
rect 4645 2125 4675 2155
rect 4165 1965 4195 1995
rect 4565 1965 4595 1995
rect 4165 1885 4195 1915
rect 2725 1805 2755 1835
rect 4565 1885 4595 1915
rect 4645 1965 4675 1995
rect 4645 1885 4675 1915
rect 4165 1805 4195 1835
rect 4645 1805 4675 1835
rect 10 1485 190 1515
rect 330 1485 510 1515
rect 650 1485 830 1515
rect 970 1485 1150 1515
rect 1450 1485 1630 1515
rect 1770 1485 1950 1515
rect 2090 1485 2270 1515
rect 2410 1485 2590 1515
rect 2890 1485 3070 1515
rect 3210 1485 3390 1515
rect 3530 1485 3710 1515
rect 3850 1485 4030 1515
rect -555 1325 -525 1355
rect -555 1245 -525 1275
rect 245 1405 275 1435
rect 245 1325 275 1355
rect 10 1085 190 1115
rect -155 845 -125 875
rect -155 685 -125 715
rect -155 525 -125 555
rect -155 365 -125 395
rect -155 205 -125 235
rect -555 45 -525 75
rect 85 765 115 795
rect 885 1405 915 1435
rect 885 1325 915 1355
rect 330 1085 510 1115
rect 650 1085 830 1115
rect 245 765 275 795
rect 405 765 435 795
rect 725 765 755 795
rect 565 445 595 475
rect -155 45 -125 75
rect -555 -35 -525 -5
rect -155 -35 -125 -5
rect -75 45 -45 75
rect 2005 1405 2035 1435
rect 2005 1325 2035 1355
rect 970 1085 1150 1115
rect 1450 1085 1630 1115
rect 1770 1085 1950 1115
rect 1285 845 1315 875
rect 885 765 915 795
rect 1045 765 1075 795
rect 1205 765 1235 795
rect 1285 685 1315 715
rect 1285 525 1315 555
rect 1285 365 1315 395
rect 1285 205 1315 235
rect 1525 765 1555 795
rect 1845 765 1875 795
rect 3445 1405 3475 1435
rect 3445 1325 3475 1355
rect 2090 1085 2270 1115
rect 2410 1085 2590 1115
rect 2890 1085 3070 1115
rect 3210 1085 3390 1115
rect 2725 845 2755 875
rect 2725 685 2755 715
rect 2005 605 2035 635
rect 2165 605 2195 635
rect 2005 445 2035 475
rect 1285 45 1315 75
rect -75 -35 -45 -5
rect 1285 -35 1315 -5
rect -155 -115 -125 -85
rect 1365 45 1395 75
rect 2485 605 2515 635
rect 2645 605 2675 635
rect 2725 525 2755 555
rect 2725 365 2755 395
rect 2725 205 2755 235
rect 2965 285 2995 315
rect 3285 285 3315 315
rect 4565 1325 4595 1355
rect 4565 1245 4595 1275
rect 3530 1085 3710 1115
rect 3850 1085 4030 1115
rect 4165 845 4195 875
rect 4165 685 4195 715
rect 4165 525 4195 555
rect 4165 365 4195 395
rect 3445 285 3475 315
rect 3605 285 3635 315
rect 3925 285 3955 315
rect 4085 285 4115 315
rect 2725 45 2755 75
rect 1365 -35 1395 -5
rect 2725 -35 2755 -5
rect 1285 -115 1315 -85
rect 2805 45 2835 75
rect 4165 205 4195 235
rect 4645 845 4675 875
rect 4645 685 4675 715
rect 4645 525 4675 555
rect 4645 365 4675 395
rect 4645 205 4675 235
rect 4165 45 4195 75
rect 2805 -35 2835 -5
rect 4565 45 4595 75
rect 4165 -35 4195 -5
rect 2725 -115 2755 -85
rect 4565 -35 4595 -5
rect 4645 45 4675 75
rect 4645 -35 4675 -5
rect 4165 -115 4195 -85
rect 4645 -115 4675 -85
<< metal2 >>
rect -1520 5595 -840 5600
rect -1520 5565 -1515 5595
rect -1485 5565 -1355 5595
rect -1325 5565 -1195 5595
rect -1165 5565 -1035 5595
rect -1005 5565 -875 5595
rect -845 5565 -840 5595
rect -1520 5560 -840 5565
rect -800 5595 5720 5600
rect -800 5565 4885 5595
rect 4915 5565 5045 5595
rect 5075 5565 5205 5595
rect 5235 5565 5365 5595
rect 5395 5565 5525 5595
rect 5555 5565 5685 5595
rect 5715 5565 5720 5595
rect -800 5560 5720 5565
rect -1520 5515 4840 5520
rect -1520 5485 -1515 5515
rect -1485 5485 -1355 5515
rect -1325 5485 -1195 5515
rect -1165 5485 -1035 5515
rect -1005 5485 -875 5515
rect -845 5485 -795 5515
rect -765 5485 -715 5515
rect -685 5485 -635 5515
rect -605 5485 -555 5515
rect -525 5485 -475 5515
rect -445 5485 -395 5515
rect -365 5485 -315 5515
rect -285 5485 -235 5515
rect -205 5485 -155 5515
rect -125 5485 -75 5515
rect -45 5485 5 5515
rect 35 5485 85 5515
rect 115 5485 165 5515
rect 195 5485 245 5515
rect 275 5485 325 5515
rect 355 5485 405 5515
rect 435 5485 485 5515
rect 515 5485 565 5515
rect 595 5485 645 5515
rect 675 5485 725 5515
rect 755 5485 805 5515
rect 835 5485 885 5515
rect 915 5485 965 5515
rect 995 5485 1045 5515
rect 1075 5485 1125 5515
rect 1155 5485 1205 5515
rect 1235 5485 1285 5515
rect 1315 5485 1365 5515
rect 1395 5485 1445 5515
rect 1475 5485 1525 5515
rect 1555 5485 1605 5515
rect 1635 5485 1685 5515
rect 1715 5485 1765 5515
rect 1795 5485 1845 5515
rect 1875 5485 1925 5515
rect 1955 5485 2005 5515
rect 2035 5485 2085 5515
rect 2115 5485 2165 5515
rect 2195 5485 2245 5515
rect 2275 5485 2325 5515
rect 2355 5485 2405 5515
rect 2435 5485 2485 5515
rect 2515 5485 2565 5515
rect 2595 5485 2645 5515
rect 2675 5485 2725 5515
rect 2755 5485 2805 5515
rect 2835 5485 2885 5515
rect 2915 5485 2965 5515
rect 2995 5485 3045 5515
rect 3075 5485 3125 5515
rect 3155 5485 3205 5515
rect 3235 5485 3285 5515
rect 3315 5485 3365 5515
rect 3395 5485 3445 5515
rect 3475 5485 3525 5515
rect 3555 5485 3605 5515
rect 3635 5485 3685 5515
rect 3715 5485 3765 5515
rect 3795 5485 3845 5515
rect 3875 5485 3925 5515
rect 3955 5485 4005 5515
rect 4035 5485 4085 5515
rect 4115 5485 4165 5515
rect 4195 5485 4245 5515
rect 4275 5485 4325 5515
rect 4355 5485 4405 5515
rect 4435 5485 4485 5515
rect 4515 5485 4565 5515
rect 4595 5485 4645 5515
rect 4675 5485 4725 5515
rect 4755 5485 4805 5515
rect 4835 5485 4840 5515
rect -1520 5480 4840 5485
rect 4880 5515 5720 5520
rect 4880 5485 4885 5515
rect 4915 5485 5045 5515
rect 5075 5485 5205 5515
rect 5235 5485 5365 5515
rect 5395 5485 5525 5515
rect 5555 5485 5685 5515
rect 5715 5485 5720 5515
rect 4880 5480 5720 5485
rect -1520 5435 4840 5440
rect -1520 5405 -1515 5435
rect -1485 5405 -1355 5435
rect -1325 5405 -1195 5435
rect -1165 5405 -1035 5435
rect -1005 5405 -875 5435
rect -845 5405 -795 5435
rect -765 5405 -715 5435
rect -685 5405 -635 5435
rect -605 5405 -555 5435
rect -525 5405 -475 5435
rect -445 5405 -395 5435
rect -365 5405 -315 5435
rect -285 5405 -235 5435
rect -205 5405 -155 5435
rect -125 5405 -75 5435
rect -45 5405 5 5435
rect 35 5405 85 5435
rect 115 5405 165 5435
rect 195 5405 245 5435
rect 275 5405 325 5435
rect 355 5405 405 5435
rect 435 5405 485 5435
rect 515 5405 565 5435
rect 595 5405 645 5435
rect 675 5405 725 5435
rect 755 5405 805 5435
rect 835 5405 885 5435
rect 915 5405 965 5435
rect 995 5405 1045 5435
rect 1075 5405 1125 5435
rect 1155 5405 1205 5435
rect 1235 5405 1285 5435
rect 1315 5405 1365 5435
rect 1395 5405 1445 5435
rect 1475 5405 1525 5435
rect 1555 5405 1605 5435
rect 1635 5405 1685 5435
rect 1715 5405 1765 5435
rect 1795 5405 1845 5435
rect 1875 5405 1925 5435
rect 1955 5405 2005 5435
rect 2035 5405 2085 5435
rect 2115 5405 2165 5435
rect 2195 5405 2245 5435
rect 2275 5405 2325 5435
rect 2355 5405 2405 5435
rect 2435 5405 2485 5435
rect 2515 5405 2565 5435
rect 2595 5405 2645 5435
rect 2675 5405 2725 5435
rect 2755 5405 2805 5435
rect 2835 5405 2885 5435
rect 2915 5405 2965 5435
rect 2995 5405 3045 5435
rect 3075 5405 3125 5435
rect 3155 5405 3205 5435
rect 3235 5405 3285 5435
rect 3315 5405 3365 5435
rect 3395 5405 3445 5435
rect 3475 5405 3525 5435
rect 3555 5405 3605 5435
rect 3635 5405 3685 5435
rect 3715 5405 3765 5435
rect 3795 5405 3845 5435
rect 3875 5405 3925 5435
rect 3955 5405 4005 5435
rect 4035 5405 4085 5435
rect 4115 5405 4165 5435
rect 4195 5405 4245 5435
rect 4275 5405 4325 5435
rect 4355 5405 4405 5435
rect 4435 5405 4485 5435
rect 4515 5405 4565 5435
rect 4595 5405 4645 5435
rect 4675 5405 4725 5435
rect 4755 5405 4805 5435
rect 4835 5405 4840 5435
rect -1520 5400 4840 5405
rect 4880 5435 5720 5440
rect 4880 5405 4885 5435
rect 4915 5405 5045 5435
rect 5075 5405 5205 5435
rect 5235 5405 5365 5435
rect 5395 5405 5525 5435
rect 5555 5405 5685 5435
rect 5715 5405 5720 5435
rect 4880 5400 5720 5405
rect -1520 5355 -1000 5360
rect -1520 5325 -1515 5355
rect -1485 5325 -1355 5355
rect -1325 5325 -1195 5355
rect -1165 5325 -1035 5355
rect -1005 5325 -1000 5355
rect -1520 5320 -1000 5325
rect -960 5355 4840 5360
rect -960 5325 -955 5355
rect -925 5325 10 5355
rect 190 5325 330 5355
rect 510 5325 650 5355
rect 830 5325 970 5355
rect 1150 5325 4840 5355
rect -960 5320 4840 5325
rect 4880 5355 5720 5360
rect 4880 5325 4885 5355
rect 4915 5325 5045 5355
rect 5075 5325 5205 5355
rect 5235 5325 5365 5355
rect 5395 5325 5525 5355
rect 5555 5325 5685 5355
rect 5715 5325 5720 5355
rect 4880 5320 5720 5325
rect -1520 5275 4840 5280
rect -1520 5245 -1515 5275
rect -1485 5245 -1355 5275
rect -1325 5245 -1195 5275
rect -1165 5245 -1035 5275
rect -1005 5245 -875 5275
rect -845 5245 -795 5275
rect -765 5245 -715 5275
rect -685 5245 -635 5275
rect -605 5245 -555 5275
rect -525 5245 -475 5275
rect -445 5245 -395 5275
rect -365 5245 -315 5275
rect -285 5245 -235 5275
rect -205 5245 -155 5275
rect -125 5245 -75 5275
rect -45 5245 5 5275
rect 35 5245 85 5275
rect 115 5245 165 5275
rect 195 5245 245 5275
rect 275 5245 325 5275
rect 355 5245 405 5275
rect 435 5245 485 5275
rect 515 5245 565 5275
rect 595 5245 645 5275
rect 675 5245 725 5275
rect 755 5245 805 5275
rect 835 5245 885 5275
rect 915 5245 965 5275
rect 995 5245 1045 5275
rect 1075 5245 1125 5275
rect 1155 5245 1205 5275
rect 1235 5245 1285 5275
rect 1315 5245 1365 5275
rect 1395 5245 1445 5275
rect 1475 5245 1525 5275
rect 1555 5245 1605 5275
rect 1635 5245 1685 5275
rect 1715 5245 1765 5275
rect 1795 5245 1845 5275
rect 1875 5245 1925 5275
rect 1955 5245 2005 5275
rect 2035 5245 2085 5275
rect 2115 5245 2165 5275
rect 2195 5245 2245 5275
rect 2275 5245 2325 5275
rect 2355 5245 2405 5275
rect 2435 5245 2485 5275
rect 2515 5245 2565 5275
rect 2595 5245 2645 5275
rect 2675 5245 2725 5275
rect 2755 5245 2805 5275
rect 2835 5245 2885 5275
rect 2915 5245 2965 5275
rect 2995 5245 3045 5275
rect 3075 5245 3125 5275
rect 3155 5245 3205 5275
rect 3235 5245 3285 5275
rect 3315 5245 3365 5275
rect 3395 5245 3445 5275
rect 3475 5245 3525 5275
rect 3555 5245 3605 5275
rect 3635 5245 3685 5275
rect 3715 5245 3765 5275
rect 3795 5245 3845 5275
rect 3875 5245 3925 5275
rect 3955 5245 4005 5275
rect 4035 5245 4085 5275
rect 4115 5245 4165 5275
rect 4195 5245 4245 5275
rect 4275 5245 4325 5275
rect 4355 5245 4405 5275
rect 4435 5245 4485 5275
rect 4515 5245 4565 5275
rect 4595 5245 4645 5275
rect 4675 5245 4725 5275
rect 4755 5245 4805 5275
rect 4835 5245 4840 5275
rect -1520 5240 4840 5245
rect 4880 5275 5720 5280
rect 4880 5245 4885 5275
rect 4915 5245 5045 5275
rect 5075 5245 5205 5275
rect 5235 5245 5365 5275
rect 5395 5245 5525 5275
rect 5555 5245 5685 5275
rect 5715 5245 5720 5275
rect 4880 5240 5720 5245
rect -1520 5195 4840 5200
rect -1520 5165 -1515 5195
rect -1485 5165 -1355 5195
rect -1325 5165 -1195 5195
rect -1165 5165 -1035 5195
rect -1005 5165 -875 5195
rect -845 5165 -795 5195
rect -765 5165 -715 5195
rect -685 5165 -635 5195
rect -605 5165 -555 5195
rect -525 5165 -475 5195
rect -445 5165 -395 5195
rect -365 5165 -315 5195
rect -285 5165 -235 5195
rect -205 5165 -155 5195
rect -125 5165 -75 5195
rect -45 5165 5 5195
rect 35 5165 85 5195
rect 115 5165 165 5195
rect 195 5165 245 5195
rect 275 5165 325 5195
rect 355 5165 405 5195
rect 435 5165 485 5195
rect 515 5165 565 5195
rect 595 5165 645 5195
rect 675 5165 725 5195
rect 755 5165 805 5195
rect 835 5165 885 5195
rect 915 5165 965 5195
rect 995 5165 1045 5195
rect 1075 5165 1125 5195
rect 1155 5165 1205 5195
rect 1235 5165 1285 5195
rect 1315 5165 1365 5195
rect 1395 5165 1445 5195
rect 1475 5165 1525 5195
rect 1555 5165 1605 5195
rect 1635 5165 1685 5195
rect 1715 5165 1765 5195
rect 1795 5165 1845 5195
rect 1875 5165 1925 5195
rect 1955 5165 2005 5195
rect 2035 5165 2085 5195
rect 2115 5165 2165 5195
rect 2195 5165 2245 5195
rect 2275 5165 2325 5195
rect 2355 5165 2405 5195
rect 2435 5165 2485 5195
rect 2515 5165 2565 5195
rect 2595 5165 2645 5195
rect 2675 5165 2725 5195
rect 2755 5165 2805 5195
rect 2835 5165 2885 5195
rect 2915 5165 2965 5195
rect 2995 5165 3045 5195
rect 3075 5165 3125 5195
rect 3155 5165 3205 5195
rect 3235 5165 3285 5195
rect 3315 5165 3365 5195
rect 3395 5165 3445 5195
rect 3475 5165 3525 5195
rect 3555 5165 3605 5195
rect 3635 5165 3685 5195
rect 3715 5165 3765 5195
rect 3795 5165 3845 5195
rect 3875 5165 3925 5195
rect 3955 5165 4005 5195
rect 4035 5165 4085 5195
rect 4115 5165 4165 5195
rect 4195 5165 4245 5195
rect 4275 5165 4325 5195
rect 4355 5165 4405 5195
rect 4435 5165 4485 5195
rect 4515 5165 4565 5195
rect 4595 5165 4645 5195
rect 4675 5165 4725 5195
rect 4755 5165 4805 5195
rect 4835 5165 4840 5195
rect -1520 5160 4840 5165
rect 4880 5195 5720 5200
rect 4880 5165 4885 5195
rect 4915 5165 5045 5195
rect 5075 5165 5205 5195
rect 5235 5165 5365 5195
rect 5395 5165 5525 5195
rect 5555 5165 5685 5195
rect 5715 5165 5720 5195
rect 4880 5160 5720 5165
rect -1520 5115 4840 5120
rect -1520 5085 -1515 5115
rect -1485 5085 -1355 5115
rect -1325 5085 -1195 5115
rect -1165 5085 -1035 5115
rect -1005 5085 -875 5115
rect -845 5085 -795 5115
rect -765 5085 -715 5115
rect -685 5085 -635 5115
rect -605 5085 -555 5115
rect -525 5085 -475 5115
rect -445 5085 -395 5115
rect -365 5085 -315 5115
rect -285 5085 -235 5115
rect -205 5085 -155 5115
rect -125 5085 -75 5115
rect -45 5085 5 5115
rect 35 5085 85 5115
rect 115 5085 165 5115
rect 195 5085 245 5115
rect 275 5085 325 5115
rect 355 5085 405 5115
rect 435 5085 485 5115
rect 515 5085 565 5115
rect 595 5085 645 5115
rect 675 5085 725 5115
rect 755 5085 805 5115
rect 835 5085 885 5115
rect 915 5085 965 5115
rect 995 5085 1045 5115
rect 1075 5085 1125 5115
rect 1155 5085 1205 5115
rect 1235 5085 1285 5115
rect 1315 5085 1365 5115
rect 1395 5085 1445 5115
rect 1475 5085 1525 5115
rect 1555 5085 1605 5115
rect 1635 5085 1685 5115
rect 1715 5085 1765 5115
rect 1795 5085 1845 5115
rect 1875 5085 1925 5115
rect 1955 5085 2005 5115
rect 2035 5085 2085 5115
rect 2115 5085 2165 5115
rect 2195 5085 2245 5115
rect 2275 5085 2325 5115
rect 2355 5085 2405 5115
rect 2435 5085 2485 5115
rect 2515 5085 2565 5115
rect 2595 5085 2645 5115
rect 2675 5085 2725 5115
rect 2755 5085 2805 5115
rect 2835 5085 2885 5115
rect 2915 5085 2965 5115
rect 2995 5085 3045 5115
rect 3075 5085 3125 5115
rect 3155 5085 3205 5115
rect 3235 5085 3285 5115
rect 3315 5085 3365 5115
rect 3395 5085 3445 5115
rect 3475 5085 3525 5115
rect 3555 5085 3605 5115
rect 3635 5085 3685 5115
rect 3715 5085 3765 5115
rect 3795 5085 3845 5115
rect 3875 5085 3925 5115
rect 3955 5085 4005 5115
rect 4035 5085 4085 5115
rect 4115 5085 4165 5115
rect 4195 5085 4245 5115
rect 4275 5085 4325 5115
rect 4355 5085 4405 5115
rect 4435 5085 4485 5115
rect 4515 5085 4565 5115
rect 4595 5085 4645 5115
rect 4675 5085 4725 5115
rect 4755 5085 4805 5115
rect 4835 5085 4840 5115
rect -1520 5080 4840 5085
rect 4880 5115 5720 5120
rect 4880 5085 4885 5115
rect 4915 5085 5045 5115
rect 5075 5085 5205 5115
rect 5235 5085 5365 5115
rect 5395 5085 5525 5115
rect 5555 5085 5685 5115
rect 5715 5085 5720 5115
rect 4880 5080 5720 5085
rect -1520 5035 4840 5040
rect -1520 5005 -1515 5035
rect -1485 5005 -1355 5035
rect -1325 5005 -1195 5035
rect -1165 5005 -1035 5035
rect -1005 5005 -875 5035
rect -845 5005 -795 5035
rect -765 5005 -715 5035
rect -685 5005 -635 5035
rect -605 5005 -555 5035
rect -525 5005 -475 5035
rect -445 5005 -395 5035
rect -365 5005 -315 5035
rect -285 5005 -235 5035
rect -205 5005 -155 5035
rect -125 5005 -75 5035
rect -45 5005 5 5035
rect 35 5005 85 5035
rect 115 5005 165 5035
rect 195 5005 245 5035
rect 275 5005 325 5035
rect 355 5005 405 5035
rect 435 5005 485 5035
rect 515 5005 565 5035
rect 595 5005 645 5035
rect 675 5005 725 5035
rect 755 5005 805 5035
rect 835 5005 885 5035
rect 915 5005 965 5035
rect 995 5005 1045 5035
rect 1075 5005 1125 5035
rect 1155 5005 1205 5035
rect 1235 5005 1285 5035
rect 1315 5005 1365 5035
rect 1395 5005 1445 5035
rect 1475 5005 1525 5035
rect 1555 5005 1605 5035
rect 1635 5005 1685 5035
rect 1715 5005 1765 5035
rect 1795 5005 1845 5035
rect 1875 5005 1925 5035
rect 1955 5005 2005 5035
rect 2035 5005 2085 5035
rect 2115 5005 2165 5035
rect 2195 5005 2245 5035
rect 2275 5005 2325 5035
rect 2355 5005 2405 5035
rect 2435 5005 2485 5035
rect 2515 5005 2565 5035
rect 2595 5005 2645 5035
rect 2675 5005 2725 5035
rect 2755 5005 2805 5035
rect 2835 5005 2885 5035
rect 2915 5005 2965 5035
rect 2995 5005 3045 5035
rect 3075 5005 3125 5035
rect 3155 5005 3205 5035
rect 3235 5005 3285 5035
rect 3315 5005 3365 5035
rect 3395 5005 3445 5035
rect 3475 5005 3525 5035
rect 3555 5005 3605 5035
rect 3635 5005 3685 5035
rect 3715 5005 3765 5035
rect 3795 5005 3845 5035
rect 3875 5005 3925 5035
rect 3955 5005 4005 5035
rect 4035 5005 4085 5035
rect 4115 5005 4165 5035
rect 4195 5005 4245 5035
rect 4275 5005 4325 5035
rect 4355 5005 4405 5035
rect 4435 5005 4485 5035
rect 4515 5005 4565 5035
rect 4595 5005 4645 5035
rect 4675 5005 4725 5035
rect 4755 5005 4805 5035
rect 4835 5005 4840 5035
rect -1520 5000 4840 5005
rect 4880 5035 5720 5040
rect 4880 5005 4885 5035
rect 4915 5005 5045 5035
rect 5075 5005 5205 5035
rect 5235 5005 5365 5035
rect 5395 5005 5525 5035
rect 5555 5005 5685 5035
rect 5715 5005 5720 5035
rect 4880 5000 5720 5005
rect -1520 4955 -1160 4960
rect -1520 4925 -1515 4955
rect -1485 4925 -1355 4955
rect -1325 4925 -1195 4955
rect -1165 4925 -1160 4955
rect -1520 4920 -1160 4925
rect -1120 4955 4840 4960
rect -1120 4925 -1115 4955
rect -1085 4925 10 4955
rect 190 4925 330 4955
rect 510 4925 650 4955
rect 830 4925 970 4955
rect 1150 4925 4840 4955
rect -1120 4920 4840 4925
rect 4880 4955 5720 4960
rect 4880 4925 4885 4955
rect 4915 4925 5045 4955
rect 5075 4925 5205 4955
rect 5235 4925 5365 4955
rect 5395 4925 5525 4955
rect 5555 4925 5685 4955
rect 5715 4925 5720 4955
rect 4880 4920 5720 4925
rect -1520 4875 4840 4880
rect -1520 4845 -1515 4875
rect -1485 4845 -1355 4875
rect -1325 4845 -1195 4875
rect -1165 4845 -1035 4875
rect -1005 4845 -875 4875
rect -845 4845 -795 4875
rect -765 4845 -715 4875
rect -685 4845 -635 4875
rect -605 4845 -555 4875
rect -525 4845 -475 4875
rect -445 4845 -395 4875
rect -365 4845 -315 4875
rect -285 4845 -235 4875
rect -205 4845 -155 4875
rect -125 4845 -75 4875
rect -45 4845 5 4875
rect 35 4845 85 4875
rect 115 4845 165 4875
rect 195 4845 245 4875
rect 275 4845 325 4875
rect 355 4845 405 4875
rect 435 4845 485 4875
rect 515 4845 565 4875
rect 595 4845 645 4875
rect 675 4845 725 4875
rect 755 4845 805 4875
rect 835 4845 885 4875
rect 915 4845 965 4875
rect 995 4845 1045 4875
rect 1075 4845 1125 4875
rect 1155 4845 1205 4875
rect 1235 4845 1285 4875
rect 1315 4845 1365 4875
rect 1395 4845 1445 4875
rect 1475 4845 1525 4875
rect 1555 4845 1605 4875
rect 1635 4845 1685 4875
rect 1715 4845 1765 4875
rect 1795 4845 1845 4875
rect 1875 4845 1925 4875
rect 1955 4845 2005 4875
rect 2035 4845 2085 4875
rect 2115 4845 2165 4875
rect 2195 4845 2245 4875
rect 2275 4845 2325 4875
rect 2355 4845 2405 4875
rect 2435 4845 2485 4875
rect 2515 4845 2565 4875
rect 2595 4845 2645 4875
rect 2675 4845 2725 4875
rect 2755 4845 2805 4875
rect 2835 4845 2885 4875
rect 2915 4845 2965 4875
rect 2995 4845 3045 4875
rect 3075 4845 3125 4875
rect 3155 4845 3205 4875
rect 3235 4845 3285 4875
rect 3315 4845 3365 4875
rect 3395 4845 3445 4875
rect 3475 4845 3525 4875
rect 3555 4845 3605 4875
rect 3635 4845 3685 4875
rect 3715 4845 3765 4875
rect 3795 4845 3845 4875
rect 3875 4845 3925 4875
rect 3955 4845 4005 4875
rect 4035 4845 4085 4875
rect 4115 4845 4165 4875
rect 4195 4845 4245 4875
rect 4275 4845 4325 4875
rect 4355 4845 4405 4875
rect 4435 4845 4485 4875
rect 4515 4845 4565 4875
rect 4595 4845 4645 4875
rect 4675 4845 4725 4875
rect 4755 4845 4805 4875
rect 4835 4845 4840 4875
rect -1520 4840 4840 4845
rect 4880 4875 5720 4880
rect 4880 4845 4885 4875
rect 4915 4845 5045 4875
rect 5075 4845 5205 4875
rect 5235 4845 5365 4875
rect 5395 4845 5525 4875
rect 5555 4845 5685 4875
rect 5715 4845 5720 4875
rect 4880 4840 5720 4845
rect -1440 4795 4840 4800
rect -1440 4765 -1435 4795
rect -1405 4765 85 4795
rect 115 4765 405 4795
rect 435 4765 725 4795
rect 755 4765 1045 4795
rect 1075 4765 1525 4795
rect 1555 4765 1845 4795
rect 1875 4765 2165 4795
rect 2195 4765 2485 4795
rect 2515 4765 2965 4795
rect 2995 4765 3285 4795
rect 3315 4765 3605 4795
rect 3635 4765 3925 4795
rect 3955 4765 4085 4795
rect 4115 4765 4840 4795
rect -1440 4760 4840 4765
rect 4880 4795 5720 4800
rect 4880 4765 4885 4795
rect 4915 4765 5045 4795
rect 5075 4765 5205 4795
rect 5235 4765 5365 4795
rect 5395 4765 5525 4795
rect 5555 4765 5685 4795
rect 5715 4765 5720 4795
rect 4880 4760 5720 4765
rect -1520 4715 4840 4720
rect -1520 4685 -1515 4715
rect -1485 4685 -1355 4715
rect -1325 4685 -1195 4715
rect -1165 4685 -1035 4715
rect -1005 4685 -875 4715
rect -845 4685 -795 4715
rect -765 4685 -715 4715
rect -685 4685 -635 4715
rect -605 4685 -555 4715
rect -525 4685 -475 4715
rect -445 4685 -395 4715
rect -365 4685 -315 4715
rect -285 4685 -235 4715
rect -205 4685 -155 4715
rect -125 4685 -75 4715
rect -45 4685 5 4715
rect 35 4685 85 4715
rect 115 4685 165 4715
rect 195 4685 245 4715
rect 275 4685 325 4715
rect 355 4685 405 4715
rect 435 4685 485 4715
rect 515 4685 565 4715
rect 595 4685 645 4715
rect 675 4685 725 4715
rect 755 4685 805 4715
rect 835 4685 885 4715
rect 915 4685 965 4715
rect 995 4685 1045 4715
rect 1075 4685 1125 4715
rect 1155 4685 1205 4715
rect 1235 4685 1285 4715
rect 1315 4685 1365 4715
rect 1395 4685 1445 4715
rect 1475 4685 1525 4715
rect 1555 4685 1605 4715
rect 1635 4685 1685 4715
rect 1715 4685 1765 4715
rect 1795 4685 1845 4715
rect 1875 4685 1925 4715
rect 1955 4685 2005 4715
rect 2035 4685 2085 4715
rect 2115 4685 2165 4715
rect 2195 4685 2245 4715
rect 2275 4685 2325 4715
rect 2355 4685 2405 4715
rect 2435 4685 2485 4715
rect 2515 4685 2565 4715
rect 2595 4685 2645 4715
rect 2675 4685 2725 4715
rect 2755 4685 2805 4715
rect 2835 4685 2885 4715
rect 2915 4685 2965 4715
rect 2995 4685 3045 4715
rect 3075 4685 3125 4715
rect 3155 4685 3205 4715
rect 3235 4685 3285 4715
rect 3315 4685 3365 4715
rect 3395 4685 3445 4715
rect 3475 4685 3525 4715
rect 3555 4685 3605 4715
rect 3635 4685 3685 4715
rect 3715 4685 3765 4715
rect 3795 4685 3845 4715
rect 3875 4685 3925 4715
rect 3955 4685 4005 4715
rect 4035 4685 4085 4715
rect 4115 4685 4165 4715
rect 4195 4685 4245 4715
rect 4275 4685 4325 4715
rect 4355 4685 4405 4715
rect 4435 4685 4485 4715
rect 4515 4685 4565 4715
rect 4595 4685 4645 4715
rect 4675 4685 4725 4715
rect 4755 4685 4805 4715
rect 4835 4685 4840 4715
rect -1520 4680 4840 4685
rect 4880 4715 5720 4720
rect 4880 4685 4885 4715
rect 4915 4685 5045 4715
rect 5075 4685 5205 4715
rect 5235 4685 5365 4715
rect 5395 4685 5525 4715
rect 5555 4685 5685 4715
rect 5715 4685 5720 4715
rect 4880 4680 5720 4685
rect -1520 4635 4840 4640
rect -1520 4605 -1515 4635
rect -1485 4605 -1355 4635
rect -1325 4605 -1195 4635
rect -1165 4605 -1035 4635
rect -1005 4605 -875 4635
rect -845 4605 -795 4635
rect -765 4605 -715 4635
rect -685 4605 -635 4635
rect -605 4605 -555 4635
rect -525 4605 -475 4635
rect -445 4605 -395 4635
rect -365 4605 -315 4635
rect -285 4605 -235 4635
rect -205 4605 -155 4635
rect -125 4605 -75 4635
rect -45 4605 5 4635
rect 35 4605 85 4635
rect 115 4605 165 4635
rect 195 4605 245 4635
rect 275 4605 325 4635
rect 355 4605 405 4635
rect 435 4605 485 4635
rect 515 4605 565 4635
rect 595 4605 645 4635
rect 675 4605 725 4635
rect 755 4605 805 4635
rect 835 4605 885 4635
rect 915 4605 965 4635
rect 995 4605 1045 4635
rect 1075 4605 1125 4635
rect 1155 4605 1205 4635
rect 1235 4605 1285 4635
rect 1315 4605 1365 4635
rect 1395 4605 1445 4635
rect 1475 4605 1525 4635
rect 1555 4605 1605 4635
rect 1635 4605 1685 4635
rect 1715 4605 1765 4635
rect 1795 4605 1845 4635
rect 1875 4605 1925 4635
rect 1955 4605 2005 4635
rect 2035 4605 2085 4635
rect 2115 4605 2165 4635
rect 2195 4605 2245 4635
rect 2275 4605 2325 4635
rect 2355 4605 2405 4635
rect 2435 4605 2485 4635
rect 2515 4605 2565 4635
rect 2595 4605 2645 4635
rect 2675 4605 2725 4635
rect 2755 4605 2805 4635
rect 2835 4605 2885 4635
rect 2915 4605 2965 4635
rect 2995 4605 3045 4635
rect 3075 4605 3125 4635
rect 3155 4605 3205 4635
rect 3235 4605 3285 4635
rect 3315 4605 3365 4635
rect 3395 4605 3445 4635
rect 3475 4605 3525 4635
rect 3555 4605 3605 4635
rect 3635 4605 3685 4635
rect 3715 4605 3765 4635
rect 3795 4605 3845 4635
rect 3875 4605 3925 4635
rect 3955 4605 4005 4635
rect 4035 4605 4085 4635
rect 4115 4605 4165 4635
rect 4195 4605 4245 4635
rect 4275 4605 4325 4635
rect 4355 4605 4405 4635
rect 4435 4605 4485 4635
rect 4515 4605 4565 4635
rect 4595 4605 4645 4635
rect 4675 4605 4725 4635
rect 4755 4605 4805 4635
rect 4835 4605 4840 4635
rect -1520 4600 4840 4605
rect 4880 4635 5720 4640
rect 4880 4605 4885 4635
rect 4915 4605 5045 4635
rect 5075 4605 5205 4635
rect 5235 4605 5365 4635
rect 5395 4605 5525 4635
rect 5555 4605 5685 4635
rect 5715 4605 5720 4635
rect 4880 4600 5720 4605
rect -1520 4555 -1000 4560
rect -1520 4525 -1515 4555
rect -1485 4525 -1355 4555
rect -1325 4525 -1195 4555
rect -1165 4525 -1035 4555
rect -1005 4525 -1000 4555
rect -1520 4520 -1000 4525
rect -960 4555 4840 4560
rect -960 4525 -955 4555
rect -925 4525 245 4555
rect 275 4525 885 4555
rect 915 4525 1685 4555
rect 1715 4525 2325 4555
rect 2355 4525 4840 4555
rect -960 4520 4840 4525
rect 4880 4555 5720 4560
rect 4880 4525 4885 4555
rect 4915 4525 5045 4555
rect 5075 4525 5205 4555
rect 5235 4525 5365 4555
rect 5395 4525 5525 4555
rect 5555 4525 5685 4555
rect 5715 4525 5720 4555
rect 4880 4520 5720 4525
rect -1520 4475 4840 4480
rect -1520 4445 -1515 4475
rect -1485 4445 -1355 4475
rect -1325 4445 -1195 4475
rect -1165 4445 -1035 4475
rect -1005 4445 -875 4475
rect -845 4445 -795 4475
rect -765 4445 -715 4475
rect -685 4445 -635 4475
rect -605 4445 -555 4475
rect -525 4445 -475 4475
rect -445 4445 -395 4475
rect -365 4445 -315 4475
rect -285 4445 -235 4475
rect -205 4445 -155 4475
rect -125 4445 -75 4475
rect -45 4445 5 4475
rect 35 4445 85 4475
rect 115 4445 165 4475
rect 195 4445 245 4475
rect 275 4445 325 4475
rect 355 4445 405 4475
rect 435 4445 485 4475
rect 515 4445 565 4475
rect 595 4445 645 4475
rect 675 4445 725 4475
rect 755 4445 805 4475
rect 835 4445 885 4475
rect 915 4445 965 4475
rect 995 4445 1045 4475
rect 1075 4445 1125 4475
rect 1155 4445 1205 4475
rect 1235 4445 1285 4475
rect 1315 4445 1365 4475
rect 1395 4445 1445 4475
rect 1475 4445 1525 4475
rect 1555 4445 1605 4475
rect 1635 4445 1685 4475
rect 1715 4445 1765 4475
rect 1795 4445 1845 4475
rect 1875 4445 1925 4475
rect 1955 4445 2005 4475
rect 2035 4445 2085 4475
rect 2115 4445 2165 4475
rect 2195 4445 2245 4475
rect 2275 4445 2325 4475
rect 2355 4445 2405 4475
rect 2435 4445 2485 4475
rect 2515 4445 2565 4475
rect 2595 4445 2645 4475
rect 2675 4445 2725 4475
rect 2755 4445 2805 4475
rect 2835 4445 2885 4475
rect 2915 4445 2965 4475
rect 2995 4445 3045 4475
rect 3075 4445 3125 4475
rect 3155 4445 3205 4475
rect 3235 4445 3285 4475
rect 3315 4445 3365 4475
rect 3395 4445 3445 4475
rect 3475 4445 3525 4475
rect 3555 4445 3605 4475
rect 3635 4445 3685 4475
rect 3715 4445 3765 4475
rect 3795 4445 3845 4475
rect 3875 4445 3925 4475
rect 3955 4445 4005 4475
rect 4035 4445 4085 4475
rect 4115 4445 4165 4475
rect 4195 4445 4245 4475
rect 4275 4445 4325 4475
rect 4355 4445 4405 4475
rect 4435 4445 4485 4475
rect 4515 4445 4565 4475
rect 4595 4445 4645 4475
rect 4675 4445 4725 4475
rect 4755 4445 4805 4475
rect 4835 4445 4840 4475
rect -1520 4440 4840 4445
rect 4880 4475 5720 4480
rect 4880 4445 4885 4475
rect 4915 4445 5045 4475
rect 5075 4445 5205 4475
rect 5235 4445 5365 4475
rect 5395 4445 5525 4475
rect 5555 4445 5685 4475
rect 5715 4445 5720 4475
rect 4880 4440 5720 4445
rect -1520 4395 -840 4400
rect -1520 4365 -1515 4395
rect -1485 4365 -1355 4395
rect -1325 4365 -1195 4395
rect -1165 4365 -1035 4395
rect -1005 4365 -875 4395
rect -845 4365 -840 4395
rect -1520 4360 -840 4365
rect -800 4395 5720 4400
rect -800 4365 -795 4395
rect -765 4365 -715 4395
rect -685 4365 -635 4395
rect -605 4365 -555 4395
rect -525 4365 -475 4395
rect -445 4365 -395 4395
rect -365 4365 -315 4395
rect -285 4365 -235 4395
rect -205 4365 -155 4395
rect -125 4365 -75 4395
rect -45 4365 5 4395
rect 35 4365 85 4395
rect 115 4365 165 4395
rect 195 4365 245 4395
rect 275 4365 325 4395
rect 355 4365 405 4395
rect 435 4365 485 4395
rect 515 4365 565 4395
rect 595 4365 645 4395
rect 675 4365 725 4395
rect 755 4365 805 4395
rect 835 4365 885 4395
rect 915 4365 965 4395
rect 995 4365 1045 4395
rect 1075 4365 1125 4395
rect 1155 4365 1205 4395
rect 1235 4365 1285 4395
rect 1315 4365 1365 4395
rect 1395 4365 1445 4395
rect 1475 4365 1525 4395
rect 1555 4365 1605 4395
rect 1635 4365 1685 4395
rect 1715 4365 1765 4395
rect 1795 4365 1845 4395
rect 1875 4365 1925 4395
rect 1955 4365 2005 4395
rect 2035 4365 2085 4395
rect 2115 4365 2165 4395
rect 2195 4365 2245 4395
rect 2275 4365 2325 4395
rect 2355 4365 2405 4395
rect 2435 4365 2485 4395
rect 2515 4365 2565 4395
rect 2595 4365 2645 4395
rect 2675 4365 2725 4395
rect 2755 4365 2805 4395
rect 2835 4365 2885 4395
rect 2915 4365 2965 4395
rect 2995 4365 3045 4395
rect 3075 4365 3125 4395
rect 3155 4365 3205 4395
rect 3235 4365 3285 4395
rect 3315 4365 3365 4395
rect 3395 4365 3445 4395
rect 3475 4365 3525 4395
rect 3555 4365 3605 4395
rect 3635 4365 3685 4395
rect 3715 4365 3765 4395
rect 3795 4365 3845 4395
rect 3875 4365 3925 4395
rect 3955 4365 4005 4395
rect 4035 4365 4085 4395
rect 4115 4365 4165 4395
rect 4195 4365 4245 4395
rect 4275 4365 4325 4395
rect 4355 4365 4405 4395
rect 4435 4365 4485 4395
rect 4515 4365 4565 4395
rect 4595 4365 4645 4395
rect 4675 4365 4725 4395
rect 4755 4365 4805 4395
rect 4835 4365 4885 4395
rect 4915 4365 5045 4395
rect 5075 4365 5205 4395
rect 5235 4365 5365 4395
rect 5395 4365 5525 4395
rect 5555 4365 5685 4395
rect 5715 4365 5720 4395
rect -800 4360 5720 4365
rect -1520 4315 -840 4320
rect -1520 4285 -1515 4315
rect -1485 4285 -1355 4315
rect -1325 4285 -1195 4315
rect -1165 4285 -1035 4315
rect -1005 4285 -875 4315
rect -845 4285 -840 4315
rect -1520 4280 -840 4285
rect -800 4315 5640 4320
rect -800 4285 565 4315
rect 595 4285 5605 4315
rect 5635 4285 5640 4315
rect -800 4280 5640 4285
rect -1520 4235 -840 4240
rect -1520 4205 -1515 4235
rect -1485 4205 -1355 4235
rect -1325 4205 -1195 4235
rect -1165 4205 -1035 4235
rect -1005 4205 -875 4235
rect -845 4205 -840 4235
rect -1520 4200 -840 4205
rect -800 4235 5720 4240
rect -800 4205 -795 4235
rect -765 4205 -715 4235
rect -685 4205 -635 4235
rect -605 4205 -555 4235
rect -525 4205 -475 4235
rect -445 4205 -395 4235
rect -365 4205 -315 4235
rect -285 4205 -235 4235
rect -205 4205 -155 4235
rect -125 4205 -75 4235
rect -45 4205 5 4235
rect 35 4205 85 4235
rect 115 4205 165 4235
rect 195 4205 245 4235
rect 275 4205 325 4235
rect 355 4205 405 4235
rect 435 4205 485 4235
rect 515 4205 565 4235
rect 595 4205 645 4235
rect 675 4205 725 4235
rect 755 4205 805 4235
rect 835 4205 885 4235
rect 915 4205 965 4235
rect 995 4205 1045 4235
rect 1075 4205 1125 4235
rect 1155 4205 1205 4235
rect 1235 4205 1285 4235
rect 1315 4205 1365 4235
rect 1395 4205 1445 4235
rect 1475 4205 1525 4235
rect 1555 4205 1605 4235
rect 1635 4205 1685 4235
rect 1715 4205 1765 4235
rect 1795 4205 1845 4235
rect 1875 4205 1925 4235
rect 1955 4205 2005 4235
rect 2035 4205 2085 4235
rect 2115 4205 2165 4235
rect 2195 4205 2245 4235
rect 2275 4205 2325 4235
rect 2355 4205 2405 4235
rect 2435 4205 2485 4235
rect 2515 4205 2565 4235
rect 2595 4205 2645 4235
rect 2675 4205 2725 4235
rect 2755 4205 2805 4235
rect 2835 4205 2885 4235
rect 2915 4205 2965 4235
rect 2995 4205 3045 4235
rect 3075 4205 3125 4235
rect 3155 4205 3205 4235
rect 3235 4205 3285 4235
rect 3315 4205 3365 4235
rect 3395 4205 3445 4235
rect 3475 4205 3525 4235
rect 3555 4205 3605 4235
rect 3635 4205 3685 4235
rect 3715 4205 3765 4235
rect 3795 4205 3845 4235
rect 3875 4205 3925 4235
rect 3955 4205 4005 4235
rect 4035 4205 4085 4235
rect 4115 4205 4165 4235
rect 4195 4205 4245 4235
rect 4275 4205 4325 4235
rect 4355 4205 4405 4235
rect 4435 4205 4485 4235
rect 4515 4205 4565 4235
rect 4595 4205 4645 4235
rect 4675 4205 4725 4235
rect 4755 4205 4805 4235
rect 4835 4205 4885 4235
rect 4915 4205 5045 4235
rect 5075 4205 5205 4235
rect 5235 4205 5365 4235
rect 5395 4205 5525 4235
rect 5555 4205 5685 4235
rect 5715 4205 5720 4235
rect -800 4200 5720 4205
rect -1520 4155 -840 4160
rect -1520 4125 -1515 4155
rect -1485 4125 -1355 4155
rect -1325 4125 -1195 4155
rect -1165 4125 -1035 4155
rect -1005 4125 -875 4155
rect -845 4125 -840 4155
rect -1520 4120 -840 4125
rect -800 4155 5000 4160
rect -800 4125 -75 4155
rect -45 4125 565 4155
rect 595 4125 1205 4155
rect 1235 4125 1365 4155
rect 1395 4125 2005 4155
rect 2035 4125 2645 4155
rect 2675 4125 2965 4155
rect 2995 4125 3285 4155
rect 3315 4125 3605 4155
rect 3635 4125 3925 4155
rect 3955 4125 4965 4155
rect 4995 4125 5000 4155
rect -800 4120 5000 4125
rect 5040 4155 5720 4160
rect 5040 4125 5045 4155
rect 5075 4125 5205 4155
rect 5235 4125 5365 4155
rect 5395 4125 5525 4155
rect 5555 4125 5685 4155
rect 5715 4125 5720 4155
rect 5040 4120 5720 4125
rect -1520 4075 -840 4080
rect -1520 4045 -1515 4075
rect -1485 4045 -1355 4075
rect -1325 4045 -1195 4075
rect -1165 4045 -1035 4075
rect -1005 4045 -875 4075
rect -845 4045 -840 4075
rect -1520 4040 -840 4045
rect -800 4075 5720 4080
rect -800 4045 -795 4075
rect -765 4045 -715 4075
rect -685 4045 -635 4075
rect -605 4045 -555 4075
rect -525 4045 -475 4075
rect -445 4045 -395 4075
rect -365 4045 -315 4075
rect -285 4045 -235 4075
rect -205 4045 -155 4075
rect -125 4045 -75 4075
rect -45 4045 5 4075
rect 35 4045 85 4075
rect 115 4045 165 4075
rect 195 4045 245 4075
rect 275 4045 325 4075
rect 355 4045 405 4075
rect 435 4045 485 4075
rect 515 4045 565 4075
rect 595 4045 645 4075
rect 675 4045 725 4075
rect 755 4045 805 4075
rect 835 4045 885 4075
rect 915 4045 965 4075
rect 995 4045 1045 4075
rect 1075 4045 1125 4075
rect 1155 4045 1205 4075
rect 1235 4045 1285 4075
rect 1315 4045 1365 4075
rect 1395 4045 1445 4075
rect 1475 4045 1525 4075
rect 1555 4045 1605 4075
rect 1635 4045 1685 4075
rect 1715 4045 1765 4075
rect 1795 4045 1845 4075
rect 1875 4045 1925 4075
rect 1955 4045 2005 4075
rect 2035 4045 2085 4075
rect 2115 4045 2165 4075
rect 2195 4045 2245 4075
rect 2275 4045 2325 4075
rect 2355 4045 2405 4075
rect 2435 4045 2485 4075
rect 2515 4045 2565 4075
rect 2595 4045 2645 4075
rect 2675 4045 2725 4075
rect 2755 4045 2805 4075
rect 2835 4045 2885 4075
rect 2915 4045 2965 4075
rect 2995 4045 3045 4075
rect 3075 4045 3125 4075
rect 3155 4045 3205 4075
rect 3235 4045 3285 4075
rect 3315 4045 3365 4075
rect 3395 4045 3445 4075
rect 3475 4045 3525 4075
rect 3555 4045 3605 4075
rect 3635 4045 3685 4075
rect 3715 4045 3765 4075
rect 3795 4045 3845 4075
rect 3875 4045 3925 4075
rect 3955 4045 4005 4075
rect 4035 4045 4085 4075
rect 4115 4045 4165 4075
rect 4195 4045 4245 4075
rect 4275 4045 4325 4075
rect 4355 4045 4405 4075
rect 4435 4045 4485 4075
rect 4515 4045 4565 4075
rect 4595 4045 4645 4075
rect 4675 4045 4725 4075
rect 4755 4045 4805 4075
rect 4835 4045 4885 4075
rect 4915 4045 5045 4075
rect 5075 4045 5205 4075
rect 5235 4045 5365 4075
rect 5395 4045 5525 4075
rect 5555 4045 5685 4075
rect 5715 4045 5720 4075
rect -800 4040 5720 4045
rect -1520 3995 -840 4000
rect -1520 3965 -1515 3995
rect -1485 3965 -1355 3995
rect -1325 3965 -1195 3995
rect -1165 3965 -1035 3995
rect -1005 3965 -875 3995
rect -845 3965 -840 3995
rect -1520 3960 -840 3965
rect -800 3995 5720 4000
rect -800 3965 -795 3995
rect -765 3965 -715 3995
rect -685 3965 -635 3995
rect -605 3965 -555 3995
rect -525 3965 -475 3995
rect -445 3965 -395 3995
rect -365 3965 -315 3995
rect -285 3965 -235 3995
rect -205 3965 -155 3995
rect -125 3965 -75 3995
rect -45 3965 5 3995
rect 35 3965 85 3995
rect 115 3965 165 3995
rect 195 3965 245 3995
rect 275 3965 325 3995
rect 355 3965 405 3995
rect 435 3965 485 3995
rect 515 3965 565 3995
rect 595 3965 645 3995
rect 675 3965 725 3995
rect 755 3965 805 3995
rect 835 3965 885 3995
rect 915 3965 965 3995
rect 995 3965 1045 3995
rect 1075 3965 1125 3995
rect 1155 3965 1205 3995
rect 1235 3965 1285 3995
rect 1315 3965 1365 3995
rect 1395 3965 1445 3995
rect 1475 3965 1525 3995
rect 1555 3965 1605 3995
rect 1635 3965 1685 3995
rect 1715 3965 1765 3995
rect 1795 3965 1845 3995
rect 1875 3965 1925 3995
rect 1955 3965 2005 3995
rect 2035 3965 2085 3995
rect 2115 3965 2165 3995
rect 2195 3965 2245 3995
rect 2275 3965 2325 3995
rect 2355 3965 2405 3995
rect 2435 3965 2485 3995
rect 2515 3965 2565 3995
rect 2595 3965 2645 3995
rect 2675 3965 2725 3995
rect 2755 3965 2805 3995
rect 2835 3965 2885 3995
rect 2915 3965 2965 3995
rect 2995 3965 3045 3995
rect 3075 3965 3125 3995
rect 3155 3965 3205 3995
rect 3235 3965 3285 3995
rect 3315 3965 3365 3995
rect 3395 3965 3445 3995
rect 3475 3965 3525 3995
rect 3555 3965 3605 3995
rect 3635 3965 3685 3995
rect 3715 3965 3765 3995
rect 3795 3965 3845 3995
rect 3875 3965 3925 3995
rect 3955 3965 4005 3995
rect 4035 3965 4085 3995
rect 4115 3965 4165 3995
rect 4195 3965 4245 3995
rect 4275 3965 4325 3995
rect 4355 3965 4405 3995
rect 4435 3965 4485 3995
rect 4515 3965 4565 3995
rect 4595 3965 4645 3995
rect 4675 3965 4725 3995
rect 4755 3965 4805 3995
rect 4835 3965 4885 3995
rect 4915 3965 5045 3995
rect 5075 3965 5205 3995
rect 5235 3965 5365 3995
rect 5395 3965 5525 3995
rect 5555 3965 5685 3995
rect 5715 3965 5720 3995
rect -800 3960 5720 3965
rect -1520 3915 -840 3920
rect -1520 3885 -1515 3915
rect -1485 3885 -1355 3915
rect -1325 3885 -1195 3915
rect -1165 3885 -1035 3915
rect -1005 3885 -875 3915
rect -845 3885 -840 3915
rect -1520 3880 -840 3885
rect -800 3915 5720 3920
rect -800 3885 -795 3915
rect -765 3885 -715 3915
rect -685 3885 -635 3915
rect -605 3885 -555 3915
rect -525 3885 -475 3915
rect -445 3885 -395 3915
rect -365 3885 -315 3915
rect -285 3885 -235 3915
rect -205 3885 -155 3915
rect -125 3885 -75 3915
rect -45 3885 5 3915
rect 35 3885 85 3915
rect 115 3885 165 3915
rect 195 3885 245 3915
rect 275 3885 325 3915
rect 355 3885 405 3915
rect 435 3885 485 3915
rect 515 3885 565 3915
rect 595 3885 645 3915
rect 675 3885 725 3915
rect 755 3885 805 3915
rect 835 3885 885 3915
rect 915 3885 965 3915
rect 995 3885 1045 3915
rect 1075 3885 1125 3915
rect 1155 3885 1205 3915
rect 1235 3885 1285 3915
rect 1315 3885 1365 3915
rect 1395 3885 1445 3915
rect 1475 3885 1525 3915
rect 1555 3885 1605 3915
rect 1635 3885 1685 3915
rect 1715 3885 1765 3915
rect 1795 3885 1845 3915
rect 1875 3885 1925 3915
rect 1955 3885 2005 3915
rect 2035 3885 2085 3915
rect 2115 3885 2165 3915
rect 2195 3885 2245 3915
rect 2275 3885 2325 3915
rect 2355 3885 2405 3915
rect 2435 3885 2485 3915
rect 2515 3885 2565 3915
rect 2595 3885 2645 3915
rect 2675 3885 2725 3915
rect 2755 3885 2805 3915
rect 2835 3885 2885 3915
rect 2915 3885 2965 3915
rect 2995 3885 3045 3915
rect 3075 3885 3125 3915
rect 3155 3885 3205 3915
rect 3235 3885 3285 3915
rect 3315 3885 3365 3915
rect 3395 3885 3445 3915
rect 3475 3885 3525 3915
rect 3555 3885 3605 3915
rect 3635 3885 3685 3915
rect 3715 3885 3765 3915
rect 3795 3885 3845 3915
rect 3875 3885 3925 3915
rect 3955 3885 4005 3915
rect 4035 3885 4085 3915
rect 4115 3885 4165 3915
rect 4195 3885 4245 3915
rect 4275 3885 4325 3915
rect 4355 3885 4405 3915
rect 4435 3885 4485 3915
rect 4515 3885 4565 3915
rect 4595 3885 4645 3915
rect 4675 3885 4725 3915
rect 4755 3885 4805 3915
rect 4835 3885 4885 3915
rect 4915 3885 5045 3915
rect 5075 3885 5205 3915
rect 5235 3885 5365 3915
rect 5395 3885 5525 3915
rect 5555 3885 5685 3915
rect 5715 3885 5720 3915
rect -800 3880 5720 3885
rect -1520 3835 -840 3840
rect -1520 3805 -1515 3835
rect -1485 3805 -1355 3835
rect -1325 3805 -1195 3835
rect -1165 3805 -1035 3835
rect -1005 3805 -875 3835
rect -845 3805 -840 3835
rect -1520 3800 -840 3805
rect -800 3835 5720 3840
rect -800 3805 -795 3835
rect -765 3805 -715 3835
rect -685 3805 -635 3835
rect -605 3805 -555 3835
rect -525 3805 -475 3835
rect -445 3805 -395 3835
rect -365 3805 -315 3835
rect -285 3805 -235 3835
rect -205 3805 -155 3835
rect -125 3805 -75 3835
rect -45 3805 5 3835
rect 35 3805 85 3835
rect 115 3805 165 3835
rect 195 3805 245 3835
rect 275 3805 325 3835
rect 355 3805 405 3835
rect 435 3805 485 3835
rect 515 3805 565 3835
rect 595 3805 645 3835
rect 675 3805 725 3835
rect 755 3805 805 3835
rect 835 3805 885 3835
rect 915 3805 965 3835
rect 995 3805 1045 3835
rect 1075 3805 1125 3835
rect 1155 3805 1205 3835
rect 1235 3805 1285 3835
rect 1315 3805 1365 3835
rect 1395 3805 1445 3835
rect 1475 3805 1525 3835
rect 1555 3805 1605 3835
rect 1635 3805 1685 3835
rect 1715 3805 1765 3835
rect 1795 3805 1845 3835
rect 1875 3805 1925 3835
rect 1955 3805 2005 3835
rect 2035 3805 2085 3835
rect 2115 3805 2165 3835
rect 2195 3805 2245 3835
rect 2275 3805 2325 3835
rect 2355 3805 2405 3835
rect 2435 3805 2485 3835
rect 2515 3805 2565 3835
rect 2595 3805 2645 3835
rect 2675 3805 2725 3835
rect 2755 3805 2805 3835
rect 2835 3805 2885 3835
rect 2915 3805 2965 3835
rect 2995 3805 3045 3835
rect 3075 3805 3125 3835
rect 3155 3805 3205 3835
rect 3235 3805 3285 3835
rect 3315 3805 3365 3835
rect 3395 3805 3445 3835
rect 3475 3805 3525 3835
rect 3555 3805 3605 3835
rect 3635 3805 3685 3835
rect 3715 3805 3765 3835
rect 3795 3805 3845 3835
rect 3875 3805 3925 3835
rect 3955 3805 4005 3835
rect 4035 3805 4085 3835
rect 4115 3805 4165 3835
rect 4195 3805 4245 3835
rect 4275 3805 4325 3835
rect 4355 3805 4405 3835
rect 4435 3805 4485 3835
rect 4515 3805 4565 3835
rect 4595 3805 4645 3835
rect 4675 3805 4725 3835
rect 4755 3805 4805 3835
rect 4835 3805 4885 3835
rect 4915 3805 5045 3835
rect 5075 3805 5205 3835
rect 5235 3805 5365 3835
rect 5395 3805 5525 3835
rect 5555 3805 5685 3835
rect 5715 3805 5720 3835
rect -800 3800 5720 3805
rect -1520 3755 -840 3760
rect -1520 3725 -1515 3755
rect -1485 3725 -1355 3755
rect -1325 3725 -1195 3755
rect -1165 3725 -1035 3755
rect -1005 3725 -875 3755
rect -845 3725 -840 3755
rect -1520 3720 -840 3725
rect -800 3755 5720 3760
rect -800 3725 -795 3755
rect -765 3725 -715 3755
rect -685 3725 -635 3755
rect -605 3725 -555 3755
rect -525 3725 -475 3755
rect -445 3725 -395 3755
rect -365 3725 -315 3755
rect -285 3725 -235 3755
rect -205 3725 -155 3755
rect -125 3725 -75 3755
rect -45 3725 5 3755
rect 35 3725 85 3755
rect 115 3725 165 3755
rect 195 3725 245 3755
rect 275 3725 325 3755
rect 355 3725 405 3755
rect 435 3725 485 3755
rect 515 3725 565 3755
rect 595 3725 645 3755
rect 675 3725 725 3755
rect 755 3725 805 3755
rect 835 3725 885 3755
rect 915 3725 965 3755
rect 995 3725 1045 3755
rect 1075 3725 1125 3755
rect 1155 3725 1205 3755
rect 1235 3725 1285 3755
rect 1315 3725 1365 3755
rect 1395 3725 1445 3755
rect 1475 3725 1525 3755
rect 1555 3725 1605 3755
rect 1635 3725 1685 3755
rect 1715 3725 1765 3755
rect 1795 3725 1845 3755
rect 1875 3725 1925 3755
rect 1955 3725 2005 3755
rect 2035 3725 2085 3755
rect 2115 3725 2165 3755
rect 2195 3725 2245 3755
rect 2275 3725 2325 3755
rect 2355 3725 2405 3755
rect 2435 3725 2485 3755
rect 2515 3725 2565 3755
rect 2595 3725 2645 3755
rect 2675 3725 2725 3755
rect 2755 3725 2805 3755
rect 2835 3725 2885 3755
rect 2915 3725 2965 3755
rect 2995 3725 3045 3755
rect 3075 3725 3125 3755
rect 3155 3725 3205 3755
rect 3235 3725 3285 3755
rect 3315 3725 3365 3755
rect 3395 3725 3445 3755
rect 3475 3725 3525 3755
rect 3555 3725 3605 3755
rect 3635 3725 3685 3755
rect 3715 3725 3765 3755
rect 3795 3725 3845 3755
rect 3875 3725 3925 3755
rect 3955 3725 4005 3755
rect 4035 3725 4085 3755
rect 4115 3725 4165 3755
rect 4195 3725 4245 3755
rect 4275 3725 4325 3755
rect 4355 3725 4405 3755
rect 4435 3725 4485 3755
rect 4515 3725 4565 3755
rect 4595 3725 4645 3755
rect 4675 3725 4725 3755
rect 4755 3725 4805 3755
rect 4835 3725 4885 3755
rect 4915 3725 5045 3755
rect 5075 3725 5205 3755
rect 5235 3725 5365 3755
rect 5395 3725 5525 3755
rect 5555 3725 5685 3755
rect 5715 3725 5720 3755
rect -800 3720 5720 3725
rect -1520 3675 -840 3680
rect -1520 3645 -1515 3675
rect -1485 3645 -1355 3675
rect -1325 3645 -1195 3675
rect -1165 3645 -1035 3675
rect -1005 3645 -875 3675
rect -845 3645 -840 3675
rect -1520 3640 -840 3645
rect -800 3675 5720 3680
rect -800 3645 -795 3675
rect -765 3645 -715 3675
rect -685 3645 -635 3675
rect -605 3645 -555 3675
rect -525 3645 -475 3675
rect -445 3645 -395 3675
rect -365 3645 -315 3675
rect -285 3645 -235 3675
rect -205 3645 -155 3675
rect -125 3645 -75 3675
rect -45 3645 5 3675
rect 35 3645 85 3675
rect 115 3645 165 3675
rect 195 3645 245 3675
rect 275 3645 325 3675
rect 355 3645 405 3675
rect 435 3645 485 3675
rect 515 3645 565 3675
rect 595 3645 645 3675
rect 675 3645 725 3675
rect 755 3645 805 3675
rect 835 3645 885 3675
rect 915 3645 965 3675
rect 995 3645 1045 3675
rect 1075 3645 1125 3675
rect 1155 3645 1205 3675
rect 1235 3645 1285 3675
rect 1315 3645 1365 3675
rect 1395 3645 1445 3675
rect 1475 3645 1525 3675
rect 1555 3645 1605 3675
rect 1635 3645 1685 3675
rect 1715 3645 1765 3675
rect 1795 3645 1845 3675
rect 1875 3645 1925 3675
rect 1955 3645 2005 3675
rect 2035 3645 2085 3675
rect 2115 3645 2165 3675
rect 2195 3645 2245 3675
rect 2275 3645 2325 3675
rect 2355 3645 2405 3675
rect 2435 3645 2485 3675
rect 2515 3645 2565 3675
rect 2595 3645 2645 3675
rect 2675 3645 2725 3675
rect 2755 3645 2805 3675
rect 2835 3645 2885 3675
rect 2915 3645 2965 3675
rect 2995 3645 3045 3675
rect 3075 3645 3125 3675
rect 3155 3645 3205 3675
rect 3235 3645 3285 3675
rect 3315 3645 3365 3675
rect 3395 3645 3445 3675
rect 3475 3645 3525 3675
rect 3555 3645 3605 3675
rect 3635 3645 3685 3675
rect 3715 3645 3765 3675
rect 3795 3645 3845 3675
rect 3875 3645 3925 3675
rect 3955 3645 4005 3675
rect 4035 3645 4085 3675
rect 4115 3645 4165 3675
rect 4195 3645 4245 3675
rect 4275 3645 4325 3675
rect 4355 3645 4405 3675
rect 4435 3645 4485 3675
rect 4515 3645 4565 3675
rect 4595 3645 4645 3675
rect 4675 3645 4725 3675
rect 4755 3645 4805 3675
rect 4835 3645 4885 3675
rect 4915 3645 5045 3675
rect 5075 3645 5205 3675
rect 5235 3645 5365 3675
rect 5395 3645 5525 3675
rect 5555 3645 5685 3675
rect 5715 3645 5720 3675
rect -800 3640 5720 3645
rect -1520 3595 4840 3600
rect -1520 3565 -1515 3595
rect -1485 3565 -1355 3595
rect -1325 3565 -1195 3595
rect -1165 3565 -1035 3595
rect -1005 3565 -875 3595
rect -845 3565 -795 3595
rect -765 3565 -715 3595
rect -685 3565 -635 3595
rect -605 3565 -555 3595
rect -525 3565 -475 3595
rect -445 3565 -395 3595
rect -365 3565 -315 3595
rect -285 3565 -235 3595
rect -205 3565 -155 3595
rect -125 3565 -75 3595
rect -45 3565 5 3595
rect 35 3565 85 3595
rect 115 3565 165 3595
rect 195 3565 245 3595
rect 275 3565 325 3595
rect 355 3565 405 3595
rect 435 3565 485 3595
rect 515 3565 565 3595
rect 595 3565 645 3595
rect 675 3565 725 3595
rect 755 3565 805 3595
rect 835 3565 885 3595
rect 915 3565 965 3595
rect 995 3565 1045 3595
rect 1075 3565 1125 3595
rect 1155 3565 1205 3595
rect 1235 3565 1285 3595
rect 1315 3565 1365 3595
rect 1395 3565 1445 3595
rect 1475 3565 1525 3595
rect 1555 3565 1605 3595
rect 1635 3565 1685 3595
rect 1715 3565 1765 3595
rect 1795 3565 1845 3595
rect 1875 3565 1925 3595
rect 1955 3565 2005 3595
rect 2035 3565 2085 3595
rect 2115 3565 2165 3595
rect 2195 3565 2245 3595
rect 2275 3565 2325 3595
rect 2355 3565 2405 3595
rect 2435 3565 2485 3595
rect 2515 3565 2565 3595
rect 2595 3565 2645 3595
rect 2675 3565 2725 3595
rect 2755 3565 2805 3595
rect 2835 3565 2885 3595
rect 2915 3565 2965 3595
rect 2995 3565 3045 3595
rect 3075 3565 3125 3595
rect 3155 3565 3205 3595
rect 3235 3565 3285 3595
rect 3315 3565 3365 3595
rect 3395 3565 3445 3595
rect 3475 3565 3525 3595
rect 3555 3565 3605 3595
rect 3635 3565 3685 3595
rect 3715 3565 3765 3595
rect 3795 3565 3845 3595
rect 3875 3565 3925 3595
rect 3955 3565 4005 3595
rect 4035 3565 4085 3595
rect 4115 3565 4165 3595
rect 4195 3565 4245 3595
rect 4275 3565 4325 3595
rect 4355 3565 4405 3595
rect 4435 3565 4485 3595
rect 4515 3565 4565 3595
rect 4595 3565 4645 3595
rect 4675 3565 4725 3595
rect 4755 3565 4805 3595
rect 4835 3565 4840 3595
rect -1520 3560 4840 3565
rect 4880 3595 5720 3600
rect 4880 3565 4885 3595
rect 4915 3565 5045 3595
rect 5075 3565 5205 3595
rect 5235 3565 5365 3595
rect 5395 3565 5525 3595
rect 5555 3565 5685 3595
rect 5715 3565 5720 3595
rect 4880 3560 5720 3565
rect -1520 3515 4840 3520
rect -1520 3485 -1515 3515
rect -1485 3485 -1355 3515
rect -1325 3485 -1195 3515
rect -1165 3485 -1035 3515
rect -1005 3485 -875 3515
rect -845 3485 -795 3515
rect -765 3485 -715 3515
rect -685 3485 -635 3515
rect -605 3485 -555 3515
rect -525 3485 -475 3515
rect -445 3485 -395 3515
rect -365 3485 -315 3515
rect -285 3485 -235 3515
rect -205 3485 -155 3515
rect -125 3485 -75 3515
rect -45 3485 5 3515
rect 35 3485 85 3515
rect 115 3485 165 3515
rect 195 3485 245 3515
rect 275 3485 325 3515
rect 355 3485 405 3515
rect 435 3485 485 3515
rect 515 3485 565 3515
rect 595 3485 645 3515
rect 675 3485 725 3515
rect 755 3485 805 3515
rect 835 3485 885 3515
rect 915 3485 965 3515
rect 995 3485 1045 3515
rect 1075 3485 1125 3515
rect 1155 3485 1205 3515
rect 1235 3485 1285 3515
rect 1315 3485 1365 3515
rect 1395 3485 1445 3515
rect 1475 3485 1525 3515
rect 1555 3485 1605 3515
rect 1635 3485 1685 3515
rect 1715 3485 1765 3515
rect 1795 3485 1845 3515
rect 1875 3485 1925 3515
rect 1955 3485 2005 3515
rect 2035 3485 2085 3515
rect 2115 3485 2165 3515
rect 2195 3485 2245 3515
rect 2275 3485 2325 3515
rect 2355 3485 2405 3515
rect 2435 3485 2485 3515
rect 2515 3485 2565 3515
rect 2595 3485 2645 3515
rect 2675 3485 2725 3515
rect 2755 3485 2805 3515
rect 2835 3485 2885 3515
rect 2915 3485 2965 3515
rect 2995 3485 3045 3515
rect 3075 3485 3125 3515
rect 3155 3485 3205 3515
rect 3235 3485 3285 3515
rect 3315 3485 3365 3515
rect 3395 3485 3445 3515
rect 3475 3485 3525 3515
rect 3555 3485 3605 3515
rect 3635 3485 3685 3515
rect 3715 3485 3765 3515
rect 3795 3485 3845 3515
rect 3875 3485 3925 3515
rect 3955 3485 4005 3515
rect 4035 3485 4085 3515
rect 4115 3485 4165 3515
rect 4195 3485 4245 3515
rect 4275 3485 4325 3515
rect 4355 3485 4405 3515
rect 4435 3485 4485 3515
rect 4515 3485 4565 3515
rect 4595 3485 4645 3515
rect 4675 3485 4725 3515
rect 4755 3485 4805 3515
rect 4835 3485 4840 3515
rect -1520 3480 4840 3485
rect 4880 3515 5720 3520
rect 4880 3485 4885 3515
rect 4915 3485 5045 3515
rect 5075 3485 5205 3515
rect 5235 3485 5365 3515
rect 5395 3485 5525 3515
rect 5555 3485 5685 3515
rect 5715 3485 5720 3515
rect 4880 3480 5720 3485
rect -1520 3435 -1320 3440
rect -1520 3405 -1515 3435
rect -1485 3405 -1355 3435
rect -1325 3405 -1320 3435
rect -1520 3400 -1320 3405
rect -1280 3435 4840 3440
rect -1280 3405 -1275 3435
rect -1245 3405 10 3435
rect 190 3405 330 3435
rect 510 3405 650 3435
rect 830 3405 970 3435
rect 1150 3405 1450 3435
rect 1630 3405 1770 3435
rect 1950 3405 2090 3435
rect 2270 3405 2410 3435
rect 2590 3405 4840 3435
rect -1280 3400 4840 3405
rect 4880 3435 5720 3440
rect 4880 3405 4885 3435
rect 4915 3405 5045 3435
rect 5075 3405 5205 3435
rect 5235 3405 5365 3435
rect 5395 3405 5525 3435
rect 5555 3405 5685 3435
rect 5715 3405 5720 3435
rect 4880 3400 5720 3405
rect -1520 3355 4840 3360
rect -1520 3325 -1515 3355
rect -1485 3325 -1355 3355
rect -1325 3325 -1195 3355
rect -1165 3325 -1035 3355
rect -1005 3325 -875 3355
rect -845 3325 -795 3355
rect -765 3325 -715 3355
rect -685 3325 -635 3355
rect -605 3325 -555 3355
rect -525 3325 -475 3355
rect -445 3325 -395 3355
rect -365 3325 -315 3355
rect -285 3325 -235 3355
rect -205 3325 -155 3355
rect -125 3325 -75 3355
rect -45 3325 5 3355
rect 35 3325 85 3355
rect 115 3325 165 3355
rect 195 3325 245 3355
rect 275 3325 325 3355
rect 355 3325 405 3355
rect 435 3325 485 3355
rect 515 3325 565 3355
rect 595 3325 645 3355
rect 675 3325 725 3355
rect 755 3325 805 3355
rect 835 3325 885 3355
rect 915 3325 965 3355
rect 995 3325 1045 3355
rect 1075 3325 1125 3355
rect 1155 3325 1205 3355
rect 1235 3325 1285 3355
rect 1315 3325 1365 3355
rect 1395 3325 1445 3355
rect 1475 3325 1525 3355
rect 1555 3325 1605 3355
rect 1635 3325 1685 3355
rect 1715 3325 1765 3355
rect 1795 3325 1845 3355
rect 1875 3325 1925 3355
rect 1955 3325 2005 3355
rect 2035 3325 2085 3355
rect 2115 3325 2165 3355
rect 2195 3325 2245 3355
rect 2275 3325 2325 3355
rect 2355 3325 2405 3355
rect 2435 3325 2485 3355
rect 2515 3325 2565 3355
rect 2595 3325 2645 3355
rect 2675 3325 2725 3355
rect 2755 3325 2805 3355
rect 2835 3325 2885 3355
rect 2915 3325 2965 3355
rect 2995 3325 3045 3355
rect 3075 3325 3125 3355
rect 3155 3325 3205 3355
rect 3235 3325 3285 3355
rect 3315 3325 3365 3355
rect 3395 3325 3445 3355
rect 3475 3325 3525 3355
rect 3555 3325 3605 3355
rect 3635 3325 3685 3355
rect 3715 3325 3765 3355
rect 3795 3325 3845 3355
rect 3875 3325 3925 3355
rect 3955 3325 4005 3355
rect 4035 3325 4085 3355
rect 4115 3325 4165 3355
rect 4195 3325 4245 3355
rect 4275 3325 4325 3355
rect 4355 3325 4405 3355
rect 4435 3325 4485 3355
rect 4515 3325 4565 3355
rect 4595 3325 4645 3355
rect 4675 3325 4725 3355
rect 4755 3325 4805 3355
rect 4835 3325 4840 3355
rect -1520 3320 4840 3325
rect 4880 3355 5720 3360
rect 4880 3325 4885 3355
rect 4915 3325 5045 3355
rect 5075 3325 5205 3355
rect 5235 3325 5365 3355
rect 5395 3325 5525 3355
rect 5555 3325 5685 3355
rect 5715 3325 5720 3355
rect 4880 3320 5720 3325
rect -1520 3275 4840 3280
rect -1520 3245 -1515 3275
rect -1485 3245 -1355 3275
rect -1325 3245 -1195 3275
rect -1165 3245 -1035 3275
rect -1005 3245 -875 3275
rect -845 3245 -795 3275
rect -765 3245 -715 3275
rect -685 3245 -635 3275
rect -605 3245 -555 3275
rect -525 3245 -475 3275
rect -445 3245 -395 3275
rect -365 3245 -315 3275
rect -285 3245 -235 3275
rect -205 3245 -155 3275
rect -125 3245 -75 3275
rect -45 3245 5 3275
rect 35 3245 85 3275
rect 115 3245 165 3275
rect 195 3245 245 3275
rect 275 3245 325 3275
rect 355 3245 405 3275
rect 435 3245 485 3275
rect 515 3245 565 3275
rect 595 3245 645 3275
rect 675 3245 725 3275
rect 755 3245 805 3275
rect 835 3245 885 3275
rect 915 3245 965 3275
rect 995 3245 1045 3275
rect 1075 3245 1125 3275
rect 1155 3245 1205 3275
rect 1235 3245 1285 3275
rect 1315 3245 1365 3275
rect 1395 3245 1445 3275
rect 1475 3245 1525 3275
rect 1555 3245 1605 3275
rect 1635 3245 1685 3275
rect 1715 3245 1765 3275
rect 1795 3245 1845 3275
rect 1875 3245 1925 3275
rect 1955 3245 2005 3275
rect 2035 3245 2085 3275
rect 2115 3245 2165 3275
rect 2195 3245 2245 3275
rect 2275 3245 2325 3275
rect 2355 3245 2405 3275
rect 2435 3245 2485 3275
rect 2515 3245 2565 3275
rect 2595 3245 2645 3275
rect 2675 3245 2725 3275
rect 2755 3245 2805 3275
rect 2835 3245 2885 3275
rect 2915 3245 2965 3275
rect 2995 3245 3045 3275
rect 3075 3245 3125 3275
rect 3155 3245 3205 3275
rect 3235 3245 3285 3275
rect 3315 3245 3365 3275
rect 3395 3245 3445 3275
rect 3475 3245 3525 3275
rect 3555 3245 3605 3275
rect 3635 3245 3685 3275
rect 3715 3245 3765 3275
rect 3795 3245 3845 3275
rect 3875 3245 3925 3275
rect 3955 3245 4005 3275
rect 4035 3245 4085 3275
rect 4115 3245 4165 3275
rect 4195 3245 4245 3275
rect 4275 3245 4325 3275
rect 4355 3245 4405 3275
rect 4435 3245 4485 3275
rect 4515 3245 4565 3275
rect 4595 3245 4645 3275
rect 4675 3245 4725 3275
rect 4755 3245 4805 3275
rect 4835 3245 4840 3275
rect -1520 3240 4840 3245
rect 4880 3275 5720 3280
rect 4880 3245 4885 3275
rect 4915 3245 5045 3275
rect 5075 3245 5205 3275
rect 5235 3245 5365 3275
rect 5395 3245 5525 3275
rect 5555 3245 5685 3275
rect 5715 3245 5720 3275
rect 4880 3240 5720 3245
rect -1520 3195 4840 3200
rect -1520 3165 -1515 3195
rect -1485 3165 -1355 3195
rect -1325 3165 -1195 3195
rect -1165 3165 -1035 3195
rect -1005 3165 -875 3195
rect -845 3165 -795 3195
rect -765 3165 -715 3195
rect -685 3165 -635 3195
rect -605 3165 -555 3195
rect -525 3165 -475 3195
rect -445 3165 -395 3195
rect -365 3165 -315 3195
rect -285 3165 -235 3195
rect -205 3165 -155 3195
rect -125 3165 -75 3195
rect -45 3165 5 3195
rect 35 3165 85 3195
rect 115 3165 165 3195
rect 195 3165 245 3195
rect 275 3165 325 3195
rect 355 3165 405 3195
rect 435 3165 485 3195
rect 515 3165 565 3195
rect 595 3165 645 3195
rect 675 3165 725 3195
rect 755 3165 805 3195
rect 835 3165 885 3195
rect 915 3165 965 3195
rect 995 3165 1045 3195
rect 1075 3165 1125 3195
rect 1155 3165 1205 3195
rect 1235 3165 1285 3195
rect 1315 3165 1365 3195
rect 1395 3165 1445 3195
rect 1475 3165 1525 3195
rect 1555 3165 1605 3195
rect 1635 3165 1685 3195
rect 1715 3165 1765 3195
rect 1795 3165 1845 3195
rect 1875 3165 1925 3195
rect 1955 3165 2005 3195
rect 2035 3165 2085 3195
rect 2115 3165 2165 3195
rect 2195 3165 2245 3195
rect 2275 3165 2325 3195
rect 2355 3165 2405 3195
rect 2435 3165 2485 3195
rect 2515 3165 2565 3195
rect 2595 3165 2645 3195
rect 2675 3165 2725 3195
rect 2755 3165 2805 3195
rect 2835 3165 2885 3195
rect 2915 3165 2965 3195
rect 2995 3165 3045 3195
rect 3075 3165 3125 3195
rect 3155 3165 3205 3195
rect 3235 3165 3285 3195
rect 3315 3165 3365 3195
rect 3395 3165 3445 3195
rect 3475 3165 3525 3195
rect 3555 3165 3605 3195
rect 3635 3165 3685 3195
rect 3715 3165 3765 3195
rect 3795 3165 3845 3195
rect 3875 3165 3925 3195
rect 3955 3165 4005 3195
rect 4035 3165 4085 3195
rect 4115 3165 4165 3195
rect 4195 3165 4245 3195
rect 4275 3165 4325 3195
rect 4355 3165 4405 3195
rect 4435 3165 4485 3195
rect 4515 3165 4565 3195
rect 4595 3165 4645 3195
rect 4675 3165 4725 3195
rect 4755 3165 4805 3195
rect 4835 3165 4840 3195
rect -1520 3160 4840 3165
rect 4880 3195 5720 3200
rect 4880 3165 4885 3195
rect 4915 3165 5045 3195
rect 5075 3165 5205 3195
rect 5235 3165 5365 3195
rect 5395 3165 5525 3195
rect 5555 3165 5685 3195
rect 5715 3165 5720 3195
rect 4880 3160 5720 3165
rect -1520 3115 4840 3120
rect -1520 3085 -1515 3115
rect -1485 3085 -1355 3115
rect -1325 3085 -1195 3115
rect -1165 3085 -1035 3115
rect -1005 3085 -875 3115
rect -845 3085 -795 3115
rect -765 3085 -715 3115
rect -685 3085 -635 3115
rect -605 3085 -555 3115
rect -525 3085 -475 3115
rect -445 3085 -395 3115
rect -365 3085 -315 3115
rect -285 3085 -235 3115
rect -205 3085 -155 3115
rect -125 3085 -75 3115
rect -45 3085 5 3115
rect 35 3085 85 3115
rect 115 3085 165 3115
rect 195 3085 245 3115
rect 275 3085 325 3115
rect 355 3085 405 3115
rect 435 3085 485 3115
rect 515 3085 565 3115
rect 595 3085 645 3115
rect 675 3085 725 3115
rect 755 3085 805 3115
rect 835 3085 885 3115
rect 915 3085 965 3115
rect 995 3085 1045 3115
rect 1075 3085 1125 3115
rect 1155 3085 1205 3115
rect 1235 3085 1285 3115
rect 1315 3085 1365 3115
rect 1395 3085 1445 3115
rect 1475 3085 1525 3115
rect 1555 3085 1605 3115
rect 1635 3085 1685 3115
rect 1715 3085 1765 3115
rect 1795 3085 1845 3115
rect 1875 3085 1925 3115
rect 1955 3085 2005 3115
rect 2035 3085 2085 3115
rect 2115 3085 2165 3115
rect 2195 3085 2245 3115
rect 2275 3085 2325 3115
rect 2355 3085 2405 3115
rect 2435 3085 2485 3115
rect 2515 3085 2565 3115
rect 2595 3085 2645 3115
rect 2675 3085 2725 3115
rect 2755 3085 2805 3115
rect 2835 3085 2885 3115
rect 2915 3085 2965 3115
rect 2995 3085 3045 3115
rect 3075 3085 3125 3115
rect 3155 3085 3205 3115
rect 3235 3085 3285 3115
rect 3315 3085 3365 3115
rect 3395 3085 3445 3115
rect 3475 3085 3525 3115
rect 3555 3085 3605 3115
rect 3635 3085 3685 3115
rect 3715 3085 3765 3115
rect 3795 3085 3845 3115
rect 3875 3085 3925 3115
rect 3955 3085 4005 3115
rect 4035 3085 4085 3115
rect 4115 3085 4165 3115
rect 4195 3085 4245 3115
rect 4275 3085 4325 3115
rect 4355 3085 4405 3115
rect 4435 3085 4485 3115
rect 4515 3085 4565 3115
rect 4595 3085 4645 3115
rect 4675 3085 4725 3115
rect 4755 3085 4805 3115
rect 4835 3085 4840 3115
rect -1520 3080 4840 3085
rect 4880 3115 5720 3120
rect 4880 3085 4885 3115
rect 4915 3085 5045 3115
rect 5075 3085 5205 3115
rect 5235 3085 5365 3115
rect 5395 3085 5525 3115
rect 5555 3085 5685 3115
rect 5715 3085 5720 3115
rect 4880 3080 5720 3085
rect -1520 3035 -1160 3040
rect -1520 3005 -1515 3035
rect -1485 3005 -1355 3035
rect -1325 3005 -1195 3035
rect -1165 3005 -1160 3035
rect -1520 3000 -1160 3005
rect -1120 3035 4840 3040
rect -1120 3005 -1115 3035
rect -1085 3005 10 3035
rect 190 3005 330 3035
rect 510 3005 650 3035
rect 830 3005 970 3035
rect 1150 3005 1450 3035
rect 1630 3005 1770 3035
rect 1950 3005 2090 3035
rect 2270 3005 2410 3035
rect 2590 3005 2890 3035
rect 3070 3005 3210 3035
rect 3390 3005 3445 3035
rect 3475 3005 3530 3035
rect 3710 3005 3850 3035
rect 4030 3005 4085 3035
rect 4115 3005 4840 3035
rect -1120 3000 4840 3005
rect 4880 3035 5720 3040
rect 4880 3005 4885 3035
rect 4915 3005 5045 3035
rect 5075 3005 5205 3035
rect 5235 3005 5365 3035
rect 5395 3005 5525 3035
rect 5555 3005 5685 3035
rect 5715 3005 5720 3035
rect 4880 3000 5720 3005
rect -1520 2955 4840 2960
rect -1520 2925 -1515 2955
rect -1485 2925 -1355 2955
rect -1325 2925 -1195 2955
rect -1165 2925 -1035 2955
rect -1005 2925 -875 2955
rect -845 2925 -795 2955
rect -765 2925 -715 2955
rect -685 2925 -635 2955
rect -605 2925 -555 2955
rect -525 2925 -475 2955
rect -445 2925 -395 2955
rect -365 2925 -315 2955
rect -285 2925 -235 2955
rect -205 2925 -155 2955
rect -125 2925 -75 2955
rect -45 2925 5 2955
rect 35 2925 85 2955
rect 115 2925 165 2955
rect 195 2925 245 2955
rect 275 2925 325 2955
rect 355 2925 405 2955
rect 435 2925 485 2955
rect 515 2925 565 2955
rect 595 2925 645 2955
rect 675 2925 725 2955
rect 755 2925 805 2955
rect 835 2925 885 2955
rect 915 2925 965 2955
rect 995 2925 1045 2955
rect 1075 2925 1125 2955
rect 1155 2925 1205 2955
rect 1235 2925 1285 2955
rect 1315 2925 1365 2955
rect 1395 2925 1445 2955
rect 1475 2925 1525 2955
rect 1555 2925 1605 2955
rect 1635 2925 1685 2955
rect 1715 2925 1765 2955
rect 1795 2925 1845 2955
rect 1875 2925 1925 2955
rect 1955 2925 2005 2955
rect 2035 2925 2085 2955
rect 2115 2925 2165 2955
rect 2195 2925 2245 2955
rect 2275 2925 2325 2955
rect 2355 2925 2405 2955
rect 2435 2925 2485 2955
rect 2515 2925 2565 2955
rect 2595 2925 2645 2955
rect 2675 2925 2725 2955
rect 2755 2925 2805 2955
rect 2835 2925 2885 2955
rect 2915 2925 2965 2955
rect 2995 2925 3045 2955
rect 3075 2925 3125 2955
rect 3155 2925 3205 2955
rect 3235 2925 3285 2955
rect 3315 2925 3365 2955
rect 3395 2925 3445 2955
rect 3475 2925 3525 2955
rect 3555 2925 3605 2955
rect 3635 2925 3685 2955
rect 3715 2925 3765 2955
rect 3795 2925 3845 2955
rect 3875 2925 3925 2955
rect 3955 2925 4005 2955
rect 4035 2925 4085 2955
rect 4115 2925 4165 2955
rect 4195 2925 4245 2955
rect 4275 2925 4325 2955
rect 4355 2925 4405 2955
rect 4435 2925 4485 2955
rect 4515 2925 4565 2955
rect 4595 2925 4645 2955
rect 4675 2925 4725 2955
rect 4755 2925 4805 2955
rect 4835 2925 4840 2955
rect -1520 2920 4840 2925
rect 4880 2955 5720 2960
rect 4880 2925 4885 2955
rect 4915 2925 5045 2955
rect 5075 2925 5205 2955
rect 5235 2925 5365 2955
rect 5395 2925 5525 2955
rect 5555 2925 5685 2955
rect 5715 2925 5720 2955
rect 4880 2920 5720 2925
rect -1520 2875 -1000 2880
rect -1520 2845 -1515 2875
rect -1485 2845 -1355 2875
rect -1325 2845 -1195 2875
rect -1165 2845 -1035 2875
rect -1005 2845 -1000 2875
rect -1520 2840 -1000 2845
rect -960 2875 4840 2880
rect -960 2845 -955 2875
rect -925 2845 2005 2875
rect 2035 2845 2645 2875
rect 2675 2845 4840 2875
rect -960 2840 4840 2845
rect 4880 2875 5720 2880
rect 4880 2845 4885 2875
rect 4915 2845 5045 2875
rect 5075 2845 5205 2875
rect 5235 2845 5365 2875
rect 5395 2845 5525 2875
rect 5555 2845 5685 2875
rect 5715 2845 5720 2875
rect 4880 2840 5720 2845
rect -1520 2795 4840 2800
rect -1520 2765 -1515 2795
rect -1485 2765 -1355 2795
rect -1325 2765 -1195 2795
rect -1165 2765 -1035 2795
rect -1005 2765 -875 2795
rect -845 2765 -795 2795
rect -765 2765 -715 2795
rect -685 2765 -635 2795
rect -605 2765 -555 2795
rect -525 2765 -475 2795
rect -445 2765 -395 2795
rect -365 2765 -315 2795
rect -285 2765 -235 2795
rect -205 2765 -155 2795
rect -125 2765 -75 2795
rect -45 2765 5 2795
rect 35 2765 85 2795
rect 115 2765 165 2795
rect 195 2765 245 2795
rect 275 2765 325 2795
rect 355 2765 405 2795
rect 435 2765 485 2795
rect 515 2765 565 2795
rect 595 2765 645 2795
rect 675 2765 725 2795
rect 755 2765 805 2795
rect 835 2765 885 2795
rect 915 2765 965 2795
rect 995 2765 1045 2795
rect 1075 2765 1125 2795
rect 1155 2765 1205 2795
rect 1235 2765 1285 2795
rect 1315 2765 1365 2795
rect 1395 2765 1445 2795
rect 1475 2765 1525 2795
rect 1555 2765 1605 2795
rect 1635 2765 1685 2795
rect 1715 2765 1765 2795
rect 1795 2765 1845 2795
rect 1875 2765 1925 2795
rect 1955 2765 2005 2795
rect 2035 2765 2085 2795
rect 2115 2765 2165 2795
rect 2195 2765 2245 2795
rect 2275 2765 2325 2795
rect 2355 2765 2405 2795
rect 2435 2765 2485 2795
rect 2515 2765 2565 2795
rect 2595 2765 2645 2795
rect 2675 2765 2725 2795
rect 2755 2765 2805 2795
rect 2835 2765 2885 2795
rect 2915 2765 2965 2795
rect 2995 2765 3045 2795
rect 3075 2765 3125 2795
rect 3155 2765 3205 2795
rect 3235 2765 3285 2795
rect 3315 2765 3365 2795
rect 3395 2765 3445 2795
rect 3475 2765 3525 2795
rect 3555 2765 3605 2795
rect 3635 2765 3685 2795
rect 3715 2765 3765 2795
rect 3795 2765 3845 2795
rect 3875 2765 3925 2795
rect 3955 2765 4005 2795
rect 4035 2765 4085 2795
rect 4115 2765 4165 2795
rect 4195 2765 4245 2795
rect 4275 2765 4325 2795
rect 4355 2765 4405 2795
rect 4435 2765 4485 2795
rect 4515 2765 4565 2795
rect 4595 2765 4645 2795
rect 4675 2765 4725 2795
rect 4755 2765 4805 2795
rect 4835 2765 4840 2795
rect -1520 2760 4840 2765
rect 4880 2795 5720 2800
rect 4880 2765 4885 2795
rect 4915 2765 5045 2795
rect 5075 2765 5205 2795
rect 5235 2765 5365 2795
rect 5395 2765 5525 2795
rect 5555 2765 5685 2795
rect 5715 2765 5720 2795
rect 4880 2760 5720 2765
rect -1520 2715 4840 2720
rect -1520 2685 -1515 2715
rect -1485 2685 -1355 2715
rect -1325 2685 -1195 2715
rect -1165 2685 -1035 2715
rect -1005 2685 -875 2715
rect -845 2685 -795 2715
rect -765 2685 -715 2715
rect -685 2685 -635 2715
rect -605 2685 -555 2715
rect -525 2685 -475 2715
rect -445 2685 -395 2715
rect -365 2685 -315 2715
rect -285 2685 -235 2715
rect -205 2685 -155 2715
rect -125 2685 -75 2715
rect -45 2685 5 2715
rect 35 2685 85 2715
rect 115 2685 165 2715
rect 195 2685 245 2715
rect 275 2685 325 2715
rect 355 2685 405 2715
rect 435 2685 485 2715
rect 515 2685 565 2715
rect 595 2685 645 2715
rect 675 2685 725 2715
rect 755 2685 805 2715
rect 835 2685 885 2715
rect 915 2685 965 2715
rect 995 2685 1045 2715
rect 1075 2685 1125 2715
rect 1155 2685 1205 2715
rect 1235 2685 1285 2715
rect 1315 2685 1365 2715
rect 1395 2685 1445 2715
rect 1475 2685 1525 2715
rect 1555 2685 1605 2715
rect 1635 2685 1685 2715
rect 1715 2685 1765 2715
rect 1795 2685 1845 2715
rect 1875 2685 1925 2715
rect 1955 2685 2005 2715
rect 2035 2685 2085 2715
rect 2115 2685 2165 2715
rect 2195 2685 2245 2715
rect 2275 2685 2325 2715
rect 2355 2685 2405 2715
rect 2435 2685 2485 2715
rect 2515 2685 2565 2715
rect 2595 2685 2645 2715
rect 2675 2685 2725 2715
rect 2755 2685 2805 2715
rect 2835 2685 2885 2715
rect 2915 2685 2965 2715
rect 2995 2685 3045 2715
rect 3075 2685 3125 2715
rect 3155 2685 3205 2715
rect 3235 2685 3285 2715
rect 3315 2685 3365 2715
rect 3395 2685 3445 2715
rect 3475 2685 3525 2715
rect 3555 2685 3605 2715
rect 3635 2685 3685 2715
rect 3715 2685 3765 2715
rect 3795 2685 3845 2715
rect 3875 2685 3925 2715
rect 3955 2685 4005 2715
rect 4035 2685 4085 2715
rect 4115 2685 4165 2715
rect 4195 2685 4245 2715
rect 4275 2685 4325 2715
rect 4355 2685 4405 2715
rect 4435 2685 4485 2715
rect 4515 2685 4565 2715
rect 4595 2685 4645 2715
rect 4675 2685 4725 2715
rect 4755 2685 4805 2715
rect 4835 2685 4840 2715
rect -1520 2680 4840 2685
rect 4880 2715 5720 2720
rect 4880 2685 4885 2715
rect 4915 2685 5045 2715
rect 5075 2685 5205 2715
rect 5235 2685 5365 2715
rect 5395 2685 5525 2715
rect 5555 2685 5685 2715
rect 5715 2685 5720 2715
rect 4880 2680 5720 2685
rect -1520 2635 -1320 2640
rect -1520 2605 -1515 2635
rect -1485 2605 -1355 2635
rect -1325 2605 -1320 2635
rect -1520 2600 -1320 2605
rect -1280 2635 4840 2640
rect -1280 2605 -1275 2635
rect -1245 2605 565 2635
rect 595 2605 1205 2635
rect 1235 2605 4840 2635
rect -1280 2600 4840 2605
rect 4880 2635 5720 2640
rect 4880 2605 4885 2635
rect 4915 2605 5045 2635
rect 5075 2605 5205 2635
rect 5235 2605 5365 2635
rect 5395 2605 5525 2635
rect 5555 2605 5685 2635
rect 5715 2605 5720 2635
rect 4880 2600 5720 2605
rect -1520 2555 4840 2560
rect -1520 2525 -1515 2555
rect -1485 2525 -1355 2555
rect -1325 2525 -1195 2555
rect -1165 2525 -1035 2555
rect -1005 2525 -875 2555
rect -845 2525 -795 2555
rect -765 2525 -715 2555
rect -685 2525 -635 2555
rect -605 2525 -555 2555
rect -525 2525 -475 2555
rect -445 2525 -395 2555
rect -365 2525 -315 2555
rect -285 2525 -235 2555
rect -205 2525 -155 2555
rect -125 2525 -75 2555
rect -45 2525 5 2555
rect 35 2525 85 2555
rect 115 2525 165 2555
rect 195 2525 245 2555
rect 275 2525 325 2555
rect 355 2525 405 2555
rect 435 2525 485 2555
rect 515 2525 565 2555
rect 595 2525 645 2555
rect 675 2525 725 2555
rect 755 2525 805 2555
rect 835 2525 885 2555
rect 915 2525 965 2555
rect 995 2525 1045 2555
rect 1075 2525 1125 2555
rect 1155 2525 1205 2555
rect 1235 2525 1285 2555
rect 1315 2525 1365 2555
rect 1395 2525 1445 2555
rect 1475 2525 1525 2555
rect 1555 2525 1605 2555
rect 1635 2525 1685 2555
rect 1715 2525 1765 2555
rect 1795 2525 1845 2555
rect 1875 2525 1925 2555
rect 1955 2525 2005 2555
rect 2035 2525 2085 2555
rect 2115 2525 2165 2555
rect 2195 2525 2245 2555
rect 2275 2525 2325 2555
rect 2355 2525 2405 2555
rect 2435 2525 2485 2555
rect 2515 2525 2565 2555
rect 2595 2525 2645 2555
rect 2675 2525 2725 2555
rect 2755 2525 2805 2555
rect 2835 2525 2885 2555
rect 2915 2525 2965 2555
rect 2995 2525 3045 2555
rect 3075 2525 3125 2555
rect 3155 2525 3205 2555
rect 3235 2525 3285 2555
rect 3315 2525 3365 2555
rect 3395 2525 3445 2555
rect 3475 2525 3525 2555
rect 3555 2525 3605 2555
rect 3635 2525 3685 2555
rect 3715 2525 3765 2555
rect 3795 2525 3845 2555
rect 3875 2525 3925 2555
rect 3955 2525 4005 2555
rect 4035 2525 4085 2555
rect 4115 2525 4165 2555
rect 4195 2525 4245 2555
rect 4275 2525 4325 2555
rect 4355 2525 4405 2555
rect 4435 2525 4485 2555
rect 4515 2525 4565 2555
rect 4595 2525 4645 2555
rect 4675 2525 4725 2555
rect 4755 2525 4805 2555
rect 4835 2525 4840 2555
rect -1520 2520 4840 2525
rect 4880 2555 5720 2560
rect 4880 2525 4885 2555
rect 4915 2525 5045 2555
rect 5075 2525 5205 2555
rect 5235 2525 5365 2555
rect 5395 2525 5525 2555
rect 5555 2525 5685 2555
rect 5715 2525 5720 2555
rect 4880 2520 5720 2525
rect -1520 2475 -840 2480
rect -1520 2445 -1515 2475
rect -1485 2445 -1355 2475
rect -1325 2445 -1195 2475
rect -1165 2445 -1035 2475
rect -1005 2445 -875 2475
rect -845 2445 -840 2475
rect -1520 2440 -840 2445
rect -800 2475 5720 2480
rect -800 2445 -795 2475
rect -765 2445 -715 2475
rect -685 2445 -635 2475
rect -605 2445 -555 2475
rect -525 2445 -475 2475
rect -445 2445 -395 2475
rect -365 2445 -315 2475
rect -285 2445 -235 2475
rect -205 2445 -155 2475
rect -125 2445 -75 2475
rect -45 2445 5 2475
rect 35 2445 85 2475
rect 115 2445 165 2475
rect 195 2445 245 2475
rect 275 2445 325 2475
rect 355 2445 405 2475
rect 435 2445 485 2475
rect 515 2445 565 2475
rect 595 2445 645 2475
rect 675 2445 725 2475
rect 755 2445 805 2475
rect 835 2445 885 2475
rect 915 2445 965 2475
rect 995 2445 1045 2475
rect 1075 2445 1125 2475
rect 1155 2445 1205 2475
rect 1235 2445 1285 2475
rect 1315 2445 1365 2475
rect 1395 2445 1445 2475
rect 1475 2445 1525 2475
rect 1555 2445 1605 2475
rect 1635 2445 1685 2475
rect 1715 2445 1765 2475
rect 1795 2445 1845 2475
rect 1875 2445 1925 2475
rect 1955 2445 2005 2475
rect 2035 2445 2085 2475
rect 2115 2445 2165 2475
rect 2195 2445 2245 2475
rect 2275 2445 2325 2475
rect 2355 2445 2405 2475
rect 2435 2445 2485 2475
rect 2515 2445 2565 2475
rect 2595 2445 2645 2475
rect 2675 2445 2725 2475
rect 2755 2445 2805 2475
rect 2835 2445 2885 2475
rect 2915 2445 2965 2475
rect 2995 2445 3045 2475
rect 3075 2445 3125 2475
rect 3155 2445 3205 2475
rect 3235 2445 3285 2475
rect 3315 2445 3365 2475
rect 3395 2445 3445 2475
rect 3475 2445 3525 2475
rect 3555 2445 3605 2475
rect 3635 2445 3685 2475
rect 3715 2445 3765 2475
rect 3795 2445 3845 2475
rect 3875 2445 3925 2475
rect 3955 2445 4005 2475
rect 4035 2445 4085 2475
rect 4115 2445 4165 2475
rect 4195 2445 4245 2475
rect 4275 2445 4325 2475
rect 4355 2445 4405 2475
rect 4435 2445 4485 2475
rect 4515 2445 4565 2475
rect 4595 2445 4645 2475
rect 4675 2445 4725 2475
rect 4755 2445 4805 2475
rect 4835 2445 4885 2475
rect 4915 2445 5045 2475
rect 5075 2445 5205 2475
rect 5235 2445 5365 2475
rect 5395 2445 5525 2475
rect 5555 2445 5685 2475
rect 5715 2445 5720 2475
rect -800 2440 5720 2445
rect -1520 2395 -840 2400
rect -1520 2365 -1515 2395
rect -1485 2365 -1355 2395
rect -1325 2365 -1195 2395
rect -1165 2365 -1035 2395
rect -1005 2365 -875 2395
rect -845 2365 -840 2395
rect -1520 2360 -840 2365
rect -800 2395 5320 2400
rect -800 2365 85 2395
rect 115 2365 405 2395
rect 435 2365 725 2395
rect 755 2365 1045 2395
rect 1075 2365 5285 2395
rect 5315 2365 5320 2395
rect -800 2360 5320 2365
rect -1520 2315 -840 2320
rect -1520 2285 -1515 2315
rect -1485 2285 -1355 2315
rect -1325 2285 -1195 2315
rect -1165 2285 -1035 2315
rect -1005 2285 -875 2315
rect -845 2285 -840 2315
rect -1520 2280 -840 2285
rect -800 2315 5720 2320
rect -800 2285 -795 2315
rect -765 2285 -715 2315
rect -685 2285 -635 2315
rect -605 2285 -555 2315
rect -525 2285 -475 2315
rect -445 2285 -395 2315
rect -365 2285 -315 2315
rect -285 2285 -235 2315
rect -205 2285 -155 2315
rect -125 2285 -75 2315
rect -45 2285 5 2315
rect 35 2285 85 2315
rect 115 2285 165 2315
rect 195 2285 245 2315
rect 275 2285 325 2315
rect 355 2285 405 2315
rect 435 2285 485 2315
rect 515 2285 565 2315
rect 595 2285 645 2315
rect 675 2285 725 2315
rect 755 2285 805 2315
rect 835 2285 885 2315
rect 915 2285 965 2315
rect 995 2285 1045 2315
rect 1075 2285 1125 2315
rect 1155 2285 1205 2315
rect 1235 2285 1285 2315
rect 1315 2285 1365 2315
rect 1395 2285 1445 2315
rect 1475 2285 1525 2315
rect 1555 2285 1605 2315
rect 1635 2285 1685 2315
rect 1715 2285 1765 2315
rect 1795 2285 1845 2315
rect 1875 2285 1925 2315
rect 1955 2285 2005 2315
rect 2035 2285 2085 2315
rect 2115 2285 2165 2315
rect 2195 2285 2245 2315
rect 2275 2285 2325 2315
rect 2355 2285 2405 2315
rect 2435 2285 2485 2315
rect 2515 2285 2565 2315
rect 2595 2285 2645 2315
rect 2675 2285 2725 2315
rect 2755 2285 2805 2315
rect 2835 2285 2885 2315
rect 2915 2285 2965 2315
rect 2995 2285 3045 2315
rect 3075 2285 3125 2315
rect 3155 2285 3205 2315
rect 3235 2285 3285 2315
rect 3315 2285 3365 2315
rect 3395 2285 3445 2315
rect 3475 2285 3525 2315
rect 3555 2285 3605 2315
rect 3635 2285 3685 2315
rect 3715 2285 3765 2315
rect 3795 2285 3845 2315
rect 3875 2285 3925 2315
rect 3955 2285 4005 2315
rect 4035 2285 4085 2315
rect 4115 2285 4165 2315
rect 4195 2285 4245 2315
rect 4275 2285 4325 2315
rect 4355 2285 4405 2315
rect 4435 2285 4485 2315
rect 4515 2285 4565 2315
rect 4595 2285 4645 2315
rect 4675 2285 4725 2315
rect 4755 2285 4805 2315
rect 4835 2285 4885 2315
rect 4915 2285 5045 2315
rect 5075 2285 5205 2315
rect 5235 2285 5365 2315
rect 5395 2285 5525 2315
rect 5555 2285 5685 2315
rect 5715 2285 5720 2315
rect -800 2280 5720 2285
rect -1520 2235 -840 2240
rect -1520 2205 -1515 2235
rect -1485 2205 -1355 2235
rect -1325 2205 -1195 2235
rect -1165 2205 -1035 2235
rect -1005 2205 -875 2235
rect -845 2205 -840 2235
rect -1520 2200 -840 2205
rect -800 2235 5000 2240
rect -800 2205 1525 2235
rect 1555 2205 1845 2235
rect 1875 2205 2165 2235
rect 2195 2205 2485 2235
rect 2515 2205 2965 2235
rect 2995 2205 3285 2235
rect 3315 2205 3605 2235
rect 3635 2205 3925 2235
rect 3955 2205 4965 2235
rect 4995 2205 5000 2235
rect -800 2200 5000 2205
rect 5040 2235 5720 2240
rect 5040 2205 5045 2235
rect 5075 2205 5205 2235
rect 5235 2205 5365 2235
rect 5395 2205 5525 2235
rect 5555 2205 5685 2235
rect 5715 2205 5720 2235
rect 5040 2200 5720 2205
rect -1520 2155 -840 2160
rect -1520 2125 -1515 2155
rect -1485 2125 -1355 2155
rect -1325 2125 -1195 2155
rect -1165 2125 -1035 2155
rect -1005 2125 -875 2155
rect -845 2125 -840 2155
rect -1520 2120 -840 2125
rect -800 2155 5720 2160
rect -800 2125 -795 2155
rect -765 2125 -715 2155
rect -685 2125 -635 2155
rect -605 2125 -555 2155
rect -525 2125 -475 2155
rect -445 2125 -395 2155
rect -365 2125 -315 2155
rect -285 2125 -235 2155
rect -205 2125 -155 2155
rect -125 2125 -75 2155
rect -45 2125 5 2155
rect 35 2125 85 2155
rect 115 2125 165 2155
rect 195 2125 245 2155
rect 275 2125 325 2155
rect 355 2125 405 2155
rect 435 2125 485 2155
rect 515 2125 565 2155
rect 595 2125 645 2155
rect 675 2125 725 2155
rect 755 2125 805 2155
rect 835 2125 885 2155
rect 915 2125 965 2155
rect 995 2125 1045 2155
rect 1075 2125 1125 2155
rect 1155 2125 1205 2155
rect 1235 2125 1285 2155
rect 1315 2125 1365 2155
rect 1395 2125 1445 2155
rect 1475 2125 1525 2155
rect 1555 2125 1605 2155
rect 1635 2125 1685 2155
rect 1715 2125 1765 2155
rect 1795 2125 1845 2155
rect 1875 2125 1925 2155
rect 1955 2125 2005 2155
rect 2035 2125 2085 2155
rect 2115 2125 2165 2155
rect 2195 2125 2245 2155
rect 2275 2125 2325 2155
rect 2355 2125 2405 2155
rect 2435 2125 2485 2155
rect 2515 2125 2565 2155
rect 2595 2125 2645 2155
rect 2675 2125 2725 2155
rect 2755 2125 2805 2155
rect 2835 2125 2885 2155
rect 2915 2125 2965 2155
rect 2995 2125 3045 2155
rect 3075 2125 3125 2155
rect 3155 2125 3205 2155
rect 3235 2125 3285 2155
rect 3315 2125 3365 2155
rect 3395 2125 3445 2155
rect 3475 2125 3525 2155
rect 3555 2125 3605 2155
rect 3635 2125 3685 2155
rect 3715 2125 3765 2155
rect 3795 2125 3845 2155
rect 3875 2125 3925 2155
rect 3955 2125 4005 2155
rect 4035 2125 4085 2155
rect 4115 2125 4165 2155
rect 4195 2125 4245 2155
rect 4275 2125 4325 2155
rect 4355 2125 4405 2155
rect 4435 2125 4485 2155
rect 4515 2125 4565 2155
rect 4595 2125 4645 2155
rect 4675 2125 4725 2155
rect 4755 2125 4805 2155
rect 4835 2125 4885 2155
rect 4915 2125 5045 2155
rect 5075 2125 5205 2155
rect 5235 2125 5365 2155
rect 5395 2125 5525 2155
rect 5555 2125 5685 2155
rect 5715 2125 5720 2155
rect -800 2120 5720 2125
rect -1520 2075 -840 2080
rect -1520 2045 -1515 2075
rect -1485 2045 -1355 2075
rect -1325 2045 -1195 2075
rect -1165 2045 -1035 2075
rect -1005 2045 -875 2075
rect -845 2045 -840 2075
rect -1520 2040 -840 2045
rect -800 2075 5720 2080
rect -800 2045 -795 2075
rect -765 2045 -715 2075
rect -685 2045 -635 2075
rect -605 2045 -555 2075
rect -525 2045 -475 2075
rect -445 2045 -395 2075
rect -365 2045 -315 2075
rect -285 2045 -235 2075
rect -205 2045 -155 2075
rect -125 2045 -75 2075
rect -45 2045 5 2075
rect 35 2045 85 2075
rect 115 2045 165 2075
rect 195 2045 245 2075
rect 275 2045 325 2075
rect 355 2045 405 2075
rect 435 2045 485 2075
rect 515 2045 565 2075
rect 595 2045 645 2075
rect 675 2045 725 2075
rect 755 2045 805 2075
rect 835 2045 885 2075
rect 915 2045 965 2075
rect 995 2045 1045 2075
rect 1075 2045 1125 2075
rect 1155 2045 1205 2075
rect 1235 2045 1285 2075
rect 1315 2045 1365 2075
rect 1395 2045 1445 2075
rect 1475 2045 1525 2075
rect 1555 2045 1605 2075
rect 1635 2045 1685 2075
rect 1715 2045 1765 2075
rect 1795 2045 1845 2075
rect 1875 2045 1925 2075
rect 1955 2045 2005 2075
rect 2035 2045 2085 2075
rect 2115 2045 2165 2075
rect 2195 2045 2245 2075
rect 2275 2045 2325 2075
rect 2355 2045 2405 2075
rect 2435 2045 2485 2075
rect 2515 2045 2565 2075
rect 2595 2045 2645 2075
rect 2675 2045 2725 2075
rect 2755 2045 2805 2075
rect 2835 2045 2885 2075
rect 2915 2045 2965 2075
rect 2995 2045 3045 2075
rect 3075 2045 3125 2075
rect 3155 2045 3205 2075
rect 3235 2045 3285 2075
rect 3315 2045 3365 2075
rect 3395 2045 3445 2075
rect 3475 2045 3525 2075
rect 3555 2045 3605 2075
rect 3635 2045 3685 2075
rect 3715 2045 3765 2075
rect 3795 2045 3845 2075
rect 3875 2045 3925 2075
rect 3955 2045 4005 2075
rect 4035 2045 4085 2075
rect 4115 2045 4165 2075
rect 4195 2045 4245 2075
rect 4275 2045 4325 2075
rect 4355 2045 4405 2075
rect 4435 2045 4485 2075
rect 4515 2045 4565 2075
rect 4595 2045 4645 2075
rect 4675 2045 4725 2075
rect 4755 2045 4805 2075
rect 4835 2045 4885 2075
rect 4915 2045 5045 2075
rect 5075 2045 5205 2075
rect 5235 2045 5365 2075
rect 5395 2045 5525 2075
rect 5555 2045 5685 2075
rect 5715 2045 5720 2075
rect -800 2040 5720 2045
rect -1520 1995 -840 2000
rect -1520 1965 -1515 1995
rect -1485 1965 -1355 1995
rect -1325 1965 -1195 1995
rect -1165 1965 -1035 1995
rect -1005 1965 -875 1995
rect -845 1965 -840 1995
rect -1520 1960 -840 1965
rect -800 1995 5720 2000
rect -800 1965 -795 1995
rect -765 1965 -715 1995
rect -685 1965 -635 1995
rect -605 1965 -555 1995
rect -525 1965 -475 1995
rect -445 1965 -395 1995
rect -365 1965 -315 1995
rect -285 1965 -235 1995
rect -205 1965 -155 1995
rect -125 1965 -75 1995
rect -45 1965 5 1995
rect 35 1965 85 1995
rect 115 1965 165 1995
rect 195 1965 245 1995
rect 275 1965 325 1995
rect 355 1965 405 1995
rect 435 1965 485 1995
rect 515 1965 565 1995
rect 595 1965 645 1995
rect 675 1965 725 1995
rect 755 1965 805 1995
rect 835 1965 885 1995
rect 915 1965 965 1995
rect 995 1965 1045 1995
rect 1075 1965 1125 1995
rect 1155 1965 1205 1995
rect 1235 1965 1285 1995
rect 1315 1965 1365 1995
rect 1395 1965 1445 1995
rect 1475 1965 1525 1995
rect 1555 1965 1605 1995
rect 1635 1965 1685 1995
rect 1715 1965 1765 1995
rect 1795 1965 1845 1995
rect 1875 1965 1925 1995
rect 1955 1965 2005 1995
rect 2035 1965 2085 1995
rect 2115 1965 2165 1995
rect 2195 1965 2245 1995
rect 2275 1965 2325 1995
rect 2355 1965 2405 1995
rect 2435 1965 2485 1995
rect 2515 1965 2565 1995
rect 2595 1965 2645 1995
rect 2675 1965 2725 1995
rect 2755 1965 2805 1995
rect 2835 1965 2885 1995
rect 2915 1965 2965 1995
rect 2995 1965 3045 1995
rect 3075 1965 3125 1995
rect 3155 1965 3205 1995
rect 3235 1965 3285 1995
rect 3315 1965 3365 1995
rect 3395 1965 3445 1995
rect 3475 1965 3525 1995
rect 3555 1965 3605 1995
rect 3635 1965 3685 1995
rect 3715 1965 3765 1995
rect 3795 1965 3845 1995
rect 3875 1965 3925 1995
rect 3955 1965 4005 1995
rect 4035 1965 4085 1995
rect 4115 1965 4165 1995
rect 4195 1965 4245 1995
rect 4275 1965 4325 1995
rect 4355 1965 4405 1995
rect 4435 1965 4485 1995
rect 4515 1965 4565 1995
rect 4595 1965 4645 1995
rect 4675 1965 4725 1995
rect 4755 1965 4805 1995
rect 4835 1965 4885 1995
rect 4915 1965 5045 1995
rect 5075 1965 5205 1995
rect 5235 1965 5365 1995
rect 5395 1965 5525 1995
rect 5555 1965 5685 1995
rect 5715 1965 5720 1995
rect -800 1960 5720 1965
rect -1520 1915 -840 1920
rect -1520 1885 -1515 1915
rect -1485 1885 -1355 1915
rect -1325 1885 -1195 1915
rect -1165 1885 -1035 1915
rect -1005 1885 -875 1915
rect -845 1885 -840 1915
rect -1520 1880 -840 1885
rect -800 1915 5720 1920
rect -800 1885 -795 1915
rect -765 1885 -715 1915
rect -685 1885 -635 1915
rect -605 1885 -555 1915
rect -525 1885 -475 1915
rect -445 1885 -395 1915
rect -365 1885 -315 1915
rect -285 1885 -235 1915
rect -205 1885 -155 1915
rect -125 1885 -75 1915
rect -45 1885 5 1915
rect 35 1885 85 1915
rect 115 1885 165 1915
rect 195 1885 245 1915
rect 275 1885 325 1915
rect 355 1885 405 1915
rect 435 1885 485 1915
rect 515 1885 565 1915
rect 595 1885 645 1915
rect 675 1885 725 1915
rect 755 1885 805 1915
rect 835 1885 885 1915
rect 915 1885 965 1915
rect 995 1885 1045 1915
rect 1075 1885 1125 1915
rect 1155 1885 1205 1915
rect 1235 1885 1285 1915
rect 1315 1885 1365 1915
rect 1395 1885 1445 1915
rect 1475 1885 1525 1915
rect 1555 1885 1605 1915
rect 1635 1885 1685 1915
rect 1715 1885 1765 1915
rect 1795 1885 1845 1915
rect 1875 1885 1925 1915
rect 1955 1885 2005 1915
rect 2035 1885 2085 1915
rect 2115 1885 2165 1915
rect 2195 1885 2245 1915
rect 2275 1885 2325 1915
rect 2355 1885 2405 1915
rect 2435 1885 2485 1915
rect 2515 1885 2565 1915
rect 2595 1885 2645 1915
rect 2675 1885 2725 1915
rect 2755 1885 2805 1915
rect 2835 1885 2885 1915
rect 2915 1885 2965 1915
rect 2995 1885 3045 1915
rect 3075 1885 3125 1915
rect 3155 1885 3205 1915
rect 3235 1885 3285 1915
rect 3315 1885 3365 1915
rect 3395 1885 3445 1915
rect 3475 1885 3525 1915
rect 3555 1885 3605 1915
rect 3635 1885 3685 1915
rect 3715 1885 3765 1915
rect 3795 1885 3845 1915
rect 3875 1885 3925 1915
rect 3955 1885 4005 1915
rect 4035 1885 4085 1915
rect 4115 1885 4165 1915
rect 4195 1885 4245 1915
rect 4275 1885 4325 1915
rect 4355 1885 4405 1915
rect 4435 1885 4485 1915
rect 4515 1885 4565 1915
rect 4595 1885 4645 1915
rect 4675 1885 4725 1915
rect 4755 1885 4805 1915
rect 4835 1885 4885 1915
rect 4915 1885 5045 1915
rect 5075 1885 5205 1915
rect 5235 1885 5365 1915
rect 5395 1885 5525 1915
rect 5555 1885 5685 1915
rect 5715 1885 5720 1915
rect -800 1880 5720 1885
rect -1520 1835 -840 1840
rect -1520 1805 -1515 1835
rect -1485 1805 -1355 1835
rect -1325 1805 -1195 1835
rect -1165 1805 -1035 1835
rect -1005 1805 -875 1835
rect -845 1805 -840 1835
rect -1520 1800 -840 1805
rect -800 1835 5720 1840
rect -800 1805 -795 1835
rect -765 1805 -715 1835
rect -685 1805 -635 1835
rect -605 1805 -555 1835
rect -525 1805 -475 1835
rect -445 1805 -395 1835
rect -365 1805 -315 1835
rect -285 1805 -235 1835
rect -205 1805 -155 1835
rect -125 1805 -75 1835
rect -45 1805 5 1835
rect 35 1805 85 1835
rect 115 1805 165 1835
rect 195 1805 245 1835
rect 275 1805 325 1835
rect 355 1805 405 1835
rect 435 1805 485 1835
rect 515 1805 565 1835
rect 595 1805 645 1835
rect 675 1805 725 1835
rect 755 1805 805 1835
rect 835 1805 885 1835
rect 915 1805 965 1835
rect 995 1805 1045 1835
rect 1075 1805 1125 1835
rect 1155 1805 1205 1835
rect 1235 1805 1285 1835
rect 1315 1805 1365 1835
rect 1395 1805 1445 1835
rect 1475 1805 1525 1835
rect 1555 1805 1605 1835
rect 1635 1805 1685 1835
rect 1715 1805 1765 1835
rect 1795 1805 1845 1835
rect 1875 1805 1925 1835
rect 1955 1805 2005 1835
rect 2035 1805 2085 1835
rect 2115 1805 2165 1835
rect 2195 1805 2245 1835
rect 2275 1805 2325 1835
rect 2355 1805 2405 1835
rect 2435 1805 2485 1835
rect 2515 1805 2565 1835
rect 2595 1805 2645 1835
rect 2675 1805 2725 1835
rect 2755 1805 2805 1835
rect 2835 1805 2885 1835
rect 2915 1805 2965 1835
rect 2995 1805 3045 1835
rect 3075 1805 3125 1835
rect 3155 1805 3205 1835
rect 3235 1805 3285 1835
rect 3315 1805 3365 1835
rect 3395 1805 3445 1835
rect 3475 1805 3525 1835
rect 3555 1805 3605 1835
rect 3635 1805 3685 1835
rect 3715 1805 3765 1835
rect 3795 1805 3845 1835
rect 3875 1805 3925 1835
rect 3955 1805 4005 1835
rect 4035 1805 4085 1835
rect 4115 1805 4165 1835
rect 4195 1805 4245 1835
rect 4275 1805 4325 1835
rect 4355 1805 4405 1835
rect 4435 1805 4485 1835
rect 4515 1805 4565 1835
rect 4595 1805 4645 1835
rect 4675 1805 4725 1835
rect 4755 1805 4805 1835
rect 4835 1805 4885 1835
rect 4915 1805 5045 1835
rect 5075 1805 5205 1835
rect 5235 1805 5365 1835
rect 5395 1805 5525 1835
rect 5555 1805 5685 1835
rect 5715 1805 5720 1835
rect -800 1800 5720 1805
rect -1520 1755 -840 1760
rect -1520 1725 -1515 1755
rect -1485 1725 -1355 1755
rect -1325 1725 -1195 1755
rect -1165 1725 -1035 1755
rect -1005 1725 -875 1755
rect -845 1725 -840 1755
rect -1520 1720 -840 1725
rect -800 1755 5720 1760
rect -800 1725 -795 1755
rect -765 1725 -715 1755
rect -685 1725 -635 1755
rect -605 1725 -555 1755
rect -525 1725 -475 1755
rect -445 1725 -395 1755
rect -365 1725 -315 1755
rect -285 1725 -235 1755
rect -205 1725 -155 1755
rect -125 1725 -75 1755
rect -45 1725 5 1755
rect 35 1725 85 1755
rect 115 1725 165 1755
rect 195 1725 245 1755
rect 275 1725 325 1755
rect 355 1725 405 1755
rect 435 1725 485 1755
rect 515 1725 565 1755
rect 595 1725 645 1755
rect 675 1725 725 1755
rect 755 1725 805 1755
rect 835 1725 885 1755
rect 915 1725 965 1755
rect 995 1725 1045 1755
rect 1075 1725 1125 1755
rect 1155 1725 1205 1755
rect 1235 1725 1285 1755
rect 1315 1725 1365 1755
rect 1395 1725 1445 1755
rect 1475 1725 1525 1755
rect 1555 1725 1605 1755
rect 1635 1725 1685 1755
rect 1715 1725 1765 1755
rect 1795 1725 1845 1755
rect 1875 1725 1925 1755
rect 1955 1725 2005 1755
rect 2035 1725 2085 1755
rect 2115 1725 2165 1755
rect 2195 1725 2245 1755
rect 2275 1725 2325 1755
rect 2355 1725 2405 1755
rect 2435 1725 2485 1755
rect 2515 1725 2565 1755
rect 2595 1725 2645 1755
rect 2675 1725 2725 1755
rect 2755 1725 2805 1755
rect 2835 1725 2885 1755
rect 2915 1725 2965 1755
rect 2995 1725 3045 1755
rect 3075 1725 3125 1755
rect 3155 1725 3205 1755
rect 3235 1725 3285 1755
rect 3315 1725 3365 1755
rect 3395 1725 3445 1755
rect 3475 1725 3525 1755
rect 3555 1725 3605 1755
rect 3635 1725 3685 1755
rect 3715 1725 3765 1755
rect 3795 1725 3845 1755
rect 3875 1725 3925 1755
rect 3955 1725 4005 1755
rect 4035 1725 4085 1755
rect 4115 1725 4165 1755
rect 4195 1725 4245 1755
rect 4275 1725 4325 1755
rect 4355 1725 4405 1755
rect 4435 1725 4485 1755
rect 4515 1725 4565 1755
rect 4595 1725 4645 1755
rect 4675 1725 4725 1755
rect 4755 1725 4805 1755
rect 4835 1725 4885 1755
rect 4915 1725 5045 1755
rect 5075 1725 5205 1755
rect 5235 1725 5365 1755
rect 5395 1725 5525 1755
rect 5555 1725 5685 1755
rect 5715 1725 5720 1755
rect -800 1720 5720 1725
rect -1520 1675 4840 1680
rect -1520 1645 -1515 1675
rect -1485 1645 -1355 1675
rect -1325 1645 -1195 1675
rect -1165 1645 -1035 1675
rect -1005 1645 -875 1675
rect -845 1645 -795 1675
rect -765 1645 -715 1675
rect -685 1645 -635 1675
rect -605 1645 -555 1675
rect -525 1645 -475 1675
rect -445 1645 -395 1675
rect -365 1645 -315 1675
rect -285 1645 -235 1675
rect -205 1645 -155 1675
rect -125 1645 -75 1675
rect -45 1645 5 1675
rect 35 1645 85 1675
rect 115 1645 165 1675
rect 195 1645 245 1675
rect 275 1645 325 1675
rect 355 1645 405 1675
rect 435 1645 485 1675
rect 515 1645 565 1675
rect 595 1645 645 1675
rect 675 1645 725 1675
rect 755 1645 805 1675
rect 835 1645 885 1675
rect 915 1645 965 1675
rect 995 1645 1045 1675
rect 1075 1645 1125 1675
rect 1155 1645 1205 1675
rect 1235 1645 1285 1675
rect 1315 1645 1365 1675
rect 1395 1645 1445 1675
rect 1475 1645 1525 1675
rect 1555 1645 1605 1675
rect 1635 1645 1685 1675
rect 1715 1645 1765 1675
rect 1795 1645 1845 1675
rect 1875 1645 1925 1675
rect 1955 1645 2005 1675
rect 2035 1645 2085 1675
rect 2115 1645 2165 1675
rect 2195 1645 2245 1675
rect 2275 1645 2325 1675
rect 2355 1645 2405 1675
rect 2435 1645 2485 1675
rect 2515 1645 2565 1675
rect 2595 1645 2645 1675
rect 2675 1645 2725 1675
rect 2755 1645 2805 1675
rect 2835 1645 2885 1675
rect 2915 1645 2965 1675
rect 2995 1645 3045 1675
rect 3075 1645 3125 1675
rect 3155 1645 3205 1675
rect 3235 1645 3285 1675
rect 3315 1645 3365 1675
rect 3395 1645 3445 1675
rect 3475 1645 3525 1675
rect 3555 1645 3605 1675
rect 3635 1645 3685 1675
rect 3715 1645 3765 1675
rect 3795 1645 3845 1675
rect 3875 1645 3925 1675
rect 3955 1645 4005 1675
rect 4035 1645 4085 1675
rect 4115 1645 4165 1675
rect 4195 1645 4245 1675
rect 4275 1645 4325 1675
rect 4355 1645 4405 1675
rect 4435 1645 4485 1675
rect 4515 1645 4565 1675
rect 4595 1645 4645 1675
rect 4675 1645 4725 1675
rect 4755 1645 4805 1675
rect 4835 1645 4840 1675
rect -1520 1640 4840 1645
rect 4880 1675 5720 1680
rect 4880 1645 4885 1675
rect 4915 1645 5045 1675
rect 5075 1645 5205 1675
rect 5235 1645 5365 1675
rect 5395 1645 5525 1675
rect 5555 1645 5685 1675
rect 5715 1645 5720 1675
rect 4880 1640 5720 1645
rect -1520 1595 4840 1600
rect -1520 1565 -1515 1595
rect -1485 1565 -1355 1595
rect -1325 1565 -1195 1595
rect -1165 1565 -1035 1595
rect -1005 1565 -875 1595
rect -845 1565 -795 1595
rect -765 1565 -715 1595
rect -685 1565 -635 1595
rect -605 1565 -555 1595
rect -525 1565 -475 1595
rect -445 1565 -395 1595
rect -365 1565 -315 1595
rect -285 1565 -235 1595
rect -205 1565 -155 1595
rect -125 1565 -75 1595
rect -45 1565 5 1595
rect 35 1565 85 1595
rect 115 1565 165 1595
rect 195 1565 245 1595
rect 275 1565 325 1595
rect 355 1565 405 1595
rect 435 1565 485 1595
rect 515 1565 565 1595
rect 595 1565 645 1595
rect 675 1565 725 1595
rect 755 1565 805 1595
rect 835 1565 885 1595
rect 915 1565 965 1595
rect 995 1565 1045 1595
rect 1075 1565 1125 1595
rect 1155 1565 1205 1595
rect 1235 1565 1285 1595
rect 1315 1565 1365 1595
rect 1395 1565 1445 1595
rect 1475 1565 1525 1595
rect 1555 1565 1605 1595
rect 1635 1565 1685 1595
rect 1715 1565 1765 1595
rect 1795 1565 1845 1595
rect 1875 1565 1925 1595
rect 1955 1565 2005 1595
rect 2035 1565 2085 1595
rect 2115 1565 2165 1595
rect 2195 1565 2245 1595
rect 2275 1565 2325 1595
rect 2355 1565 2405 1595
rect 2435 1565 2485 1595
rect 2515 1565 2565 1595
rect 2595 1565 2645 1595
rect 2675 1565 2725 1595
rect 2755 1565 2805 1595
rect 2835 1565 2885 1595
rect 2915 1565 2965 1595
rect 2995 1565 3045 1595
rect 3075 1565 3125 1595
rect 3155 1565 3205 1595
rect 3235 1565 3285 1595
rect 3315 1565 3365 1595
rect 3395 1565 3445 1595
rect 3475 1565 3525 1595
rect 3555 1565 3605 1595
rect 3635 1565 3685 1595
rect 3715 1565 3765 1595
rect 3795 1565 3845 1595
rect 3875 1565 3925 1595
rect 3955 1565 4005 1595
rect 4035 1565 4085 1595
rect 4115 1565 4165 1595
rect 4195 1565 4245 1595
rect 4275 1565 4325 1595
rect 4355 1565 4405 1595
rect 4435 1565 4485 1595
rect 4515 1565 4565 1595
rect 4595 1565 4645 1595
rect 4675 1565 4725 1595
rect 4755 1565 4805 1595
rect 4835 1565 4840 1595
rect -1520 1560 4840 1565
rect 4880 1595 5720 1600
rect 4880 1565 4885 1595
rect 4915 1565 5045 1595
rect 5075 1565 5205 1595
rect 5235 1565 5365 1595
rect 5395 1565 5525 1595
rect 5555 1565 5685 1595
rect 5715 1565 5720 1595
rect 4880 1560 5720 1565
rect -1520 1515 -1000 1520
rect -1520 1485 -1515 1515
rect -1485 1485 -1355 1515
rect -1325 1485 -1195 1515
rect -1165 1485 -1035 1515
rect -1005 1485 -1000 1515
rect -1520 1480 -1000 1485
rect -960 1515 4840 1520
rect -960 1485 -955 1515
rect -925 1485 10 1515
rect 190 1485 330 1515
rect 510 1485 650 1515
rect 830 1485 970 1515
rect 1150 1485 1450 1515
rect 1630 1485 1770 1515
rect 1950 1485 2090 1515
rect 2270 1485 2410 1515
rect 2590 1485 2890 1515
rect 3070 1485 3210 1515
rect 3390 1485 3530 1515
rect 3710 1485 3850 1515
rect 4030 1485 4840 1515
rect -960 1480 4840 1485
rect 4880 1515 5720 1520
rect 4880 1485 4885 1515
rect 4915 1485 5045 1515
rect 5075 1485 5205 1515
rect 5235 1485 5365 1515
rect 5395 1485 5525 1515
rect 5555 1485 5685 1515
rect 5715 1485 5720 1515
rect 4880 1480 5720 1485
rect -1520 1435 4840 1440
rect -1520 1405 -1515 1435
rect -1485 1405 -1355 1435
rect -1325 1405 -1195 1435
rect -1165 1405 -1035 1435
rect -1005 1405 -875 1435
rect -845 1405 -795 1435
rect -765 1405 -715 1435
rect -685 1405 -635 1435
rect -605 1405 -555 1435
rect -525 1405 -475 1435
rect -445 1405 -395 1435
rect -365 1405 -315 1435
rect -285 1405 -235 1435
rect -205 1405 -155 1435
rect -125 1405 -75 1435
rect -45 1405 5 1435
rect 35 1405 85 1435
rect 115 1405 165 1435
rect 195 1405 245 1435
rect 275 1405 325 1435
rect 355 1405 405 1435
rect 435 1405 485 1435
rect 515 1405 565 1435
rect 595 1405 645 1435
rect 675 1405 725 1435
rect 755 1405 805 1435
rect 835 1405 885 1435
rect 915 1405 965 1435
rect 995 1405 1045 1435
rect 1075 1405 1125 1435
rect 1155 1405 1205 1435
rect 1235 1405 1285 1435
rect 1315 1405 1365 1435
rect 1395 1405 1445 1435
rect 1475 1405 1525 1435
rect 1555 1405 1605 1435
rect 1635 1405 1685 1435
rect 1715 1405 1765 1435
rect 1795 1405 1845 1435
rect 1875 1405 1925 1435
rect 1955 1405 2005 1435
rect 2035 1405 2085 1435
rect 2115 1405 2165 1435
rect 2195 1405 2245 1435
rect 2275 1405 2325 1435
rect 2355 1405 2405 1435
rect 2435 1405 2485 1435
rect 2515 1405 2565 1435
rect 2595 1405 2645 1435
rect 2675 1405 2725 1435
rect 2755 1405 2805 1435
rect 2835 1405 2885 1435
rect 2915 1405 2965 1435
rect 2995 1405 3045 1435
rect 3075 1405 3125 1435
rect 3155 1405 3205 1435
rect 3235 1405 3285 1435
rect 3315 1405 3365 1435
rect 3395 1405 3445 1435
rect 3475 1405 3525 1435
rect 3555 1405 3605 1435
rect 3635 1405 3685 1435
rect 3715 1405 3765 1435
rect 3795 1405 3845 1435
rect 3875 1405 3925 1435
rect 3955 1405 4005 1435
rect 4035 1405 4085 1435
rect 4115 1405 4165 1435
rect 4195 1405 4245 1435
rect 4275 1405 4325 1435
rect 4355 1405 4405 1435
rect 4435 1405 4485 1435
rect 4515 1405 4565 1435
rect 4595 1405 4645 1435
rect 4675 1405 4725 1435
rect 4755 1405 4805 1435
rect 4835 1405 4840 1435
rect -1520 1400 4840 1405
rect 4880 1435 5720 1440
rect 4880 1405 4885 1435
rect 4915 1405 5045 1435
rect 5075 1405 5205 1435
rect 5235 1405 5365 1435
rect 5395 1405 5525 1435
rect 5555 1405 5685 1435
rect 5715 1405 5720 1435
rect 4880 1400 5720 1405
rect -1520 1355 4840 1360
rect -1520 1325 -1515 1355
rect -1485 1325 -1355 1355
rect -1325 1325 -1195 1355
rect -1165 1325 -1035 1355
rect -1005 1325 -875 1355
rect -845 1325 -795 1355
rect -765 1325 -715 1355
rect -685 1325 -635 1355
rect -605 1325 -555 1355
rect -525 1325 -475 1355
rect -445 1325 -395 1355
rect -365 1325 -315 1355
rect -285 1325 -235 1355
rect -205 1325 -155 1355
rect -125 1325 -75 1355
rect -45 1325 5 1355
rect 35 1325 85 1355
rect 115 1325 165 1355
rect 195 1325 245 1355
rect 275 1325 325 1355
rect 355 1325 405 1355
rect 435 1325 485 1355
rect 515 1325 565 1355
rect 595 1325 645 1355
rect 675 1325 725 1355
rect 755 1325 805 1355
rect 835 1325 885 1355
rect 915 1325 965 1355
rect 995 1325 1045 1355
rect 1075 1325 1125 1355
rect 1155 1325 1205 1355
rect 1235 1325 1285 1355
rect 1315 1325 1365 1355
rect 1395 1325 1445 1355
rect 1475 1325 1525 1355
rect 1555 1325 1605 1355
rect 1635 1325 1685 1355
rect 1715 1325 1765 1355
rect 1795 1325 1845 1355
rect 1875 1325 1925 1355
rect 1955 1325 2005 1355
rect 2035 1325 2085 1355
rect 2115 1325 2165 1355
rect 2195 1325 2245 1355
rect 2275 1325 2325 1355
rect 2355 1325 2405 1355
rect 2435 1325 2485 1355
rect 2515 1325 2565 1355
rect 2595 1325 2645 1355
rect 2675 1325 2725 1355
rect 2755 1325 2805 1355
rect 2835 1325 2885 1355
rect 2915 1325 2965 1355
rect 2995 1325 3045 1355
rect 3075 1325 3125 1355
rect 3155 1325 3205 1355
rect 3235 1325 3285 1355
rect 3315 1325 3365 1355
rect 3395 1325 3445 1355
rect 3475 1325 3525 1355
rect 3555 1325 3605 1355
rect 3635 1325 3685 1355
rect 3715 1325 3765 1355
rect 3795 1325 3845 1355
rect 3875 1325 3925 1355
rect 3955 1325 4005 1355
rect 4035 1325 4085 1355
rect 4115 1325 4165 1355
rect 4195 1325 4245 1355
rect 4275 1325 4325 1355
rect 4355 1325 4405 1355
rect 4435 1325 4485 1355
rect 4515 1325 4565 1355
rect 4595 1325 4645 1355
rect 4675 1325 4725 1355
rect 4755 1325 4805 1355
rect 4835 1325 4840 1355
rect -1520 1320 4840 1325
rect 4880 1355 5720 1360
rect 4880 1325 4885 1355
rect 4915 1325 5045 1355
rect 5075 1325 5205 1355
rect 5235 1325 5365 1355
rect 5395 1325 5525 1355
rect 5555 1325 5685 1355
rect 5715 1325 5720 1355
rect 4880 1320 5720 1325
rect -1520 1275 4840 1280
rect -1520 1245 -1515 1275
rect -1485 1245 -1355 1275
rect -1325 1245 -1195 1275
rect -1165 1245 -1035 1275
rect -1005 1245 -875 1275
rect -845 1245 -795 1275
rect -765 1245 -715 1275
rect -685 1245 -635 1275
rect -605 1245 -555 1275
rect -525 1245 -475 1275
rect -445 1245 -395 1275
rect -365 1245 -315 1275
rect -285 1245 -235 1275
rect -205 1245 -155 1275
rect -125 1245 -75 1275
rect -45 1245 5 1275
rect 35 1245 85 1275
rect 115 1245 165 1275
rect 195 1245 245 1275
rect 275 1245 325 1275
rect 355 1245 405 1275
rect 435 1245 485 1275
rect 515 1245 565 1275
rect 595 1245 645 1275
rect 675 1245 725 1275
rect 755 1245 805 1275
rect 835 1245 885 1275
rect 915 1245 965 1275
rect 995 1245 1045 1275
rect 1075 1245 1125 1275
rect 1155 1245 1205 1275
rect 1235 1245 1285 1275
rect 1315 1245 1365 1275
rect 1395 1245 1445 1275
rect 1475 1245 1525 1275
rect 1555 1245 1605 1275
rect 1635 1245 1685 1275
rect 1715 1245 1765 1275
rect 1795 1245 1845 1275
rect 1875 1245 1925 1275
rect 1955 1245 2005 1275
rect 2035 1245 2085 1275
rect 2115 1245 2165 1275
rect 2195 1245 2245 1275
rect 2275 1245 2325 1275
rect 2355 1245 2405 1275
rect 2435 1245 2485 1275
rect 2515 1245 2565 1275
rect 2595 1245 2645 1275
rect 2675 1245 2725 1275
rect 2755 1245 2805 1275
rect 2835 1245 2885 1275
rect 2915 1245 2965 1275
rect 2995 1245 3045 1275
rect 3075 1245 3125 1275
rect 3155 1245 3205 1275
rect 3235 1245 3285 1275
rect 3315 1245 3365 1275
rect 3395 1245 3445 1275
rect 3475 1245 3525 1275
rect 3555 1245 3605 1275
rect 3635 1245 3685 1275
rect 3715 1245 3765 1275
rect 3795 1245 3845 1275
rect 3875 1245 3925 1275
rect 3955 1245 4005 1275
rect 4035 1245 4085 1275
rect 4115 1245 4165 1275
rect 4195 1245 4245 1275
rect 4275 1245 4325 1275
rect 4355 1245 4405 1275
rect 4435 1245 4485 1275
rect 4515 1245 4565 1275
rect 4595 1245 4645 1275
rect 4675 1245 4725 1275
rect 4755 1245 4805 1275
rect 4835 1245 4840 1275
rect -1520 1240 4840 1245
rect 4880 1275 5720 1280
rect 4880 1245 4885 1275
rect 4915 1245 5045 1275
rect 5075 1245 5205 1275
rect 5235 1245 5365 1275
rect 5395 1245 5525 1275
rect 5555 1245 5685 1275
rect 5715 1245 5720 1275
rect 4880 1240 5720 1245
rect -1520 1195 4840 1200
rect -1520 1165 -1515 1195
rect -1485 1165 -1355 1195
rect -1325 1165 -1195 1195
rect -1165 1165 -1035 1195
rect -1005 1165 -875 1195
rect -845 1165 -795 1195
rect -765 1165 -715 1195
rect -685 1165 -635 1195
rect -605 1165 -555 1195
rect -525 1165 -475 1195
rect -445 1165 -395 1195
rect -365 1165 -315 1195
rect -285 1165 -235 1195
rect -205 1165 -155 1195
rect -125 1165 -75 1195
rect -45 1165 5 1195
rect 35 1165 85 1195
rect 115 1165 165 1195
rect 195 1165 245 1195
rect 275 1165 325 1195
rect 355 1165 405 1195
rect 435 1165 485 1195
rect 515 1165 565 1195
rect 595 1165 645 1195
rect 675 1165 725 1195
rect 755 1165 805 1195
rect 835 1165 885 1195
rect 915 1165 965 1195
rect 995 1165 1045 1195
rect 1075 1165 1125 1195
rect 1155 1165 1205 1195
rect 1235 1165 1285 1195
rect 1315 1165 1365 1195
rect 1395 1165 1445 1195
rect 1475 1165 1525 1195
rect 1555 1165 1605 1195
rect 1635 1165 1685 1195
rect 1715 1165 1765 1195
rect 1795 1165 1845 1195
rect 1875 1165 1925 1195
rect 1955 1165 2005 1195
rect 2035 1165 2085 1195
rect 2115 1165 2165 1195
rect 2195 1165 2245 1195
rect 2275 1165 2325 1195
rect 2355 1165 2405 1195
rect 2435 1165 2485 1195
rect 2515 1165 2565 1195
rect 2595 1165 2645 1195
rect 2675 1165 2725 1195
rect 2755 1165 2805 1195
rect 2835 1165 2885 1195
rect 2915 1165 2965 1195
rect 2995 1165 3045 1195
rect 3075 1165 3125 1195
rect 3155 1165 3205 1195
rect 3235 1165 3285 1195
rect 3315 1165 3365 1195
rect 3395 1165 3445 1195
rect 3475 1165 3525 1195
rect 3555 1165 3605 1195
rect 3635 1165 3685 1195
rect 3715 1165 3765 1195
rect 3795 1165 3845 1195
rect 3875 1165 3925 1195
rect 3955 1165 4005 1195
rect 4035 1165 4085 1195
rect 4115 1165 4165 1195
rect 4195 1165 4245 1195
rect 4275 1165 4325 1195
rect 4355 1165 4405 1195
rect 4435 1165 4485 1195
rect 4515 1165 4565 1195
rect 4595 1165 4645 1195
rect 4675 1165 4725 1195
rect 4755 1165 4805 1195
rect 4835 1165 4840 1195
rect -1520 1160 4840 1165
rect 4880 1195 5720 1200
rect 4880 1165 4885 1195
rect 4915 1165 5045 1195
rect 5075 1165 5205 1195
rect 5235 1165 5365 1195
rect 5395 1165 5525 1195
rect 5555 1165 5685 1195
rect 5715 1165 5720 1195
rect 4880 1160 5720 1165
rect -1520 1115 -1160 1120
rect -1520 1085 -1515 1115
rect -1485 1085 -1355 1115
rect -1325 1085 -1195 1115
rect -1165 1085 -1160 1115
rect -1520 1080 -1160 1085
rect -1120 1115 4840 1120
rect -1120 1085 -1115 1115
rect -1085 1085 10 1115
rect 190 1085 330 1115
rect 510 1085 650 1115
rect 830 1085 970 1115
rect 1150 1085 1450 1115
rect 1630 1085 1770 1115
rect 1950 1085 2090 1115
rect 2270 1085 2410 1115
rect 2590 1085 2890 1115
rect 3070 1085 3210 1115
rect 3390 1085 3530 1115
rect 3710 1085 3850 1115
rect 4030 1085 4840 1115
rect -1120 1080 4840 1085
rect 4880 1115 5720 1120
rect 4880 1085 4885 1115
rect 4915 1085 5045 1115
rect 5075 1085 5205 1115
rect 5235 1085 5365 1115
rect 5395 1085 5525 1115
rect 5555 1085 5685 1115
rect 5715 1085 5720 1115
rect 4880 1080 5720 1085
rect -1520 1035 4840 1040
rect -1520 1005 -1515 1035
rect -1485 1005 -1355 1035
rect -1325 1005 -1195 1035
rect -1165 1005 -1035 1035
rect -1005 1005 -875 1035
rect -845 1005 -795 1035
rect -765 1005 -715 1035
rect -685 1005 -635 1035
rect -605 1005 -555 1035
rect -525 1005 -475 1035
rect -445 1005 -395 1035
rect -365 1005 -315 1035
rect -285 1005 -235 1035
rect -205 1005 -155 1035
rect -125 1005 -75 1035
rect -45 1005 5 1035
rect 35 1005 85 1035
rect 115 1005 165 1035
rect 195 1005 245 1035
rect 275 1005 325 1035
rect 355 1005 405 1035
rect 435 1005 485 1035
rect 515 1005 565 1035
rect 595 1005 645 1035
rect 675 1005 725 1035
rect 755 1005 805 1035
rect 835 1005 885 1035
rect 915 1005 965 1035
rect 995 1005 1045 1035
rect 1075 1005 1125 1035
rect 1155 1005 1205 1035
rect 1235 1005 1285 1035
rect 1315 1005 1365 1035
rect 1395 1005 1445 1035
rect 1475 1005 1525 1035
rect 1555 1005 1605 1035
rect 1635 1005 1685 1035
rect 1715 1005 1765 1035
rect 1795 1005 1845 1035
rect 1875 1005 1925 1035
rect 1955 1005 2005 1035
rect 2035 1005 2085 1035
rect 2115 1005 2165 1035
rect 2195 1005 2245 1035
rect 2275 1005 2325 1035
rect 2355 1005 2405 1035
rect 2435 1005 2485 1035
rect 2515 1005 2565 1035
rect 2595 1005 2645 1035
rect 2675 1005 2725 1035
rect 2755 1005 2805 1035
rect 2835 1005 2885 1035
rect 2915 1005 2965 1035
rect 2995 1005 3045 1035
rect 3075 1005 3125 1035
rect 3155 1005 3205 1035
rect 3235 1005 3285 1035
rect 3315 1005 3365 1035
rect 3395 1005 3445 1035
rect 3475 1005 3525 1035
rect 3555 1005 3605 1035
rect 3635 1005 3685 1035
rect 3715 1005 3765 1035
rect 3795 1005 3845 1035
rect 3875 1005 3925 1035
rect 3955 1005 4005 1035
rect 4035 1005 4085 1035
rect 4115 1005 4165 1035
rect 4195 1005 4245 1035
rect 4275 1005 4325 1035
rect 4355 1005 4405 1035
rect 4435 1005 4485 1035
rect 4515 1005 4565 1035
rect 4595 1005 4645 1035
rect 4675 1005 4725 1035
rect 4755 1005 4805 1035
rect 4835 1005 4840 1035
rect -1520 1000 4840 1005
rect 4880 1035 5720 1040
rect 4880 1005 4885 1035
rect 4915 1005 5045 1035
rect 5075 1005 5205 1035
rect 5235 1005 5365 1035
rect 5395 1005 5525 1035
rect 5555 1005 5685 1035
rect 5715 1005 5720 1035
rect 4880 1000 5720 1005
rect -1520 955 4840 960
rect -1520 925 -1515 955
rect -1485 925 -1355 955
rect -1325 925 -1195 955
rect -1165 925 -1035 955
rect -1005 925 -875 955
rect -845 925 -795 955
rect -765 925 -715 955
rect -685 925 -635 955
rect -605 925 -555 955
rect -525 925 -475 955
rect -445 925 -395 955
rect -365 925 -315 955
rect -285 925 -235 955
rect -205 925 -155 955
rect -125 925 -75 955
rect -45 925 5 955
rect 35 925 85 955
rect 115 925 165 955
rect 195 925 245 955
rect 275 925 325 955
rect 355 925 405 955
rect 435 925 485 955
rect 515 925 565 955
rect 595 925 645 955
rect 675 925 725 955
rect 755 925 805 955
rect 835 925 885 955
rect 915 925 965 955
rect 995 925 1045 955
rect 1075 925 1125 955
rect 1155 925 1205 955
rect 1235 925 1285 955
rect 1315 925 1365 955
rect 1395 925 1445 955
rect 1475 925 1525 955
rect 1555 925 1605 955
rect 1635 925 1685 955
rect 1715 925 1765 955
rect 1795 925 1845 955
rect 1875 925 1925 955
rect 1955 925 2005 955
rect 2035 925 2085 955
rect 2115 925 2165 955
rect 2195 925 2245 955
rect 2275 925 2325 955
rect 2355 925 2405 955
rect 2435 925 2485 955
rect 2515 925 2565 955
rect 2595 925 2645 955
rect 2675 925 2725 955
rect 2755 925 2805 955
rect 2835 925 2885 955
rect 2915 925 2965 955
rect 2995 925 3045 955
rect 3075 925 3125 955
rect 3155 925 3205 955
rect 3235 925 3285 955
rect 3315 925 3365 955
rect 3395 925 3445 955
rect 3475 925 3525 955
rect 3555 925 3605 955
rect 3635 925 3685 955
rect 3715 925 3765 955
rect 3795 925 3845 955
rect 3875 925 3925 955
rect 3955 925 4005 955
rect 4035 925 4085 955
rect 4115 925 4165 955
rect 4195 925 4245 955
rect 4275 925 4325 955
rect 4355 925 4405 955
rect 4435 925 4485 955
rect 4515 925 4565 955
rect 4595 925 4645 955
rect 4675 925 4725 955
rect 4755 925 4805 955
rect 4835 925 4840 955
rect -1520 920 4840 925
rect 4880 955 5720 960
rect 4880 925 4885 955
rect 4915 925 5045 955
rect 5075 925 5205 955
rect 5235 925 5365 955
rect 5395 925 5525 955
rect 5555 925 5685 955
rect 5715 925 5720 955
rect 4880 920 5720 925
rect -1520 875 -840 880
rect -1520 845 -1515 875
rect -1485 845 -1355 875
rect -1325 845 -1195 875
rect -1165 845 -1035 875
rect -1005 845 -875 875
rect -845 845 -840 875
rect -1520 840 -840 845
rect -800 875 5720 880
rect -800 845 -795 875
rect -765 845 -715 875
rect -685 845 -635 875
rect -605 845 -555 875
rect -525 845 -475 875
rect -445 845 -395 875
rect -365 845 -315 875
rect -285 845 -235 875
rect -205 845 -155 875
rect -125 845 -75 875
rect -45 845 5 875
rect 35 845 85 875
rect 115 845 165 875
rect 195 845 245 875
rect 275 845 325 875
rect 355 845 405 875
rect 435 845 485 875
rect 515 845 565 875
rect 595 845 645 875
rect 675 845 725 875
rect 755 845 805 875
rect 835 845 885 875
rect 915 845 965 875
rect 995 845 1045 875
rect 1075 845 1125 875
rect 1155 845 1205 875
rect 1235 845 1285 875
rect 1315 845 1365 875
rect 1395 845 1445 875
rect 1475 845 1525 875
rect 1555 845 1605 875
rect 1635 845 1685 875
rect 1715 845 1765 875
rect 1795 845 1845 875
rect 1875 845 1925 875
rect 1955 845 2005 875
rect 2035 845 2085 875
rect 2115 845 2165 875
rect 2195 845 2245 875
rect 2275 845 2325 875
rect 2355 845 2405 875
rect 2435 845 2485 875
rect 2515 845 2565 875
rect 2595 845 2645 875
rect 2675 845 2725 875
rect 2755 845 2805 875
rect 2835 845 2885 875
rect 2915 845 2965 875
rect 2995 845 3045 875
rect 3075 845 3125 875
rect 3155 845 3205 875
rect 3235 845 3285 875
rect 3315 845 3365 875
rect 3395 845 3445 875
rect 3475 845 3525 875
rect 3555 845 3605 875
rect 3635 845 3685 875
rect 3715 845 3765 875
rect 3795 845 3845 875
rect 3875 845 3925 875
rect 3955 845 4005 875
rect 4035 845 4085 875
rect 4115 845 4165 875
rect 4195 845 4245 875
rect 4275 845 4325 875
rect 4355 845 4405 875
rect 4435 845 4485 875
rect 4515 845 4565 875
rect 4595 845 4645 875
rect 4675 845 4725 875
rect 4755 845 4805 875
rect 4835 845 4885 875
rect 4915 845 5045 875
rect 5075 845 5205 875
rect 5235 845 5365 875
rect 5395 845 5525 875
rect 5555 845 5685 875
rect 5715 845 5720 875
rect -800 840 5720 845
rect -1520 795 -840 800
rect -1520 765 -1515 795
rect -1485 765 -1355 795
rect -1325 765 -1195 795
rect -1165 765 -1035 795
rect -1005 765 -875 795
rect -845 765 -840 795
rect -1520 760 -840 765
rect -800 795 5480 800
rect -800 765 85 795
rect 115 765 245 795
rect 275 765 405 795
rect 435 765 725 795
rect 755 765 885 795
rect 915 765 1045 795
rect 1075 765 1205 795
rect 1235 765 1525 795
rect 1555 765 1845 795
rect 1875 765 5445 795
rect 5475 765 5480 795
rect -800 760 5480 765
rect 5520 795 5720 800
rect 5520 765 5525 795
rect 5555 765 5685 795
rect 5715 765 5720 795
rect 5520 760 5720 765
rect -1520 715 -840 720
rect -1520 685 -1515 715
rect -1485 685 -1355 715
rect -1325 685 -1195 715
rect -1165 685 -1035 715
rect -1005 685 -875 715
rect -845 685 -840 715
rect -1520 680 -840 685
rect -800 715 5720 720
rect -800 685 -795 715
rect -765 685 -715 715
rect -685 685 -635 715
rect -605 685 -555 715
rect -525 685 -475 715
rect -445 685 -395 715
rect -365 685 -315 715
rect -285 685 -235 715
rect -205 685 -155 715
rect -125 685 -75 715
rect -45 685 5 715
rect 35 685 85 715
rect 115 685 165 715
rect 195 685 245 715
rect 275 685 325 715
rect 355 685 405 715
rect 435 685 485 715
rect 515 685 565 715
rect 595 685 645 715
rect 675 685 725 715
rect 755 685 805 715
rect 835 685 885 715
rect 915 685 965 715
rect 995 685 1045 715
rect 1075 685 1125 715
rect 1155 685 1205 715
rect 1235 685 1285 715
rect 1315 685 1365 715
rect 1395 685 1445 715
rect 1475 685 1525 715
rect 1555 685 1605 715
rect 1635 685 1685 715
rect 1715 685 1765 715
rect 1795 685 1845 715
rect 1875 685 1925 715
rect 1955 685 2005 715
rect 2035 685 2085 715
rect 2115 685 2165 715
rect 2195 685 2245 715
rect 2275 685 2325 715
rect 2355 685 2405 715
rect 2435 685 2485 715
rect 2515 685 2565 715
rect 2595 685 2645 715
rect 2675 685 2725 715
rect 2755 685 2805 715
rect 2835 685 2885 715
rect 2915 685 2965 715
rect 2995 685 3045 715
rect 3075 685 3125 715
rect 3155 685 3205 715
rect 3235 685 3285 715
rect 3315 685 3365 715
rect 3395 685 3445 715
rect 3475 685 3525 715
rect 3555 685 3605 715
rect 3635 685 3685 715
rect 3715 685 3765 715
rect 3795 685 3845 715
rect 3875 685 3925 715
rect 3955 685 4005 715
rect 4035 685 4085 715
rect 4115 685 4165 715
rect 4195 685 4245 715
rect 4275 685 4325 715
rect 4355 685 4405 715
rect 4435 685 4485 715
rect 4515 685 4565 715
rect 4595 685 4645 715
rect 4675 685 4725 715
rect 4755 685 4805 715
rect 4835 685 4885 715
rect 4915 685 5045 715
rect 5075 685 5205 715
rect 5235 685 5365 715
rect 5395 685 5525 715
rect 5555 685 5685 715
rect 5715 685 5720 715
rect -800 680 5720 685
rect -1520 635 -840 640
rect -1520 605 -1515 635
rect -1485 605 -1355 635
rect -1325 605 -1195 635
rect -1165 605 -1035 635
rect -1005 605 -875 635
rect -845 605 -840 635
rect -1520 600 -840 605
rect -800 635 5320 640
rect -800 605 2005 635
rect 2035 605 2165 635
rect 2195 605 2485 635
rect 2515 605 2645 635
rect 2675 605 5285 635
rect 5315 605 5320 635
rect -800 600 5320 605
rect 5360 635 5720 640
rect 5360 605 5365 635
rect 5395 605 5525 635
rect 5555 605 5685 635
rect 5715 605 5720 635
rect 5360 600 5720 605
rect -1520 555 -840 560
rect -1520 525 -1515 555
rect -1485 525 -1355 555
rect -1325 525 -1195 555
rect -1165 525 -1035 555
rect -1005 525 -875 555
rect -845 525 -840 555
rect -1520 520 -840 525
rect -800 555 5720 560
rect -800 525 -795 555
rect -765 525 -715 555
rect -685 525 -635 555
rect -605 525 -555 555
rect -525 525 -475 555
rect -445 525 -395 555
rect -365 525 -315 555
rect -285 525 -235 555
rect -205 525 -155 555
rect -125 525 -75 555
rect -45 525 5 555
rect 35 525 85 555
rect 115 525 165 555
rect 195 525 245 555
rect 275 525 325 555
rect 355 525 405 555
rect 435 525 485 555
rect 515 525 565 555
rect 595 525 645 555
rect 675 525 725 555
rect 755 525 805 555
rect 835 525 885 555
rect 915 525 965 555
rect 995 525 1045 555
rect 1075 525 1125 555
rect 1155 525 1205 555
rect 1235 525 1285 555
rect 1315 525 1365 555
rect 1395 525 1445 555
rect 1475 525 1525 555
rect 1555 525 1605 555
rect 1635 525 1685 555
rect 1715 525 1765 555
rect 1795 525 1845 555
rect 1875 525 1925 555
rect 1955 525 2005 555
rect 2035 525 2085 555
rect 2115 525 2165 555
rect 2195 525 2245 555
rect 2275 525 2325 555
rect 2355 525 2405 555
rect 2435 525 2485 555
rect 2515 525 2565 555
rect 2595 525 2645 555
rect 2675 525 2725 555
rect 2755 525 2805 555
rect 2835 525 2885 555
rect 2915 525 2965 555
rect 2995 525 3045 555
rect 3075 525 3125 555
rect 3155 525 3205 555
rect 3235 525 3285 555
rect 3315 525 3365 555
rect 3395 525 3445 555
rect 3475 525 3525 555
rect 3555 525 3605 555
rect 3635 525 3685 555
rect 3715 525 3765 555
rect 3795 525 3845 555
rect 3875 525 3925 555
rect 3955 525 4005 555
rect 4035 525 4085 555
rect 4115 525 4165 555
rect 4195 525 4245 555
rect 4275 525 4325 555
rect 4355 525 4405 555
rect 4435 525 4485 555
rect 4515 525 4565 555
rect 4595 525 4645 555
rect 4675 525 4725 555
rect 4755 525 4805 555
rect 4835 525 4885 555
rect 4915 525 5045 555
rect 5075 525 5205 555
rect 5235 525 5365 555
rect 5395 525 5525 555
rect 5555 525 5685 555
rect 5715 525 5720 555
rect -800 520 5720 525
rect -1520 475 -840 480
rect -1520 445 -1515 475
rect -1485 445 -1355 475
rect -1325 445 -1195 475
rect -1165 445 -1035 475
rect -1005 445 -875 475
rect -845 445 -840 475
rect -1520 440 -840 445
rect -800 475 5160 480
rect -800 445 565 475
rect 595 445 2005 475
rect 2035 445 5125 475
rect 5155 445 5160 475
rect -800 440 5160 445
rect 5200 475 5720 480
rect 5200 445 5205 475
rect 5235 445 5365 475
rect 5395 445 5525 475
rect 5555 445 5685 475
rect 5715 445 5720 475
rect 5200 440 5720 445
rect -1520 395 -840 400
rect -1520 365 -1515 395
rect -1485 365 -1355 395
rect -1325 365 -1195 395
rect -1165 365 -1035 395
rect -1005 365 -875 395
rect -845 365 -840 395
rect -1520 360 -840 365
rect -800 395 5720 400
rect -800 365 -795 395
rect -765 365 -715 395
rect -685 365 -635 395
rect -605 365 -555 395
rect -525 365 -475 395
rect -445 365 -395 395
rect -365 365 -315 395
rect -285 365 -235 395
rect -205 365 -155 395
rect -125 365 -75 395
rect -45 365 5 395
rect 35 365 85 395
rect 115 365 165 395
rect 195 365 245 395
rect 275 365 325 395
rect 355 365 405 395
rect 435 365 485 395
rect 515 365 565 395
rect 595 365 645 395
rect 675 365 725 395
rect 755 365 805 395
rect 835 365 885 395
rect 915 365 965 395
rect 995 365 1045 395
rect 1075 365 1125 395
rect 1155 365 1205 395
rect 1235 365 1285 395
rect 1315 365 1365 395
rect 1395 365 1445 395
rect 1475 365 1525 395
rect 1555 365 1605 395
rect 1635 365 1685 395
rect 1715 365 1765 395
rect 1795 365 1845 395
rect 1875 365 1925 395
rect 1955 365 2005 395
rect 2035 365 2085 395
rect 2115 365 2165 395
rect 2195 365 2245 395
rect 2275 365 2325 395
rect 2355 365 2405 395
rect 2435 365 2485 395
rect 2515 365 2565 395
rect 2595 365 2645 395
rect 2675 365 2725 395
rect 2755 365 2805 395
rect 2835 365 2885 395
rect 2915 365 2965 395
rect 2995 365 3045 395
rect 3075 365 3125 395
rect 3155 365 3205 395
rect 3235 365 3285 395
rect 3315 365 3365 395
rect 3395 365 3445 395
rect 3475 365 3525 395
rect 3555 365 3605 395
rect 3635 365 3685 395
rect 3715 365 3765 395
rect 3795 365 3845 395
rect 3875 365 3925 395
rect 3955 365 4005 395
rect 4035 365 4085 395
rect 4115 365 4165 395
rect 4195 365 4245 395
rect 4275 365 4325 395
rect 4355 365 4405 395
rect 4435 365 4485 395
rect 4515 365 4565 395
rect 4595 365 4645 395
rect 4675 365 4725 395
rect 4755 365 4805 395
rect 4835 365 4885 395
rect 4915 365 5045 395
rect 5075 365 5205 395
rect 5235 365 5365 395
rect 5395 365 5525 395
rect 5555 365 5685 395
rect 5715 365 5720 395
rect -800 360 5720 365
rect -1520 315 -840 320
rect -1520 285 -1515 315
rect -1485 285 -1355 315
rect -1325 285 -1195 315
rect -1165 285 -1035 315
rect -1005 285 -875 315
rect -845 285 -840 315
rect -1520 280 -840 285
rect -800 315 5000 320
rect -800 285 2965 315
rect 2995 285 3285 315
rect 3315 285 3445 315
rect 3475 285 3605 315
rect 3635 285 3925 315
rect 3955 285 4085 315
rect 4115 285 4965 315
rect 4995 285 5000 315
rect -800 280 5000 285
rect 5040 315 5720 320
rect 5040 285 5045 315
rect 5075 285 5205 315
rect 5235 285 5365 315
rect 5395 285 5525 315
rect 5555 285 5685 315
rect 5715 285 5720 315
rect 5040 280 5720 285
rect -1520 235 -840 240
rect -1520 205 -1515 235
rect -1485 205 -1355 235
rect -1325 205 -1195 235
rect -1165 205 -1035 235
rect -1005 205 -875 235
rect -845 205 -840 235
rect -1520 200 -840 205
rect -800 235 5720 240
rect -800 205 -795 235
rect -765 205 -715 235
rect -685 205 -635 235
rect -605 205 -555 235
rect -525 205 -475 235
rect -445 205 -395 235
rect -365 205 -315 235
rect -285 205 -235 235
rect -205 205 -155 235
rect -125 205 -75 235
rect -45 205 5 235
rect 35 205 85 235
rect 115 205 165 235
rect 195 205 245 235
rect 275 205 325 235
rect 355 205 405 235
rect 435 205 485 235
rect 515 205 565 235
rect 595 205 645 235
rect 675 205 725 235
rect 755 205 805 235
rect 835 205 885 235
rect 915 205 965 235
rect 995 205 1045 235
rect 1075 205 1125 235
rect 1155 205 1205 235
rect 1235 205 1285 235
rect 1315 205 1365 235
rect 1395 205 1445 235
rect 1475 205 1525 235
rect 1555 205 1605 235
rect 1635 205 1685 235
rect 1715 205 1765 235
rect 1795 205 1845 235
rect 1875 205 1925 235
rect 1955 205 2005 235
rect 2035 205 2085 235
rect 2115 205 2165 235
rect 2195 205 2245 235
rect 2275 205 2325 235
rect 2355 205 2405 235
rect 2435 205 2485 235
rect 2515 205 2565 235
rect 2595 205 2645 235
rect 2675 205 2725 235
rect 2755 205 2805 235
rect 2835 205 2885 235
rect 2915 205 2965 235
rect 2995 205 3045 235
rect 3075 205 3125 235
rect 3155 205 3205 235
rect 3235 205 3285 235
rect 3315 205 3365 235
rect 3395 205 3445 235
rect 3475 205 3525 235
rect 3555 205 3605 235
rect 3635 205 3685 235
rect 3715 205 3765 235
rect 3795 205 3845 235
rect 3875 205 3925 235
rect 3955 205 4005 235
rect 4035 205 4085 235
rect 4115 205 4165 235
rect 4195 205 4245 235
rect 4275 205 4325 235
rect 4355 205 4405 235
rect 4435 205 4485 235
rect 4515 205 4565 235
rect 4595 205 4645 235
rect 4675 205 4725 235
rect 4755 205 4805 235
rect 4835 205 4885 235
rect 4915 205 5045 235
rect 5075 205 5205 235
rect 5235 205 5365 235
rect 5395 205 5525 235
rect 5555 205 5685 235
rect 5715 205 5720 235
rect -800 200 5720 205
rect -1520 155 -840 160
rect -1520 125 -1515 155
rect -1485 125 -1355 155
rect -1325 125 -1195 155
rect -1165 125 -1035 155
rect -1005 125 -875 155
rect -845 125 -840 155
rect -1520 120 -840 125
rect -800 155 5720 160
rect -800 125 -795 155
rect -765 125 -715 155
rect -685 125 -635 155
rect -605 125 -555 155
rect -525 125 -475 155
rect -445 125 -395 155
rect -365 125 -315 155
rect -285 125 -235 155
rect -205 125 -155 155
rect -125 125 -75 155
rect -45 125 5 155
rect 35 125 85 155
rect 115 125 165 155
rect 195 125 245 155
rect 275 125 325 155
rect 355 125 405 155
rect 435 125 485 155
rect 515 125 565 155
rect 595 125 645 155
rect 675 125 725 155
rect 755 125 805 155
rect 835 125 885 155
rect 915 125 965 155
rect 995 125 1045 155
rect 1075 125 1125 155
rect 1155 125 1205 155
rect 1235 125 1285 155
rect 1315 125 1365 155
rect 1395 125 1445 155
rect 1475 125 1525 155
rect 1555 125 1605 155
rect 1635 125 1685 155
rect 1715 125 1765 155
rect 1795 125 1845 155
rect 1875 125 1925 155
rect 1955 125 2005 155
rect 2035 125 2085 155
rect 2115 125 2165 155
rect 2195 125 2245 155
rect 2275 125 2325 155
rect 2355 125 2405 155
rect 2435 125 2485 155
rect 2515 125 2565 155
rect 2595 125 2645 155
rect 2675 125 2725 155
rect 2755 125 2805 155
rect 2835 125 2885 155
rect 2915 125 2965 155
rect 2995 125 3045 155
rect 3075 125 3125 155
rect 3155 125 3205 155
rect 3235 125 3285 155
rect 3315 125 3365 155
rect 3395 125 3445 155
rect 3475 125 3525 155
rect 3555 125 3605 155
rect 3635 125 3685 155
rect 3715 125 3765 155
rect 3795 125 3845 155
rect 3875 125 3925 155
rect 3955 125 4005 155
rect 4035 125 4085 155
rect 4115 125 4165 155
rect 4195 125 4245 155
rect 4275 125 4325 155
rect 4355 125 4405 155
rect 4435 125 4485 155
rect 4515 125 4565 155
rect 4595 125 4645 155
rect 4675 125 4725 155
rect 4755 125 4805 155
rect 4835 125 4885 155
rect 4915 125 5045 155
rect 5075 125 5205 155
rect 5235 125 5365 155
rect 5395 125 5525 155
rect 5555 125 5685 155
rect 5715 125 5720 155
rect -800 120 5720 125
rect -1520 75 -840 80
rect -1520 45 -1515 75
rect -1485 45 -1355 75
rect -1325 45 -1195 75
rect -1165 45 -1035 75
rect -1005 45 -875 75
rect -845 45 -840 75
rect -1520 40 -840 45
rect -800 75 5720 80
rect -800 45 -795 75
rect -765 45 -715 75
rect -685 45 -635 75
rect -605 45 -555 75
rect -525 45 -475 75
rect -445 45 -395 75
rect -365 45 -315 75
rect -285 45 -235 75
rect -205 45 -155 75
rect -125 45 -75 75
rect -45 45 5 75
rect 35 45 85 75
rect 115 45 165 75
rect 195 45 245 75
rect 275 45 325 75
rect 355 45 405 75
rect 435 45 485 75
rect 515 45 565 75
rect 595 45 645 75
rect 675 45 725 75
rect 755 45 805 75
rect 835 45 885 75
rect 915 45 965 75
rect 995 45 1045 75
rect 1075 45 1125 75
rect 1155 45 1205 75
rect 1235 45 1285 75
rect 1315 45 1365 75
rect 1395 45 1445 75
rect 1475 45 1525 75
rect 1555 45 1605 75
rect 1635 45 1685 75
rect 1715 45 1765 75
rect 1795 45 1845 75
rect 1875 45 1925 75
rect 1955 45 2005 75
rect 2035 45 2085 75
rect 2115 45 2165 75
rect 2195 45 2245 75
rect 2275 45 2325 75
rect 2355 45 2405 75
rect 2435 45 2485 75
rect 2515 45 2565 75
rect 2595 45 2645 75
rect 2675 45 2725 75
rect 2755 45 2805 75
rect 2835 45 2885 75
rect 2915 45 2965 75
rect 2995 45 3045 75
rect 3075 45 3125 75
rect 3155 45 3205 75
rect 3235 45 3285 75
rect 3315 45 3365 75
rect 3395 45 3445 75
rect 3475 45 3525 75
rect 3555 45 3605 75
rect 3635 45 3685 75
rect 3715 45 3765 75
rect 3795 45 3845 75
rect 3875 45 3925 75
rect 3955 45 4005 75
rect 4035 45 4085 75
rect 4115 45 4165 75
rect 4195 45 4245 75
rect 4275 45 4325 75
rect 4355 45 4405 75
rect 4435 45 4485 75
rect 4515 45 4565 75
rect 4595 45 4645 75
rect 4675 45 4725 75
rect 4755 45 4805 75
rect 4835 45 4885 75
rect 4915 45 5045 75
rect 5075 45 5205 75
rect 5235 45 5365 75
rect 5395 45 5525 75
rect 5555 45 5685 75
rect 5715 45 5720 75
rect -800 40 5720 45
rect -1520 -5 -840 0
rect -1520 -35 -1515 -5
rect -1485 -35 -1355 -5
rect -1325 -35 -1195 -5
rect -1165 -35 -1035 -5
rect -1005 -35 -875 -5
rect -845 -35 -840 -5
rect -1520 -40 -840 -35
rect -800 -5 5720 0
rect -800 -35 -795 -5
rect -765 -35 -715 -5
rect -685 -35 -635 -5
rect -605 -35 -555 -5
rect -525 -35 -475 -5
rect -445 -35 -395 -5
rect -365 -35 -315 -5
rect -285 -35 -235 -5
rect -205 -35 -155 -5
rect -125 -35 -75 -5
rect -45 -35 5 -5
rect 35 -35 85 -5
rect 115 -35 165 -5
rect 195 -35 245 -5
rect 275 -35 325 -5
rect 355 -35 405 -5
rect 435 -35 485 -5
rect 515 -35 565 -5
rect 595 -35 645 -5
rect 675 -35 725 -5
rect 755 -35 805 -5
rect 835 -35 885 -5
rect 915 -35 965 -5
rect 995 -35 1045 -5
rect 1075 -35 1125 -5
rect 1155 -35 1205 -5
rect 1235 -35 1285 -5
rect 1315 -35 1365 -5
rect 1395 -35 1445 -5
rect 1475 -35 1525 -5
rect 1555 -35 1605 -5
rect 1635 -35 1685 -5
rect 1715 -35 1765 -5
rect 1795 -35 1845 -5
rect 1875 -35 1925 -5
rect 1955 -35 2005 -5
rect 2035 -35 2085 -5
rect 2115 -35 2165 -5
rect 2195 -35 2245 -5
rect 2275 -35 2325 -5
rect 2355 -35 2405 -5
rect 2435 -35 2485 -5
rect 2515 -35 2565 -5
rect 2595 -35 2645 -5
rect 2675 -35 2725 -5
rect 2755 -35 2805 -5
rect 2835 -35 2885 -5
rect 2915 -35 2965 -5
rect 2995 -35 3045 -5
rect 3075 -35 3125 -5
rect 3155 -35 3205 -5
rect 3235 -35 3285 -5
rect 3315 -35 3365 -5
rect 3395 -35 3445 -5
rect 3475 -35 3525 -5
rect 3555 -35 3605 -5
rect 3635 -35 3685 -5
rect 3715 -35 3765 -5
rect 3795 -35 3845 -5
rect 3875 -35 3925 -5
rect 3955 -35 4005 -5
rect 4035 -35 4085 -5
rect 4115 -35 4165 -5
rect 4195 -35 4245 -5
rect 4275 -35 4325 -5
rect 4355 -35 4405 -5
rect 4435 -35 4485 -5
rect 4515 -35 4565 -5
rect 4595 -35 4645 -5
rect 4675 -35 4725 -5
rect 4755 -35 4805 -5
rect 4835 -35 4885 -5
rect 4915 -35 5045 -5
rect 5075 -35 5205 -5
rect 5235 -35 5365 -5
rect 5395 -35 5525 -5
rect 5555 -35 5685 -5
rect 5715 -35 5720 -5
rect -800 -40 5720 -35
rect -1520 -85 -840 -80
rect -1520 -115 -1515 -85
rect -1485 -115 -1355 -85
rect -1325 -115 -1195 -85
rect -1165 -115 -1035 -85
rect -1005 -115 -875 -85
rect -845 -115 -840 -85
rect -1520 -120 -840 -115
rect -800 -85 5720 -80
rect -800 -115 -795 -85
rect -765 -115 -715 -85
rect -685 -115 -635 -85
rect -605 -115 -555 -85
rect -525 -115 -475 -85
rect -445 -115 -395 -85
rect -365 -115 -315 -85
rect -285 -115 -235 -85
rect -205 -115 -155 -85
rect -125 -115 -75 -85
rect -45 -115 5 -85
rect 35 -115 85 -85
rect 115 -115 165 -85
rect 195 -115 245 -85
rect 275 -115 325 -85
rect 355 -115 405 -85
rect 435 -115 485 -85
rect 515 -115 565 -85
rect 595 -115 645 -85
rect 675 -115 725 -85
rect 755 -115 805 -85
rect 835 -115 885 -85
rect 915 -115 965 -85
rect 995 -115 1045 -85
rect 1075 -115 1125 -85
rect 1155 -115 1205 -85
rect 1235 -115 1285 -85
rect 1315 -115 1365 -85
rect 1395 -115 1445 -85
rect 1475 -115 1525 -85
rect 1555 -115 1605 -85
rect 1635 -115 1685 -85
rect 1715 -115 1765 -85
rect 1795 -115 1845 -85
rect 1875 -115 1925 -85
rect 1955 -115 2005 -85
rect 2035 -115 2085 -85
rect 2115 -115 2165 -85
rect 2195 -115 2245 -85
rect 2275 -115 2325 -85
rect 2355 -115 2405 -85
rect 2435 -115 2485 -85
rect 2515 -115 2565 -85
rect 2595 -115 2645 -85
rect 2675 -115 2725 -85
rect 2755 -115 2805 -85
rect 2835 -115 2885 -85
rect 2915 -115 2965 -85
rect 2995 -115 3045 -85
rect 3075 -115 3125 -85
rect 3155 -115 3205 -85
rect 3235 -115 3285 -85
rect 3315 -115 3365 -85
rect 3395 -115 3445 -85
rect 3475 -115 3525 -85
rect 3555 -115 3605 -85
rect 3635 -115 3685 -85
rect 3715 -115 3765 -85
rect 3795 -115 3845 -85
rect 3875 -115 3925 -85
rect 3955 -115 4005 -85
rect 4035 -115 4085 -85
rect 4115 -115 4165 -85
rect 4195 -115 4245 -85
rect 4275 -115 4325 -85
rect 4355 -115 4405 -85
rect 4435 -115 4485 -85
rect 4515 -115 4565 -85
rect 4595 -115 4645 -85
rect 4675 -115 4725 -85
rect 4755 -115 4805 -85
rect 4835 -115 4885 -85
rect 4915 -115 5045 -85
rect 5075 -115 5205 -85
rect 5235 -115 5365 -85
rect 5395 -115 5525 -85
rect 5555 -115 5685 -85
rect 5715 -115 5720 -85
rect -800 -120 5720 -115
<< via2 >>
rect -1515 5565 -1485 5595
rect -1355 5565 -1325 5595
rect -1195 5565 -1165 5595
rect -1035 5565 -1005 5595
rect -875 5565 -845 5595
rect 4885 5565 4915 5595
rect 5045 5565 5075 5595
rect 5205 5565 5235 5595
rect 5365 5565 5395 5595
rect 5525 5565 5555 5595
rect 5685 5565 5715 5595
rect -1515 5485 -1485 5515
rect -1355 5485 -1325 5515
rect -1195 5485 -1165 5515
rect -1035 5485 -1005 5515
rect -875 5485 -845 5515
rect -795 5485 -765 5515
rect -715 5485 -685 5515
rect -635 5485 -605 5515
rect -555 5485 -525 5515
rect -475 5485 -445 5515
rect -395 5485 -365 5515
rect -315 5485 -285 5515
rect -235 5485 -205 5515
rect -155 5485 -125 5515
rect -75 5485 -45 5515
rect 5 5485 35 5515
rect 85 5485 115 5515
rect 165 5485 195 5515
rect 245 5485 275 5515
rect 325 5485 355 5515
rect 405 5485 435 5515
rect 485 5485 515 5515
rect 565 5485 595 5515
rect 645 5485 675 5515
rect 725 5485 755 5515
rect 805 5485 835 5515
rect 885 5485 915 5515
rect 965 5485 995 5515
rect 1045 5485 1075 5515
rect 1125 5485 1155 5515
rect 1205 5485 1235 5515
rect 1285 5485 1315 5515
rect 1365 5485 1395 5515
rect 1445 5485 1475 5515
rect 1525 5485 1555 5515
rect 1605 5485 1635 5515
rect 1685 5485 1715 5515
rect 1765 5485 1795 5515
rect 1845 5485 1875 5515
rect 1925 5485 1955 5515
rect 2005 5485 2035 5515
rect 2085 5485 2115 5515
rect 2165 5485 2195 5515
rect 2245 5485 2275 5515
rect 2325 5485 2355 5515
rect 2405 5485 2435 5515
rect 2485 5485 2515 5515
rect 2565 5485 2595 5515
rect 2645 5485 2675 5515
rect 2725 5485 2755 5515
rect 2805 5485 2835 5515
rect 2885 5485 2915 5515
rect 2965 5485 2995 5515
rect 3045 5485 3075 5515
rect 3125 5485 3155 5515
rect 3205 5485 3235 5515
rect 3285 5485 3315 5515
rect 3365 5485 3395 5515
rect 3445 5485 3475 5515
rect 3525 5485 3555 5515
rect 3605 5485 3635 5515
rect 3685 5485 3715 5515
rect 3765 5485 3795 5515
rect 3845 5485 3875 5515
rect 3925 5485 3955 5515
rect 4005 5485 4035 5515
rect 4085 5485 4115 5515
rect 4165 5485 4195 5515
rect 4245 5485 4275 5515
rect 4325 5485 4355 5515
rect 4405 5485 4435 5515
rect 4485 5485 4515 5515
rect 4565 5485 4595 5515
rect 4645 5485 4675 5515
rect 4725 5485 4755 5515
rect 4805 5485 4835 5515
rect 4885 5485 4915 5515
rect 5045 5485 5075 5515
rect 5205 5485 5235 5515
rect 5365 5485 5395 5515
rect 5525 5485 5555 5515
rect 5685 5485 5715 5515
rect -1515 5405 -1485 5435
rect -1355 5405 -1325 5435
rect -1195 5405 -1165 5435
rect -1035 5405 -1005 5435
rect -875 5405 -845 5435
rect -795 5405 -765 5435
rect -715 5405 -685 5435
rect -635 5405 -605 5435
rect -555 5405 -525 5435
rect -475 5405 -445 5435
rect -395 5405 -365 5435
rect -315 5405 -285 5435
rect -235 5405 -205 5435
rect -155 5405 -125 5435
rect -75 5405 -45 5435
rect 5 5405 35 5435
rect 85 5405 115 5435
rect 165 5405 195 5435
rect 245 5405 275 5435
rect 325 5405 355 5435
rect 405 5405 435 5435
rect 485 5405 515 5435
rect 565 5405 595 5435
rect 645 5405 675 5435
rect 725 5405 755 5435
rect 805 5405 835 5435
rect 885 5405 915 5435
rect 965 5405 995 5435
rect 1045 5405 1075 5435
rect 1125 5405 1155 5435
rect 1205 5405 1235 5435
rect 1285 5405 1315 5435
rect 1365 5405 1395 5435
rect 1445 5405 1475 5435
rect 1525 5405 1555 5435
rect 1605 5405 1635 5435
rect 1685 5405 1715 5435
rect 1765 5405 1795 5435
rect 1845 5405 1875 5435
rect 1925 5405 1955 5435
rect 2005 5405 2035 5435
rect 2085 5405 2115 5435
rect 2165 5405 2195 5435
rect 2245 5405 2275 5435
rect 2325 5405 2355 5435
rect 2405 5405 2435 5435
rect 2485 5405 2515 5435
rect 2565 5405 2595 5435
rect 2645 5405 2675 5435
rect 2725 5405 2755 5435
rect 2805 5405 2835 5435
rect 2885 5405 2915 5435
rect 2965 5405 2995 5435
rect 3045 5405 3075 5435
rect 3125 5405 3155 5435
rect 3205 5405 3235 5435
rect 3285 5405 3315 5435
rect 3365 5405 3395 5435
rect 3445 5405 3475 5435
rect 3525 5405 3555 5435
rect 3605 5405 3635 5435
rect 3685 5405 3715 5435
rect 3765 5405 3795 5435
rect 3845 5405 3875 5435
rect 3925 5405 3955 5435
rect 4005 5405 4035 5435
rect 4085 5405 4115 5435
rect 4165 5405 4195 5435
rect 4245 5405 4275 5435
rect 4325 5405 4355 5435
rect 4405 5405 4435 5435
rect 4485 5405 4515 5435
rect 4565 5405 4595 5435
rect 4645 5405 4675 5435
rect 4725 5405 4755 5435
rect 4805 5405 4835 5435
rect 4885 5405 4915 5435
rect 5045 5405 5075 5435
rect 5205 5405 5235 5435
rect 5365 5405 5395 5435
rect 5525 5405 5555 5435
rect 5685 5405 5715 5435
rect -1515 5325 -1485 5355
rect -1355 5325 -1325 5355
rect -1195 5325 -1165 5355
rect -1035 5325 -1005 5355
rect -955 5325 -925 5355
rect 4885 5325 4915 5355
rect 5045 5325 5075 5355
rect 5205 5325 5235 5355
rect 5365 5325 5395 5355
rect 5525 5325 5555 5355
rect 5685 5325 5715 5355
rect -1515 5245 -1485 5275
rect -1355 5245 -1325 5275
rect -1195 5245 -1165 5275
rect -1035 5245 -1005 5275
rect -875 5245 -845 5275
rect -795 5245 -765 5275
rect -715 5245 -685 5275
rect -635 5245 -605 5275
rect -555 5245 -525 5275
rect -475 5245 -445 5275
rect -395 5245 -365 5275
rect -315 5245 -285 5275
rect -235 5245 -205 5275
rect -155 5245 -125 5275
rect -75 5245 -45 5275
rect 5 5245 35 5275
rect 85 5245 115 5275
rect 165 5245 195 5275
rect 245 5245 275 5275
rect 325 5245 355 5275
rect 405 5245 435 5275
rect 485 5245 515 5275
rect 565 5245 595 5275
rect 645 5245 675 5275
rect 725 5245 755 5275
rect 805 5245 835 5275
rect 885 5245 915 5275
rect 965 5245 995 5275
rect 1045 5245 1075 5275
rect 1125 5245 1155 5275
rect 1205 5245 1235 5275
rect 1285 5245 1315 5275
rect 1365 5245 1395 5275
rect 1445 5245 1475 5275
rect 1525 5245 1555 5275
rect 1605 5245 1635 5275
rect 1685 5245 1715 5275
rect 1765 5245 1795 5275
rect 1845 5245 1875 5275
rect 1925 5245 1955 5275
rect 2005 5245 2035 5275
rect 2085 5245 2115 5275
rect 2165 5245 2195 5275
rect 2245 5245 2275 5275
rect 2325 5245 2355 5275
rect 2405 5245 2435 5275
rect 2485 5245 2515 5275
rect 2565 5245 2595 5275
rect 2645 5245 2675 5275
rect 2725 5245 2755 5275
rect 2805 5245 2835 5275
rect 2885 5245 2915 5275
rect 2965 5245 2995 5275
rect 3045 5245 3075 5275
rect 3125 5245 3155 5275
rect 3205 5245 3235 5275
rect 3285 5245 3315 5275
rect 3365 5245 3395 5275
rect 3445 5245 3475 5275
rect 3525 5245 3555 5275
rect 3605 5245 3635 5275
rect 3685 5245 3715 5275
rect 3765 5245 3795 5275
rect 3845 5245 3875 5275
rect 3925 5245 3955 5275
rect 4005 5245 4035 5275
rect 4085 5245 4115 5275
rect 4165 5245 4195 5275
rect 4245 5245 4275 5275
rect 4325 5245 4355 5275
rect 4405 5245 4435 5275
rect 4485 5245 4515 5275
rect 4565 5245 4595 5275
rect 4645 5245 4675 5275
rect 4725 5245 4755 5275
rect 4805 5245 4835 5275
rect 4885 5245 4915 5275
rect 5045 5245 5075 5275
rect 5205 5245 5235 5275
rect 5365 5245 5395 5275
rect 5525 5245 5555 5275
rect 5685 5245 5715 5275
rect -1515 5165 -1485 5195
rect -1355 5165 -1325 5195
rect -1195 5165 -1165 5195
rect -1035 5165 -1005 5195
rect -875 5165 -845 5195
rect -795 5165 -765 5195
rect -715 5165 -685 5195
rect -635 5165 -605 5195
rect -555 5165 -525 5195
rect -475 5165 -445 5195
rect -395 5165 -365 5195
rect -315 5165 -285 5195
rect -235 5165 -205 5195
rect -155 5165 -125 5195
rect -75 5165 -45 5195
rect 5 5165 35 5195
rect 85 5165 115 5195
rect 165 5165 195 5195
rect 245 5165 275 5195
rect 325 5165 355 5195
rect 405 5165 435 5195
rect 485 5165 515 5195
rect 565 5165 595 5195
rect 645 5165 675 5195
rect 725 5165 755 5195
rect 805 5165 835 5195
rect 885 5165 915 5195
rect 965 5165 995 5195
rect 1045 5165 1075 5195
rect 1125 5165 1155 5195
rect 1205 5165 1235 5195
rect 1285 5165 1315 5195
rect 1365 5165 1395 5195
rect 1445 5165 1475 5195
rect 1525 5165 1555 5195
rect 1605 5165 1635 5195
rect 1685 5165 1715 5195
rect 1765 5165 1795 5195
rect 1845 5165 1875 5195
rect 1925 5165 1955 5195
rect 2005 5165 2035 5195
rect 2085 5165 2115 5195
rect 2165 5165 2195 5195
rect 2245 5165 2275 5195
rect 2325 5165 2355 5195
rect 2405 5165 2435 5195
rect 2485 5165 2515 5195
rect 2565 5165 2595 5195
rect 2645 5165 2675 5195
rect 2725 5165 2755 5195
rect 2805 5165 2835 5195
rect 2885 5165 2915 5195
rect 2965 5165 2995 5195
rect 3045 5165 3075 5195
rect 3125 5165 3155 5195
rect 3205 5165 3235 5195
rect 3285 5165 3315 5195
rect 3365 5165 3395 5195
rect 3445 5165 3475 5195
rect 3525 5165 3555 5195
rect 3605 5165 3635 5195
rect 3685 5165 3715 5195
rect 3765 5165 3795 5195
rect 3845 5165 3875 5195
rect 3925 5165 3955 5195
rect 4005 5165 4035 5195
rect 4085 5165 4115 5195
rect 4165 5165 4195 5195
rect 4245 5165 4275 5195
rect 4325 5165 4355 5195
rect 4405 5165 4435 5195
rect 4485 5165 4515 5195
rect 4565 5165 4595 5195
rect 4645 5165 4675 5195
rect 4725 5165 4755 5195
rect 4805 5165 4835 5195
rect 4885 5165 4915 5195
rect 5045 5165 5075 5195
rect 5205 5165 5235 5195
rect 5365 5165 5395 5195
rect 5525 5165 5555 5195
rect 5685 5165 5715 5195
rect -1515 5085 -1485 5115
rect -1355 5085 -1325 5115
rect -1195 5085 -1165 5115
rect -1035 5085 -1005 5115
rect -875 5085 -845 5115
rect -795 5085 -765 5115
rect -715 5085 -685 5115
rect -635 5085 -605 5115
rect -555 5085 -525 5115
rect -475 5085 -445 5115
rect -395 5085 -365 5115
rect -315 5085 -285 5115
rect -235 5085 -205 5115
rect -155 5085 -125 5115
rect -75 5085 -45 5115
rect 5 5085 35 5115
rect 85 5085 115 5115
rect 165 5085 195 5115
rect 245 5085 275 5115
rect 325 5085 355 5115
rect 405 5085 435 5115
rect 485 5085 515 5115
rect 565 5085 595 5115
rect 645 5085 675 5115
rect 725 5085 755 5115
rect 805 5085 835 5115
rect 885 5085 915 5115
rect 965 5085 995 5115
rect 1045 5085 1075 5115
rect 1125 5085 1155 5115
rect 1205 5085 1235 5115
rect 1285 5085 1315 5115
rect 1365 5085 1395 5115
rect 1445 5085 1475 5115
rect 1525 5085 1555 5115
rect 1605 5085 1635 5115
rect 1685 5085 1715 5115
rect 1765 5085 1795 5115
rect 1845 5085 1875 5115
rect 1925 5085 1955 5115
rect 2005 5085 2035 5115
rect 2085 5085 2115 5115
rect 2165 5085 2195 5115
rect 2245 5085 2275 5115
rect 2325 5085 2355 5115
rect 2405 5085 2435 5115
rect 2485 5085 2515 5115
rect 2565 5085 2595 5115
rect 2645 5085 2675 5115
rect 2725 5085 2755 5115
rect 2805 5085 2835 5115
rect 2885 5085 2915 5115
rect 2965 5085 2995 5115
rect 3045 5085 3075 5115
rect 3125 5085 3155 5115
rect 3205 5085 3235 5115
rect 3285 5085 3315 5115
rect 3365 5085 3395 5115
rect 3445 5085 3475 5115
rect 3525 5085 3555 5115
rect 3605 5085 3635 5115
rect 3685 5085 3715 5115
rect 3765 5085 3795 5115
rect 3845 5085 3875 5115
rect 3925 5085 3955 5115
rect 4005 5085 4035 5115
rect 4085 5085 4115 5115
rect 4165 5085 4195 5115
rect 4245 5085 4275 5115
rect 4325 5085 4355 5115
rect 4405 5085 4435 5115
rect 4485 5085 4515 5115
rect 4565 5085 4595 5115
rect 4645 5085 4675 5115
rect 4725 5085 4755 5115
rect 4805 5085 4835 5115
rect 4885 5085 4915 5115
rect 5045 5085 5075 5115
rect 5205 5085 5235 5115
rect 5365 5085 5395 5115
rect 5525 5085 5555 5115
rect 5685 5085 5715 5115
rect -1515 5005 -1485 5035
rect -1355 5005 -1325 5035
rect -1195 5005 -1165 5035
rect -1035 5005 -1005 5035
rect -875 5005 -845 5035
rect -795 5005 -765 5035
rect -715 5005 -685 5035
rect -635 5005 -605 5035
rect -555 5005 -525 5035
rect -475 5005 -445 5035
rect -395 5005 -365 5035
rect -315 5005 -285 5035
rect -235 5005 -205 5035
rect -155 5005 -125 5035
rect -75 5005 -45 5035
rect 5 5005 35 5035
rect 85 5005 115 5035
rect 165 5005 195 5035
rect 245 5005 275 5035
rect 325 5005 355 5035
rect 405 5005 435 5035
rect 485 5005 515 5035
rect 565 5005 595 5035
rect 645 5005 675 5035
rect 725 5005 755 5035
rect 805 5005 835 5035
rect 885 5005 915 5035
rect 965 5005 995 5035
rect 1045 5005 1075 5035
rect 1125 5005 1155 5035
rect 1205 5005 1235 5035
rect 1285 5005 1315 5035
rect 1365 5005 1395 5035
rect 1445 5005 1475 5035
rect 1525 5005 1555 5035
rect 1605 5005 1635 5035
rect 1685 5005 1715 5035
rect 1765 5005 1795 5035
rect 1845 5005 1875 5035
rect 1925 5005 1955 5035
rect 2005 5005 2035 5035
rect 2085 5005 2115 5035
rect 2165 5005 2195 5035
rect 2245 5005 2275 5035
rect 2325 5005 2355 5035
rect 2405 5005 2435 5035
rect 2485 5005 2515 5035
rect 2565 5005 2595 5035
rect 2645 5005 2675 5035
rect 2725 5005 2755 5035
rect 2805 5005 2835 5035
rect 2885 5005 2915 5035
rect 2965 5005 2995 5035
rect 3045 5005 3075 5035
rect 3125 5005 3155 5035
rect 3205 5005 3235 5035
rect 3285 5005 3315 5035
rect 3365 5005 3395 5035
rect 3445 5005 3475 5035
rect 3525 5005 3555 5035
rect 3605 5005 3635 5035
rect 3685 5005 3715 5035
rect 3765 5005 3795 5035
rect 3845 5005 3875 5035
rect 3925 5005 3955 5035
rect 4005 5005 4035 5035
rect 4085 5005 4115 5035
rect 4165 5005 4195 5035
rect 4245 5005 4275 5035
rect 4325 5005 4355 5035
rect 4405 5005 4435 5035
rect 4485 5005 4515 5035
rect 4565 5005 4595 5035
rect 4645 5005 4675 5035
rect 4725 5005 4755 5035
rect 4805 5005 4835 5035
rect 4885 5005 4915 5035
rect 5045 5005 5075 5035
rect 5205 5005 5235 5035
rect 5365 5005 5395 5035
rect 5525 5005 5555 5035
rect 5685 5005 5715 5035
rect -1515 4925 -1485 4955
rect -1355 4925 -1325 4955
rect -1195 4925 -1165 4955
rect -1115 4925 -1085 4955
rect 4885 4925 4915 4955
rect 5045 4925 5075 4955
rect 5205 4925 5235 4955
rect 5365 4925 5395 4955
rect 5525 4925 5555 4955
rect 5685 4925 5715 4955
rect -1515 4845 -1485 4875
rect -1355 4845 -1325 4875
rect -1195 4845 -1165 4875
rect -1035 4845 -1005 4875
rect -875 4845 -845 4875
rect -795 4845 -765 4875
rect -715 4845 -685 4875
rect -635 4845 -605 4875
rect -555 4845 -525 4875
rect -475 4845 -445 4875
rect -395 4845 -365 4875
rect -315 4845 -285 4875
rect -235 4845 -205 4875
rect -155 4845 -125 4875
rect -75 4845 -45 4875
rect 5 4845 35 4875
rect 85 4845 115 4875
rect 165 4845 195 4875
rect 245 4845 275 4875
rect 325 4845 355 4875
rect 405 4845 435 4875
rect 485 4845 515 4875
rect 565 4845 595 4875
rect 645 4845 675 4875
rect 725 4845 755 4875
rect 805 4845 835 4875
rect 885 4845 915 4875
rect 965 4845 995 4875
rect 1045 4845 1075 4875
rect 1125 4845 1155 4875
rect 1205 4845 1235 4875
rect 1285 4845 1315 4875
rect 1365 4845 1395 4875
rect 1445 4845 1475 4875
rect 1525 4845 1555 4875
rect 1605 4845 1635 4875
rect 1685 4845 1715 4875
rect 1765 4845 1795 4875
rect 1845 4845 1875 4875
rect 1925 4845 1955 4875
rect 2005 4845 2035 4875
rect 2085 4845 2115 4875
rect 2165 4845 2195 4875
rect 2245 4845 2275 4875
rect 2325 4845 2355 4875
rect 2405 4845 2435 4875
rect 2485 4845 2515 4875
rect 2565 4845 2595 4875
rect 2645 4845 2675 4875
rect 2725 4845 2755 4875
rect 2805 4845 2835 4875
rect 2885 4845 2915 4875
rect 2965 4845 2995 4875
rect 3045 4845 3075 4875
rect 3125 4845 3155 4875
rect 3205 4845 3235 4875
rect 3285 4845 3315 4875
rect 3365 4845 3395 4875
rect 3445 4845 3475 4875
rect 3525 4845 3555 4875
rect 3605 4845 3635 4875
rect 3685 4845 3715 4875
rect 3765 4845 3795 4875
rect 3845 4845 3875 4875
rect 3925 4845 3955 4875
rect 4005 4845 4035 4875
rect 4085 4845 4115 4875
rect 4165 4845 4195 4875
rect 4245 4845 4275 4875
rect 4325 4845 4355 4875
rect 4405 4845 4435 4875
rect 4485 4845 4515 4875
rect 4565 4845 4595 4875
rect 4645 4845 4675 4875
rect 4725 4845 4755 4875
rect 4805 4845 4835 4875
rect 4885 4845 4915 4875
rect 5045 4845 5075 4875
rect 5205 4845 5235 4875
rect 5365 4845 5395 4875
rect 5525 4845 5555 4875
rect 5685 4845 5715 4875
rect -1435 4765 -1405 4795
rect 4885 4765 4915 4795
rect 5045 4765 5075 4795
rect 5205 4765 5235 4795
rect 5365 4765 5395 4795
rect 5525 4765 5555 4795
rect 5685 4765 5715 4795
rect -1515 4685 -1485 4715
rect -1355 4685 -1325 4715
rect -1195 4685 -1165 4715
rect -1035 4685 -1005 4715
rect -875 4685 -845 4715
rect -795 4685 -765 4715
rect -715 4685 -685 4715
rect -635 4685 -605 4715
rect -555 4685 -525 4715
rect -475 4685 -445 4715
rect -395 4685 -365 4715
rect -315 4685 -285 4715
rect -235 4685 -205 4715
rect -155 4685 -125 4715
rect -75 4685 -45 4715
rect 5 4685 35 4715
rect 85 4685 115 4715
rect 165 4685 195 4715
rect 245 4685 275 4715
rect 325 4685 355 4715
rect 405 4685 435 4715
rect 485 4685 515 4715
rect 565 4685 595 4715
rect 645 4685 675 4715
rect 725 4685 755 4715
rect 805 4685 835 4715
rect 885 4685 915 4715
rect 965 4685 995 4715
rect 1045 4685 1075 4715
rect 1125 4685 1155 4715
rect 1205 4685 1235 4715
rect 1285 4685 1315 4715
rect 1365 4685 1395 4715
rect 1445 4685 1475 4715
rect 1525 4685 1555 4715
rect 1605 4685 1635 4715
rect 1685 4685 1715 4715
rect 1765 4685 1795 4715
rect 1845 4685 1875 4715
rect 1925 4685 1955 4715
rect 2005 4685 2035 4715
rect 2085 4685 2115 4715
rect 2165 4685 2195 4715
rect 2245 4685 2275 4715
rect 2325 4685 2355 4715
rect 2405 4685 2435 4715
rect 2485 4685 2515 4715
rect 2565 4685 2595 4715
rect 2645 4685 2675 4715
rect 2725 4685 2755 4715
rect 2805 4685 2835 4715
rect 2885 4685 2915 4715
rect 2965 4685 2995 4715
rect 3045 4685 3075 4715
rect 3125 4685 3155 4715
rect 3205 4685 3235 4715
rect 3285 4685 3315 4715
rect 3365 4685 3395 4715
rect 3445 4685 3475 4715
rect 3525 4685 3555 4715
rect 3605 4685 3635 4715
rect 3685 4685 3715 4715
rect 3765 4685 3795 4715
rect 3845 4685 3875 4715
rect 3925 4685 3955 4715
rect 4005 4685 4035 4715
rect 4085 4685 4115 4715
rect 4165 4685 4195 4715
rect 4245 4685 4275 4715
rect 4325 4685 4355 4715
rect 4405 4685 4435 4715
rect 4485 4685 4515 4715
rect 4565 4685 4595 4715
rect 4645 4685 4675 4715
rect 4725 4685 4755 4715
rect 4805 4685 4835 4715
rect 4885 4685 4915 4715
rect 5045 4685 5075 4715
rect 5205 4685 5235 4715
rect 5365 4685 5395 4715
rect 5525 4685 5555 4715
rect 5685 4685 5715 4715
rect -1515 4605 -1485 4635
rect -1355 4605 -1325 4635
rect -1195 4605 -1165 4635
rect -1035 4605 -1005 4635
rect -875 4605 -845 4635
rect -795 4605 -765 4635
rect -715 4605 -685 4635
rect -635 4605 -605 4635
rect -555 4605 -525 4635
rect -475 4605 -445 4635
rect -395 4605 -365 4635
rect -315 4605 -285 4635
rect -235 4605 -205 4635
rect -155 4605 -125 4635
rect -75 4605 -45 4635
rect 5 4605 35 4635
rect 85 4605 115 4635
rect 165 4605 195 4635
rect 245 4605 275 4635
rect 325 4605 355 4635
rect 405 4605 435 4635
rect 485 4605 515 4635
rect 565 4605 595 4635
rect 645 4605 675 4635
rect 725 4605 755 4635
rect 805 4605 835 4635
rect 885 4605 915 4635
rect 965 4605 995 4635
rect 1045 4605 1075 4635
rect 1125 4605 1155 4635
rect 1205 4605 1235 4635
rect 1285 4605 1315 4635
rect 1365 4605 1395 4635
rect 1445 4605 1475 4635
rect 1525 4605 1555 4635
rect 1605 4605 1635 4635
rect 1685 4605 1715 4635
rect 1765 4605 1795 4635
rect 1845 4605 1875 4635
rect 1925 4605 1955 4635
rect 2005 4605 2035 4635
rect 2085 4605 2115 4635
rect 2165 4605 2195 4635
rect 2245 4605 2275 4635
rect 2325 4605 2355 4635
rect 2405 4605 2435 4635
rect 2485 4605 2515 4635
rect 2565 4605 2595 4635
rect 2645 4605 2675 4635
rect 2725 4605 2755 4635
rect 2805 4605 2835 4635
rect 2885 4605 2915 4635
rect 2965 4605 2995 4635
rect 3045 4605 3075 4635
rect 3125 4605 3155 4635
rect 3205 4605 3235 4635
rect 3285 4605 3315 4635
rect 3365 4605 3395 4635
rect 3445 4605 3475 4635
rect 3525 4605 3555 4635
rect 3605 4605 3635 4635
rect 3685 4605 3715 4635
rect 3765 4605 3795 4635
rect 3845 4605 3875 4635
rect 3925 4605 3955 4635
rect 4005 4605 4035 4635
rect 4085 4605 4115 4635
rect 4165 4605 4195 4635
rect 4245 4605 4275 4635
rect 4325 4605 4355 4635
rect 4405 4605 4435 4635
rect 4485 4605 4515 4635
rect 4565 4605 4595 4635
rect 4645 4605 4675 4635
rect 4725 4605 4755 4635
rect 4805 4605 4835 4635
rect 4885 4605 4915 4635
rect 5045 4605 5075 4635
rect 5205 4605 5235 4635
rect 5365 4605 5395 4635
rect 5525 4605 5555 4635
rect 5685 4605 5715 4635
rect -1515 4525 -1485 4555
rect -1355 4525 -1325 4555
rect -1195 4525 -1165 4555
rect -1035 4525 -1005 4555
rect -955 4525 -925 4555
rect 4885 4525 4915 4555
rect 5045 4525 5075 4555
rect 5205 4525 5235 4555
rect 5365 4525 5395 4555
rect 5525 4525 5555 4555
rect 5685 4525 5715 4555
rect -1515 4445 -1485 4475
rect -1355 4445 -1325 4475
rect -1195 4445 -1165 4475
rect -1035 4445 -1005 4475
rect -875 4445 -845 4475
rect -795 4445 -765 4475
rect -715 4445 -685 4475
rect -635 4445 -605 4475
rect -555 4445 -525 4475
rect -475 4445 -445 4475
rect -395 4445 -365 4475
rect -315 4445 -285 4475
rect -235 4445 -205 4475
rect -155 4445 -125 4475
rect -75 4445 -45 4475
rect 5 4445 35 4475
rect 85 4445 115 4475
rect 165 4445 195 4475
rect 245 4445 275 4475
rect 325 4445 355 4475
rect 405 4445 435 4475
rect 485 4445 515 4475
rect 565 4445 595 4475
rect 645 4445 675 4475
rect 725 4445 755 4475
rect 805 4445 835 4475
rect 885 4445 915 4475
rect 965 4445 995 4475
rect 1045 4445 1075 4475
rect 1125 4445 1155 4475
rect 1205 4445 1235 4475
rect 1285 4445 1315 4475
rect 1365 4445 1395 4475
rect 1445 4445 1475 4475
rect 1525 4445 1555 4475
rect 1605 4445 1635 4475
rect 1685 4445 1715 4475
rect 1765 4445 1795 4475
rect 1845 4445 1875 4475
rect 1925 4445 1955 4475
rect 2005 4445 2035 4475
rect 2085 4445 2115 4475
rect 2165 4445 2195 4475
rect 2245 4445 2275 4475
rect 2325 4445 2355 4475
rect 2405 4445 2435 4475
rect 2485 4445 2515 4475
rect 2565 4445 2595 4475
rect 2645 4445 2675 4475
rect 2725 4445 2755 4475
rect 2805 4445 2835 4475
rect 2885 4445 2915 4475
rect 2965 4445 2995 4475
rect 3045 4445 3075 4475
rect 3125 4445 3155 4475
rect 3205 4445 3235 4475
rect 3285 4445 3315 4475
rect 3365 4445 3395 4475
rect 3445 4445 3475 4475
rect 3525 4445 3555 4475
rect 3605 4445 3635 4475
rect 3685 4445 3715 4475
rect 3765 4445 3795 4475
rect 3845 4445 3875 4475
rect 3925 4445 3955 4475
rect 4005 4445 4035 4475
rect 4085 4445 4115 4475
rect 4165 4445 4195 4475
rect 4245 4445 4275 4475
rect 4325 4445 4355 4475
rect 4405 4445 4435 4475
rect 4485 4445 4515 4475
rect 4565 4445 4595 4475
rect 4645 4445 4675 4475
rect 4725 4445 4755 4475
rect 4805 4445 4835 4475
rect 4885 4445 4915 4475
rect 5045 4445 5075 4475
rect 5205 4445 5235 4475
rect 5365 4445 5395 4475
rect 5525 4445 5555 4475
rect 5685 4445 5715 4475
rect -1515 4365 -1485 4395
rect -1355 4365 -1325 4395
rect -1195 4365 -1165 4395
rect -1035 4365 -1005 4395
rect -875 4365 -845 4395
rect -795 4365 -765 4395
rect -715 4365 -685 4395
rect -635 4365 -605 4395
rect -555 4365 -525 4395
rect -475 4365 -445 4395
rect -395 4365 -365 4395
rect -315 4365 -285 4395
rect -235 4365 -205 4395
rect -155 4365 -125 4395
rect -75 4365 -45 4395
rect 5 4365 35 4395
rect 85 4365 115 4395
rect 165 4365 195 4395
rect 245 4365 275 4395
rect 325 4365 355 4395
rect 405 4365 435 4395
rect 485 4365 515 4395
rect 565 4365 595 4395
rect 645 4365 675 4395
rect 725 4365 755 4395
rect 805 4365 835 4395
rect 885 4365 915 4395
rect 965 4365 995 4395
rect 1045 4365 1075 4395
rect 1125 4365 1155 4395
rect 1205 4365 1235 4395
rect 1285 4365 1315 4395
rect 1365 4365 1395 4395
rect 1445 4365 1475 4395
rect 1525 4365 1555 4395
rect 1605 4365 1635 4395
rect 1685 4365 1715 4395
rect 1765 4365 1795 4395
rect 1845 4365 1875 4395
rect 1925 4365 1955 4395
rect 2005 4365 2035 4395
rect 2085 4365 2115 4395
rect 2165 4365 2195 4395
rect 2245 4365 2275 4395
rect 2325 4365 2355 4395
rect 2405 4365 2435 4395
rect 2485 4365 2515 4395
rect 2565 4365 2595 4395
rect 2645 4365 2675 4395
rect 2725 4365 2755 4395
rect 2805 4365 2835 4395
rect 2885 4365 2915 4395
rect 2965 4365 2995 4395
rect 3045 4365 3075 4395
rect 3125 4365 3155 4395
rect 3205 4365 3235 4395
rect 3285 4365 3315 4395
rect 3365 4365 3395 4395
rect 3445 4365 3475 4395
rect 3525 4365 3555 4395
rect 3605 4365 3635 4395
rect 3685 4365 3715 4395
rect 3765 4365 3795 4395
rect 3845 4365 3875 4395
rect 3925 4365 3955 4395
rect 4005 4365 4035 4395
rect 4085 4365 4115 4395
rect 4165 4365 4195 4395
rect 4245 4365 4275 4395
rect 4325 4365 4355 4395
rect 4405 4365 4435 4395
rect 4485 4365 4515 4395
rect 4565 4365 4595 4395
rect 4645 4365 4675 4395
rect 4725 4365 4755 4395
rect 4805 4365 4835 4395
rect 4885 4365 4915 4395
rect 5045 4365 5075 4395
rect 5205 4365 5235 4395
rect 5365 4365 5395 4395
rect 5525 4365 5555 4395
rect 5685 4365 5715 4395
rect -1515 4285 -1485 4315
rect -1355 4285 -1325 4315
rect -1195 4285 -1165 4315
rect -1035 4285 -1005 4315
rect -875 4285 -845 4315
rect 5605 4285 5635 4315
rect -1515 4205 -1485 4235
rect -1355 4205 -1325 4235
rect -1195 4205 -1165 4235
rect -1035 4205 -1005 4235
rect -875 4205 -845 4235
rect -795 4205 -765 4235
rect -715 4205 -685 4235
rect -635 4205 -605 4235
rect -555 4205 -525 4235
rect -475 4205 -445 4235
rect -395 4205 -365 4235
rect -315 4205 -285 4235
rect -235 4205 -205 4235
rect -155 4205 -125 4235
rect -75 4205 -45 4235
rect 5 4205 35 4235
rect 85 4205 115 4235
rect 165 4205 195 4235
rect 245 4205 275 4235
rect 325 4205 355 4235
rect 405 4205 435 4235
rect 485 4205 515 4235
rect 565 4205 595 4235
rect 645 4205 675 4235
rect 725 4205 755 4235
rect 805 4205 835 4235
rect 885 4205 915 4235
rect 965 4205 995 4235
rect 1045 4205 1075 4235
rect 1125 4205 1155 4235
rect 1205 4205 1235 4235
rect 1285 4205 1315 4235
rect 1365 4205 1395 4235
rect 1445 4205 1475 4235
rect 1525 4205 1555 4235
rect 1605 4205 1635 4235
rect 1685 4205 1715 4235
rect 1765 4205 1795 4235
rect 1845 4205 1875 4235
rect 1925 4205 1955 4235
rect 2005 4205 2035 4235
rect 2085 4205 2115 4235
rect 2165 4205 2195 4235
rect 2245 4205 2275 4235
rect 2325 4205 2355 4235
rect 2405 4205 2435 4235
rect 2485 4205 2515 4235
rect 2565 4205 2595 4235
rect 2645 4205 2675 4235
rect 2725 4205 2755 4235
rect 2805 4205 2835 4235
rect 2885 4205 2915 4235
rect 2965 4205 2995 4235
rect 3045 4205 3075 4235
rect 3125 4205 3155 4235
rect 3205 4205 3235 4235
rect 3285 4205 3315 4235
rect 3365 4205 3395 4235
rect 3445 4205 3475 4235
rect 3525 4205 3555 4235
rect 3605 4205 3635 4235
rect 3685 4205 3715 4235
rect 3765 4205 3795 4235
rect 3845 4205 3875 4235
rect 3925 4205 3955 4235
rect 4005 4205 4035 4235
rect 4085 4205 4115 4235
rect 4165 4205 4195 4235
rect 4245 4205 4275 4235
rect 4325 4205 4355 4235
rect 4405 4205 4435 4235
rect 4485 4205 4515 4235
rect 4565 4205 4595 4235
rect 4645 4205 4675 4235
rect 4725 4205 4755 4235
rect 4805 4205 4835 4235
rect 4885 4205 4915 4235
rect 5045 4205 5075 4235
rect 5205 4205 5235 4235
rect 5365 4205 5395 4235
rect 5525 4205 5555 4235
rect 5685 4205 5715 4235
rect -1515 4125 -1485 4155
rect -1355 4125 -1325 4155
rect -1195 4125 -1165 4155
rect -1035 4125 -1005 4155
rect -875 4125 -845 4155
rect 4965 4125 4995 4155
rect 5045 4125 5075 4155
rect 5205 4125 5235 4155
rect 5365 4125 5395 4155
rect 5525 4125 5555 4155
rect 5685 4125 5715 4155
rect -1515 4045 -1485 4075
rect -1355 4045 -1325 4075
rect -1195 4045 -1165 4075
rect -1035 4045 -1005 4075
rect -875 4045 -845 4075
rect -795 4045 -765 4075
rect -715 4045 -685 4075
rect -635 4045 -605 4075
rect -555 4045 -525 4075
rect -475 4045 -445 4075
rect -395 4045 -365 4075
rect -315 4045 -285 4075
rect -235 4045 -205 4075
rect -155 4045 -125 4075
rect -75 4045 -45 4075
rect 5 4045 35 4075
rect 85 4045 115 4075
rect 165 4045 195 4075
rect 245 4045 275 4075
rect 325 4045 355 4075
rect 405 4045 435 4075
rect 485 4045 515 4075
rect 565 4045 595 4075
rect 645 4045 675 4075
rect 725 4045 755 4075
rect 805 4045 835 4075
rect 885 4045 915 4075
rect 965 4045 995 4075
rect 1045 4045 1075 4075
rect 1125 4045 1155 4075
rect 1205 4045 1235 4075
rect 1285 4045 1315 4075
rect 1365 4045 1395 4075
rect 1445 4045 1475 4075
rect 1525 4045 1555 4075
rect 1605 4045 1635 4075
rect 1685 4045 1715 4075
rect 1765 4045 1795 4075
rect 1845 4045 1875 4075
rect 1925 4045 1955 4075
rect 2005 4045 2035 4075
rect 2085 4045 2115 4075
rect 2165 4045 2195 4075
rect 2245 4045 2275 4075
rect 2325 4045 2355 4075
rect 2405 4045 2435 4075
rect 2485 4045 2515 4075
rect 2565 4045 2595 4075
rect 2645 4045 2675 4075
rect 2725 4045 2755 4075
rect 2805 4045 2835 4075
rect 2885 4045 2915 4075
rect 2965 4045 2995 4075
rect 3045 4045 3075 4075
rect 3125 4045 3155 4075
rect 3205 4045 3235 4075
rect 3285 4045 3315 4075
rect 3365 4045 3395 4075
rect 3445 4045 3475 4075
rect 3525 4045 3555 4075
rect 3605 4045 3635 4075
rect 3685 4045 3715 4075
rect 3765 4045 3795 4075
rect 3845 4045 3875 4075
rect 3925 4045 3955 4075
rect 4005 4045 4035 4075
rect 4085 4045 4115 4075
rect 4165 4045 4195 4075
rect 4245 4045 4275 4075
rect 4325 4045 4355 4075
rect 4405 4045 4435 4075
rect 4485 4045 4515 4075
rect 4565 4045 4595 4075
rect 4645 4045 4675 4075
rect 4725 4045 4755 4075
rect 4805 4045 4835 4075
rect 4885 4045 4915 4075
rect 5045 4045 5075 4075
rect 5205 4045 5235 4075
rect 5365 4045 5395 4075
rect 5525 4045 5555 4075
rect 5685 4045 5715 4075
rect -1515 3965 -1485 3995
rect -1355 3965 -1325 3995
rect -1195 3965 -1165 3995
rect -1035 3965 -1005 3995
rect -875 3965 -845 3995
rect -795 3965 -765 3995
rect -715 3965 -685 3995
rect -635 3965 -605 3995
rect -555 3965 -525 3995
rect -475 3965 -445 3995
rect -395 3965 -365 3995
rect -315 3965 -285 3995
rect -235 3965 -205 3995
rect -155 3965 -125 3995
rect -75 3965 -45 3995
rect 5 3965 35 3995
rect 85 3965 115 3995
rect 165 3965 195 3995
rect 245 3965 275 3995
rect 325 3965 355 3995
rect 405 3965 435 3995
rect 485 3965 515 3995
rect 565 3965 595 3995
rect 645 3965 675 3995
rect 725 3965 755 3995
rect 805 3965 835 3995
rect 885 3965 915 3995
rect 965 3965 995 3995
rect 1045 3965 1075 3995
rect 1125 3965 1155 3995
rect 1205 3965 1235 3995
rect 1285 3965 1315 3995
rect 1365 3965 1395 3995
rect 1445 3965 1475 3995
rect 1525 3965 1555 3995
rect 1605 3965 1635 3995
rect 1685 3965 1715 3995
rect 1765 3965 1795 3995
rect 1845 3965 1875 3995
rect 1925 3965 1955 3995
rect 2005 3965 2035 3995
rect 2085 3965 2115 3995
rect 2165 3965 2195 3995
rect 2245 3965 2275 3995
rect 2325 3965 2355 3995
rect 2405 3965 2435 3995
rect 2485 3965 2515 3995
rect 2565 3965 2595 3995
rect 2645 3965 2675 3995
rect 2725 3965 2755 3995
rect 2805 3965 2835 3995
rect 2885 3965 2915 3995
rect 2965 3965 2995 3995
rect 3045 3965 3075 3995
rect 3125 3965 3155 3995
rect 3205 3965 3235 3995
rect 3285 3965 3315 3995
rect 3365 3965 3395 3995
rect 3445 3965 3475 3995
rect 3525 3965 3555 3995
rect 3605 3965 3635 3995
rect 3685 3965 3715 3995
rect 3765 3965 3795 3995
rect 3845 3965 3875 3995
rect 3925 3965 3955 3995
rect 4005 3965 4035 3995
rect 4085 3965 4115 3995
rect 4165 3965 4195 3995
rect 4245 3965 4275 3995
rect 4325 3965 4355 3995
rect 4405 3965 4435 3995
rect 4485 3965 4515 3995
rect 4565 3965 4595 3995
rect 4645 3965 4675 3995
rect 4725 3965 4755 3995
rect 4805 3965 4835 3995
rect 4885 3965 4915 3995
rect 5045 3965 5075 3995
rect 5205 3965 5235 3995
rect 5365 3965 5395 3995
rect 5525 3965 5555 3995
rect 5685 3965 5715 3995
rect -1515 3885 -1485 3915
rect -1355 3885 -1325 3915
rect -1195 3885 -1165 3915
rect -1035 3885 -1005 3915
rect -875 3885 -845 3915
rect -795 3885 -765 3915
rect -715 3885 -685 3915
rect -635 3885 -605 3915
rect -555 3885 -525 3915
rect -475 3885 -445 3915
rect -395 3885 -365 3915
rect -315 3885 -285 3915
rect -235 3885 -205 3915
rect -155 3885 -125 3915
rect -75 3885 -45 3915
rect 5 3885 35 3915
rect 85 3885 115 3915
rect 165 3885 195 3915
rect 245 3885 275 3915
rect 325 3885 355 3915
rect 405 3885 435 3915
rect 485 3885 515 3915
rect 565 3885 595 3915
rect 645 3885 675 3915
rect 725 3885 755 3915
rect 805 3885 835 3915
rect 885 3885 915 3915
rect 965 3885 995 3915
rect 1045 3885 1075 3915
rect 1125 3885 1155 3915
rect 1205 3885 1235 3915
rect 1285 3885 1315 3915
rect 1365 3885 1395 3915
rect 1445 3885 1475 3915
rect 1525 3885 1555 3915
rect 1605 3885 1635 3915
rect 1685 3885 1715 3915
rect 1765 3885 1795 3915
rect 1845 3885 1875 3915
rect 1925 3885 1955 3915
rect 2005 3885 2035 3915
rect 2085 3885 2115 3915
rect 2165 3885 2195 3915
rect 2245 3885 2275 3915
rect 2325 3885 2355 3915
rect 2405 3885 2435 3915
rect 2485 3885 2515 3915
rect 2565 3885 2595 3915
rect 2645 3885 2675 3915
rect 2725 3885 2755 3915
rect 2805 3885 2835 3915
rect 2885 3885 2915 3915
rect 2965 3885 2995 3915
rect 3045 3885 3075 3915
rect 3125 3885 3155 3915
rect 3205 3885 3235 3915
rect 3285 3885 3315 3915
rect 3365 3885 3395 3915
rect 3445 3885 3475 3915
rect 3525 3885 3555 3915
rect 3605 3885 3635 3915
rect 3685 3885 3715 3915
rect 3765 3885 3795 3915
rect 3845 3885 3875 3915
rect 3925 3885 3955 3915
rect 4005 3885 4035 3915
rect 4085 3885 4115 3915
rect 4165 3885 4195 3915
rect 4245 3885 4275 3915
rect 4325 3885 4355 3915
rect 4405 3885 4435 3915
rect 4485 3885 4515 3915
rect 4565 3885 4595 3915
rect 4645 3885 4675 3915
rect 4725 3885 4755 3915
rect 4805 3885 4835 3915
rect 4885 3885 4915 3915
rect 5045 3885 5075 3915
rect 5205 3885 5235 3915
rect 5365 3885 5395 3915
rect 5525 3885 5555 3915
rect 5685 3885 5715 3915
rect -1515 3805 -1485 3835
rect -1355 3805 -1325 3835
rect -1195 3805 -1165 3835
rect -1035 3805 -1005 3835
rect -875 3805 -845 3835
rect -795 3805 -765 3835
rect -715 3805 -685 3835
rect -635 3805 -605 3835
rect -555 3805 -525 3835
rect -475 3805 -445 3835
rect -395 3805 -365 3835
rect -315 3805 -285 3835
rect -235 3805 -205 3835
rect -155 3805 -125 3835
rect -75 3805 -45 3835
rect 5 3805 35 3835
rect 85 3805 115 3835
rect 165 3805 195 3835
rect 245 3805 275 3835
rect 325 3805 355 3835
rect 405 3805 435 3835
rect 485 3805 515 3835
rect 565 3805 595 3835
rect 645 3805 675 3835
rect 725 3805 755 3835
rect 805 3805 835 3835
rect 885 3805 915 3835
rect 965 3805 995 3835
rect 1045 3805 1075 3835
rect 1125 3805 1155 3835
rect 1205 3805 1235 3835
rect 1285 3805 1315 3835
rect 1365 3805 1395 3835
rect 1445 3805 1475 3835
rect 1525 3805 1555 3835
rect 1605 3805 1635 3835
rect 1685 3805 1715 3835
rect 1765 3805 1795 3835
rect 1845 3805 1875 3835
rect 1925 3805 1955 3835
rect 2005 3805 2035 3835
rect 2085 3805 2115 3835
rect 2165 3805 2195 3835
rect 2245 3805 2275 3835
rect 2325 3805 2355 3835
rect 2405 3805 2435 3835
rect 2485 3805 2515 3835
rect 2565 3805 2595 3835
rect 2645 3805 2675 3835
rect 2725 3805 2755 3835
rect 2805 3805 2835 3835
rect 2885 3805 2915 3835
rect 2965 3805 2995 3835
rect 3045 3805 3075 3835
rect 3125 3805 3155 3835
rect 3205 3805 3235 3835
rect 3285 3805 3315 3835
rect 3365 3805 3395 3835
rect 3445 3805 3475 3835
rect 3525 3805 3555 3835
rect 3605 3805 3635 3835
rect 3685 3805 3715 3835
rect 3765 3805 3795 3835
rect 3845 3805 3875 3835
rect 3925 3805 3955 3835
rect 4005 3805 4035 3835
rect 4085 3805 4115 3835
rect 4165 3805 4195 3835
rect 4245 3805 4275 3835
rect 4325 3805 4355 3835
rect 4405 3805 4435 3835
rect 4485 3805 4515 3835
rect 4565 3805 4595 3835
rect 4645 3805 4675 3835
rect 4725 3805 4755 3835
rect 4805 3805 4835 3835
rect 4885 3805 4915 3835
rect 5045 3805 5075 3835
rect 5205 3805 5235 3835
rect 5365 3805 5395 3835
rect 5525 3805 5555 3835
rect 5685 3805 5715 3835
rect -1515 3725 -1485 3755
rect -1355 3725 -1325 3755
rect -1195 3725 -1165 3755
rect -1035 3725 -1005 3755
rect -875 3725 -845 3755
rect -795 3725 -765 3755
rect -715 3725 -685 3755
rect -635 3725 -605 3755
rect -555 3725 -525 3755
rect -475 3725 -445 3755
rect -395 3725 -365 3755
rect -315 3725 -285 3755
rect -235 3725 -205 3755
rect -155 3725 -125 3755
rect -75 3725 -45 3755
rect 5 3725 35 3755
rect 85 3725 115 3755
rect 165 3725 195 3755
rect 245 3725 275 3755
rect 325 3725 355 3755
rect 405 3725 435 3755
rect 485 3725 515 3755
rect 565 3725 595 3755
rect 645 3725 675 3755
rect 725 3725 755 3755
rect 805 3725 835 3755
rect 885 3725 915 3755
rect 965 3725 995 3755
rect 1045 3725 1075 3755
rect 1125 3725 1155 3755
rect 1205 3725 1235 3755
rect 1285 3725 1315 3755
rect 1365 3725 1395 3755
rect 1445 3725 1475 3755
rect 1525 3725 1555 3755
rect 1605 3725 1635 3755
rect 1685 3725 1715 3755
rect 1765 3725 1795 3755
rect 1845 3725 1875 3755
rect 1925 3725 1955 3755
rect 2005 3725 2035 3755
rect 2085 3725 2115 3755
rect 2165 3725 2195 3755
rect 2245 3725 2275 3755
rect 2325 3725 2355 3755
rect 2405 3725 2435 3755
rect 2485 3725 2515 3755
rect 2565 3725 2595 3755
rect 2645 3725 2675 3755
rect 2725 3725 2755 3755
rect 2805 3725 2835 3755
rect 2885 3725 2915 3755
rect 2965 3725 2995 3755
rect 3045 3725 3075 3755
rect 3125 3725 3155 3755
rect 3205 3725 3235 3755
rect 3285 3725 3315 3755
rect 3365 3725 3395 3755
rect 3445 3725 3475 3755
rect 3525 3725 3555 3755
rect 3605 3725 3635 3755
rect 3685 3725 3715 3755
rect 3765 3725 3795 3755
rect 3845 3725 3875 3755
rect 3925 3725 3955 3755
rect 4005 3725 4035 3755
rect 4085 3725 4115 3755
rect 4165 3725 4195 3755
rect 4245 3725 4275 3755
rect 4325 3725 4355 3755
rect 4405 3725 4435 3755
rect 4485 3725 4515 3755
rect 4565 3725 4595 3755
rect 4645 3725 4675 3755
rect 4725 3725 4755 3755
rect 4805 3725 4835 3755
rect 4885 3725 4915 3755
rect 5045 3725 5075 3755
rect 5205 3725 5235 3755
rect 5365 3725 5395 3755
rect 5525 3725 5555 3755
rect 5685 3725 5715 3755
rect -1515 3645 -1485 3675
rect -1355 3645 -1325 3675
rect -1195 3645 -1165 3675
rect -1035 3645 -1005 3675
rect -875 3645 -845 3675
rect -795 3645 -765 3675
rect -715 3645 -685 3675
rect -635 3645 -605 3675
rect -555 3645 -525 3675
rect -475 3645 -445 3675
rect -395 3645 -365 3675
rect -315 3645 -285 3675
rect -235 3645 -205 3675
rect -155 3645 -125 3675
rect -75 3645 -45 3675
rect 5 3645 35 3675
rect 85 3645 115 3675
rect 165 3645 195 3675
rect 245 3645 275 3675
rect 325 3645 355 3675
rect 405 3645 435 3675
rect 485 3645 515 3675
rect 565 3645 595 3675
rect 645 3645 675 3675
rect 725 3645 755 3675
rect 805 3645 835 3675
rect 885 3645 915 3675
rect 965 3645 995 3675
rect 1045 3645 1075 3675
rect 1125 3645 1155 3675
rect 1205 3645 1235 3675
rect 1285 3645 1315 3675
rect 1365 3645 1395 3675
rect 1445 3645 1475 3675
rect 1525 3645 1555 3675
rect 1605 3645 1635 3675
rect 1685 3645 1715 3675
rect 1765 3645 1795 3675
rect 1845 3645 1875 3675
rect 1925 3645 1955 3675
rect 2005 3645 2035 3675
rect 2085 3645 2115 3675
rect 2165 3645 2195 3675
rect 2245 3645 2275 3675
rect 2325 3645 2355 3675
rect 2405 3645 2435 3675
rect 2485 3645 2515 3675
rect 2565 3645 2595 3675
rect 2645 3645 2675 3675
rect 2725 3645 2755 3675
rect 2805 3645 2835 3675
rect 2885 3645 2915 3675
rect 2965 3645 2995 3675
rect 3045 3645 3075 3675
rect 3125 3645 3155 3675
rect 3205 3645 3235 3675
rect 3285 3645 3315 3675
rect 3365 3645 3395 3675
rect 3445 3645 3475 3675
rect 3525 3645 3555 3675
rect 3605 3645 3635 3675
rect 3685 3645 3715 3675
rect 3765 3645 3795 3675
rect 3845 3645 3875 3675
rect 3925 3645 3955 3675
rect 4005 3645 4035 3675
rect 4085 3645 4115 3675
rect 4165 3645 4195 3675
rect 4245 3645 4275 3675
rect 4325 3645 4355 3675
rect 4405 3645 4435 3675
rect 4485 3645 4515 3675
rect 4565 3645 4595 3675
rect 4645 3645 4675 3675
rect 4725 3645 4755 3675
rect 4805 3645 4835 3675
rect 4885 3645 4915 3675
rect 5045 3645 5075 3675
rect 5205 3645 5235 3675
rect 5365 3645 5395 3675
rect 5525 3645 5555 3675
rect 5685 3645 5715 3675
rect -1515 3565 -1485 3595
rect -1355 3565 -1325 3595
rect -1195 3565 -1165 3595
rect -1035 3565 -1005 3595
rect -875 3565 -845 3595
rect -795 3565 -765 3595
rect -715 3565 -685 3595
rect -635 3565 -605 3595
rect -555 3565 -525 3595
rect -475 3565 -445 3595
rect -395 3565 -365 3595
rect -315 3565 -285 3595
rect -235 3565 -205 3595
rect -155 3565 -125 3595
rect -75 3565 -45 3595
rect 5 3565 35 3595
rect 85 3565 115 3595
rect 165 3565 195 3595
rect 245 3565 275 3595
rect 325 3565 355 3595
rect 405 3565 435 3595
rect 485 3565 515 3595
rect 565 3565 595 3595
rect 645 3565 675 3595
rect 725 3565 755 3595
rect 805 3565 835 3595
rect 885 3565 915 3595
rect 965 3565 995 3595
rect 1045 3565 1075 3595
rect 1125 3565 1155 3595
rect 1205 3565 1235 3595
rect 1285 3565 1315 3595
rect 1365 3565 1395 3595
rect 1445 3565 1475 3595
rect 1525 3565 1555 3595
rect 1605 3565 1635 3595
rect 1685 3565 1715 3595
rect 1765 3565 1795 3595
rect 1845 3565 1875 3595
rect 1925 3565 1955 3595
rect 2005 3565 2035 3595
rect 2085 3565 2115 3595
rect 2165 3565 2195 3595
rect 2245 3565 2275 3595
rect 2325 3565 2355 3595
rect 2405 3565 2435 3595
rect 2485 3565 2515 3595
rect 2565 3565 2595 3595
rect 2645 3565 2675 3595
rect 2725 3565 2755 3595
rect 2805 3565 2835 3595
rect 2885 3565 2915 3595
rect 2965 3565 2995 3595
rect 3045 3565 3075 3595
rect 3125 3565 3155 3595
rect 3205 3565 3235 3595
rect 3285 3565 3315 3595
rect 3365 3565 3395 3595
rect 3445 3565 3475 3595
rect 3525 3565 3555 3595
rect 3605 3565 3635 3595
rect 3685 3565 3715 3595
rect 3765 3565 3795 3595
rect 3845 3565 3875 3595
rect 3925 3565 3955 3595
rect 4005 3565 4035 3595
rect 4085 3565 4115 3595
rect 4165 3565 4195 3595
rect 4245 3565 4275 3595
rect 4325 3565 4355 3595
rect 4405 3565 4435 3595
rect 4485 3565 4515 3595
rect 4565 3565 4595 3595
rect 4645 3565 4675 3595
rect 4725 3565 4755 3595
rect 4805 3565 4835 3595
rect 4885 3565 4915 3595
rect 5045 3565 5075 3595
rect 5205 3565 5235 3595
rect 5365 3565 5395 3595
rect 5525 3565 5555 3595
rect 5685 3565 5715 3595
rect -1515 3485 -1485 3515
rect -1355 3485 -1325 3515
rect -1195 3485 -1165 3515
rect -1035 3485 -1005 3515
rect -875 3485 -845 3515
rect -795 3485 -765 3515
rect -715 3485 -685 3515
rect -635 3485 -605 3515
rect -555 3485 -525 3515
rect -475 3485 -445 3515
rect -395 3485 -365 3515
rect -315 3485 -285 3515
rect -235 3485 -205 3515
rect -155 3485 -125 3515
rect -75 3485 -45 3515
rect 5 3485 35 3515
rect 85 3485 115 3515
rect 165 3485 195 3515
rect 245 3485 275 3515
rect 325 3485 355 3515
rect 405 3485 435 3515
rect 485 3485 515 3515
rect 565 3485 595 3515
rect 645 3485 675 3515
rect 725 3485 755 3515
rect 805 3485 835 3515
rect 885 3485 915 3515
rect 965 3485 995 3515
rect 1045 3485 1075 3515
rect 1125 3485 1155 3515
rect 1205 3485 1235 3515
rect 1285 3485 1315 3515
rect 1365 3485 1395 3515
rect 1445 3485 1475 3515
rect 1525 3485 1555 3515
rect 1605 3485 1635 3515
rect 1685 3485 1715 3515
rect 1765 3485 1795 3515
rect 1845 3485 1875 3515
rect 1925 3485 1955 3515
rect 2005 3485 2035 3515
rect 2085 3485 2115 3515
rect 2165 3485 2195 3515
rect 2245 3485 2275 3515
rect 2325 3485 2355 3515
rect 2405 3485 2435 3515
rect 2485 3485 2515 3515
rect 2565 3485 2595 3515
rect 2645 3485 2675 3515
rect 2725 3485 2755 3515
rect 2805 3485 2835 3515
rect 2885 3485 2915 3515
rect 2965 3485 2995 3515
rect 3045 3485 3075 3515
rect 3125 3485 3155 3515
rect 3205 3485 3235 3515
rect 3285 3485 3315 3515
rect 3365 3485 3395 3515
rect 3445 3485 3475 3515
rect 3525 3485 3555 3515
rect 3605 3485 3635 3515
rect 3685 3485 3715 3515
rect 3765 3485 3795 3515
rect 3845 3485 3875 3515
rect 3925 3485 3955 3515
rect 4005 3485 4035 3515
rect 4085 3485 4115 3515
rect 4165 3485 4195 3515
rect 4245 3485 4275 3515
rect 4325 3485 4355 3515
rect 4405 3485 4435 3515
rect 4485 3485 4515 3515
rect 4565 3485 4595 3515
rect 4645 3485 4675 3515
rect 4725 3485 4755 3515
rect 4805 3485 4835 3515
rect 4885 3485 4915 3515
rect 5045 3485 5075 3515
rect 5205 3485 5235 3515
rect 5365 3485 5395 3515
rect 5525 3485 5555 3515
rect 5685 3485 5715 3515
rect -1515 3405 -1485 3435
rect -1355 3405 -1325 3435
rect -1275 3405 -1245 3435
rect 4885 3405 4915 3435
rect 5045 3405 5075 3435
rect 5205 3405 5235 3435
rect 5365 3405 5395 3435
rect 5525 3405 5555 3435
rect 5685 3405 5715 3435
rect -1515 3325 -1485 3355
rect -1355 3325 -1325 3355
rect -1195 3325 -1165 3355
rect -1035 3325 -1005 3355
rect -875 3325 -845 3355
rect -795 3325 -765 3355
rect -715 3325 -685 3355
rect -635 3325 -605 3355
rect -555 3325 -525 3355
rect -475 3325 -445 3355
rect -395 3325 -365 3355
rect -315 3325 -285 3355
rect -235 3325 -205 3355
rect -155 3325 -125 3355
rect -75 3325 -45 3355
rect 5 3325 35 3355
rect 85 3325 115 3355
rect 165 3325 195 3355
rect 245 3325 275 3355
rect 325 3325 355 3355
rect 405 3325 435 3355
rect 485 3325 515 3355
rect 565 3325 595 3355
rect 645 3325 675 3355
rect 725 3325 755 3355
rect 805 3325 835 3355
rect 885 3325 915 3355
rect 965 3325 995 3355
rect 1045 3325 1075 3355
rect 1125 3325 1155 3355
rect 1205 3325 1235 3355
rect 1285 3325 1315 3355
rect 1365 3325 1395 3355
rect 1445 3325 1475 3355
rect 1525 3325 1555 3355
rect 1605 3325 1635 3355
rect 1685 3325 1715 3355
rect 1765 3325 1795 3355
rect 1845 3325 1875 3355
rect 1925 3325 1955 3355
rect 2005 3325 2035 3355
rect 2085 3325 2115 3355
rect 2165 3325 2195 3355
rect 2245 3325 2275 3355
rect 2325 3325 2355 3355
rect 2405 3325 2435 3355
rect 2485 3325 2515 3355
rect 2565 3325 2595 3355
rect 2645 3325 2675 3355
rect 2725 3325 2755 3355
rect 2805 3325 2835 3355
rect 2885 3325 2915 3355
rect 2965 3325 2995 3355
rect 3045 3325 3075 3355
rect 3125 3325 3155 3355
rect 3205 3325 3235 3355
rect 3285 3325 3315 3355
rect 3365 3325 3395 3355
rect 3445 3325 3475 3355
rect 3525 3325 3555 3355
rect 3605 3325 3635 3355
rect 3685 3325 3715 3355
rect 3765 3325 3795 3355
rect 3845 3325 3875 3355
rect 3925 3325 3955 3355
rect 4005 3325 4035 3355
rect 4085 3325 4115 3355
rect 4165 3325 4195 3355
rect 4245 3325 4275 3355
rect 4325 3325 4355 3355
rect 4405 3325 4435 3355
rect 4485 3325 4515 3355
rect 4565 3325 4595 3355
rect 4645 3325 4675 3355
rect 4725 3325 4755 3355
rect 4805 3325 4835 3355
rect 4885 3325 4915 3355
rect 5045 3325 5075 3355
rect 5205 3325 5235 3355
rect 5365 3325 5395 3355
rect 5525 3325 5555 3355
rect 5685 3325 5715 3355
rect -1515 3245 -1485 3275
rect -1355 3245 -1325 3275
rect -1195 3245 -1165 3275
rect -1035 3245 -1005 3275
rect -875 3245 -845 3275
rect -795 3245 -765 3275
rect -715 3245 -685 3275
rect -635 3245 -605 3275
rect -555 3245 -525 3275
rect -475 3245 -445 3275
rect -395 3245 -365 3275
rect -315 3245 -285 3275
rect -235 3245 -205 3275
rect -155 3245 -125 3275
rect -75 3245 -45 3275
rect 5 3245 35 3275
rect 85 3245 115 3275
rect 165 3245 195 3275
rect 245 3245 275 3275
rect 325 3245 355 3275
rect 405 3245 435 3275
rect 485 3245 515 3275
rect 565 3245 595 3275
rect 645 3245 675 3275
rect 725 3245 755 3275
rect 805 3245 835 3275
rect 885 3245 915 3275
rect 965 3245 995 3275
rect 1045 3245 1075 3275
rect 1125 3245 1155 3275
rect 1205 3245 1235 3275
rect 1285 3245 1315 3275
rect 1365 3245 1395 3275
rect 1445 3245 1475 3275
rect 1525 3245 1555 3275
rect 1605 3245 1635 3275
rect 1685 3245 1715 3275
rect 1765 3245 1795 3275
rect 1845 3245 1875 3275
rect 1925 3245 1955 3275
rect 2005 3245 2035 3275
rect 2085 3245 2115 3275
rect 2165 3245 2195 3275
rect 2245 3245 2275 3275
rect 2325 3245 2355 3275
rect 2405 3245 2435 3275
rect 2485 3245 2515 3275
rect 2565 3245 2595 3275
rect 2645 3245 2675 3275
rect 2725 3245 2755 3275
rect 2805 3245 2835 3275
rect 2885 3245 2915 3275
rect 2965 3245 2995 3275
rect 3045 3245 3075 3275
rect 3125 3245 3155 3275
rect 3205 3245 3235 3275
rect 3285 3245 3315 3275
rect 3365 3245 3395 3275
rect 3445 3245 3475 3275
rect 3525 3245 3555 3275
rect 3605 3245 3635 3275
rect 3685 3245 3715 3275
rect 3765 3245 3795 3275
rect 3845 3245 3875 3275
rect 3925 3245 3955 3275
rect 4005 3245 4035 3275
rect 4085 3245 4115 3275
rect 4165 3245 4195 3275
rect 4245 3245 4275 3275
rect 4325 3245 4355 3275
rect 4405 3245 4435 3275
rect 4485 3245 4515 3275
rect 4565 3245 4595 3275
rect 4645 3245 4675 3275
rect 4725 3245 4755 3275
rect 4805 3245 4835 3275
rect 4885 3245 4915 3275
rect 5045 3245 5075 3275
rect 5205 3245 5235 3275
rect 5365 3245 5395 3275
rect 5525 3245 5555 3275
rect 5685 3245 5715 3275
rect -1515 3165 -1485 3195
rect -1355 3165 -1325 3195
rect -1195 3165 -1165 3195
rect -1035 3165 -1005 3195
rect -875 3165 -845 3195
rect -795 3165 -765 3195
rect -715 3165 -685 3195
rect -635 3165 -605 3195
rect -555 3165 -525 3195
rect -475 3165 -445 3195
rect -395 3165 -365 3195
rect -315 3165 -285 3195
rect -235 3165 -205 3195
rect -155 3165 -125 3195
rect -75 3165 -45 3195
rect 5 3165 35 3195
rect 85 3165 115 3195
rect 165 3165 195 3195
rect 245 3165 275 3195
rect 325 3165 355 3195
rect 405 3165 435 3195
rect 485 3165 515 3195
rect 565 3165 595 3195
rect 645 3165 675 3195
rect 725 3165 755 3195
rect 805 3165 835 3195
rect 885 3165 915 3195
rect 965 3165 995 3195
rect 1045 3165 1075 3195
rect 1125 3165 1155 3195
rect 1205 3165 1235 3195
rect 1285 3165 1315 3195
rect 1365 3165 1395 3195
rect 1445 3165 1475 3195
rect 1525 3165 1555 3195
rect 1605 3165 1635 3195
rect 1685 3165 1715 3195
rect 1765 3165 1795 3195
rect 1845 3165 1875 3195
rect 1925 3165 1955 3195
rect 2005 3165 2035 3195
rect 2085 3165 2115 3195
rect 2165 3165 2195 3195
rect 2245 3165 2275 3195
rect 2325 3165 2355 3195
rect 2405 3165 2435 3195
rect 2485 3165 2515 3195
rect 2565 3165 2595 3195
rect 2645 3165 2675 3195
rect 2725 3165 2755 3195
rect 2805 3165 2835 3195
rect 2885 3165 2915 3195
rect 2965 3165 2995 3195
rect 3045 3165 3075 3195
rect 3125 3165 3155 3195
rect 3205 3165 3235 3195
rect 3285 3165 3315 3195
rect 3365 3165 3395 3195
rect 3445 3165 3475 3195
rect 3525 3165 3555 3195
rect 3605 3165 3635 3195
rect 3685 3165 3715 3195
rect 3765 3165 3795 3195
rect 3845 3165 3875 3195
rect 3925 3165 3955 3195
rect 4005 3165 4035 3195
rect 4085 3165 4115 3195
rect 4165 3165 4195 3195
rect 4245 3165 4275 3195
rect 4325 3165 4355 3195
rect 4405 3165 4435 3195
rect 4485 3165 4515 3195
rect 4565 3165 4595 3195
rect 4645 3165 4675 3195
rect 4725 3165 4755 3195
rect 4805 3165 4835 3195
rect 4885 3165 4915 3195
rect 5045 3165 5075 3195
rect 5205 3165 5235 3195
rect 5365 3165 5395 3195
rect 5525 3165 5555 3195
rect 5685 3165 5715 3195
rect -1515 3085 -1485 3115
rect -1355 3085 -1325 3115
rect -1195 3085 -1165 3115
rect -1035 3085 -1005 3115
rect -875 3085 -845 3115
rect -795 3085 -765 3115
rect -715 3085 -685 3115
rect -635 3085 -605 3115
rect -555 3085 -525 3115
rect -475 3085 -445 3115
rect -395 3085 -365 3115
rect -315 3085 -285 3115
rect -235 3085 -205 3115
rect -155 3085 -125 3115
rect -75 3085 -45 3115
rect 5 3085 35 3115
rect 85 3085 115 3115
rect 165 3085 195 3115
rect 245 3085 275 3115
rect 325 3085 355 3115
rect 405 3085 435 3115
rect 485 3085 515 3115
rect 565 3085 595 3115
rect 645 3085 675 3115
rect 725 3085 755 3115
rect 805 3085 835 3115
rect 885 3085 915 3115
rect 965 3085 995 3115
rect 1045 3085 1075 3115
rect 1125 3085 1155 3115
rect 1205 3085 1235 3115
rect 1285 3085 1315 3115
rect 1365 3085 1395 3115
rect 1445 3085 1475 3115
rect 1525 3085 1555 3115
rect 1605 3085 1635 3115
rect 1685 3085 1715 3115
rect 1765 3085 1795 3115
rect 1845 3085 1875 3115
rect 1925 3085 1955 3115
rect 2005 3085 2035 3115
rect 2085 3085 2115 3115
rect 2165 3085 2195 3115
rect 2245 3085 2275 3115
rect 2325 3085 2355 3115
rect 2405 3085 2435 3115
rect 2485 3085 2515 3115
rect 2565 3085 2595 3115
rect 2645 3085 2675 3115
rect 2725 3085 2755 3115
rect 2805 3085 2835 3115
rect 2885 3085 2915 3115
rect 2965 3085 2995 3115
rect 3045 3085 3075 3115
rect 3125 3085 3155 3115
rect 3205 3085 3235 3115
rect 3285 3085 3315 3115
rect 3365 3085 3395 3115
rect 3445 3085 3475 3115
rect 3525 3085 3555 3115
rect 3605 3085 3635 3115
rect 3685 3085 3715 3115
rect 3765 3085 3795 3115
rect 3845 3085 3875 3115
rect 3925 3085 3955 3115
rect 4005 3085 4035 3115
rect 4085 3085 4115 3115
rect 4165 3085 4195 3115
rect 4245 3085 4275 3115
rect 4325 3085 4355 3115
rect 4405 3085 4435 3115
rect 4485 3085 4515 3115
rect 4565 3085 4595 3115
rect 4645 3085 4675 3115
rect 4725 3085 4755 3115
rect 4805 3085 4835 3115
rect 4885 3085 4915 3115
rect 5045 3085 5075 3115
rect 5205 3085 5235 3115
rect 5365 3085 5395 3115
rect 5525 3085 5555 3115
rect 5685 3085 5715 3115
rect -1515 3005 -1485 3035
rect -1355 3005 -1325 3035
rect -1195 3005 -1165 3035
rect -1115 3005 -1085 3035
rect 4885 3005 4915 3035
rect 5045 3005 5075 3035
rect 5205 3005 5235 3035
rect 5365 3005 5395 3035
rect 5525 3005 5555 3035
rect 5685 3005 5715 3035
rect -1515 2925 -1485 2955
rect -1355 2925 -1325 2955
rect -1195 2925 -1165 2955
rect -1035 2925 -1005 2955
rect -875 2925 -845 2955
rect -795 2925 -765 2955
rect -715 2925 -685 2955
rect -635 2925 -605 2955
rect -555 2925 -525 2955
rect -475 2925 -445 2955
rect -395 2925 -365 2955
rect -315 2925 -285 2955
rect -235 2925 -205 2955
rect -155 2925 -125 2955
rect -75 2925 -45 2955
rect 5 2925 35 2955
rect 85 2925 115 2955
rect 165 2925 195 2955
rect 245 2925 275 2955
rect 325 2925 355 2955
rect 405 2925 435 2955
rect 485 2925 515 2955
rect 565 2925 595 2955
rect 645 2925 675 2955
rect 725 2925 755 2955
rect 805 2925 835 2955
rect 885 2925 915 2955
rect 965 2925 995 2955
rect 1045 2925 1075 2955
rect 1125 2925 1155 2955
rect 1205 2925 1235 2955
rect 1285 2925 1315 2955
rect 1365 2925 1395 2955
rect 1445 2925 1475 2955
rect 1525 2925 1555 2955
rect 1605 2925 1635 2955
rect 1685 2925 1715 2955
rect 1765 2925 1795 2955
rect 1845 2925 1875 2955
rect 1925 2925 1955 2955
rect 2005 2925 2035 2955
rect 2085 2925 2115 2955
rect 2165 2925 2195 2955
rect 2245 2925 2275 2955
rect 2325 2925 2355 2955
rect 2405 2925 2435 2955
rect 2485 2925 2515 2955
rect 2565 2925 2595 2955
rect 2645 2925 2675 2955
rect 2725 2925 2755 2955
rect 2805 2925 2835 2955
rect 2885 2925 2915 2955
rect 2965 2925 2995 2955
rect 3045 2925 3075 2955
rect 3125 2925 3155 2955
rect 3205 2925 3235 2955
rect 3285 2925 3315 2955
rect 3365 2925 3395 2955
rect 3445 2925 3475 2955
rect 3525 2925 3555 2955
rect 3605 2925 3635 2955
rect 3685 2925 3715 2955
rect 3765 2925 3795 2955
rect 3845 2925 3875 2955
rect 3925 2925 3955 2955
rect 4005 2925 4035 2955
rect 4085 2925 4115 2955
rect 4165 2925 4195 2955
rect 4245 2925 4275 2955
rect 4325 2925 4355 2955
rect 4405 2925 4435 2955
rect 4485 2925 4515 2955
rect 4565 2925 4595 2955
rect 4645 2925 4675 2955
rect 4725 2925 4755 2955
rect 4805 2925 4835 2955
rect 4885 2925 4915 2955
rect 5045 2925 5075 2955
rect 5205 2925 5235 2955
rect 5365 2925 5395 2955
rect 5525 2925 5555 2955
rect 5685 2925 5715 2955
rect -1515 2845 -1485 2875
rect -1355 2845 -1325 2875
rect -1195 2845 -1165 2875
rect -1035 2845 -1005 2875
rect -955 2845 -925 2875
rect 4885 2845 4915 2875
rect 5045 2845 5075 2875
rect 5205 2845 5235 2875
rect 5365 2845 5395 2875
rect 5525 2845 5555 2875
rect 5685 2845 5715 2875
rect -1515 2765 -1485 2795
rect -1355 2765 -1325 2795
rect -1195 2765 -1165 2795
rect -1035 2765 -1005 2795
rect -875 2765 -845 2795
rect -795 2765 -765 2795
rect -715 2765 -685 2795
rect -635 2765 -605 2795
rect -555 2765 -525 2795
rect -475 2765 -445 2795
rect -395 2765 -365 2795
rect -315 2765 -285 2795
rect -235 2765 -205 2795
rect -155 2765 -125 2795
rect -75 2765 -45 2795
rect 5 2765 35 2795
rect 85 2765 115 2795
rect 165 2765 195 2795
rect 245 2765 275 2795
rect 325 2765 355 2795
rect 405 2765 435 2795
rect 485 2765 515 2795
rect 565 2765 595 2795
rect 645 2765 675 2795
rect 725 2765 755 2795
rect 805 2765 835 2795
rect 885 2765 915 2795
rect 965 2765 995 2795
rect 1045 2765 1075 2795
rect 1125 2765 1155 2795
rect 1205 2765 1235 2795
rect 1285 2765 1315 2795
rect 1365 2765 1395 2795
rect 1445 2765 1475 2795
rect 1525 2765 1555 2795
rect 1605 2765 1635 2795
rect 1685 2765 1715 2795
rect 1765 2765 1795 2795
rect 1845 2765 1875 2795
rect 1925 2765 1955 2795
rect 2005 2765 2035 2795
rect 2085 2765 2115 2795
rect 2165 2765 2195 2795
rect 2245 2765 2275 2795
rect 2325 2765 2355 2795
rect 2405 2765 2435 2795
rect 2485 2765 2515 2795
rect 2565 2765 2595 2795
rect 2645 2765 2675 2795
rect 2725 2765 2755 2795
rect 2805 2765 2835 2795
rect 2885 2765 2915 2795
rect 2965 2765 2995 2795
rect 3045 2765 3075 2795
rect 3125 2765 3155 2795
rect 3205 2765 3235 2795
rect 3285 2765 3315 2795
rect 3365 2765 3395 2795
rect 3445 2765 3475 2795
rect 3525 2765 3555 2795
rect 3605 2765 3635 2795
rect 3685 2765 3715 2795
rect 3765 2765 3795 2795
rect 3845 2765 3875 2795
rect 3925 2765 3955 2795
rect 4005 2765 4035 2795
rect 4085 2765 4115 2795
rect 4165 2765 4195 2795
rect 4245 2765 4275 2795
rect 4325 2765 4355 2795
rect 4405 2765 4435 2795
rect 4485 2765 4515 2795
rect 4565 2765 4595 2795
rect 4645 2765 4675 2795
rect 4725 2765 4755 2795
rect 4805 2765 4835 2795
rect 4885 2765 4915 2795
rect 5045 2765 5075 2795
rect 5205 2765 5235 2795
rect 5365 2765 5395 2795
rect 5525 2765 5555 2795
rect 5685 2765 5715 2795
rect -1515 2685 -1485 2715
rect -1355 2685 -1325 2715
rect -1195 2685 -1165 2715
rect -1035 2685 -1005 2715
rect -875 2685 -845 2715
rect -795 2685 -765 2715
rect -715 2685 -685 2715
rect -635 2685 -605 2715
rect -555 2685 -525 2715
rect -475 2685 -445 2715
rect -395 2685 -365 2715
rect -315 2685 -285 2715
rect -235 2685 -205 2715
rect -155 2685 -125 2715
rect -75 2685 -45 2715
rect 5 2685 35 2715
rect 85 2685 115 2715
rect 165 2685 195 2715
rect 245 2685 275 2715
rect 325 2685 355 2715
rect 405 2685 435 2715
rect 485 2685 515 2715
rect 565 2685 595 2715
rect 645 2685 675 2715
rect 725 2685 755 2715
rect 805 2685 835 2715
rect 885 2685 915 2715
rect 965 2685 995 2715
rect 1045 2685 1075 2715
rect 1125 2685 1155 2715
rect 1205 2685 1235 2715
rect 1285 2685 1315 2715
rect 1365 2685 1395 2715
rect 1445 2685 1475 2715
rect 1525 2685 1555 2715
rect 1605 2685 1635 2715
rect 1685 2685 1715 2715
rect 1765 2685 1795 2715
rect 1845 2685 1875 2715
rect 1925 2685 1955 2715
rect 2005 2685 2035 2715
rect 2085 2685 2115 2715
rect 2165 2685 2195 2715
rect 2245 2685 2275 2715
rect 2325 2685 2355 2715
rect 2405 2685 2435 2715
rect 2485 2685 2515 2715
rect 2565 2685 2595 2715
rect 2645 2685 2675 2715
rect 2725 2685 2755 2715
rect 2805 2685 2835 2715
rect 2885 2685 2915 2715
rect 2965 2685 2995 2715
rect 3045 2685 3075 2715
rect 3125 2685 3155 2715
rect 3205 2685 3235 2715
rect 3285 2685 3315 2715
rect 3365 2685 3395 2715
rect 3445 2685 3475 2715
rect 3525 2685 3555 2715
rect 3605 2685 3635 2715
rect 3685 2685 3715 2715
rect 3765 2685 3795 2715
rect 3845 2685 3875 2715
rect 3925 2685 3955 2715
rect 4005 2685 4035 2715
rect 4085 2685 4115 2715
rect 4165 2685 4195 2715
rect 4245 2685 4275 2715
rect 4325 2685 4355 2715
rect 4405 2685 4435 2715
rect 4485 2685 4515 2715
rect 4565 2685 4595 2715
rect 4645 2685 4675 2715
rect 4725 2685 4755 2715
rect 4805 2685 4835 2715
rect 4885 2685 4915 2715
rect 5045 2685 5075 2715
rect 5205 2685 5235 2715
rect 5365 2685 5395 2715
rect 5525 2685 5555 2715
rect 5685 2685 5715 2715
rect -1515 2605 -1485 2635
rect -1355 2605 -1325 2635
rect -1275 2605 -1245 2635
rect 4885 2605 4915 2635
rect 5045 2605 5075 2635
rect 5205 2605 5235 2635
rect 5365 2605 5395 2635
rect 5525 2605 5555 2635
rect 5685 2605 5715 2635
rect -1515 2525 -1485 2555
rect -1355 2525 -1325 2555
rect -1195 2525 -1165 2555
rect -1035 2525 -1005 2555
rect -875 2525 -845 2555
rect -795 2525 -765 2555
rect -715 2525 -685 2555
rect -635 2525 -605 2555
rect -555 2525 -525 2555
rect -475 2525 -445 2555
rect -395 2525 -365 2555
rect -315 2525 -285 2555
rect -235 2525 -205 2555
rect -155 2525 -125 2555
rect -75 2525 -45 2555
rect 5 2525 35 2555
rect 85 2525 115 2555
rect 165 2525 195 2555
rect 245 2525 275 2555
rect 325 2525 355 2555
rect 405 2525 435 2555
rect 485 2525 515 2555
rect 565 2525 595 2555
rect 645 2525 675 2555
rect 725 2525 755 2555
rect 805 2525 835 2555
rect 885 2525 915 2555
rect 965 2525 995 2555
rect 1045 2525 1075 2555
rect 1125 2525 1155 2555
rect 1205 2525 1235 2555
rect 1285 2525 1315 2555
rect 1365 2525 1395 2555
rect 1445 2525 1475 2555
rect 1525 2525 1555 2555
rect 1605 2525 1635 2555
rect 1685 2525 1715 2555
rect 1765 2525 1795 2555
rect 1845 2525 1875 2555
rect 1925 2525 1955 2555
rect 2005 2525 2035 2555
rect 2085 2525 2115 2555
rect 2165 2525 2195 2555
rect 2245 2525 2275 2555
rect 2325 2525 2355 2555
rect 2405 2525 2435 2555
rect 2485 2525 2515 2555
rect 2565 2525 2595 2555
rect 2645 2525 2675 2555
rect 2725 2525 2755 2555
rect 2805 2525 2835 2555
rect 2885 2525 2915 2555
rect 2965 2525 2995 2555
rect 3045 2525 3075 2555
rect 3125 2525 3155 2555
rect 3205 2525 3235 2555
rect 3285 2525 3315 2555
rect 3365 2525 3395 2555
rect 3445 2525 3475 2555
rect 3525 2525 3555 2555
rect 3605 2525 3635 2555
rect 3685 2525 3715 2555
rect 3765 2525 3795 2555
rect 3845 2525 3875 2555
rect 3925 2525 3955 2555
rect 4005 2525 4035 2555
rect 4085 2525 4115 2555
rect 4165 2525 4195 2555
rect 4245 2525 4275 2555
rect 4325 2525 4355 2555
rect 4405 2525 4435 2555
rect 4485 2525 4515 2555
rect 4565 2525 4595 2555
rect 4645 2525 4675 2555
rect 4725 2525 4755 2555
rect 4805 2525 4835 2555
rect 4885 2525 4915 2555
rect 5045 2525 5075 2555
rect 5205 2525 5235 2555
rect 5365 2525 5395 2555
rect 5525 2525 5555 2555
rect 5685 2525 5715 2555
rect -1515 2445 -1485 2475
rect -1355 2445 -1325 2475
rect -1195 2445 -1165 2475
rect -1035 2445 -1005 2475
rect -875 2445 -845 2475
rect -795 2445 -765 2475
rect -715 2445 -685 2475
rect -635 2445 -605 2475
rect -555 2445 -525 2475
rect -475 2445 -445 2475
rect -395 2445 -365 2475
rect -315 2445 -285 2475
rect -235 2445 -205 2475
rect -155 2445 -125 2475
rect -75 2445 -45 2475
rect 5 2445 35 2475
rect 85 2445 115 2475
rect 165 2445 195 2475
rect 245 2445 275 2475
rect 325 2445 355 2475
rect 405 2445 435 2475
rect 485 2445 515 2475
rect 565 2445 595 2475
rect 645 2445 675 2475
rect 725 2445 755 2475
rect 805 2445 835 2475
rect 885 2445 915 2475
rect 965 2445 995 2475
rect 1045 2445 1075 2475
rect 1125 2445 1155 2475
rect 1205 2445 1235 2475
rect 1285 2445 1315 2475
rect 1365 2445 1395 2475
rect 1445 2445 1475 2475
rect 1525 2445 1555 2475
rect 1605 2445 1635 2475
rect 1685 2445 1715 2475
rect 1765 2445 1795 2475
rect 1845 2445 1875 2475
rect 1925 2445 1955 2475
rect 2005 2445 2035 2475
rect 2085 2445 2115 2475
rect 2165 2445 2195 2475
rect 2245 2445 2275 2475
rect 2325 2445 2355 2475
rect 2405 2445 2435 2475
rect 2485 2445 2515 2475
rect 2565 2445 2595 2475
rect 2645 2445 2675 2475
rect 2725 2445 2755 2475
rect 2805 2445 2835 2475
rect 2885 2445 2915 2475
rect 2965 2445 2995 2475
rect 3045 2445 3075 2475
rect 3125 2445 3155 2475
rect 3205 2445 3235 2475
rect 3285 2445 3315 2475
rect 3365 2445 3395 2475
rect 3445 2445 3475 2475
rect 3525 2445 3555 2475
rect 3605 2445 3635 2475
rect 3685 2445 3715 2475
rect 3765 2445 3795 2475
rect 3845 2445 3875 2475
rect 3925 2445 3955 2475
rect 4005 2445 4035 2475
rect 4085 2445 4115 2475
rect 4165 2445 4195 2475
rect 4245 2445 4275 2475
rect 4325 2445 4355 2475
rect 4405 2445 4435 2475
rect 4485 2445 4515 2475
rect 4565 2445 4595 2475
rect 4645 2445 4675 2475
rect 4725 2445 4755 2475
rect 4805 2445 4835 2475
rect 4885 2445 4915 2475
rect 5045 2445 5075 2475
rect 5205 2445 5235 2475
rect 5365 2445 5395 2475
rect 5525 2445 5555 2475
rect 5685 2445 5715 2475
rect -1515 2365 -1485 2395
rect -1355 2365 -1325 2395
rect -1195 2365 -1165 2395
rect -1035 2365 -1005 2395
rect -875 2365 -845 2395
rect 5285 2365 5315 2395
rect -1515 2285 -1485 2315
rect -1355 2285 -1325 2315
rect -1195 2285 -1165 2315
rect -1035 2285 -1005 2315
rect -875 2285 -845 2315
rect -795 2285 -765 2315
rect -715 2285 -685 2315
rect -635 2285 -605 2315
rect -555 2285 -525 2315
rect -475 2285 -445 2315
rect -395 2285 -365 2315
rect -315 2285 -285 2315
rect -235 2285 -205 2315
rect -155 2285 -125 2315
rect -75 2285 -45 2315
rect 5 2285 35 2315
rect 85 2285 115 2315
rect 165 2285 195 2315
rect 245 2285 275 2315
rect 325 2285 355 2315
rect 405 2285 435 2315
rect 485 2285 515 2315
rect 565 2285 595 2315
rect 645 2285 675 2315
rect 725 2285 755 2315
rect 805 2285 835 2315
rect 885 2285 915 2315
rect 965 2285 995 2315
rect 1045 2285 1075 2315
rect 1125 2285 1155 2315
rect 1205 2285 1235 2315
rect 1285 2285 1315 2315
rect 1365 2285 1395 2315
rect 1445 2285 1475 2315
rect 1525 2285 1555 2315
rect 1605 2285 1635 2315
rect 1685 2285 1715 2315
rect 1765 2285 1795 2315
rect 1845 2285 1875 2315
rect 1925 2285 1955 2315
rect 2005 2285 2035 2315
rect 2085 2285 2115 2315
rect 2165 2285 2195 2315
rect 2245 2285 2275 2315
rect 2325 2285 2355 2315
rect 2405 2285 2435 2315
rect 2485 2285 2515 2315
rect 2565 2285 2595 2315
rect 2645 2285 2675 2315
rect 2725 2285 2755 2315
rect 2805 2285 2835 2315
rect 2885 2285 2915 2315
rect 2965 2285 2995 2315
rect 3045 2285 3075 2315
rect 3125 2285 3155 2315
rect 3205 2285 3235 2315
rect 3285 2285 3315 2315
rect 3365 2285 3395 2315
rect 3445 2285 3475 2315
rect 3525 2285 3555 2315
rect 3605 2285 3635 2315
rect 3685 2285 3715 2315
rect 3765 2285 3795 2315
rect 3845 2285 3875 2315
rect 3925 2285 3955 2315
rect 4005 2285 4035 2315
rect 4085 2285 4115 2315
rect 4165 2285 4195 2315
rect 4245 2285 4275 2315
rect 4325 2285 4355 2315
rect 4405 2285 4435 2315
rect 4485 2285 4515 2315
rect 4565 2285 4595 2315
rect 4645 2285 4675 2315
rect 4725 2285 4755 2315
rect 4805 2285 4835 2315
rect 4885 2285 4915 2315
rect 5045 2285 5075 2315
rect 5205 2285 5235 2315
rect 5365 2285 5395 2315
rect 5525 2285 5555 2315
rect 5685 2285 5715 2315
rect -1515 2205 -1485 2235
rect -1355 2205 -1325 2235
rect -1195 2205 -1165 2235
rect -1035 2205 -1005 2235
rect -875 2205 -845 2235
rect 4965 2205 4995 2235
rect 5045 2205 5075 2235
rect 5205 2205 5235 2235
rect 5365 2205 5395 2235
rect 5525 2205 5555 2235
rect 5685 2205 5715 2235
rect -1515 2125 -1485 2155
rect -1355 2125 -1325 2155
rect -1195 2125 -1165 2155
rect -1035 2125 -1005 2155
rect -875 2125 -845 2155
rect -795 2125 -765 2155
rect -715 2125 -685 2155
rect -635 2125 -605 2155
rect -555 2125 -525 2155
rect -475 2125 -445 2155
rect -395 2125 -365 2155
rect -315 2125 -285 2155
rect -235 2125 -205 2155
rect -155 2125 -125 2155
rect -75 2125 -45 2155
rect 5 2125 35 2155
rect 85 2125 115 2155
rect 165 2125 195 2155
rect 245 2125 275 2155
rect 325 2125 355 2155
rect 405 2125 435 2155
rect 485 2125 515 2155
rect 565 2125 595 2155
rect 645 2125 675 2155
rect 725 2125 755 2155
rect 805 2125 835 2155
rect 885 2125 915 2155
rect 965 2125 995 2155
rect 1045 2125 1075 2155
rect 1125 2125 1155 2155
rect 1205 2125 1235 2155
rect 1285 2125 1315 2155
rect 1365 2125 1395 2155
rect 1445 2125 1475 2155
rect 1525 2125 1555 2155
rect 1605 2125 1635 2155
rect 1685 2125 1715 2155
rect 1765 2125 1795 2155
rect 1845 2125 1875 2155
rect 1925 2125 1955 2155
rect 2005 2125 2035 2155
rect 2085 2125 2115 2155
rect 2165 2125 2195 2155
rect 2245 2125 2275 2155
rect 2325 2125 2355 2155
rect 2405 2125 2435 2155
rect 2485 2125 2515 2155
rect 2565 2125 2595 2155
rect 2645 2125 2675 2155
rect 2725 2125 2755 2155
rect 2805 2125 2835 2155
rect 2885 2125 2915 2155
rect 2965 2125 2995 2155
rect 3045 2125 3075 2155
rect 3125 2125 3155 2155
rect 3205 2125 3235 2155
rect 3285 2125 3315 2155
rect 3365 2125 3395 2155
rect 3445 2125 3475 2155
rect 3525 2125 3555 2155
rect 3605 2125 3635 2155
rect 3685 2125 3715 2155
rect 3765 2125 3795 2155
rect 3845 2125 3875 2155
rect 3925 2125 3955 2155
rect 4005 2125 4035 2155
rect 4085 2125 4115 2155
rect 4165 2125 4195 2155
rect 4245 2125 4275 2155
rect 4325 2125 4355 2155
rect 4405 2125 4435 2155
rect 4485 2125 4515 2155
rect 4565 2125 4595 2155
rect 4645 2125 4675 2155
rect 4725 2125 4755 2155
rect 4805 2125 4835 2155
rect 4885 2125 4915 2155
rect 5045 2125 5075 2155
rect 5205 2125 5235 2155
rect 5365 2125 5395 2155
rect 5525 2125 5555 2155
rect 5685 2125 5715 2155
rect -1515 2045 -1485 2075
rect -1355 2045 -1325 2075
rect -1195 2045 -1165 2075
rect -1035 2045 -1005 2075
rect -875 2045 -845 2075
rect -795 2045 -765 2075
rect -715 2045 -685 2075
rect -635 2045 -605 2075
rect -555 2045 -525 2075
rect -475 2045 -445 2075
rect -395 2045 -365 2075
rect -315 2045 -285 2075
rect -235 2045 -205 2075
rect -155 2045 -125 2075
rect -75 2045 -45 2075
rect 5 2045 35 2075
rect 85 2045 115 2075
rect 165 2045 195 2075
rect 245 2045 275 2075
rect 325 2045 355 2075
rect 405 2045 435 2075
rect 485 2045 515 2075
rect 565 2045 595 2075
rect 645 2045 675 2075
rect 725 2045 755 2075
rect 805 2045 835 2075
rect 885 2045 915 2075
rect 965 2045 995 2075
rect 1045 2045 1075 2075
rect 1125 2045 1155 2075
rect 1205 2045 1235 2075
rect 1285 2045 1315 2075
rect 1365 2045 1395 2075
rect 1445 2045 1475 2075
rect 1525 2045 1555 2075
rect 1605 2045 1635 2075
rect 1685 2045 1715 2075
rect 1765 2045 1795 2075
rect 1845 2045 1875 2075
rect 1925 2045 1955 2075
rect 2005 2045 2035 2075
rect 2085 2045 2115 2075
rect 2165 2045 2195 2075
rect 2245 2045 2275 2075
rect 2325 2045 2355 2075
rect 2405 2045 2435 2075
rect 2485 2045 2515 2075
rect 2565 2045 2595 2075
rect 2645 2045 2675 2075
rect 2725 2045 2755 2075
rect 2805 2045 2835 2075
rect 2885 2045 2915 2075
rect 2965 2045 2995 2075
rect 3045 2045 3075 2075
rect 3125 2045 3155 2075
rect 3205 2045 3235 2075
rect 3285 2045 3315 2075
rect 3365 2045 3395 2075
rect 3445 2045 3475 2075
rect 3525 2045 3555 2075
rect 3605 2045 3635 2075
rect 3685 2045 3715 2075
rect 3765 2045 3795 2075
rect 3845 2045 3875 2075
rect 3925 2045 3955 2075
rect 4005 2045 4035 2075
rect 4085 2045 4115 2075
rect 4165 2045 4195 2075
rect 4245 2045 4275 2075
rect 4325 2045 4355 2075
rect 4405 2045 4435 2075
rect 4485 2045 4515 2075
rect 4565 2045 4595 2075
rect 4645 2045 4675 2075
rect 4725 2045 4755 2075
rect 4805 2045 4835 2075
rect 4885 2045 4915 2075
rect 5045 2045 5075 2075
rect 5205 2045 5235 2075
rect 5365 2045 5395 2075
rect 5525 2045 5555 2075
rect 5685 2045 5715 2075
rect -1515 1965 -1485 1995
rect -1355 1965 -1325 1995
rect -1195 1965 -1165 1995
rect -1035 1965 -1005 1995
rect -875 1965 -845 1995
rect -795 1965 -765 1995
rect -715 1965 -685 1995
rect -635 1965 -605 1995
rect -555 1965 -525 1995
rect -475 1965 -445 1995
rect -395 1965 -365 1995
rect -315 1965 -285 1995
rect -235 1965 -205 1995
rect -155 1965 -125 1995
rect -75 1965 -45 1995
rect 5 1965 35 1995
rect 85 1965 115 1995
rect 165 1965 195 1995
rect 245 1965 275 1995
rect 325 1965 355 1995
rect 405 1965 435 1995
rect 485 1965 515 1995
rect 565 1965 595 1995
rect 645 1965 675 1995
rect 725 1965 755 1995
rect 805 1965 835 1995
rect 885 1965 915 1995
rect 965 1965 995 1995
rect 1045 1965 1075 1995
rect 1125 1965 1155 1995
rect 1205 1965 1235 1995
rect 1285 1965 1315 1995
rect 1365 1965 1395 1995
rect 1445 1965 1475 1995
rect 1525 1965 1555 1995
rect 1605 1965 1635 1995
rect 1685 1965 1715 1995
rect 1765 1965 1795 1995
rect 1845 1965 1875 1995
rect 1925 1965 1955 1995
rect 2005 1965 2035 1995
rect 2085 1965 2115 1995
rect 2165 1965 2195 1995
rect 2245 1965 2275 1995
rect 2325 1965 2355 1995
rect 2405 1965 2435 1995
rect 2485 1965 2515 1995
rect 2565 1965 2595 1995
rect 2645 1965 2675 1995
rect 2725 1965 2755 1995
rect 2805 1965 2835 1995
rect 2885 1965 2915 1995
rect 2965 1965 2995 1995
rect 3045 1965 3075 1995
rect 3125 1965 3155 1995
rect 3205 1965 3235 1995
rect 3285 1965 3315 1995
rect 3365 1965 3395 1995
rect 3445 1965 3475 1995
rect 3525 1965 3555 1995
rect 3605 1965 3635 1995
rect 3685 1965 3715 1995
rect 3765 1965 3795 1995
rect 3845 1965 3875 1995
rect 3925 1965 3955 1995
rect 4005 1965 4035 1995
rect 4085 1965 4115 1995
rect 4165 1965 4195 1995
rect 4245 1965 4275 1995
rect 4325 1965 4355 1995
rect 4405 1965 4435 1995
rect 4485 1965 4515 1995
rect 4565 1965 4595 1995
rect 4645 1965 4675 1995
rect 4725 1965 4755 1995
rect 4805 1965 4835 1995
rect 4885 1965 4915 1995
rect 5045 1965 5075 1995
rect 5205 1965 5235 1995
rect 5365 1965 5395 1995
rect 5525 1965 5555 1995
rect 5685 1965 5715 1995
rect -1515 1885 -1485 1915
rect -1355 1885 -1325 1915
rect -1195 1885 -1165 1915
rect -1035 1885 -1005 1915
rect -875 1885 -845 1915
rect -795 1885 -765 1915
rect -715 1885 -685 1915
rect -635 1885 -605 1915
rect -555 1885 -525 1915
rect -475 1885 -445 1915
rect -395 1885 -365 1915
rect -315 1885 -285 1915
rect -235 1885 -205 1915
rect -155 1885 -125 1915
rect -75 1885 -45 1915
rect 5 1885 35 1915
rect 85 1885 115 1915
rect 165 1885 195 1915
rect 245 1885 275 1915
rect 325 1885 355 1915
rect 405 1885 435 1915
rect 485 1885 515 1915
rect 565 1885 595 1915
rect 645 1885 675 1915
rect 725 1885 755 1915
rect 805 1885 835 1915
rect 885 1885 915 1915
rect 965 1885 995 1915
rect 1045 1885 1075 1915
rect 1125 1885 1155 1915
rect 1205 1885 1235 1915
rect 1285 1885 1315 1915
rect 1365 1885 1395 1915
rect 1445 1885 1475 1915
rect 1525 1885 1555 1915
rect 1605 1885 1635 1915
rect 1685 1885 1715 1915
rect 1765 1885 1795 1915
rect 1845 1885 1875 1915
rect 1925 1885 1955 1915
rect 2005 1885 2035 1915
rect 2085 1885 2115 1915
rect 2165 1885 2195 1915
rect 2245 1885 2275 1915
rect 2325 1885 2355 1915
rect 2405 1885 2435 1915
rect 2485 1885 2515 1915
rect 2565 1885 2595 1915
rect 2645 1885 2675 1915
rect 2725 1885 2755 1915
rect 2805 1885 2835 1915
rect 2885 1885 2915 1915
rect 2965 1885 2995 1915
rect 3045 1885 3075 1915
rect 3125 1885 3155 1915
rect 3205 1885 3235 1915
rect 3285 1885 3315 1915
rect 3365 1885 3395 1915
rect 3445 1885 3475 1915
rect 3525 1885 3555 1915
rect 3605 1885 3635 1915
rect 3685 1885 3715 1915
rect 3765 1885 3795 1915
rect 3845 1885 3875 1915
rect 3925 1885 3955 1915
rect 4005 1885 4035 1915
rect 4085 1885 4115 1915
rect 4165 1885 4195 1915
rect 4245 1885 4275 1915
rect 4325 1885 4355 1915
rect 4405 1885 4435 1915
rect 4485 1885 4515 1915
rect 4565 1885 4595 1915
rect 4645 1885 4675 1915
rect 4725 1885 4755 1915
rect 4805 1885 4835 1915
rect 4885 1885 4915 1915
rect 5045 1885 5075 1915
rect 5205 1885 5235 1915
rect 5365 1885 5395 1915
rect 5525 1885 5555 1915
rect 5685 1885 5715 1915
rect -1515 1805 -1485 1835
rect -1355 1805 -1325 1835
rect -1195 1805 -1165 1835
rect -1035 1805 -1005 1835
rect -875 1805 -845 1835
rect -795 1805 -765 1835
rect -715 1805 -685 1835
rect -635 1805 -605 1835
rect -555 1805 -525 1835
rect -475 1805 -445 1835
rect -395 1805 -365 1835
rect -315 1805 -285 1835
rect -235 1805 -205 1835
rect -155 1805 -125 1835
rect -75 1805 -45 1835
rect 5 1805 35 1835
rect 85 1805 115 1835
rect 165 1805 195 1835
rect 245 1805 275 1835
rect 325 1805 355 1835
rect 405 1805 435 1835
rect 485 1805 515 1835
rect 565 1805 595 1835
rect 645 1805 675 1835
rect 725 1805 755 1835
rect 805 1805 835 1835
rect 885 1805 915 1835
rect 965 1805 995 1835
rect 1045 1805 1075 1835
rect 1125 1805 1155 1835
rect 1205 1805 1235 1835
rect 1285 1805 1315 1835
rect 1365 1805 1395 1835
rect 1445 1805 1475 1835
rect 1525 1805 1555 1835
rect 1605 1805 1635 1835
rect 1685 1805 1715 1835
rect 1765 1805 1795 1835
rect 1845 1805 1875 1835
rect 1925 1805 1955 1835
rect 2005 1805 2035 1835
rect 2085 1805 2115 1835
rect 2165 1805 2195 1835
rect 2245 1805 2275 1835
rect 2325 1805 2355 1835
rect 2405 1805 2435 1835
rect 2485 1805 2515 1835
rect 2565 1805 2595 1835
rect 2645 1805 2675 1835
rect 2725 1805 2755 1835
rect 2805 1805 2835 1835
rect 2885 1805 2915 1835
rect 2965 1805 2995 1835
rect 3045 1805 3075 1835
rect 3125 1805 3155 1835
rect 3205 1805 3235 1835
rect 3285 1805 3315 1835
rect 3365 1805 3395 1835
rect 3445 1805 3475 1835
rect 3525 1805 3555 1835
rect 3605 1805 3635 1835
rect 3685 1805 3715 1835
rect 3765 1805 3795 1835
rect 3845 1805 3875 1835
rect 3925 1805 3955 1835
rect 4005 1805 4035 1835
rect 4085 1805 4115 1835
rect 4165 1805 4195 1835
rect 4245 1805 4275 1835
rect 4325 1805 4355 1835
rect 4405 1805 4435 1835
rect 4485 1805 4515 1835
rect 4565 1805 4595 1835
rect 4645 1805 4675 1835
rect 4725 1805 4755 1835
rect 4805 1805 4835 1835
rect 4885 1805 4915 1835
rect 5045 1805 5075 1835
rect 5205 1805 5235 1835
rect 5365 1805 5395 1835
rect 5525 1805 5555 1835
rect 5685 1805 5715 1835
rect -1515 1725 -1485 1755
rect -1355 1725 -1325 1755
rect -1195 1725 -1165 1755
rect -1035 1725 -1005 1755
rect -875 1725 -845 1755
rect -795 1725 -765 1755
rect -715 1725 -685 1755
rect -635 1725 -605 1755
rect -555 1725 -525 1755
rect -475 1725 -445 1755
rect -395 1725 -365 1755
rect -315 1725 -285 1755
rect -235 1725 -205 1755
rect -155 1725 -125 1755
rect -75 1725 -45 1755
rect 5 1725 35 1755
rect 85 1725 115 1755
rect 165 1725 195 1755
rect 245 1725 275 1755
rect 325 1725 355 1755
rect 405 1725 435 1755
rect 485 1725 515 1755
rect 565 1725 595 1755
rect 645 1725 675 1755
rect 725 1725 755 1755
rect 805 1725 835 1755
rect 885 1725 915 1755
rect 965 1725 995 1755
rect 1045 1725 1075 1755
rect 1125 1725 1155 1755
rect 1205 1725 1235 1755
rect 1285 1725 1315 1755
rect 1365 1725 1395 1755
rect 1445 1725 1475 1755
rect 1525 1725 1555 1755
rect 1605 1725 1635 1755
rect 1685 1725 1715 1755
rect 1765 1725 1795 1755
rect 1845 1725 1875 1755
rect 1925 1725 1955 1755
rect 2005 1725 2035 1755
rect 2085 1725 2115 1755
rect 2165 1725 2195 1755
rect 2245 1725 2275 1755
rect 2325 1725 2355 1755
rect 2405 1725 2435 1755
rect 2485 1725 2515 1755
rect 2565 1725 2595 1755
rect 2645 1725 2675 1755
rect 2725 1725 2755 1755
rect 2805 1725 2835 1755
rect 2885 1725 2915 1755
rect 2965 1725 2995 1755
rect 3045 1725 3075 1755
rect 3125 1725 3155 1755
rect 3205 1725 3235 1755
rect 3285 1725 3315 1755
rect 3365 1725 3395 1755
rect 3445 1725 3475 1755
rect 3525 1725 3555 1755
rect 3605 1725 3635 1755
rect 3685 1725 3715 1755
rect 3765 1725 3795 1755
rect 3845 1725 3875 1755
rect 3925 1725 3955 1755
rect 4005 1725 4035 1755
rect 4085 1725 4115 1755
rect 4165 1725 4195 1755
rect 4245 1725 4275 1755
rect 4325 1725 4355 1755
rect 4405 1725 4435 1755
rect 4485 1725 4515 1755
rect 4565 1725 4595 1755
rect 4645 1725 4675 1755
rect 4725 1725 4755 1755
rect 4805 1725 4835 1755
rect 4885 1725 4915 1755
rect 5045 1725 5075 1755
rect 5205 1725 5235 1755
rect 5365 1725 5395 1755
rect 5525 1725 5555 1755
rect 5685 1725 5715 1755
rect -1515 1645 -1485 1675
rect -1355 1645 -1325 1675
rect -1195 1645 -1165 1675
rect -1035 1645 -1005 1675
rect -875 1645 -845 1675
rect -795 1645 -765 1675
rect -715 1645 -685 1675
rect -635 1645 -605 1675
rect -555 1645 -525 1675
rect -475 1645 -445 1675
rect -395 1645 -365 1675
rect -315 1645 -285 1675
rect -235 1645 -205 1675
rect -155 1645 -125 1675
rect -75 1645 -45 1675
rect 5 1645 35 1675
rect 85 1645 115 1675
rect 165 1645 195 1675
rect 245 1645 275 1675
rect 325 1645 355 1675
rect 405 1645 435 1675
rect 485 1645 515 1675
rect 565 1645 595 1675
rect 645 1645 675 1675
rect 725 1645 755 1675
rect 805 1645 835 1675
rect 885 1645 915 1675
rect 965 1645 995 1675
rect 1045 1645 1075 1675
rect 1125 1645 1155 1675
rect 1205 1645 1235 1675
rect 1285 1645 1315 1675
rect 1365 1645 1395 1675
rect 1445 1645 1475 1675
rect 1525 1645 1555 1675
rect 1605 1645 1635 1675
rect 1685 1645 1715 1675
rect 1765 1645 1795 1675
rect 1845 1645 1875 1675
rect 1925 1645 1955 1675
rect 2005 1645 2035 1675
rect 2085 1645 2115 1675
rect 2165 1645 2195 1675
rect 2245 1645 2275 1675
rect 2325 1645 2355 1675
rect 2405 1645 2435 1675
rect 2485 1645 2515 1675
rect 2565 1645 2595 1675
rect 2645 1645 2675 1675
rect 2725 1645 2755 1675
rect 2805 1645 2835 1675
rect 2885 1645 2915 1675
rect 2965 1645 2995 1675
rect 3045 1645 3075 1675
rect 3125 1645 3155 1675
rect 3205 1645 3235 1675
rect 3285 1645 3315 1675
rect 3365 1645 3395 1675
rect 3445 1645 3475 1675
rect 3525 1645 3555 1675
rect 3605 1645 3635 1675
rect 3685 1645 3715 1675
rect 3765 1645 3795 1675
rect 3845 1645 3875 1675
rect 3925 1645 3955 1675
rect 4005 1645 4035 1675
rect 4085 1645 4115 1675
rect 4165 1645 4195 1675
rect 4245 1645 4275 1675
rect 4325 1645 4355 1675
rect 4405 1645 4435 1675
rect 4485 1645 4515 1675
rect 4565 1645 4595 1675
rect 4645 1645 4675 1675
rect 4725 1645 4755 1675
rect 4805 1645 4835 1675
rect 4885 1645 4915 1675
rect 5045 1645 5075 1675
rect 5205 1645 5235 1675
rect 5365 1645 5395 1675
rect 5525 1645 5555 1675
rect 5685 1645 5715 1675
rect -1515 1565 -1485 1595
rect -1355 1565 -1325 1595
rect -1195 1565 -1165 1595
rect -1035 1565 -1005 1595
rect -875 1565 -845 1595
rect -795 1565 -765 1595
rect -715 1565 -685 1595
rect -635 1565 -605 1595
rect -555 1565 -525 1595
rect -475 1565 -445 1595
rect -395 1565 -365 1595
rect -315 1565 -285 1595
rect -235 1565 -205 1595
rect -155 1565 -125 1595
rect -75 1565 -45 1595
rect 5 1565 35 1595
rect 85 1565 115 1595
rect 165 1565 195 1595
rect 245 1565 275 1595
rect 325 1565 355 1595
rect 405 1565 435 1595
rect 485 1565 515 1595
rect 565 1565 595 1595
rect 645 1565 675 1595
rect 725 1565 755 1595
rect 805 1565 835 1595
rect 885 1565 915 1595
rect 965 1565 995 1595
rect 1045 1565 1075 1595
rect 1125 1565 1155 1595
rect 1205 1565 1235 1595
rect 1285 1565 1315 1595
rect 1365 1565 1395 1595
rect 1445 1565 1475 1595
rect 1525 1565 1555 1595
rect 1605 1565 1635 1595
rect 1685 1565 1715 1595
rect 1765 1565 1795 1595
rect 1845 1565 1875 1595
rect 1925 1565 1955 1595
rect 2005 1565 2035 1595
rect 2085 1565 2115 1595
rect 2165 1565 2195 1595
rect 2245 1565 2275 1595
rect 2325 1565 2355 1595
rect 2405 1565 2435 1595
rect 2485 1565 2515 1595
rect 2565 1565 2595 1595
rect 2645 1565 2675 1595
rect 2725 1565 2755 1595
rect 2805 1565 2835 1595
rect 2885 1565 2915 1595
rect 2965 1565 2995 1595
rect 3045 1565 3075 1595
rect 3125 1565 3155 1595
rect 3205 1565 3235 1595
rect 3285 1565 3315 1595
rect 3365 1565 3395 1595
rect 3445 1565 3475 1595
rect 3525 1565 3555 1595
rect 3605 1565 3635 1595
rect 3685 1565 3715 1595
rect 3765 1565 3795 1595
rect 3845 1565 3875 1595
rect 3925 1565 3955 1595
rect 4005 1565 4035 1595
rect 4085 1565 4115 1595
rect 4165 1565 4195 1595
rect 4245 1565 4275 1595
rect 4325 1565 4355 1595
rect 4405 1565 4435 1595
rect 4485 1565 4515 1595
rect 4565 1565 4595 1595
rect 4645 1565 4675 1595
rect 4725 1565 4755 1595
rect 4805 1565 4835 1595
rect 4885 1565 4915 1595
rect 5045 1565 5075 1595
rect 5205 1565 5235 1595
rect 5365 1565 5395 1595
rect 5525 1565 5555 1595
rect 5685 1565 5715 1595
rect -1515 1485 -1485 1515
rect -1355 1485 -1325 1515
rect -1195 1485 -1165 1515
rect -1035 1485 -1005 1515
rect -955 1485 -925 1515
rect 4885 1485 4915 1515
rect 5045 1485 5075 1515
rect 5205 1485 5235 1515
rect 5365 1485 5395 1515
rect 5525 1485 5555 1515
rect 5685 1485 5715 1515
rect -1515 1405 -1485 1435
rect -1355 1405 -1325 1435
rect -1195 1405 -1165 1435
rect -1035 1405 -1005 1435
rect -875 1405 -845 1435
rect -795 1405 -765 1435
rect -715 1405 -685 1435
rect -635 1405 -605 1435
rect -555 1405 -525 1435
rect -475 1405 -445 1435
rect -395 1405 -365 1435
rect -315 1405 -285 1435
rect -235 1405 -205 1435
rect -155 1405 -125 1435
rect -75 1405 -45 1435
rect 5 1405 35 1435
rect 85 1405 115 1435
rect 165 1405 195 1435
rect 245 1405 275 1435
rect 325 1405 355 1435
rect 405 1405 435 1435
rect 485 1405 515 1435
rect 565 1405 595 1435
rect 645 1405 675 1435
rect 725 1405 755 1435
rect 805 1405 835 1435
rect 885 1405 915 1435
rect 965 1405 995 1435
rect 1045 1405 1075 1435
rect 1125 1405 1155 1435
rect 1205 1405 1235 1435
rect 1285 1405 1315 1435
rect 1365 1405 1395 1435
rect 1445 1405 1475 1435
rect 1525 1405 1555 1435
rect 1605 1405 1635 1435
rect 1685 1405 1715 1435
rect 1765 1405 1795 1435
rect 1845 1405 1875 1435
rect 1925 1405 1955 1435
rect 2005 1405 2035 1435
rect 2085 1405 2115 1435
rect 2165 1405 2195 1435
rect 2245 1405 2275 1435
rect 2325 1405 2355 1435
rect 2405 1405 2435 1435
rect 2485 1405 2515 1435
rect 2565 1405 2595 1435
rect 2645 1405 2675 1435
rect 2725 1405 2755 1435
rect 2805 1405 2835 1435
rect 2885 1405 2915 1435
rect 2965 1405 2995 1435
rect 3045 1405 3075 1435
rect 3125 1405 3155 1435
rect 3205 1405 3235 1435
rect 3285 1405 3315 1435
rect 3365 1405 3395 1435
rect 3445 1405 3475 1435
rect 3525 1405 3555 1435
rect 3605 1405 3635 1435
rect 3685 1405 3715 1435
rect 3765 1405 3795 1435
rect 3845 1405 3875 1435
rect 3925 1405 3955 1435
rect 4005 1405 4035 1435
rect 4085 1405 4115 1435
rect 4165 1405 4195 1435
rect 4245 1405 4275 1435
rect 4325 1405 4355 1435
rect 4405 1405 4435 1435
rect 4485 1405 4515 1435
rect 4565 1405 4595 1435
rect 4645 1405 4675 1435
rect 4725 1405 4755 1435
rect 4805 1405 4835 1435
rect 4885 1405 4915 1435
rect 5045 1405 5075 1435
rect 5205 1405 5235 1435
rect 5365 1405 5395 1435
rect 5525 1405 5555 1435
rect 5685 1405 5715 1435
rect -1515 1325 -1485 1355
rect -1355 1325 -1325 1355
rect -1195 1325 -1165 1355
rect -1035 1325 -1005 1355
rect -875 1325 -845 1355
rect -795 1325 -765 1355
rect -715 1325 -685 1355
rect -635 1325 -605 1355
rect -555 1325 -525 1355
rect -475 1325 -445 1355
rect -395 1325 -365 1355
rect -315 1325 -285 1355
rect -235 1325 -205 1355
rect -155 1325 -125 1355
rect -75 1325 -45 1355
rect 5 1325 35 1355
rect 85 1325 115 1355
rect 165 1325 195 1355
rect 245 1325 275 1355
rect 325 1325 355 1355
rect 405 1325 435 1355
rect 485 1325 515 1355
rect 565 1325 595 1355
rect 645 1325 675 1355
rect 725 1325 755 1355
rect 805 1325 835 1355
rect 885 1325 915 1355
rect 965 1325 995 1355
rect 1045 1325 1075 1355
rect 1125 1325 1155 1355
rect 1205 1325 1235 1355
rect 1285 1325 1315 1355
rect 1365 1325 1395 1355
rect 1445 1325 1475 1355
rect 1525 1325 1555 1355
rect 1605 1325 1635 1355
rect 1685 1325 1715 1355
rect 1765 1325 1795 1355
rect 1845 1325 1875 1355
rect 1925 1325 1955 1355
rect 2005 1325 2035 1355
rect 2085 1325 2115 1355
rect 2165 1325 2195 1355
rect 2245 1325 2275 1355
rect 2325 1325 2355 1355
rect 2405 1325 2435 1355
rect 2485 1325 2515 1355
rect 2565 1325 2595 1355
rect 2645 1325 2675 1355
rect 2725 1325 2755 1355
rect 2805 1325 2835 1355
rect 2885 1325 2915 1355
rect 2965 1325 2995 1355
rect 3045 1325 3075 1355
rect 3125 1325 3155 1355
rect 3205 1325 3235 1355
rect 3285 1325 3315 1355
rect 3365 1325 3395 1355
rect 3445 1325 3475 1355
rect 3525 1325 3555 1355
rect 3605 1325 3635 1355
rect 3685 1325 3715 1355
rect 3765 1325 3795 1355
rect 3845 1325 3875 1355
rect 3925 1325 3955 1355
rect 4005 1325 4035 1355
rect 4085 1325 4115 1355
rect 4165 1325 4195 1355
rect 4245 1325 4275 1355
rect 4325 1325 4355 1355
rect 4405 1325 4435 1355
rect 4485 1325 4515 1355
rect 4565 1325 4595 1355
rect 4645 1325 4675 1355
rect 4725 1325 4755 1355
rect 4805 1325 4835 1355
rect 4885 1325 4915 1355
rect 5045 1325 5075 1355
rect 5205 1325 5235 1355
rect 5365 1325 5395 1355
rect 5525 1325 5555 1355
rect 5685 1325 5715 1355
rect -1515 1245 -1485 1275
rect -1355 1245 -1325 1275
rect -1195 1245 -1165 1275
rect -1035 1245 -1005 1275
rect -875 1245 -845 1275
rect -795 1245 -765 1275
rect -715 1245 -685 1275
rect -635 1245 -605 1275
rect -555 1245 -525 1275
rect -475 1245 -445 1275
rect -395 1245 -365 1275
rect -315 1245 -285 1275
rect -235 1245 -205 1275
rect -155 1245 -125 1275
rect -75 1245 -45 1275
rect 5 1245 35 1275
rect 85 1245 115 1275
rect 165 1245 195 1275
rect 245 1245 275 1275
rect 325 1245 355 1275
rect 405 1245 435 1275
rect 485 1245 515 1275
rect 565 1245 595 1275
rect 645 1245 675 1275
rect 725 1245 755 1275
rect 805 1245 835 1275
rect 885 1245 915 1275
rect 965 1245 995 1275
rect 1045 1245 1075 1275
rect 1125 1245 1155 1275
rect 1205 1245 1235 1275
rect 1285 1245 1315 1275
rect 1365 1245 1395 1275
rect 1445 1245 1475 1275
rect 1525 1245 1555 1275
rect 1605 1245 1635 1275
rect 1685 1245 1715 1275
rect 1765 1245 1795 1275
rect 1845 1245 1875 1275
rect 1925 1245 1955 1275
rect 2005 1245 2035 1275
rect 2085 1245 2115 1275
rect 2165 1245 2195 1275
rect 2245 1245 2275 1275
rect 2325 1245 2355 1275
rect 2405 1245 2435 1275
rect 2485 1245 2515 1275
rect 2565 1245 2595 1275
rect 2645 1245 2675 1275
rect 2725 1245 2755 1275
rect 2805 1245 2835 1275
rect 2885 1245 2915 1275
rect 2965 1245 2995 1275
rect 3045 1245 3075 1275
rect 3125 1245 3155 1275
rect 3205 1245 3235 1275
rect 3285 1245 3315 1275
rect 3365 1245 3395 1275
rect 3445 1245 3475 1275
rect 3525 1245 3555 1275
rect 3605 1245 3635 1275
rect 3685 1245 3715 1275
rect 3765 1245 3795 1275
rect 3845 1245 3875 1275
rect 3925 1245 3955 1275
rect 4005 1245 4035 1275
rect 4085 1245 4115 1275
rect 4165 1245 4195 1275
rect 4245 1245 4275 1275
rect 4325 1245 4355 1275
rect 4405 1245 4435 1275
rect 4485 1245 4515 1275
rect 4565 1245 4595 1275
rect 4645 1245 4675 1275
rect 4725 1245 4755 1275
rect 4805 1245 4835 1275
rect 4885 1245 4915 1275
rect 5045 1245 5075 1275
rect 5205 1245 5235 1275
rect 5365 1245 5395 1275
rect 5525 1245 5555 1275
rect 5685 1245 5715 1275
rect -1515 1165 -1485 1195
rect -1355 1165 -1325 1195
rect -1195 1165 -1165 1195
rect -1035 1165 -1005 1195
rect -875 1165 -845 1195
rect -795 1165 -765 1195
rect -715 1165 -685 1195
rect -635 1165 -605 1195
rect -555 1165 -525 1195
rect -475 1165 -445 1195
rect -395 1165 -365 1195
rect -315 1165 -285 1195
rect -235 1165 -205 1195
rect -155 1165 -125 1195
rect -75 1165 -45 1195
rect 5 1165 35 1195
rect 85 1165 115 1195
rect 165 1165 195 1195
rect 245 1165 275 1195
rect 325 1165 355 1195
rect 405 1165 435 1195
rect 485 1165 515 1195
rect 565 1165 595 1195
rect 645 1165 675 1195
rect 725 1165 755 1195
rect 805 1165 835 1195
rect 885 1165 915 1195
rect 965 1165 995 1195
rect 1045 1165 1075 1195
rect 1125 1165 1155 1195
rect 1205 1165 1235 1195
rect 1285 1165 1315 1195
rect 1365 1165 1395 1195
rect 1445 1165 1475 1195
rect 1525 1165 1555 1195
rect 1605 1165 1635 1195
rect 1685 1165 1715 1195
rect 1765 1165 1795 1195
rect 1845 1165 1875 1195
rect 1925 1165 1955 1195
rect 2005 1165 2035 1195
rect 2085 1165 2115 1195
rect 2165 1165 2195 1195
rect 2245 1165 2275 1195
rect 2325 1165 2355 1195
rect 2405 1165 2435 1195
rect 2485 1165 2515 1195
rect 2565 1165 2595 1195
rect 2645 1165 2675 1195
rect 2725 1165 2755 1195
rect 2805 1165 2835 1195
rect 2885 1165 2915 1195
rect 2965 1165 2995 1195
rect 3045 1165 3075 1195
rect 3125 1165 3155 1195
rect 3205 1165 3235 1195
rect 3285 1165 3315 1195
rect 3365 1165 3395 1195
rect 3445 1165 3475 1195
rect 3525 1165 3555 1195
rect 3605 1165 3635 1195
rect 3685 1165 3715 1195
rect 3765 1165 3795 1195
rect 3845 1165 3875 1195
rect 3925 1165 3955 1195
rect 4005 1165 4035 1195
rect 4085 1165 4115 1195
rect 4165 1165 4195 1195
rect 4245 1165 4275 1195
rect 4325 1165 4355 1195
rect 4405 1165 4435 1195
rect 4485 1165 4515 1195
rect 4565 1165 4595 1195
rect 4645 1165 4675 1195
rect 4725 1165 4755 1195
rect 4805 1165 4835 1195
rect 4885 1165 4915 1195
rect 5045 1165 5075 1195
rect 5205 1165 5235 1195
rect 5365 1165 5395 1195
rect 5525 1165 5555 1195
rect 5685 1165 5715 1195
rect -1515 1085 -1485 1115
rect -1355 1085 -1325 1115
rect -1195 1085 -1165 1115
rect -1115 1085 -1085 1115
rect 4885 1085 4915 1115
rect 5045 1085 5075 1115
rect 5205 1085 5235 1115
rect 5365 1085 5395 1115
rect 5525 1085 5555 1115
rect 5685 1085 5715 1115
rect -1515 1005 -1485 1035
rect -1355 1005 -1325 1035
rect -1195 1005 -1165 1035
rect -1035 1005 -1005 1035
rect -875 1005 -845 1035
rect -795 1005 -765 1035
rect -715 1005 -685 1035
rect -635 1005 -605 1035
rect -555 1005 -525 1035
rect -475 1005 -445 1035
rect -395 1005 -365 1035
rect -315 1005 -285 1035
rect -235 1005 -205 1035
rect -155 1005 -125 1035
rect -75 1005 -45 1035
rect 5 1005 35 1035
rect 85 1005 115 1035
rect 165 1005 195 1035
rect 245 1005 275 1035
rect 325 1005 355 1035
rect 405 1005 435 1035
rect 485 1005 515 1035
rect 565 1005 595 1035
rect 645 1005 675 1035
rect 725 1005 755 1035
rect 805 1005 835 1035
rect 885 1005 915 1035
rect 965 1005 995 1035
rect 1045 1005 1075 1035
rect 1125 1005 1155 1035
rect 1205 1005 1235 1035
rect 1285 1005 1315 1035
rect 1365 1005 1395 1035
rect 1445 1005 1475 1035
rect 1525 1005 1555 1035
rect 1605 1005 1635 1035
rect 1685 1005 1715 1035
rect 1765 1005 1795 1035
rect 1845 1005 1875 1035
rect 1925 1005 1955 1035
rect 2005 1005 2035 1035
rect 2085 1005 2115 1035
rect 2165 1005 2195 1035
rect 2245 1005 2275 1035
rect 2325 1005 2355 1035
rect 2405 1005 2435 1035
rect 2485 1005 2515 1035
rect 2565 1005 2595 1035
rect 2645 1005 2675 1035
rect 2725 1005 2755 1035
rect 2805 1005 2835 1035
rect 2885 1005 2915 1035
rect 2965 1005 2995 1035
rect 3045 1005 3075 1035
rect 3125 1005 3155 1035
rect 3205 1005 3235 1035
rect 3285 1005 3315 1035
rect 3365 1005 3395 1035
rect 3445 1005 3475 1035
rect 3525 1005 3555 1035
rect 3605 1005 3635 1035
rect 3685 1005 3715 1035
rect 3765 1005 3795 1035
rect 3845 1005 3875 1035
rect 3925 1005 3955 1035
rect 4005 1005 4035 1035
rect 4085 1005 4115 1035
rect 4165 1005 4195 1035
rect 4245 1005 4275 1035
rect 4325 1005 4355 1035
rect 4405 1005 4435 1035
rect 4485 1005 4515 1035
rect 4565 1005 4595 1035
rect 4645 1005 4675 1035
rect 4725 1005 4755 1035
rect 4805 1005 4835 1035
rect 4885 1005 4915 1035
rect 5045 1005 5075 1035
rect 5205 1005 5235 1035
rect 5365 1005 5395 1035
rect 5525 1005 5555 1035
rect 5685 1005 5715 1035
rect -1515 925 -1485 955
rect -1355 925 -1325 955
rect -1195 925 -1165 955
rect -1035 925 -1005 955
rect -875 925 -845 955
rect -795 925 -765 955
rect -715 925 -685 955
rect -635 925 -605 955
rect -555 925 -525 955
rect -475 925 -445 955
rect -395 925 -365 955
rect -315 925 -285 955
rect -235 925 -205 955
rect -155 925 -125 955
rect -75 925 -45 955
rect 5 925 35 955
rect 85 925 115 955
rect 165 925 195 955
rect 245 925 275 955
rect 325 925 355 955
rect 405 925 435 955
rect 485 925 515 955
rect 565 925 595 955
rect 645 925 675 955
rect 725 925 755 955
rect 805 925 835 955
rect 885 925 915 955
rect 965 925 995 955
rect 1045 925 1075 955
rect 1125 925 1155 955
rect 1205 925 1235 955
rect 1285 925 1315 955
rect 1365 925 1395 955
rect 1445 925 1475 955
rect 1525 925 1555 955
rect 1605 925 1635 955
rect 1685 925 1715 955
rect 1765 925 1795 955
rect 1845 925 1875 955
rect 1925 925 1955 955
rect 2005 925 2035 955
rect 2085 925 2115 955
rect 2165 925 2195 955
rect 2245 925 2275 955
rect 2325 925 2355 955
rect 2405 925 2435 955
rect 2485 925 2515 955
rect 2565 925 2595 955
rect 2645 925 2675 955
rect 2725 925 2755 955
rect 2805 925 2835 955
rect 2885 925 2915 955
rect 2965 925 2995 955
rect 3045 925 3075 955
rect 3125 925 3155 955
rect 3205 925 3235 955
rect 3285 925 3315 955
rect 3365 925 3395 955
rect 3445 925 3475 955
rect 3525 925 3555 955
rect 3605 925 3635 955
rect 3685 925 3715 955
rect 3765 925 3795 955
rect 3845 925 3875 955
rect 3925 925 3955 955
rect 4005 925 4035 955
rect 4085 925 4115 955
rect 4165 925 4195 955
rect 4245 925 4275 955
rect 4325 925 4355 955
rect 4405 925 4435 955
rect 4485 925 4515 955
rect 4565 925 4595 955
rect 4645 925 4675 955
rect 4725 925 4755 955
rect 4805 925 4835 955
rect 4885 925 4915 955
rect 5045 925 5075 955
rect 5205 925 5235 955
rect 5365 925 5395 955
rect 5525 925 5555 955
rect 5685 925 5715 955
rect -1515 845 -1485 875
rect -1355 845 -1325 875
rect -1195 845 -1165 875
rect -1035 845 -1005 875
rect -875 845 -845 875
rect -795 845 -765 875
rect -715 845 -685 875
rect -635 845 -605 875
rect -555 845 -525 875
rect -475 845 -445 875
rect -395 845 -365 875
rect -315 845 -285 875
rect -235 845 -205 875
rect -155 845 -125 875
rect -75 845 -45 875
rect 5 845 35 875
rect 85 845 115 875
rect 165 845 195 875
rect 245 845 275 875
rect 325 845 355 875
rect 405 845 435 875
rect 485 845 515 875
rect 565 845 595 875
rect 645 845 675 875
rect 725 845 755 875
rect 805 845 835 875
rect 885 845 915 875
rect 965 845 995 875
rect 1045 845 1075 875
rect 1125 845 1155 875
rect 1205 845 1235 875
rect 1285 845 1315 875
rect 1365 845 1395 875
rect 1445 845 1475 875
rect 1525 845 1555 875
rect 1605 845 1635 875
rect 1685 845 1715 875
rect 1765 845 1795 875
rect 1845 845 1875 875
rect 1925 845 1955 875
rect 2005 845 2035 875
rect 2085 845 2115 875
rect 2165 845 2195 875
rect 2245 845 2275 875
rect 2325 845 2355 875
rect 2405 845 2435 875
rect 2485 845 2515 875
rect 2565 845 2595 875
rect 2645 845 2675 875
rect 2725 845 2755 875
rect 2805 845 2835 875
rect 2885 845 2915 875
rect 2965 845 2995 875
rect 3045 845 3075 875
rect 3125 845 3155 875
rect 3205 845 3235 875
rect 3285 845 3315 875
rect 3365 845 3395 875
rect 3445 845 3475 875
rect 3525 845 3555 875
rect 3605 845 3635 875
rect 3685 845 3715 875
rect 3765 845 3795 875
rect 3845 845 3875 875
rect 3925 845 3955 875
rect 4005 845 4035 875
rect 4085 845 4115 875
rect 4165 845 4195 875
rect 4245 845 4275 875
rect 4325 845 4355 875
rect 4405 845 4435 875
rect 4485 845 4515 875
rect 4565 845 4595 875
rect 4645 845 4675 875
rect 4725 845 4755 875
rect 4805 845 4835 875
rect 4885 845 4915 875
rect 5045 845 5075 875
rect 5205 845 5235 875
rect 5365 845 5395 875
rect 5525 845 5555 875
rect 5685 845 5715 875
rect -1515 765 -1485 795
rect -1355 765 -1325 795
rect -1195 765 -1165 795
rect -1035 765 -1005 795
rect -875 765 -845 795
rect 5445 765 5475 795
rect 5525 765 5555 795
rect 5685 765 5715 795
rect -1515 685 -1485 715
rect -1355 685 -1325 715
rect -1195 685 -1165 715
rect -1035 685 -1005 715
rect -875 685 -845 715
rect -795 685 -765 715
rect -715 685 -685 715
rect -635 685 -605 715
rect -555 685 -525 715
rect -475 685 -445 715
rect -395 685 -365 715
rect -315 685 -285 715
rect -235 685 -205 715
rect -155 685 -125 715
rect -75 685 -45 715
rect 5 685 35 715
rect 85 685 115 715
rect 165 685 195 715
rect 245 685 275 715
rect 325 685 355 715
rect 405 685 435 715
rect 485 685 515 715
rect 565 685 595 715
rect 645 685 675 715
rect 725 685 755 715
rect 805 685 835 715
rect 885 685 915 715
rect 965 685 995 715
rect 1045 685 1075 715
rect 1125 685 1155 715
rect 1205 685 1235 715
rect 1285 685 1315 715
rect 1365 685 1395 715
rect 1445 685 1475 715
rect 1525 685 1555 715
rect 1605 685 1635 715
rect 1685 685 1715 715
rect 1765 685 1795 715
rect 1845 685 1875 715
rect 1925 685 1955 715
rect 2005 685 2035 715
rect 2085 685 2115 715
rect 2165 685 2195 715
rect 2245 685 2275 715
rect 2325 685 2355 715
rect 2405 685 2435 715
rect 2485 685 2515 715
rect 2565 685 2595 715
rect 2645 685 2675 715
rect 2725 685 2755 715
rect 2805 685 2835 715
rect 2885 685 2915 715
rect 2965 685 2995 715
rect 3045 685 3075 715
rect 3125 685 3155 715
rect 3205 685 3235 715
rect 3285 685 3315 715
rect 3365 685 3395 715
rect 3445 685 3475 715
rect 3525 685 3555 715
rect 3605 685 3635 715
rect 3685 685 3715 715
rect 3765 685 3795 715
rect 3845 685 3875 715
rect 3925 685 3955 715
rect 4005 685 4035 715
rect 4085 685 4115 715
rect 4165 685 4195 715
rect 4245 685 4275 715
rect 4325 685 4355 715
rect 4405 685 4435 715
rect 4485 685 4515 715
rect 4565 685 4595 715
rect 4645 685 4675 715
rect 4725 685 4755 715
rect 4805 685 4835 715
rect 4885 685 4915 715
rect 5045 685 5075 715
rect 5205 685 5235 715
rect 5365 685 5395 715
rect 5525 685 5555 715
rect 5685 685 5715 715
rect -1515 605 -1485 635
rect -1355 605 -1325 635
rect -1195 605 -1165 635
rect -1035 605 -1005 635
rect -875 605 -845 635
rect 5285 605 5315 635
rect 5365 605 5395 635
rect 5525 605 5555 635
rect 5685 605 5715 635
rect -1515 525 -1485 555
rect -1355 525 -1325 555
rect -1195 525 -1165 555
rect -1035 525 -1005 555
rect -875 525 -845 555
rect -795 525 -765 555
rect -715 525 -685 555
rect -635 525 -605 555
rect -555 525 -525 555
rect -475 525 -445 555
rect -395 525 -365 555
rect -315 525 -285 555
rect -235 525 -205 555
rect -155 525 -125 555
rect -75 525 -45 555
rect 5 525 35 555
rect 85 525 115 555
rect 165 525 195 555
rect 245 525 275 555
rect 325 525 355 555
rect 405 525 435 555
rect 485 525 515 555
rect 565 525 595 555
rect 645 525 675 555
rect 725 525 755 555
rect 805 525 835 555
rect 885 525 915 555
rect 965 525 995 555
rect 1045 525 1075 555
rect 1125 525 1155 555
rect 1205 525 1235 555
rect 1285 525 1315 555
rect 1365 525 1395 555
rect 1445 525 1475 555
rect 1525 525 1555 555
rect 1605 525 1635 555
rect 1685 525 1715 555
rect 1765 525 1795 555
rect 1845 525 1875 555
rect 1925 525 1955 555
rect 2005 525 2035 555
rect 2085 525 2115 555
rect 2165 525 2195 555
rect 2245 525 2275 555
rect 2325 525 2355 555
rect 2405 525 2435 555
rect 2485 525 2515 555
rect 2565 525 2595 555
rect 2645 525 2675 555
rect 2725 525 2755 555
rect 2805 525 2835 555
rect 2885 525 2915 555
rect 2965 525 2995 555
rect 3045 525 3075 555
rect 3125 525 3155 555
rect 3205 525 3235 555
rect 3285 525 3315 555
rect 3365 525 3395 555
rect 3445 525 3475 555
rect 3525 525 3555 555
rect 3605 525 3635 555
rect 3685 525 3715 555
rect 3765 525 3795 555
rect 3845 525 3875 555
rect 3925 525 3955 555
rect 4005 525 4035 555
rect 4085 525 4115 555
rect 4165 525 4195 555
rect 4245 525 4275 555
rect 4325 525 4355 555
rect 4405 525 4435 555
rect 4485 525 4515 555
rect 4565 525 4595 555
rect 4645 525 4675 555
rect 4725 525 4755 555
rect 4805 525 4835 555
rect 4885 525 4915 555
rect 5045 525 5075 555
rect 5205 525 5235 555
rect 5365 525 5395 555
rect 5525 525 5555 555
rect 5685 525 5715 555
rect -1515 445 -1485 475
rect -1355 445 -1325 475
rect -1195 445 -1165 475
rect -1035 445 -1005 475
rect -875 445 -845 475
rect 5125 445 5155 475
rect 5205 445 5235 475
rect 5365 445 5395 475
rect 5525 445 5555 475
rect 5685 445 5715 475
rect -1515 365 -1485 395
rect -1355 365 -1325 395
rect -1195 365 -1165 395
rect -1035 365 -1005 395
rect -875 365 -845 395
rect -795 365 -765 395
rect -715 365 -685 395
rect -635 365 -605 395
rect -555 365 -525 395
rect -475 365 -445 395
rect -395 365 -365 395
rect -315 365 -285 395
rect -235 365 -205 395
rect -155 365 -125 395
rect -75 365 -45 395
rect 5 365 35 395
rect 85 365 115 395
rect 165 365 195 395
rect 245 365 275 395
rect 325 365 355 395
rect 405 365 435 395
rect 485 365 515 395
rect 565 365 595 395
rect 645 365 675 395
rect 725 365 755 395
rect 805 365 835 395
rect 885 365 915 395
rect 965 365 995 395
rect 1045 365 1075 395
rect 1125 365 1155 395
rect 1205 365 1235 395
rect 1285 365 1315 395
rect 1365 365 1395 395
rect 1445 365 1475 395
rect 1525 365 1555 395
rect 1605 365 1635 395
rect 1685 365 1715 395
rect 1765 365 1795 395
rect 1845 365 1875 395
rect 1925 365 1955 395
rect 2005 365 2035 395
rect 2085 365 2115 395
rect 2165 365 2195 395
rect 2245 365 2275 395
rect 2325 365 2355 395
rect 2405 365 2435 395
rect 2485 365 2515 395
rect 2565 365 2595 395
rect 2645 365 2675 395
rect 2725 365 2755 395
rect 2805 365 2835 395
rect 2885 365 2915 395
rect 2965 365 2995 395
rect 3045 365 3075 395
rect 3125 365 3155 395
rect 3205 365 3235 395
rect 3285 365 3315 395
rect 3365 365 3395 395
rect 3445 365 3475 395
rect 3525 365 3555 395
rect 3605 365 3635 395
rect 3685 365 3715 395
rect 3765 365 3795 395
rect 3845 365 3875 395
rect 3925 365 3955 395
rect 4005 365 4035 395
rect 4085 365 4115 395
rect 4165 365 4195 395
rect 4245 365 4275 395
rect 4325 365 4355 395
rect 4405 365 4435 395
rect 4485 365 4515 395
rect 4565 365 4595 395
rect 4645 365 4675 395
rect 4725 365 4755 395
rect 4805 365 4835 395
rect 4885 365 4915 395
rect 5045 365 5075 395
rect 5205 365 5235 395
rect 5365 365 5395 395
rect 5525 365 5555 395
rect 5685 365 5715 395
rect -1515 285 -1485 315
rect -1355 285 -1325 315
rect -1195 285 -1165 315
rect -1035 285 -1005 315
rect -875 285 -845 315
rect 4965 285 4995 315
rect 5045 285 5075 315
rect 5205 285 5235 315
rect 5365 285 5395 315
rect 5525 285 5555 315
rect 5685 285 5715 315
rect -1515 205 -1485 235
rect -1355 205 -1325 235
rect -1195 205 -1165 235
rect -1035 205 -1005 235
rect -875 205 -845 235
rect -795 205 -765 235
rect -715 205 -685 235
rect -635 205 -605 235
rect -555 205 -525 235
rect -475 205 -445 235
rect -395 205 -365 235
rect -315 205 -285 235
rect -235 205 -205 235
rect -155 205 -125 235
rect -75 205 -45 235
rect 5 205 35 235
rect 85 205 115 235
rect 165 205 195 235
rect 245 205 275 235
rect 325 205 355 235
rect 405 205 435 235
rect 485 205 515 235
rect 565 205 595 235
rect 645 205 675 235
rect 725 205 755 235
rect 805 205 835 235
rect 885 205 915 235
rect 965 205 995 235
rect 1045 205 1075 235
rect 1125 205 1155 235
rect 1205 205 1235 235
rect 1285 205 1315 235
rect 1365 205 1395 235
rect 1445 205 1475 235
rect 1525 205 1555 235
rect 1605 205 1635 235
rect 1685 205 1715 235
rect 1765 205 1795 235
rect 1845 205 1875 235
rect 1925 205 1955 235
rect 2005 205 2035 235
rect 2085 205 2115 235
rect 2165 205 2195 235
rect 2245 205 2275 235
rect 2325 205 2355 235
rect 2405 205 2435 235
rect 2485 205 2515 235
rect 2565 205 2595 235
rect 2645 205 2675 235
rect 2725 205 2755 235
rect 2805 205 2835 235
rect 2885 205 2915 235
rect 2965 205 2995 235
rect 3045 205 3075 235
rect 3125 205 3155 235
rect 3205 205 3235 235
rect 3285 205 3315 235
rect 3365 205 3395 235
rect 3445 205 3475 235
rect 3525 205 3555 235
rect 3605 205 3635 235
rect 3685 205 3715 235
rect 3765 205 3795 235
rect 3845 205 3875 235
rect 3925 205 3955 235
rect 4005 205 4035 235
rect 4085 205 4115 235
rect 4165 205 4195 235
rect 4245 205 4275 235
rect 4325 205 4355 235
rect 4405 205 4435 235
rect 4485 205 4515 235
rect 4565 205 4595 235
rect 4645 205 4675 235
rect 4725 205 4755 235
rect 4805 205 4835 235
rect 4885 205 4915 235
rect 5045 205 5075 235
rect 5205 205 5235 235
rect 5365 205 5395 235
rect 5525 205 5555 235
rect 5685 205 5715 235
rect -1515 125 -1485 155
rect -1355 125 -1325 155
rect -1195 125 -1165 155
rect -1035 125 -1005 155
rect -875 125 -845 155
rect -795 125 -765 155
rect -715 125 -685 155
rect -635 125 -605 155
rect -555 125 -525 155
rect -475 125 -445 155
rect -395 125 -365 155
rect -315 125 -285 155
rect -235 125 -205 155
rect -155 125 -125 155
rect -75 125 -45 155
rect 5 125 35 155
rect 85 125 115 155
rect 165 125 195 155
rect 245 125 275 155
rect 325 125 355 155
rect 405 125 435 155
rect 485 125 515 155
rect 565 125 595 155
rect 645 125 675 155
rect 725 125 755 155
rect 805 125 835 155
rect 885 125 915 155
rect 965 125 995 155
rect 1045 125 1075 155
rect 1125 125 1155 155
rect 1205 125 1235 155
rect 1285 125 1315 155
rect 1365 125 1395 155
rect 1445 125 1475 155
rect 1525 125 1555 155
rect 1605 125 1635 155
rect 1685 125 1715 155
rect 1765 125 1795 155
rect 1845 125 1875 155
rect 1925 125 1955 155
rect 2005 125 2035 155
rect 2085 125 2115 155
rect 2165 125 2195 155
rect 2245 125 2275 155
rect 2325 125 2355 155
rect 2405 125 2435 155
rect 2485 125 2515 155
rect 2565 125 2595 155
rect 2645 125 2675 155
rect 2725 125 2755 155
rect 2805 125 2835 155
rect 2885 125 2915 155
rect 2965 125 2995 155
rect 3045 125 3075 155
rect 3125 125 3155 155
rect 3205 125 3235 155
rect 3285 125 3315 155
rect 3365 125 3395 155
rect 3445 125 3475 155
rect 3525 125 3555 155
rect 3605 125 3635 155
rect 3685 125 3715 155
rect 3765 125 3795 155
rect 3845 125 3875 155
rect 3925 125 3955 155
rect 4005 125 4035 155
rect 4085 125 4115 155
rect 4165 125 4195 155
rect 4245 125 4275 155
rect 4325 125 4355 155
rect 4405 125 4435 155
rect 4485 125 4515 155
rect 4565 125 4595 155
rect 4645 125 4675 155
rect 4725 125 4755 155
rect 4805 125 4835 155
rect 4885 125 4915 155
rect 5045 125 5075 155
rect 5205 125 5235 155
rect 5365 125 5395 155
rect 5525 125 5555 155
rect 5685 125 5715 155
rect -1515 45 -1485 75
rect -1355 45 -1325 75
rect -1195 45 -1165 75
rect -1035 45 -1005 75
rect -875 45 -845 75
rect -795 45 -765 75
rect -715 45 -685 75
rect -635 45 -605 75
rect -555 45 -525 75
rect -475 45 -445 75
rect -395 45 -365 75
rect -315 45 -285 75
rect -235 45 -205 75
rect -155 45 -125 75
rect -75 45 -45 75
rect 5 45 35 75
rect 85 45 115 75
rect 165 45 195 75
rect 245 45 275 75
rect 325 45 355 75
rect 405 45 435 75
rect 485 45 515 75
rect 565 45 595 75
rect 645 45 675 75
rect 725 45 755 75
rect 805 45 835 75
rect 885 45 915 75
rect 965 45 995 75
rect 1045 45 1075 75
rect 1125 45 1155 75
rect 1205 45 1235 75
rect 1285 45 1315 75
rect 1365 45 1395 75
rect 1445 45 1475 75
rect 1525 45 1555 75
rect 1605 45 1635 75
rect 1685 45 1715 75
rect 1765 45 1795 75
rect 1845 45 1875 75
rect 1925 45 1955 75
rect 2005 45 2035 75
rect 2085 45 2115 75
rect 2165 45 2195 75
rect 2245 45 2275 75
rect 2325 45 2355 75
rect 2405 45 2435 75
rect 2485 45 2515 75
rect 2565 45 2595 75
rect 2645 45 2675 75
rect 2725 45 2755 75
rect 2805 45 2835 75
rect 2885 45 2915 75
rect 2965 45 2995 75
rect 3045 45 3075 75
rect 3125 45 3155 75
rect 3205 45 3235 75
rect 3285 45 3315 75
rect 3365 45 3395 75
rect 3445 45 3475 75
rect 3525 45 3555 75
rect 3605 45 3635 75
rect 3685 45 3715 75
rect 3765 45 3795 75
rect 3845 45 3875 75
rect 3925 45 3955 75
rect 4005 45 4035 75
rect 4085 45 4115 75
rect 4165 45 4195 75
rect 4245 45 4275 75
rect 4325 45 4355 75
rect 4405 45 4435 75
rect 4485 45 4515 75
rect 4565 45 4595 75
rect 4645 45 4675 75
rect 4725 45 4755 75
rect 4805 45 4835 75
rect 4885 45 4915 75
rect 5045 45 5075 75
rect 5205 45 5235 75
rect 5365 45 5395 75
rect 5525 45 5555 75
rect 5685 45 5715 75
rect -1515 -35 -1485 -5
rect -1355 -35 -1325 -5
rect -1195 -35 -1165 -5
rect -1035 -35 -1005 -5
rect -875 -35 -845 -5
rect -795 -35 -765 -5
rect -715 -35 -685 -5
rect -635 -35 -605 -5
rect -555 -35 -525 -5
rect -475 -35 -445 -5
rect -395 -35 -365 -5
rect -315 -35 -285 -5
rect -235 -35 -205 -5
rect -155 -35 -125 -5
rect -75 -35 -45 -5
rect 5 -35 35 -5
rect 85 -35 115 -5
rect 165 -35 195 -5
rect 245 -35 275 -5
rect 325 -35 355 -5
rect 405 -35 435 -5
rect 485 -35 515 -5
rect 565 -35 595 -5
rect 645 -35 675 -5
rect 725 -35 755 -5
rect 805 -35 835 -5
rect 885 -35 915 -5
rect 965 -35 995 -5
rect 1045 -35 1075 -5
rect 1125 -35 1155 -5
rect 1205 -35 1235 -5
rect 1285 -35 1315 -5
rect 1365 -35 1395 -5
rect 1445 -35 1475 -5
rect 1525 -35 1555 -5
rect 1605 -35 1635 -5
rect 1685 -35 1715 -5
rect 1765 -35 1795 -5
rect 1845 -35 1875 -5
rect 1925 -35 1955 -5
rect 2005 -35 2035 -5
rect 2085 -35 2115 -5
rect 2165 -35 2195 -5
rect 2245 -35 2275 -5
rect 2325 -35 2355 -5
rect 2405 -35 2435 -5
rect 2485 -35 2515 -5
rect 2565 -35 2595 -5
rect 2645 -35 2675 -5
rect 2725 -35 2755 -5
rect 2805 -35 2835 -5
rect 2885 -35 2915 -5
rect 2965 -35 2995 -5
rect 3045 -35 3075 -5
rect 3125 -35 3155 -5
rect 3205 -35 3235 -5
rect 3285 -35 3315 -5
rect 3365 -35 3395 -5
rect 3445 -35 3475 -5
rect 3525 -35 3555 -5
rect 3605 -35 3635 -5
rect 3685 -35 3715 -5
rect 3765 -35 3795 -5
rect 3845 -35 3875 -5
rect 3925 -35 3955 -5
rect 4005 -35 4035 -5
rect 4085 -35 4115 -5
rect 4165 -35 4195 -5
rect 4245 -35 4275 -5
rect 4325 -35 4355 -5
rect 4405 -35 4435 -5
rect 4485 -35 4515 -5
rect 4565 -35 4595 -5
rect 4645 -35 4675 -5
rect 4725 -35 4755 -5
rect 4805 -35 4835 -5
rect 4885 -35 4915 -5
rect 5045 -35 5075 -5
rect 5205 -35 5235 -5
rect 5365 -35 5395 -5
rect 5525 -35 5555 -5
rect 5685 -35 5715 -5
rect -1515 -115 -1485 -85
rect -1355 -115 -1325 -85
rect -1195 -115 -1165 -85
rect -1035 -115 -1005 -85
rect -875 -115 -845 -85
rect -795 -115 -765 -85
rect -715 -115 -685 -85
rect -635 -115 -605 -85
rect -555 -115 -525 -85
rect -475 -115 -445 -85
rect -395 -115 -365 -85
rect -315 -115 -285 -85
rect -235 -115 -205 -85
rect -155 -115 -125 -85
rect -75 -115 -45 -85
rect 5 -115 35 -85
rect 85 -115 115 -85
rect 165 -115 195 -85
rect 245 -115 275 -85
rect 325 -115 355 -85
rect 405 -115 435 -85
rect 485 -115 515 -85
rect 565 -115 595 -85
rect 645 -115 675 -85
rect 725 -115 755 -85
rect 805 -115 835 -85
rect 885 -115 915 -85
rect 965 -115 995 -85
rect 1045 -115 1075 -85
rect 1125 -115 1155 -85
rect 1205 -115 1235 -85
rect 1285 -115 1315 -85
rect 1365 -115 1395 -85
rect 1445 -115 1475 -85
rect 1525 -115 1555 -85
rect 1605 -115 1635 -85
rect 1685 -115 1715 -85
rect 1765 -115 1795 -85
rect 1845 -115 1875 -85
rect 1925 -115 1955 -85
rect 2005 -115 2035 -85
rect 2085 -115 2115 -85
rect 2165 -115 2195 -85
rect 2245 -115 2275 -85
rect 2325 -115 2355 -85
rect 2405 -115 2435 -85
rect 2485 -115 2515 -85
rect 2565 -115 2595 -85
rect 2645 -115 2675 -85
rect 2725 -115 2755 -85
rect 2805 -115 2835 -85
rect 2885 -115 2915 -85
rect 2965 -115 2995 -85
rect 3045 -115 3075 -85
rect 3125 -115 3155 -85
rect 3205 -115 3235 -85
rect 3285 -115 3315 -85
rect 3365 -115 3395 -85
rect 3445 -115 3475 -85
rect 3525 -115 3555 -85
rect 3605 -115 3635 -85
rect 3685 -115 3715 -85
rect 3765 -115 3795 -85
rect 3845 -115 3875 -85
rect 3925 -115 3955 -85
rect 4005 -115 4035 -85
rect 4085 -115 4115 -85
rect 4165 -115 4195 -85
rect 4245 -115 4275 -85
rect 4325 -115 4355 -85
rect 4405 -115 4435 -85
rect 4485 -115 4515 -85
rect 4565 -115 4595 -85
rect 4645 -115 4675 -85
rect 4725 -115 4755 -85
rect 4805 -115 4835 -85
rect 4885 -115 4915 -85
rect 5045 -115 5075 -85
rect 5205 -115 5235 -85
rect 5365 -115 5395 -85
rect 5525 -115 5555 -85
rect 5685 -115 5715 -85
<< metal3 >>
rect -1520 5596 -1480 5640
rect -1520 5564 -1516 5596
rect -1484 5564 -1480 5596
rect -1520 5516 -1480 5564
rect -1520 5484 -1516 5516
rect -1484 5484 -1480 5516
rect -1520 5436 -1480 5484
rect -1520 5404 -1516 5436
rect -1484 5404 -1480 5436
rect -1520 5356 -1480 5404
rect -1520 5324 -1516 5356
rect -1484 5324 -1480 5356
rect -1520 5276 -1480 5324
rect -1520 5244 -1516 5276
rect -1484 5244 -1480 5276
rect -1520 5196 -1480 5244
rect -1520 5164 -1516 5196
rect -1484 5164 -1480 5196
rect -1520 5116 -1480 5164
rect -1520 5084 -1516 5116
rect -1484 5084 -1480 5116
rect -1520 5036 -1480 5084
rect -1520 5004 -1516 5036
rect -1484 5004 -1480 5036
rect -1520 4956 -1480 5004
rect -1520 4924 -1516 4956
rect -1484 4924 -1480 4956
rect -1520 4876 -1480 4924
rect -1520 4844 -1516 4876
rect -1484 4844 -1480 4876
rect -1520 4796 -1480 4844
rect -1520 4764 -1516 4796
rect -1484 4764 -1480 4796
rect -1520 4716 -1480 4764
rect -1520 4684 -1516 4716
rect -1484 4684 -1480 4716
rect -1520 4636 -1480 4684
rect -1520 4604 -1516 4636
rect -1484 4604 -1480 4636
rect -1520 4556 -1480 4604
rect -1520 4524 -1516 4556
rect -1484 4524 -1480 4556
rect -1520 4476 -1480 4524
rect -1520 4444 -1516 4476
rect -1484 4444 -1480 4476
rect -1520 4396 -1480 4444
rect -1520 4364 -1516 4396
rect -1484 4364 -1480 4396
rect -1520 4316 -1480 4364
rect -1520 4284 -1516 4316
rect -1484 4284 -1480 4316
rect -1520 4236 -1480 4284
rect -1520 4204 -1516 4236
rect -1484 4204 -1480 4236
rect -1520 4156 -1480 4204
rect -1520 4124 -1516 4156
rect -1484 4124 -1480 4156
rect -1520 4076 -1480 4124
rect -1520 4044 -1516 4076
rect -1484 4044 -1480 4076
rect -1520 3996 -1480 4044
rect -1520 3964 -1516 3996
rect -1484 3964 -1480 3996
rect -1520 3916 -1480 3964
rect -1520 3884 -1516 3916
rect -1484 3884 -1480 3916
rect -1520 3836 -1480 3884
rect -1520 3804 -1516 3836
rect -1484 3804 -1480 3836
rect -1520 3756 -1480 3804
rect -1520 3724 -1516 3756
rect -1484 3724 -1480 3756
rect -1520 3676 -1480 3724
rect -1520 3644 -1516 3676
rect -1484 3644 -1480 3676
rect -1520 3596 -1480 3644
rect -1520 3564 -1516 3596
rect -1484 3564 -1480 3596
rect -1520 3516 -1480 3564
rect -1520 3484 -1516 3516
rect -1484 3484 -1480 3516
rect -1520 3436 -1480 3484
rect -1520 3404 -1516 3436
rect -1484 3404 -1480 3436
rect -1520 3356 -1480 3404
rect -1520 3324 -1516 3356
rect -1484 3324 -1480 3356
rect -1520 3276 -1480 3324
rect -1520 3244 -1516 3276
rect -1484 3244 -1480 3276
rect -1520 3196 -1480 3244
rect -1520 3164 -1516 3196
rect -1484 3164 -1480 3196
rect -1520 3116 -1480 3164
rect -1520 3084 -1516 3116
rect -1484 3084 -1480 3116
rect -1520 3036 -1480 3084
rect -1520 3004 -1516 3036
rect -1484 3004 -1480 3036
rect -1520 2956 -1480 3004
rect -1520 2924 -1516 2956
rect -1484 2924 -1480 2956
rect -1520 2876 -1480 2924
rect -1520 2844 -1516 2876
rect -1484 2844 -1480 2876
rect -1520 2796 -1480 2844
rect -1520 2764 -1516 2796
rect -1484 2764 -1480 2796
rect -1520 2716 -1480 2764
rect -1520 2684 -1516 2716
rect -1484 2684 -1480 2716
rect -1520 2636 -1480 2684
rect -1520 2604 -1516 2636
rect -1484 2604 -1480 2636
rect -1520 2556 -1480 2604
rect -1520 2524 -1516 2556
rect -1484 2524 -1480 2556
rect -1520 2476 -1480 2524
rect -1520 2444 -1516 2476
rect -1484 2444 -1480 2476
rect -1520 2396 -1480 2444
rect -1520 2364 -1516 2396
rect -1484 2364 -1480 2396
rect -1520 2316 -1480 2364
rect -1520 2284 -1516 2316
rect -1484 2284 -1480 2316
rect -1520 2236 -1480 2284
rect -1520 2204 -1516 2236
rect -1484 2204 -1480 2236
rect -1520 2156 -1480 2204
rect -1520 2124 -1516 2156
rect -1484 2124 -1480 2156
rect -1520 2076 -1480 2124
rect -1520 2044 -1516 2076
rect -1484 2044 -1480 2076
rect -1520 1996 -1480 2044
rect -1520 1964 -1516 1996
rect -1484 1964 -1480 1996
rect -1520 1916 -1480 1964
rect -1520 1884 -1516 1916
rect -1484 1884 -1480 1916
rect -1520 1836 -1480 1884
rect -1520 1804 -1516 1836
rect -1484 1804 -1480 1836
rect -1520 1756 -1480 1804
rect -1520 1724 -1516 1756
rect -1484 1724 -1480 1756
rect -1520 1676 -1480 1724
rect -1520 1644 -1516 1676
rect -1484 1644 -1480 1676
rect -1520 1596 -1480 1644
rect -1520 1564 -1516 1596
rect -1484 1564 -1480 1596
rect -1520 1516 -1480 1564
rect -1520 1484 -1516 1516
rect -1484 1484 -1480 1516
rect -1520 1436 -1480 1484
rect -1520 1404 -1516 1436
rect -1484 1404 -1480 1436
rect -1520 1356 -1480 1404
rect -1520 1324 -1516 1356
rect -1484 1324 -1480 1356
rect -1520 1276 -1480 1324
rect -1520 1244 -1516 1276
rect -1484 1244 -1480 1276
rect -1520 1196 -1480 1244
rect -1520 1164 -1516 1196
rect -1484 1164 -1480 1196
rect -1520 1116 -1480 1164
rect -1520 1084 -1516 1116
rect -1484 1084 -1480 1116
rect -1520 1036 -1480 1084
rect -1520 1004 -1516 1036
rect -1484 1004 -1480 1036
rect -1520 956 -1480 1004
rect -1520 924 -1516 956
rect -1484 924 -1480 956
rect -1520 876 -1480 924
rect -1520 844 -1516 876
rect -1484 844 -1480 876
rect -1520 796 -1480 844
rect -1520 764 -1516 796
rect -1484 764 -1480 796
rect -1520 716 -1480 764
rect -1520 684 -1516 716
rect -1484 684 -1480 716
rect -1520 636 -1480 684
rect -1520 604 -1516 636
rect -1484 604 -1480 636
rect -1520 556 -1480 604
rect -1520 524 -1516 556
rect -1484 524 -1480 556
rect -1520 476 -1480 524
rect -1520 444 -1516 476
rect -1484 444 -1480 476
rect -1520 396 -1480 444
rect -1520 364 -1516 396
rect -1484 364 -1480 396
rect -1520 316 -1480 364
rect -1520 284 -1516 316
rect -1484 284 -1480 316
rect -1520 236 -1480 284
rect -1520 204 -1516 236
rect -1484 204 -1480 236
rect -1520 156 -1480 204
rect -1520 124 -1516 156
rect -1484 124 -1480 156
rect -1520 76 -1480 124
rect -1520 44 -1516 76
rect -1484 44 -1480 76
rect -1520 -4 -1480 44
rect -1520 -36 -1516 -4
rect -1484 -36 -1480 -4
rect -1520 -84 -1480 -36
rect -1520 -116 -1516 -84
rect -1484 -116 -1480 -84
rect -1520 -120 -1480 -116
rect -1440 4795 -1400 5640
rect -1440 4765 -1435 4795
rect -1405 4765 -1400 4795
rect -1440 -120 -1400 4765
rect -1360 5596 -1320 5640
rect -1360 5564 -1356 5596
rect -1324 5564 -1320 5596
rect -1360 5516 -1320 5564
rect -1360 5484 -1356 5516
rect -1324 5484 -1320 5516
rect -1360 5436 -1320 5484
rect -1360 5404 -1356 5436
rect -1324 5404 -1320 5436
rect -1360 5356 -1320 5404
rect -1360 5324 -1356 5356
rect -1324 5324 -1320 5356
rect -1360 5276 -1320 5324
rect -1360 5244 -1356 5276
rect -1324 5244 -1320 5276
rect -1360 5196 -1320 5244
rect -1360 5164 -1356 5196
rect -1324 5164 -1320 5196
rect -1360 5116 -1320 5164
rect -1360 5084 -1356 5116
rect -1324 5084 -1320 5116
rect -1360 5036 -1320 5084
rect -1360 5004 -1356 5036
rect -1324 5004 -1320 5036
rect -1360 4956 -1320 5004
rect -1360 4924 -1356 4956
rect -1324 4924 -1320 4956
rect -1360 4876 -1320 4924
rect -1360 4844 -1356 4876
rect -1324 4844 -1320 4876
rect -1360 4796 -1320 4844
rect -1360 4764 -1356 4796
rect -1324 4764 -1320 4796
rect -1360 4716 -1320 4764
rect -1360 4684 -1356 4716
rect -1324 4684 -1320 4716
rect -1360 4636 -1320 4684
rect -1360 4604 -1356 4636
rect -1324 4604 -1320 4636
rect -1360 4556 -1320 4604
rect -1360 4524 -1356 4556
rect -1324 4524 -1320 4556
rect -1360 4476 -1320 4524
rect -1360 4444 -1356 4476
rect -1324 4444 -1320 4476
rect -1360 4396 -1320 4444
rect -1360 4364 -1356 4396
rect -1324 4364 -1320 4396
rect -1360 4316 -1320 4364
rect -1360 4284 -1356 4316
rect -1324 4284 -1320 4316
rect -1360 4236 -1320 4284
rect -1360 4204 -1356 4236
rect -1324 4204 -1320 4236
rect -1360 4156 -1320 4204
rect -1360 4124 -1356 4156
rect -1324 4124 -1320 4156
rect -1360 4076 -1320 4124
rect -1360 4044 -1356 4076
rect -1324 4044 -1320 4076
rect -1360 3996 -1320 4044
rect -1360 3964 -1356 3996
rect -1324 3964 -1320 3996
rect -1360 3916 -1320 3964
rect -1360 3884 -1356 3916
rect -1324 3884 -1320 3916
rect -1360 3836 -1320 3884
rect -1360 3804 -1356 3836
rect -1324 3804 -1320 3836
rect -1360 3756 -1320 3804
rect -1360 3724 -1356 3756
rect -1324 3724 -1320 3756
rect -1360 3676 -1320 3724
rect -1360 3644 -1356 3676
rect -1324 3644 -1320 3676
rect -1360 3596 -1320 3644
rect -1360 3564 -1356 3596
rect -1324 3564 -1320 3596
rect -1360 3516 -1320 3564
rect -1360 3484 -1356 3516
rect -1324 3484 -1320 3516
rect -1360 3436 -1320 3484
rect -1360 3404 -1356 3436
rect -1324 3404 -1320 3436
rect -1360 3356 -1320 3404
rect -1360 3324 -1356 3356
rect -1324 3324 -1320 3356
rect -1360 3276 -1320 3324
rect -1360 3244 -1356 3276
rect -1324 3244 -1320 3276
rect -1360 3196 -1320 3244
rect -1360 3164 -1356 3196
rect -1324 3164 -1320 3196
rect -1360 3116 -1320 3164
rect -1360 3084 -1356 3116
rect -1324 3084 -1320 3116
rect -1360 3036 -1320 3084
rect -1360 3004 -1356 3036
rect -1324 3004 -1320 3036
rect -1360 2956 -1320 3004
rect -1360 2924 -1356 2956
rect -1324 2924 -1320 2956
rect -1360 2876 -1320 2924
rect -1360 2844 -1356 2876
rect -1324 2844 -1320 2876
rect -1360 2796 -1320 2844
rect -1360 2764 -1356 2796
rect -1324 2764 -1320 2796
rect -1360 2716 -1320 2764
rect -1360 2684 -1356 2716
rect -1324 2684 -1320 2716
rect -1360 2636 -1320 2684
rect -1360 2604 -1356 2636
rect -1324 2604 -1320 2636
rect -1360 2556 -1320 2604
rect -1360 2524 -1356 2556
rect -1324 2524 -1320 2556
rect -1360 2476 -1320 2524
rect -1360 2444 -1356 2476
rect -1324 2444 -1320 2476
rect -1360 2396 -1320 2444
rect -1360 2364 -1356 2396
rect -1324 2364 -1320 2396
rect -1360 2316 -1320 2364
rect -1360 2284 -1356 2316
rect -1324 2284 -1320 2316
rect -1360 2236 -1320 2284
rect -1360 2204 -1356 2236
rect -1324 2204 -1320 2236
rect -1360 2156 -1320 2204
rect -1360 2124 -1356 2156
rect -1324 2124 -1320 2156
rect -1360 2076 -1320 2124
rect -1360 2044 -1356 2076
rect -1324 2044 -1320 2076
rect -1360 1996 -1320 2044
rect -1360 1964 -1356 1996
rect -1324 1964 -1320 1996
rect -1360 1916 -1320 1964
rect -1360 1884 -1356 1916
rect -1324 1884 -1320 1916
rect -1360 1836 -1320 1884
rect -1360 1804 -1356 1836
rect -1324 1804 -1320 1836
rect -1360 1756 -1320 1804
rect -1360 1724 -1356 1756
rect -1324 1724 -1320 1756
rect -1360 1676 -1320 1724
rect -1360 1644 -1356 1676
rect -1324 1644 -1320 1676
rect -1360 1596 -1320 1644
rect -1360 1564 -1356 1596
rect -1324 1564 -1320 1596
rect -1360 1516 -1320 1564
rect -1360 1484 -1356 1516
rect -1324 1484 -1320 1516
rect -1360 1436 -1320 1484
rect -1360 1404 -1356 1436
rect -1324 1404 -1320 1436
rect -1360 1356 -1320 1404
rect -1360 1324 -1356 1356
rect -1324 1324 -1320 1356
rect -1360 1276 -1320 1324
rect -1360 1244 -1356 1276
rect -1324 1244 -1320 1276
rect -1360 1196 -1320 1244
rect -1360 1164 -1356 1196
rect -1324 1164 -1320 1196
rect -1360 1116 -1320 1164
rect -1360 1084 -1356 1116
rect -1324 1084 -1320 1116
rect -1360 1036 -1320 1084
rect -1360 1004 -1356 1036
rect -1324 1004 -1320 1036
rect -1360 956 -1320 1004
rect -1360 924 -1356 956
rect -1324 924 -1320 956
rect -1360 876 -1320 924
rect -1360 844 -1356 876
rect -1324 844 -1320 876
rect -1360 796 -1320 844
rect -1360 764 -1356 796
rect -1324 764 -1320 796
rect -1360 716 -1320 764
rect -1360 684 -1356 716
rect -1324 684 -1320 716
rect -1360 636 -1320 684
rect -1360 604 -1356 636
rect -1324 604 -1320 636
rect -1360 556 -1320 604
rect -1360 524 -1356 556
rect -1324 524 -1320 556
rect -1360 476 -1320 524
rect -1360 444 -1356 476
rect -1324 444 -1320 476
rect -1360 396 -1320 444
rect -1360 364 -1356 396
rect -1324 364 -1320 396
rect -1360 316 -1320 364
rect -1360 284 -1356 316
rect -1324 284 -1320 316
rect -1360 236 -1320 284
rect -1360 204 -1356 236
rect -1324 204 -1320 236
rect -1360 156 -1320 204
rect -1360 124 -1356 156
rect -1324 124 -1320 156
rect -1360 76 -1320 124
rect -1360 44 -1356 76
rect -1324 44 -1320 76
rect -1360 -4 -1320 44
rect -1360 -36 -1356 -4
rect -1324 -36 -1320 -4
rect -1360 -84 -1320 -36
rect -1360 -116 -1356 -84
rect -1324 -116 -1320 -84
rect -1360 -120 -1320 -116
rect -1280 3435 -1240 5640
rect -1280 3405 -1275 3435
rect -1245 3405 -1240 3435
rect -1280 2635 -1240 3405
rect -1280 2605 -1275 2635
rect -1245 2605 -1240 2635
rect -1280 -120 -1240 2605
rect -1200 5596 -1160 5640
rect -1200 5564 -1196 5596
rect -1164 5564 -1160 5596
rect -1200 5516 -1160 5564
rect -1200 5484 -1196 5516
rect -1164 5484 -1160 5516
rect -1200 5436 -1160 5484
rect -1200 5404 -1196 5436
rect -1164 5404 -1160 5436
rect -1200 5356 -1160 5404
rect -1200 5324 -1196 5356
rect -1164 5324 -1160 5356
rect -1200 5276 -1160 5324
rect -1200 5244 -1196 5276
rect -1164 5244 -1160 5276
rect -1200 5196 -1160 5244
rect -1200 5164 -1196 5196
rect -1164 5164 -1160 5196
rect -1200 5116 -1160 5164
rect -1200 5084 -1196 5116
rect -1164 5084 -1160 5116
rect -1200 5036 -1160 5084
rect -1200 5004 -1196 5036
rect -1164 5004 -1160 5036
rect -1200 4956 -1160 5004
rect -1200 4924 -1196 4956
rect -1164 4924 -1160 4956
rect -1200 4876 -1160 4924
rect -1200 4844 -1196 4876
rect -1164 4844 -1160 4876
rect -1200 4796 -1160 4844
rect -1200 4764 -1196 4796
rect -1164 4764 -1160 4796
rect -1200 4716 -1160 4764
rect -1200 4684 -1196 4716
rect -1164 4684 -1160 4716
rect -1200 4636 -1160 4684
rect -1200 4604 -1196 4636
rect -1164 4604 -1160 4636
rect -1200 4556 -1160 4604
rect -1200 4524 -1196 4556
rect -1164 4524 -1160 4556
rect -1200 4476 -1160 4524
rect -1200 4444 -1196 4476
rect -1164 4444 -1160 4476
rect -1200 4396 -1160 4444
rect -1200 4364 -1196 4396
rect -1164 4364 -1160 4396
rect -1200 4316 -1160 4364
rect -1200 4284 -1196 4316
rect -1164 4284 -1160 4316
rect -1200 4236 -1160 4284
rect -1200 4204 -1196 4236
rect -1164 4204 -1160 4236
rect -1200 4156 -1160 4204
rect -1200 4124 -1196 4156
rect -1164 4124 -1160 4156
rect -1200 4076 -1160 4124
rect -1200 4044 -1196 4076
rect -1164 4044 -1160 4076
rect -1200 3996 -1160 4044
rect -1200 3964 -1196 3996
rect -1164 3964 -1160 3996
rect -1200 3916 -1160 3964
rect -1200 3884 -1196 3916
rect -1164 3884 -1160 3916
rect -1200 3836 -1160 3884
rect -1200 3804 -1196 3836
rect -1164 3804 -1160 3836
rect -1200 3756 -1160 3804
rect -1200 3724 -1196 3756
rect -1164 3724 -1160 3756
rect -1200 3676 -1160 3724
rect -1200 3644 -1196 3676
rect -1164 3644 -1160 3676
rect -1200 3596 -1160 3644
rect -1200 3564 -1196 3596
rect -1164 3564 -1160 3596
rect -1200 3516 -1160 3564
rect -1200 3484 -1196 3516
rect -1164 3484 -1160 3516
rect -1200 3436 -1160 3484
rect -1200 3404 -1196 3436
rect -1164 3404 -1160 3436
rect -1200 3356 -1160 3404
rect -1200 3324 -1196 3356
rect -1164 3324 -1160 3356
rect -1200 3276 -1160 3324
rect -1200 3244 -1196 3276
rect -1164 3244 -1160 3276
rect -1200 3196 -1160 3244
rect -1200 3164 -1196 3196
rect -1164 3164 -1160 3196
rect -1200 3116 -1160 3164
rect -1200 3084 -1196 3116
rect -1164 3084 -1160 3116
rect -1200 3036 -1160 3084
rect -1200 3004 -1196 3036
rect -1164 3004 -1160 3036
rect -1200 2956 -1160 3004
rect -1200 2924 -1196 2956
rect -1164 2924 -1160 2956
rect -1200 2876 -1160 2924
rect -1200 2844 -1196 2876
rect -1164 2844 -1160 2876
rect -1200 2796 -1160 2844
rect -1200 2764 -1196 2796
rect -1164 2764 -1160 2796
rect -1200 2716 -1160 2764
rect -1200 2684 -1196 2716
rect -1164 2684 -1160 2716
rect -1200 2636 -1160 2684
rect -1200 2604 -1196 2636
rect -1164 2604 -1160 2636
rect -1200 2556 -1160 2604
rect -1200 2524 -1196 2556
rect -1164 2524 -1160 2556
rect -1200 2476 -1160 2524
rect -1200 2444 -1196 2476
rect -1164 2444 -1160 2476
rect -1200 2396 -1160 2444
rect -1200 2364 -1196 2396
rect -1164 2364 -1160 2396
rect -1200 2316 -1160 2364
rect -1200 2284 -1196 2316
rect -1164 2284 -1160 2316
rect -1200 2236 -1160 2284
rect -1200 2204 -1196 2236
rect -1164 2204 -1160 2236
rect -1200 2156 -1160 2204
rect -1200 2124 -1196 2156
rect -1164 2124 -1160 2156
rect -1200 2076 -1160 2124
rect -1200 2044 -1196 2076
rect -1164 2044 -1160 2076
rect -1200 1996 -1160 2044
rect -1200 1964 -1196 1996
rect -1164 1964 -1160 1996
rect -1200 1916 -1160 1964
rect -1200 1884 -1196 1916
rect -1164 1884 -1160 1916
rect -1200 1836 -1160 1884
rect -1200 1804 -1196 1836
rect -1164 1804 -1160 1836
rect -1200 1756 -1160 1804
rect -1200 1724 -1196 1756
rect -1164 1724 -1160 1756
rect -1200 1676 -1160 1724
rect -1200 1644 -1196 1676
rect -1164 1644 -1160 1676
rect -1200 1596 -1160 1644
rect -1200 1564 -1196 1596
rect -1164 1564 -1160 1596
rect -1200 1516 -1160 1564
rect -1200 1484 -1196 1516
rect -1164 1484 -1160 1516
rect -1200 1436 -1160 1484
rect -1200 1404 -1196 1436
rect -1164 1404 -1160 1436
rect -1200 1356 -1160 1404
rect -1200 1324 -1196 1356
rect -1164 1324 -1160 1356
rect -1200 1276 -1160 1324
rect -1200 1244 -1196 1276
rect -1164 1244 -1160 1276
rect -1200 1196 -1160 1244
rect -1200 1164 -1196 1196
rect -1164 1164 -1160 1196
rect -1200 1116 -1160 1164
rect -1200 1084 -1196 1116
rect -1164 1084 -1160 1116
rect -1200 1036 -1160 1084
rect -1200 1004 -1196 1036
rect -1164 1004 -1160 1036
rect -1200 956 -1160 1004
rect -1200 924 -1196 956
rect -1164 924 -1160 956
rect -1200 876 -1160 924
rect -1200 844 -1196 876
rect -1164 844 -1160 876
rect -1200 796 -1160 844
rect -1200 764 -1196 796
rect -1164 764 -1160 796
rect -1200 716 -1160 764
rect -1200 684 -1196 716
rect -1164 684 -1160 716
rect -1200 636 -1160 684
rect -1200 604 -1196 636
rect -1164 604 -1160 636
rect -1200 556 -1160 604
rect -1200 524 -1196 556
rect -1164 524 -1160 556
rect -1200 476 -1160 524
rect -1200 444 -1196 476
rect -1164 444 -1160 476
rect -1200 396 -1160 444
rect -1200 364 -1196 396
rect -1164 364 -1160 396
rect -1200 316 -1160 364
rect -1200 284 -1196 316
rect -1164 284 -1160 316
rect -1200 236 -1160 284
rect -1200 204 -1196 236
rect -1164 204 -1160 236
rect -1200 156 -1160 204
rect -1200 124 -1196 156
rect -1164 124 -1160 156
rect -1200 76 -1160 124
rect -1200 44 -1196 76
rect -1164 44 -1160 76
rect -1200 -4 -1160 44
rect -1200 -36 -1196 -4
rect -1164 -36 -1160 -4
rect -1200 -84 -1160 -36
rect -1200 -116 -1196 -84
rect -1164 -116 -1160 -84
rect -1200 -120 -1160 -116
rect -1120 4955 -1080 5640
rect -1120 4925 -1115 4955
rect -1085 4925 -1080 4955
rect -1120 3035 -1080 4925
rect -1120 3005 -1115 3035
rect -1085 3005 -1080 3035
rect -1120 1115 -1080 3005
rect -1120 1085 -1115 1115
rect -1085 1085 -1080 1115
rect -1120 -120 -1080 1085
rect -1040 5596 -1000 5640
rect -1040 5564 -1036 5596
rect -1004 5564 -1000 5596
rect -1040 5516 -1000 5564
rect -1040 5484 -1036 5516
rect -1004 5484 -1000 5516
rect -1040 5436 -1000 5484
rect -1040 5404 -1036 5436
rect -1004 5404 -1000 5436
rect -1040 5356 -1000 5404
rect -1040 5324 -1036 5356
rect -1004 5324 -1000 5356
rect -1040 5276 -1000 5324
rect -1040 5244 -1036 5276
rect -1004 5244 -1000 5276
rect -1040 5196 -1000 5244
rect -1040 5164 -1036 5196
rect -1004 5164 -1000 5196
rect -1040 5116 -1000 5164
rect -1040 5084 -1036 5116
rect -1004 5084 -1000 5116
rect -1040 5036 -1000 5084
rect -1040 5004 -1036 5036
rect -1004 5004 -1000 5036
rect -1040 4956 -1000 5004
rect -1040 4924 -1036 4956
rect -1004 4924 -1000 4956
rect -1040 4876 -1000 4924
rect -1040 4844 -1036 4876
rect -1004 4844 -1000 4876
rect -1040 4796 -1000 4844
rect -1040 4764 -1036 4796
rect -1004 4764 -1000 4796
rect -1040 4716 -1000 4764
rect -1040 4684 -1036 4716
rect -1004 4684 -1000 4716
rect -1040 4636 -1000 4684
rect -1040 4604 -1036 4636
rect -1004 4604 -1000 4636
rect -1040 4556 -1000 4604
rect -1040 4524 -1036 4556
rect -1004 4524 -1000 4556
rect -1040 4476 -1000 4524
rect -1040 4444 -1036 4476
rect -1004 4444 -1000 4476
rect -1040 4396 -1000 4444
rect -1040 4364 -1036 4396
rect -1004 4364 -1000 4396
rect -1040 4316 -1000 4364
rect -1040 4284 -1036 4316
rect -1004 4284 -1000 4316
rect -1040 4236 -1000 4284
rect -1040 4204 -1036 4236
rect -1004 4204 -1000 4236
rect -1040 4156 -1000 4204
rect -1040 4124 -1036 4156
rect -1004 4124 -1000 4156
rect -1040 4076 -1000 4124
rect -1040 4044 -1036 4076
rect -1004 4044 -1000 4076
rect -1040 3996 -1000 4044
rect -1040 3964 -1036 3996
rect -1004 3964 -1000 3996
rect -1040 3916 -1000 3964
rect -1040 3884 -1036 3916
rect -1004 3884 -1000 3916
rect -1040 3836 -1000 3884
rect -1040 3804 -1036 3836
rect -1004 3804 -1000 3836
rect -1040 3756 -1000 3804
rect -1040 3724 -1036 3756
rect -1004 3724 -1000 3756
rect -1040 3676 -1000 3724
rect -1040 3644 -1036 3676
rect -1004 3644 -1000 3676
rect -1040 3596 -1000 3644
rect -1040 3564 -1036 3596
rect -1004 3564 -1000 3596
rect -1040 3516 -1000 3564
rect -1040 3484 -1036 3516
rect -1004 3484 -1000 3516
rect -1040 3436 -1000 3484
rect -1040 3404 -1036 3436
rect -1004 3404 -1000 3436
rect -1040 3356 -1000 3404
rect -1040 3324 -1036 3356
rect -1004 3324 -1000 3356
rect -1040 3276 -1000 3324
rect -1040 3244 -1036 3276
rect -1004 3244 -1000 3276
rect -1040 3196 -1000 3244
rect -1040 3164 -1036 3196
rect -1004 3164 -1000 3196
rect -1040 3116 -1000 3164
rect -1040 3084 -1036 3116
rect -1004 3084 -1000 3116
rect -1040 3036 -1000 3084
rect -1040 3004 -1036 3036
rect -1004 3004 -1000 3036
rect -1040 2956 -1000 3004
rect -1040 2924 -1036 2956
rect -1004 2924 -1000 2956
rect -1040 2876 -1000 2924
rect -1040 2844 -1036 2876
rect -1004 2844 -1000 2876
rect -1040 2796 -1000 2844
rect -1040 2764 -1036 2796
rect -1004 2764 -1000 2796
rect -1040 2716 -1000 2764
rect -1040 2684 -1036 2716
rect -1004 2684 -1000 2716
rect -1040 2636 -1000 2684
rect -1040 2604 -1036 2636
rect -1004 2604 -1000 2636
rect -1040 2556 -1000 2604
rect -1040 2524 -1036 2556
rect -1004 2524 -1000 2556
rect -1040 2476 -1000 2524
rect -1040 2444 -1036 2476
rect -1004 2444 -1000 2476
rect -1040 2396 -1000 2444
rect -1040 2364 -1036 2396
rect -1004 2364 -1000 2396
rect -1040 2316 -1000 2364
rect -1040 2284 -1036 2316
rect -1004 2284 -1000 2316
rect -1040 2236 -1000 2284
rect -1040 2204 -1036 2236
rect -1004 2204 -1000 2236
rect -1040 2156 -1000 2204
rect -1040 2124 -1036 2156
rect -1004 2124 -1000 2156
rect -1040 2076 -1000 2124
rect -1040 2044 -1036 2076
rect -1004 2044 -1000 2076
rect -1040 1996 -1000 2044
rect -1040 1964 -1036 1996
rect -1004 1964 -1000 1996
rect -1040 1916 -1000 1964
rect -1040 1884 -1036 1916
rect -1004 1884 -1000 1916
rect -1040 1836 -1000 1884
rect -1040 1804 -1036 1836
rect -1004 1804 -1000 1836
rect -1040 1756 -1000 1804
rect -1040 1724 -1036 1756
rect -1004 1724 -1000 1756
rect -1040 1676 -1000 1724
rect -1040 1644 -1036 1676
rect -1004 1644 -1000 1676
rect -1040 1596 -1000 1644
rect -1040 1564 -1036 1596
rect -1004 1564 -1000 1596
rect -1040 1516 -1000 1564
rect -1040 1484 -1036 1516
rect -1004 1484 -1000 1516
rect -1040 1436 -1000 1484
rect -1040 1404 -1036 1436
rect -1004 1404 -1000 1436
rect -1040 1356 -1000 1404
rect -1040 1324 -1036 1356
rect -1004 1324 -1000 1356
rect -1040 1276 -1000 1324
rect -1040 1244 -1036 1276
rect -1004 1244 -1000 1276
rect -1040 1196 -1000 1244
rect -1040 1164 -1036 1196
rect -1004 1164 -1000 1196
rect -1040 1116 -1000 1164
rect -1040 1084 -1036 1116
rect -1004 1084 -1000 1116
rect -1040 1036 -1000 1084
rect -1040 1004 -1036 1036
rect -1004 1004 -1000 1036
rect -1040 956 -1000 1004
rect -1040 924 -1036 956
rect -1004 924 -1000 956
rect -1040 876 -1000 924
rect -1040 844 -1036 876
rect -1004 844 -1000 876
rect -1040 796 -1000 844
rect -1040 764 -1036 796
rect -1004 764 -1000 796
rect -1040 716 -1000 764
rect -1040 684 -1036 716
rect -1004 684 -1000 716
rect -1040 636 -1000 684
rect -1040 604 -1036 636
rect -1004 604 -1000 636
rect -1040 556 -1000 604
rect -1040 524 -1036 556
rect -1004 524 -1000 556
rect -1040 476 -1000 524
rect -1040 444 -1036 476
rect -1004 444 -1000 476
rect -1040 396 -1000 444
rect -1040 364 -1036 396
rect -1004 364 -1000 396
rect -1040 316 -1000 364
rect -1040 284 -1036 316
rect -1004 284 -1000 316
rect -1040 236 -1000 284
rect -1040 204 -1036 236
rect -1004 204 -1000 236
rect -1040 156 -1000 204
rect -1040 124 -1036 156
rect -1004 124 -1000 156
rect -1040 76 -1000 124
rect -1040 44 -1036 76
rect -1004 44 -1000 76
rect -1040 -4 -1000 44
rect -1040 -36 -1036 -4
rect -1004 -36 -1000 -4
rect -1040 -84 -1000 -36
rect -1040 -116 -1036 -84
rect -1004 -116 -1000 -84
rect -1040 -120 -1000 -116
rect -960 5355 -920 5640
rect -960 5325 -955 5355
rect -925 5325 -920 5355
rect -960 4555 -920 5325
rect -960 4525 -955 4555
rect -925 4525 -920 4555
rect -960 2875 -920 4525
rect -960 2845 -955 2875
rect -925 2845 -920 2875
rect -960 1515 -920 2845
rect -960 1485 -955 1515
rect -925 1485 -920 1515
rect -960 -120 -920 1485
rect -880 5596 -840 5640
rect -880 5564 -876 5596
rect -844 5564 -840 5596
rect -880 5516 -840 5564
rect 4880 5596 4920 5600
rect 4880 5564 4884 5596
rect 4916 5564 4920 5596
rect -880 5484 -876 5516
rect -844 5484 -840 5516
rect -880 5436 -840 5484
rect -880 5404 -876 5436
rect -844 5404 -840 5436
rect -880 5356 -840 5404
rect -880 5324 -876 5356
rect -844 5324 -840 5356
rect -880 5276 -840 5324
rect -880 5244 -876 5276
rect -844 5244 -840 5276
rect -880 5196 -840 5244
rect -880 5164 -876 5196
rect -844 5164 -840 5196
rect -880 5116 -840 5164
rect -880 5084 -876 5116
rect -844 5084 -840 5116
rect -880 5036 -840 5084
rect -880 5004 -876 5036
rect -844 5004 -840 5036
rect -880 4956 -840 5004
rect -880 4924 -876 4956
rect -844 4924 -840 4956
rect -880 4876 -840 4924
rect -880 4844 -876 4876
rect -844 4844 -840 4876
rect -880 4796 -840 4844
rect -880 4764 -876 4796
rect -844 4764 -840 4796
rect -880 4716 -840 4764
rect -880 4684 -876 4716
rect -844 4684 -840 4716
rect -880 4636 -840 4684
rect -880 4604 -876 4636
rect -844 4604 -840 4636
rect -880 4556 -840 4604
rect -880 4524 -876 4556
rect -844 4524 -840 4556
rect -880 4476 -840 4524
rect -880 4444 -876 4476
rect -844 4444 -840 4476
rect -880 4396 -840 4444
rect -800 5516 -760 5520
rect -800 5484 -796 5516
rect -764 5484 -760 5516
rect -800 5436 -760 5484
rect -800 5404 -796 5436
rect -764 5404 -760 5436
rect -800 5356 -760 5404
rect -800 5324 -796 5356
rect -764 5324 -760 5356
rect -800 5276 -760 5324
rect -800 5244 -796 5276
rect -764 5244 -760 5276
rect -800 5196 -760 5244
rect -800 5164 -796 5196
rect -764 5164 -760 5196
rect -800 5116 -760 5164
rect -800 5084 -796 5116
rect -764 5084 -760 5116
rect -800 5036 -760 5084
rect -800 5004 -796 5036
rect -764 5004 -760 5036
rect -800 4956 -760 5004
rect -800 4924 -796 4956
rect -764 4924 -760 4956
rect -800 4876 -760 4924
rect -800 4844 -796 4876
rect -764 4844 -760 4876
rect -800 4796 -760 4844
rect -800 4764 -796 4796
rect -764 4764 -760 4796
rect -800 4716 -760 4764
rect -800 4684 -796 4716
rect -764 4684 -760 4716
rect -800 4636 -760 4684
rect -800 4604 -796 4636
rect -764 4604 -760 4636
rect -800 4556 -760 4604
rect -800 4524 -796 4556
rect -764 4524 -760 4556
rect -800 4476 -760 4524
rect -800 4444 -796 4476
rect -764 4444 -760 4476
rect -800 4440 -760 4444
rect -720 5516 -680 5520
rect -720 5484 -716 5516
rect -684 5484 -680 5516
rect -720 5436 -680 5484
rect -720 5404 -716 5436
rect -684 5404 -680 5436
rect -720 5356 -680 5404
rect -720 5324 -716 5356
rect -684 5324 -680 5356
rect -720 5276 -680 5324
rect -720 5244 -716 5276
rect -684 5244 -680 5276
rect -720 5196 -680 5244
rect -720 5164 -716 5196
rect -684 5164 -680 5196
rect -720 5116 -680 5164
rect -720 5084 -716 5116
rect -684 5084 -680 5116
rect -720 5036 -680 5084
rect -720 5004 -716 5036
rect -684 5004 -680 5036
rect -720 4956 -680 5004
rect -720 4924 -716 4956
rect -684 4924 -680 4956
rect -720 4876 -680 4924
rect -720 4844 -716 4876
rect -684 4844 -680 4876
rect -720 4796 -680 4844
rect -720 4764 -716 4796
rect -684 4764 -680 4796
rect -720 4716 -680 4764
rect -720 4684 -716 4716
rect -684 4684 -680 4716
rect -720 4636 -680 4684
rect -720 4604 -716 4636
rect -684 4604 -680 4636
rect -720 4556 -680 4604
rect -720 4524 -716 4556
rect -684 4524 -680 4556
rect -720 4476 -680 4524
rect -720 4444 -716 4476
rect -684 4444 -680 4476
rect -720 4440 -680 4444
rect -640 5516 -600 5520
rect -640 5484 -636 5516
rect -604 5484 -600 5516
rect -640 5436 -600 5484
rect -640 5404 -636 5436
rect -604 5404 -600 5436
rect -640 5356 -600 5404
rect -640 5324 -636 5356
rect -604 5324 -600 5356
rect -640 5276 -600 5324
rect -640 5244 -636 5276
rect -604 5244 -600 5276
rect -640 5196 -600 5244
rect -640 5164 -636 5196
rect -604 5164 -600 5196
rect -640 5116 -600 5164
rect -640 5084 -636 5116
rect -604 5084 -600 5116
rect -640 5036 -600 5084
rect -640 5004 -636 5036
rect -604 5004 -600 5036
rect -640 4956 -600 5004
rect -640 4924 -636 4956
rect -604 4924 -600 4956
rect -640 4876 -600 4924
rect -640 4844 -636 4876
rect -604 4844 -600 4876
rect -640 4796 -600 4844
rect -640 4764 -636 4796
rect -604 4764 -600 4796
rect -640 4716 -600 4764
rect -640 4684 -636 4716
rect -604 4684 -600 4716
rect -640 4636 -600 4684
rect -640 4604 -636 4636
rect -604 4604 -600 4636
rect -640 4556 -600 4604
rect -640 4524 -636 4556
rect -604 4524 -600 4556
rect -640 4476 -600 4524
rect -640 4444 -636 4476
rect -604 4444 -600 4476
rect -640 4440 -600 4444
rect -560 5516 -520 5520
rect -560 5484 -556 5516
rect -524 5484 -520 5516
rect -560 5436 -520 5484
rect -560 5404 -556 5436
rect -524 5404 -520 5436
rect -560 5356 -520 5404
rect -560 5324 -556 5356
rect -524 5324 -520 5356
rect -560 5276 -520 5324
rect -560 5244 -556 5276
rect -524 5244 -520 5276
rect -560 5196 -520 5244
rect -560 5164 -556 5196
rect -524 5164 -520 5196
rect -560 5116 -520 5164
rect -560 5084 -556 5116
rect -524 5084 -520 5116
rect -560 5036 -520 5084
rect -560 5004 -556 5036
rect -524 5004 -520 5036
rect -560 4956 -520 5004
rect -560 4924 -556 4956
rect -524 4924 -520 4956
rect -560 4876 -520 4924
rect -560 4844 -556 4876
rect -524 4844 -520 4876
rect -560 4796 -520 4844
rect -560 4764 -556 4796
rect -524 4764 -520 4796
rect -560 4716 -520 4764
rect -560 4684 -556 4716
rect -524 4684 -520 4716
rect -560 4636 -520 4684
rect -560 4604 -556 4636
rect -524 4604 -520 4636
rect -560 4556 -520 4604
rect -560 4524 -556 4556
rect -524 4524 -520 4556
rect -560 4476 -520 4524
rect -560 4444 -556 4476
rect -524 4444 -520 4476
rect -560 4440 -520 4444
rect -480 5516 -440 5520
rect -480 5484 -476 5516
rect -444 5484 -440 5516
rect -480 5436 -440 5484
rect -480 5404 -476 5436
rect -444 5404 -440 5436
rect -480 5356 -440 5404
rect -480 5324 -476 5356
rect -444 5324 -440 5356
rect -480 5276 -440 5324
rect -480 5244 -476 5276
rect -444 5244 -440 5276
rect -480 5196 -440 5244
rect -480 5164 -476 5196
rect -444 5164 -440 5196
rect -480 5116 -440 5164
rect -480 5084 -476 5116
rect -444 5084 -440 5116
rect -480 5036 -440 5084
rect -480 5004 -476 5036
rect -444 5004 -440 5036
rect -480 4956 -440 5004
rect -480 4924 -476 4956
rect -444 4924 -440 4956
rect -480 4876 -440 4924
rect -480 4844 -476 4876
rect -444 4844 -440 4876
rect -480 4796 -440 4844
rect -480 4764 -476 4796
rect -444 4764 -440 4796
rect -480 4716 -440 4764
rect -480 4684 -476 4716
rect -444 4684 -440 4716
rect -480 4636 -440 4684
rect -480 4604 -476 4636
rect -444 4604 -440 4636
rect -480 4556 -440 4604
rect -480 4524 -476 4556
rect -444 4524 -440 4556
rect -480 4476 -440 4524
rect -480 4444 -476 4476
rect -444 4444 -440 4476
rect -480 4440 -440 4444
rect -400 5516 -360 5520
rect -400 5484 -396 5516
rect -364 5484 -360 5516
rect -400 5436 -360 5484
rect -400 5404 -396 5436
rect -364 5404 -360 5436
rect -400 5356 -360 5404
rect -400 5324 -396 5356
rect -364 5324 -360 5356
rect -400 5276 -360 5324
rect -400 5244 -396 5276
rect -364 5244 -360 5276
rect -400 5196 -360 5244
rect -400 5164 -396 5196
rect -364 5164 -360 5196
rect -400 5116 -360 5164
rect -400 5084 -396 5116
rect -364 5084 -360 5116
rect -400 5036 -360 5084
rect -400 5004 -396 5036
rect -364 5004 -360 5036
rect -400 4956 -360 5004
rect -400 4924 -396 4956
rect -364 4924 -360 4956
rect -400 4876 -360 4924
rect -400 4844 -396 4876
rect -364 4844 -360 4876
rect -400 4796 -360 4844
rect -400 4764 -396 4796
rect -364 4764 -360 4796
rect -400 4716 -360 4764
rect -400 4684 -396 4716
rect -364 4684 -360 4716
rect -400 4636 -360 4684
rect -400 4604 -396 4636
rect -364 4604 -360 4636
rect -400 4556 -360 4604
rect -400 4524 -396 4556
rect -364 4524 -360 4556
rect -400 4476 -360 4524
rect -400 4444 -396 4476
rect -364 4444 -360 4476
rect -400 4440 -360 4444
rect -320 5516 -280 5520
rect -320 5484 -316 5516
rect -284 5484 -280 5516
rect -320 5436 -280 5484
rect -320 5404 -316 5436
rect -284 5404 -280 5436
rect -320 5356 -280 5404
rect -320 5324 -316 5356
rect -284 5324 -280 5356
rect -320 5276 -280 5324
rect -320 5244 -316 5276
rect -284 5244 -280 5276
rect -320 5196 -280 5244
rect -320 5164 -316 5196
rect -284 5164 -280 5196
rect -320 5116 -280 5164
rect -320 5084 -316 5116
rect -284 5084 -280 5116
rect -320 5036 -280 5084
rect -320 5004 -316 5036
rect -284 5004 -280 5036
rect -320 4956 -280 5004
rect -320 4924 -316 4956
rect -284 4924 -280 4956
rect -320 4876 -280 4924
rect -320 4844 -316 4876
rect -284 4844 -280 4876
rect -320 4796 -280 4844
rect -320 4764 -316 4796
rect -284 4764 -280 4796
rect -320 4716 -280 4764
rect -320 4684 -316 4716
rect -284 4684 -280 4716
rect -320 4636 -280 4684
rect -320 4604 -316 4636
rect -284 4604 -280 4636
rect -320 4556 -280 4604
rect -320 4524 -316 4556
rect -284 4524 -280 4556
rect -320 4476 -280 4524
rect -320 4444 -316 4476
rect -284 4444 -280 4476
rect -320 4440 -280 4444
rect -240 5516 -200 5520
rect -240 5484 -236 5516
rect -204 5484 -200 5516
rect -240 5436 -200 5484
rect -240 5404 -236 5436
rect -204 5404 -200 5436
rect -240 5356 -200 5404
rect -240 5324 -236 5356
rect -204 5324 -200 5356
rect -240 5276 -200 5324
rect -240 5244 -236 5276
rect -204 5244 -200 5276
rect -240 5196 -200 5244
rect -240 5164 -236 5196
rect -204 5164 -200 5196
rect -240 5116 -200 5164
rect -240 5084 -236 5116
rect -204 5084 -200 5116
rect -240 5036 -200 5084
rect -240 5004 -236 5036
rect -204 5004 -200 5036
rect -240 4956 -200 5004
rect -240 4924 -236 4956
rect -204 4924 -200 4956
rect -240 4876 -200 4924
rect -240 4844 -236 4876
rect -204 4844 -200 4876
rect -240 4796 -200 4844
rect -240 4764 -236 4796
rect -204 4764 -200 4796
rect -240 4716 -200 4764
rect -240 4684 -236 4716
rect -204 4684 -200 4716
rect -240 4636 -200 4684
rect -240 4604 -236 4636
rect -204 4604 -200 4636
rect -240 4556 -200 4604
rect -240 4524 -236 4556
rect -204 4524 -200 4556
rect -240 4476 -200 4524
rect -240 4444 -236 4476
rect -204 4444 -200 4476
rect -240 4440 -200 4444
rect -160 5516 -120 5520
rect -160 5484 -156 5516
rect -124 5484 -120 5516
rect -160 5436 -120 5484
rect -160 5404 -156 5436
rect -124 5404 -120 5436
rect -160 5356 -120 5404
rect -160 5324 -156 5356
rect -124 5324 -120 5356
rect -160 5276 -120 5324
rect -160 5244 -156 5276
rect -124 5244 -120 5276
rect -160 5196 -120 5244
rect -160 5164 -156 5196
rect -124 5164 -120 5196
rect -160 5116 -120 5164
rect -160 5084 -156 5116
rect -124 5084 -120 5116
rect -160 5036 -120 5084
rect -160 5004 -156 5036
rect -124 5004 -120 5036
rect -160 4956 -120 5004
rect -160 4924 -156 4956
rect -124 4924 -120 4956
rect -160 4876 -120 4924
rect -160 4844 -156 4876
rect -124 4844 -120 4876
rect -160 4796 -120 4844
rect -160 4764 -156 4796
rect -124 4764 -120 4796
rect -160 4716 -120 4764
rect -160 4684 -156 4716
rect -124 4684 -120 4716
rect -160 4636 -120 4684
rect -160 4604 -156 4636
rect -124 4604 -120 4636
rect -160 4556 -120 4604
rect -160 4524 -156 4556
rect -124 4524 -120 4556
rect -160 4476 -120 4524
rect -160 4444 -156 4476
rect -124 4444 -120 4476
rect -160 4440 -120 4444
rect -80 5516 -40 5520
rect -80 5484 -76 5516
rect -44 5484 -40 5516
rect -80 5436 -40 5484
rect -80 5404 -76 5436
rect -44 5404 -40 5436
rect -80 5356 -40 5404
rect -80 5324 -76 5356
rect -44 5324 -40 5356
rect -80 5276 -40 5324
rect -80 5244 -76 5276
rect -44 5244 -40 5276
rect -80 5196 -40 5244
rect -80 5164 -76 5196
rect -44 5164 -40 5196
rect -80 5116 -40 5164
rect -80 5084 -76 5116
rect -44 5084 -40 5116
rect -80 5036 -40 5084
rect -80 5004 -76 5036
rect -44 5004 -40 5036
rect -80 4956 -40 5004
rect -80 4924 -76 4956
rect -44 4924 -40 4956
rect -80 4876 -40 4924
rect -80 4844 -76 4876
rect -44 4844 -40 4876
rect -80 4796 -40 4844
rect -80 4764 -76 4796
rect -44 4764 -40 4796
rect -80 4716 -40 4764
rect -80 4684 -76 4716
rect -44 4684 -40 4716
rect -80 4636 -40 4684
rect -80 4604 -76 4636
rect -44 4604 -40 4636
rect -80 4556 -40 4604
rect -80 4524 -76 4556
rect -44 4524 -40 4556
rect -80 4476 -40 4524
rect -80 4444 -76 4476
rect -44 4444 -40 4476
rect -80 4440 -40 4444
rect 0 5516 40 5520
rect 0 5484 4 5516
rect 36 5484 40 5516
rect 0 5436 40 5484
rect 0 5404 4 5436
rect 36 5404 40 5436
rect 0 5356 40 5404
rect 0 5324 4 5356
rect 36 5324 40 5356
rect 0 5276 40 5324
rect 0 5244 4 5276
rect 36 5244 40 5276
rect 0 5196 40 5244
rect 0 5164 4 5196
rect 36 5164 40 5196
rect 0 5116 40 5164
rect 0 5084 4 5116
rect 36 5084 40 5116
rect 0 5036 40 5084
rect 0 5004 4 5036
rect 36 5004 40 5036
rect 0 4956 40 5004
rect 0 4924 4 4956
rect 36 4924 40 4956
rect 0 4876 40 4924
rect 0 4844 4 4876
rect 36 4844 40 4876
rect 0 4796 40 4844
rect 0 4764 4 4796
rect 36 4764 40 4796
rect 0 4716 40 4764
rect 0 4684 4 4716
rect 36 4684 40 4716
rect 0 4636 40 4684
rect 0 4604 4 4636
rect 36 4604 40 4636
rect 0 4556 40 4604
rect 0 4524 4 4556
rect 36 4524 40 4556
rect 0 4476 40 4524
rect 0 4444 4 4476
rect 36 4444 40 4476
rect 0 4440 40 4444
rect 80 5516 120 5520
rect 80 5484 84 5516
rect 116 5484 120 5516
rect 80 5436 120 5484
rect 80 5404 84 5436
rect 116 5404 120 5436
rect 80 5356 120 5404
rect 80 5324 84 5356
rect 116 5324 120 5356
rect 80 5276 120 5324
rect 80 5244 84 5276
rect 116 5244 120 5276
rect 80 5196 120 5244
rect 80 5164 84 5196
rect 116 5164 120 5196
rect 80 5116 120 5164
rect 80 5084 84 5116
rect 116 5084 120 5116
rect 80 5036 120 5084
rect 80 5004 84 5036
rect 116 5004 120 5036
rect 80 4956 120 5004
rect 80 4924 84 4956
rect 116 4924 120 4956
rect 80 4876 120 4924
rect 80 4844 84 4876
rect 116 4844 120 4876
rect 80 4796 120 4844
rect 80 4764 84 4796
rect 116 4764 120 4796
rect 80 4716 120 4764
rect 80 4684 84 4716
rect 116 4684 120 4716
rect 80 4636 120 4684
rect 80 4604 84 4636
rect 116 4604 120 4636
rect 80 4556 120 4604
rect 80 4524 84 4556
rect 116 4524 120 4556
rect 80 4476 120 4524
rect 80 4444 84 4476
rect 116 4444 120 4476
rect 80 4440 120 4444
rect 160 5516 200 5520
rect 160 5484 164 5516
rect 196 5484 200 5516
rect 160 5436 200 5484
rect 160 5404 164 5436
rect 196 5404 200 5436
rect 160 5356 200 5404
rect 160 5324 164 5356
rect 196 5324 200 5356
rect 160 5276 200 5324
rect 160 5244 164 5276
rect 196 5244 200 5276
rect 160 5196 200 5244
rect 160 5164 164 5196
rect 196 5164 200 5196
rect 160 5116 200 5164
rect 160 5084 164 5116
rect 196 5084 200 5116
rect 160 5036 200 5084
rect 160 5004 164 5036
rect 196 5004 200 5036
rect 160 4956 200 5004
rect 160 4924 164 4956
rect 196 4924 200 4956
rect 160 4876 200 4924
rect 160 4844 164 4876
rect 196 4844 200 4876
rect 160 4796 200 4844
rect 160 4764 164 4796
rect 196 4764 200 4796
rect 160 4716 200 4764
rect 160 4684 164 4716
rect 196 4684 200 4716
rect 160 4636 200 4684
rect 160 4604 164 4636
rect 196 4604 200 4636
rect 160 4556 200 4604
rect 160 4524 164 4556
rect 196 4524 200 4556
rect 160 4476 200 4524
rect 160 4444 164 4476
rect 196 4444 200 4476
rect 160 4440 200 4444
rect 240 5516 280 5520
rect 240 5484 244 5516
rect 276 5484 280 5516
rect 240 5436 280 5484
rect 240 5404 244 5436
rect 276 5404 280 5436
rect 240 5356 280 5404
rect 240 5324 244 5356
rect 276 5324 280 5356
rect 240 5276 280 5324
rect 240 5244 244 5276
rect 276 5244 280 5276
rect 240 5196 280 5244
rect 240 5164 244 5196
rect 276 5164 280 5196
rect 240 5116 280 5164
rect 240 5084 244 5116
rect 276 5084 280 5116
rect 240 5036 280 5084
rect 240 5004 244 5036
rect 276 5004 280 5036
rect 240 4956 280 5004
rect 240 4924 244 4956
rect 276 4924 280 4956
rect 240 4876 280 4924
rect 240 4844 244 4876
rect 276 4844 280 4876
rect 240 4796 280 4844
rect 240 4764 244 4796
rect 276 4764 280 4796
rect 240 4716 280 4764
rect 240 4684 244 4716
rect 276 4684 280 4716
rect 240 4636 280 4684
rect 240 4604 244 4636
rect 276 4604 280 4636
rect 240 4556 280 4604
rect 240 4524 244 4556
rect 276 4524 280 4556
rect 240 4476 280 4524
rect 240 4444 244 4476
rect 276 4444 280 4476
rect 240 4440 280 4444
rect 320 5516 360 5520
rect 320 5484 324 5516
rect 356 5484 360 5516
rect 320 5436 360 5484
rect 320 5404 324 5436
rect 356 5404 360 5436
rect 320 5356 360 5404
rect 320 5324 324 5356
rect 356 5324 360 5356
rect 320 5276 360 5324
rect 320 5244 324 5276
rect 356 5244 360 5276
rect 320 5196 360 5244
rect 320 5164 324 5196
rect 356 5164 360 5196
rect 320 5116 360 5164
rect 320 5084 324 5116
rect 356 5084 360 5116
rect 320 5036 360 5084
rect 320 5004 324 5036
rect 356 5004 360 5036
rect 320 4956 360 5004
rect 320 4924 324 4956
rect 356 4924 360 4956
rect 320 4876 360 4924
rect 320 4844 324 4876
rect 356 4844 360 4876
rect 320 4796 360 4844
rect 320 4764 324 4796
rect 356 4764 360 4796
rect 320 4716 360 4764
rect 320 4684 324 4716
rect 356 4684 360 4716
rect 320 4636 360 4684
rect 320 4604 324 4636
rect 356 4604 360 4636
rect 320 4556 360 4604
rect 320 4524 324 4556
rect 356 4524 360 4556
rect 320 4476 360 4524
rect 320 4444 324 4476
rect 356 4444 360 4476
rect 320 4440 360 4444
rect 400 5516 440 5520
rect 400 5484 404 5516
rect 436 5484 440 5516
rect 400 5436 440 5484
rect 400 5404 404 5436
rect 436 5404 440 5436
rect 400 5356 440 5404
rect 400 5324 404 5356
rect 436 5324 440 5356
rect 400 5276 440 5324
rect 400 5244 404 5276
rect 436 5244 440 5276
rect 400 5196 440 5244
rect 400 5164 404 5196
rect 436 5164 440 5196
rect 400 5116 440 5164
rect 400 5084 404 5116
rect 436 5084 440 5116
rect 400 5036 440 5084
rect 400 5004 404 5036
rect 436 5004 440 5036
rect 400 4956 440 5004
rect 400 4924 404 4956
rect 436 4924 440 4956
rect 400 4876 440 4924
rect 400 4844 404 4876
rect 436 4844 440 4876
rect 400 4796 440 4844
rect 400 4764 404 4796
rect 436 4764 440 4796
rect 400 4716 440 4764
rect 400 4684 404 4716
rect 436 4684 440 4716
rect 400 4636 440 4684
rect 400 4604 404 4636
rect 436 4604 440 4636
rect 400 4556 440 4604
rect 400 4524 404 4556
rect 436 4524 440 4556
rect 400 4476 440 4524
rect 400 4444 404 4476
rect 436 4444 440 4476
rect 400 4440 440 4444
rect 480 5516 520 5520
rect 480 5484 484 5516
rect 516 5484 520 5516
rect 480 5436 520 5484
rect 480 5404 484 5436
rect 516 5404 520 5436
rect 480 5356 520 5404
rect 480 5324 484 5356
rect 516 5324 520 5356
rect 480 5276 520 5324
rect 480 5244 484 5276
rect 516 5244 520 5276
rect 480 5196 520 5244
rect 480 5164 484 5196
rect 516 5164 520 5196
rect 480 5116 520 5164
rect 480 5084 484 5116
rect 516 5084 520 5116
rect 480 5036 520 5084
rect 480 5004 484 5036
rect 516 5004 520 5036
rect 480 4956 520 5004
rect 480 4924 484 4956
rect 516 4924 520 4956
rect 480 4876 520 4924
rect 480 4844 484 4876
rect 516 4844 520 4876
rect 480 4796 520 4844
rect 480 4764 484 4796
rect 516 4764 520 4796
rect 480 4716 520 4764
rect 480 4684 484 4716
rect 516 4684 520 4716
rect 480 4636 520 4684
rect 480 4604 484 4636
rect 516 4604 520 4636
rect 480 4556 520 4604
rect 480 4524 484 4556
rect 516 4524 520 4556
rect 480 4476 520 4524
rect 480 4444 484 4476
rect 516 4444 520 4476
rect 480 4440 520 4444
rect 560 5516 600 5520
rect 560 5484 564 5516
rect 596 5484 600 5516
rect 560 5436 600 5484
rect 560 5404 564 5436
rect 596 5404 600 5436
rect 560 5356 600 5404
rect 560 5324 564 5356
rect 596 5324 600 5356
rect 560 5276 600 5324
rect 560 5244 564 5276
rect 596 5244 600 5276
rect 560 5196 600 5244
rect 560 5164 564 5196
rect 596 5164 600 5196
rect 560 5116 600 5164
rect 560 5084 564 5116
rect 596 5084 600 5116
rect 560 5036 600 5084
rect 560 5004 564 5036
rect 596 5004 600 5036
rect 560 4956 600 5004
rect 560 4924 564 4956
rect 596 4924 600 4956
rect 560 4876 600 4924
rect 560 4844 564 4876
rect 596 4844 600 4876
rect 560 4796 600 4844
rect 560 4764 564 4796
rect 596 4764 600 4796
rect 560 4716 600 4764
rect 560 4684 564 4716
rect 596 4684 600 4716
rect 560 4636 600 4684
rect 560 4604 564 4636
rect 596 4604 600 4636
rect 560 4556 600 4604
rect 560 4524 564 4556
rect 596 4524 600 4556
rect 560 4476 600 4524
rect 560 4444 564 4476
rect 596 4444 600 4476
rect 560 4440 600 4444
rect 640 5516 680 5520
rect 640 5484 644 5516
rect 676 5484 680 5516
rect 640 5436 680 5484
rect 640 5404 644 5436
rect 676 5404 680 5436
rect 640 5356 680 5404
rect 640 5324 644 5356
rect 676 5324 680 5356
rect 640 5276 680 5324
rect 640 5244 644 5276
rect 676 5244 680 5276
rect 640 5196 680 5244
rect 640 5164 644 5196
rect 676 5164 680 5196
rect 640 5116 680 5164
rect 640 5084 644 5116
rect 676 5084 680 5116
rect 640 5036 680 5084
rect 640 5004 644 5036
rect 676 5004 680 5036
rect 640 4956 680 5004
rect 640 4924 644 4956
rect 676 4924 680 4956
rect 640 4876 680 4924
rect 640 4844 644 4876
rect 676 4844 680 4876
rect 640 4796 680 4844
rect 640 4764 644 4796
rect 676 4764 680 4796
rect 640 4716 680 4764
rect 640 4684 644 4716
rect 676 4684 680 4716
rect 640 4636 680 4684
rect 640 4604 644 4636
rect 676 4604 680 4636
rect 640 4556 680 4604
rect 640 4524 644 4556
rect 676 4524 680 4556
rect 640 4476 680 4524
rect 640 4444 644 4476
rect 676 4444 680 4476
rect 640 4440 680 4444
rect 720 5516 760 5520
rect 720 5484 724 5516
rect 756 5484 760 5516
rect 720 5436 760 5484
rect 720 5404 724 5436
rect 756 5404 760 5436
rect 720 5356 760 5404
rect 720 5324 724 5356
rect 756 5324 760 5356
rect 720 5276 760 5324
rect 720 5244 724 5276
rect 756 5244 760 5276
rect 720 5196 760 5244
rect 720 5164 724 5196
rect 756 5164 760 5196
rect 720 5116 760 5164
rect 720 5084 724 5116
rect 756 5084 760 5116
rect 720 5036 760 5084
rect 720 5004 724 5036
rect 756 5004 760 5036
rect 720 4956 760 5004
rect 720 4924 724 4956
rect 756 4924 760 4956
rect 720 4876 760 4924
rect 720 4844 724 4876
rect 756 4844 760 4876
rect 720 4796 760 4844
rect 720 4764 724 4796
rect 756 4764 760 4796
rect 720 4716 760 4764
rect 720 4684 724 4716
rect 756 4684 760 4716
rect 720 4636 760 4684
rect 720 4604 724 4636
rect 756 4604 760 4636
rect 720 4556 760 4604
rect 720 4524 724 4556
rect 756 4524 760 4556
rect 720 4476 760 4524
rect 720 4444 724 4476
rect 756 4444 760 4476
rect 720 4440 760 4444
rect 800 5516 840 5520
rect 800 5484 804 5516
rect 836 5484 840 5516
rect 800 5436 840 5484
rect 800 5404 804 5436
rect 836 5404 840 5436
rect 800 5356 840 5404
rect 800 5324 804 5356
rect 836 5324 840 5356
rect 800 5276 840 5324
rect 800 5244 804 5276
rect 836 5244 840 5276
rect 800 5196 840 5244
rect 800 5164 804 5196
rect 836 5164 840 5196
rect 800 5116 840 5164
rect 800 5084 804 5116
rect 836 5084 840 5116
rect 800 5036 840 5084
rect 800 5004 804 5036
rect 836 5004 840 5036
rect 800 4956 840 5004
rect 800 4924 804 4956
rect 836 4924 840 4956
rect 800 4876 840 4924
rect 800 4844 804 4876
rect 836 4844 840 4876
rect 800 4796 840 4844
rect 800 4764 804 4796
rect 836 4764 840 4796
rect 800 4716 840 4764
rect 800 4684 804 4716
rect 836 4684 840 4716
rect 800 4636 840 4684
rect 800 4604 804 4636
rect 836 4604 840 4636
rect 800 4556 840 4604
rect 800 4524 804 4556
rect 836 4524 840 4556
rect 800 4476 840 4524
rect 800 4444 804 4476
rect 836 4444 840 4476
rect 800 4440 840 4444
rect 880 5516 920 5520
rect 880 5484 884 5516
rect 916 5484 920 5516
rect 880 5436 920 5484
rect 880 5404 884 5436
rect 916 5404 920 5436
rect 880 5356 920 5404
rect 880 5324 884 5356
rect 916 5324 920 5356
rect 880 5276 920 5324
rect 880 5244 884 5276
rect 916 5244 920 5276
rect 880 5196 920 5244
rect 880 5164 884 5196
rect 916 5164 920 5196
rect 880 5116 920 5164
rect 880 5084 884 5116
rect 916 5084 920 5116
rect 880 5036 920 5084
rect 880 5004 884 5036
rect 916 5004 920 5036
rect 880 4956 920 5004
rect 880 4924 884 4956
rect 916 4924 920 4956
rect 880 4876 920 4924
rect 880 4844 884 4876
rect 916 4844 920 4876
rect 880 4796 920 4844
rect 880 4764 884 4796
rect 916 4764 920 4796
rect 880 4716 920 4764
rect 880 4684 884 4716
rect 916 4684 920 4716
rect 880 4636 920 4684
rect 880 4604 884 4636
rect 916 4604 920 4636
rect 880 4556 920 4604
rect 880 4524 884 4556
rect 916 4524 920 4556
rect 880 4476 920 4524
rect 880 4444 884 4476
rect 916 4444 920 4476
rect 880 4440 920 4444
rect 960 5516 1000 5520
rect 960 5484 964 5516
rect 996 5484 1000 5516
rect 960 5436 1000 5484
rect 960 5404 964 5436
rect 996 5404 1000 5436
rect 960 5356 1000 5404
rect 960 5324 964 5356
rect 996 5324 1000 5356
rect 960 5276 1000 5324
rect 960 5244 964 5276
rect 996 5244 1000 5276
rect 960 5196 1000 5244
rect 960 5164 964 5196
rect 996 5164 1000 5196
rect 960 5116 1000 5164
rect 960 5084 964 5116
rect 996 5084 1000 5116
rect 960 5036 1000 5084
rect 960 5004 964 5036
rect 996 5004 1000 5036
rect 960 4956 1000 5004
rect 960 4924 964 4956
rect 996 4924 1000 4956
rect 960 4876 1000 4924
rect 960 4844 964 4876
rect 996 4844 1000 4876
rect 960 4796 1000 4844
rect 960 4764 964 4796
rect 996 4764 1000 4796
rect 960 4716 1000 4764
rect 960 4684 964 4716
rect 996 4684 1000 4716
rect 960 4636 1000 4684
rect 960 4604 964 4636
rect 996 4604 1000 4636
rect 960 4556 1000 4604
rect 960 4524 964 4556
rect 996 4524 1000 4556
rect 960 4476 1000 4524
rect 960 4444 964 4476
rect 996 4444 1000 4476
rect 960 4440 1000 4444
rect 1040 5516 1080 5520
rect 1040 5484 1044 5516
rect 1076 5484 1080 5516
rect 1040 5436 1080 5484
rect 1040 5404 1044 5436
rect 1076 5404 1080 5436
rect 1040 5356 1080 5404
rect 1040 5324 1044 5356
rect 1076 5324 1080 5356
rect 1040 5276 1080 5324
rect 1040 5244 1044 5276
rect 1076 5244 1080 5276
rect 1040 5196 1080 5244
rect 1040 5164 1044 5196
rect 1076 5164 1080 5196
rect 1040 5116 1080 5164
rect 1040 5084 1044 5116
rect 1076 5084 1080 5116
rect 1040 5036 1080 5084
rect 1040 5004 1044 5036
rect 1076 5004 1080 5036
rect 1040 4956 1080 5004
rect 1040 4924 1044 4956
rect 1076 4924 1080 4956
rect 1040 4876 1080 4924
rect 1040 4844 1044 4876
rect 1076 4844 1080 4876
rect 1040 4796 1080 4844
rect 1040 4764 1044 4796
rect 1076 4764 1080 4796
rect 1040 4716 1080 4764
rect 1040 4684 1044 4716
rect 1076 4684 1080 4716
rect 1040 4636 1080 4684
rect 1040 4604 1044 4636
rect 1076 4604 1080 4636
rect 1040 4556 1080 4604
rect 1040 4524 1044 4556
rect 1076 4524 1080 4556
rect 1040 4476 1080 4524
rect 1040 4444 1044 4476
rect 1076 4444 1080 4476
rect 1040 4440 1080 4444
rect 1120 5516 1160 5520
rect 1120 5484 1124 5516
rect 1156 5484 1160 5516
rect 1120 5436 1160 5484
rect 1120 5404 1124 5436
rect 1156 5404 1160 5436
rect 1120 5356 1160 5404
rect 1120 5324 1124 5356
rect 1156 5324 1160 5356
rect 1120 5276 1160 5324
rect 1120 5244 1124 5276
rect 1156 5244 1160 5276
rect 1120 5196 1160 5244
rect 1120 5164 1124 5196
rect 1156 5164 1160 5196
rect 1120 5116 1160 5164
rect 1120 5084 1124 5116
rect 1156 5084 1160 5116
rect 1120 5036 1160 5084
rect 1120 5004 1124 5036
rect 1156 5004 1160 5036
rect 1120 4956 1160 5004
rect 1120 4924 1124 4956
rect 1156 4924 1160 4956
rect 1120 4876 1160 4924
rect 1120 4844 1124 4876
rect 1156 4844 1160 4876
rect 1120 4796 1160 4844
rect 1120 4764 1124 4796
rect 1156 4764 1160 4796
rect 1120 4716 1160 4764
rect 1120 4684 1124 4716
rect 1156 4684 1160 4716
rect 1120 4636 1160 4684
rect 1120 4604 1124 4636
rect 1156 4604 1160 4636
rect 1120 4556 1160 4604
rect 1120 4524 1124 4556
rect 1156 4524 1160 4556
rect 1120 4476 1160 4524
rect 1120 4444 1124 4476
rect 1156 4444 1160 4476
rect 1120 4440 1160 4444
rect 1200 5516 1240 5520
rect 1200 5484 1204 5516
rect 1236 5484 1240 5516
rect 1200 5436 1240 5484
rect 1200 5404 1204 5436
rect 1236 5404 1240 5436
rect 1200 5356 1240 5404
rect 1200 5324 1204 5356
rect 1236 5324 1240 5356
rect 1200 5276 1240 5324
rect 1200 5244 1204 5276
rect 1236 5244 1240 5276
rect 1200 5196 1240 5244
rect 1200 5164 1204 5196
rect 1236 5164 1240 5196
rect 1200 5116 1240 5164
rect 1200 5084 1204 5116
rect 1236 5084 1240 5116
rect 1200 5036 1240 5084
rect 1200 5004 1204 5036
rect 1236 5004 1240 5036
rect 1200 4956 1240 5004
rect 1200 4924 1204 4956
rect 1236 4924 1240 4956
rect 1200 4876 1240 4924
rect 1200 4844 1204 4876
rect 1236 4844 1240 4876
rect 1200 4796 1240 4844
rect 1200 4764 1204 4796
rect 1236 4764 1240 4796
rect 1200 4716 1240 4764
rect 1200 4684 1204 4716
rect 1236 4684 1240 4716
rect 1200 4636 1240 4684
rect 1200 4604 1204 4636
rect 1236 4604 1240 4636
rect 1200 4556 1240 4604
rect 1200 4524 1204 4556
rect 1236 4524 1240 4556
rect 1200 4476 1240 4524
rect 1200 4444 1204 4476
rect 1236 4444 1240 4476
rect 1200 4440 1240 4444
rect 1280 5516 1320 5520
rect 1280 5484 1284 5516
rect 1316 5484 1320 5516
rect 1280 5436 1320 5484
rect 1280 5404 1284 5436
rect 1316 5404 1320 5436
rect 1280 5356 1320 5404
rect 1280 5324 1284 5356
rect 1316 5324 1320 5356
rect 1280 5276 1320 5324
rect 1280 5244 1284 5276
rect 1316 5244 1320 5276
rect 1280 5196 1320 5244
rect 1280 5164 1284 5196
rect 1316 5164 1320 5196
rect 1280 5116 1320 5164
rect 1280 5084 1284 5116
rect 1316 5084 1320 5116
rect 1280 5036 1320 5084
rect 1280 5004 1284 5036
rect 1316 5004 1320 5036
rect 1280 4956 1320 5004
rect 1280 4924 1284 4956
rect 1316 4924 1320 4956
rect 1280 4876 1320 4924
rect 1280 4844 1284 4876
rect 1316 4844 1320 4876
rect 1280 4796 1320 4844
rect 1280 4764 1284 4796
rect 1316 4764 1320 4796
rect 1280 4716 1320 4764
rect 1280 4684 1284 4716
rect 1316 4684 1320 4716
rect 1280 4636 1320 4684
rect 1280 4604 1284 4636
rect 1316 4604 1320 4636
rect 1280 4556 1320 4604
rect 1280 4524 1284 4556
rect 1316 4524 1320 4556
rect 1280 4476 1320 4524
rect 1280 4444 1284 4476
rect 1316 4444 1320 4476
rect 1280 4440 1320 4444
rect 1360 5516 1400 5520
rect 1360 5484 1364 5516
rect 1396 5484 1400 5516
rect 1360 5436 1400 5484
rect 1360 5404 1364 5436
rect 1396 5404 1400 5436
rect 1360 5356 1400 5404
rect 1360 5324 1364 5356
rect 1396 5324 1400 5356
rect 1360 5276 1400 5324
rect 1360 5244 1364 5276
rect 1396 5244 1400 5276
rect 1360 5196 1400 5244
rect 1360 5164 1364 5196
rect 1396 5164 1400 5196
rect 1360 5116 1400 5164
rect 1360 5084 1364 5116
rect 1396 5084 1400 5116
rect 1360 5036 1400 5084
rect 1360 5004 1364 5036
rect 1396 5004 1400 5036
rect 1360 4956 1400 5004
rect 1360 4924 1364 4956
rect 1396 4924 1400 4956
rect 1360 4876 1400 4924
rect 1360 4844 1364 4876
rect 1396 4844 1400 4876
rect 1360 4796 1400 4844
rect 1360 4764 1364 4796
rect 1396 4764 1400 4796
rect 1360 4716 1400 4764
rect 1360 4684 1364 4716
rect 1396 4684 1400 4716
rect 1360 4636 1400 4684
rect 1360 4604 1364 4636
rect 1396 4604 1400 4636
rect 1360 4556 1400 4604
rect 1360 4524 1364 4556
rect 1396 4524 1400 4556
rect 1360 4476 1400 4524
rect 1360 4444 1364 4476
rect 1396 4444 1400 4476
rect 1360 4440 1400 4444
rect 1440 5516 1480 5520
rect 1440 5484 1444 5516
rect 1476 5484 1480 5516
rect 1440 5436 1480 5484
rect 1440 5404 1444 5436
rect 1476 5404 1480 5436
rect 1440 5356 1480 5404
rect 1440 5324 1444 5356
rect 1476 5324 1480 5356
rect 1440 5276 1480 5324
rect 1440 5244 1444 5276
rect 1476 5244 1480 5276
rect 1440 5196 1480 5244
rect 1440 5164 1444 5196
rect 1476 5164 1480 5196
rect 1440 5116 1480 5164
rect 1440 5084 1444 5116
rect 1476 5084 1480 5116
rect 1440 5036 1480 5084
rect 1440 5004 1444 5036
rect 1476 5004 1480 5036
rect 1440 4956 1480 5004
rect 1440 4924 1444 4956
rect 1476 4924 1480 4956
rect 1440 4876 1480 4924
rect 1440 4844 1444 4876
rect 1476 4844 1480 4876
rect 1440 4796 1480 4844
rect 1440 4764 1444 4796
rect 1476 4764 1480 4796
rect 1440 4716 1480 4764
rect 1440 4684 1444 4716
rect 1476 4684 1480 4716
rect 1440 4636 1480 4684
rect 1440 4604 1444 4636
rect 1476 4604 1480 4636
rect 1440 4556 1480 4604
rect 1440 4524 1444 4556
rect 1476 4524 1480 4556
rect 1440 4476 1480 4524
rect 1440 4444 1444 4476
rect 1476 4444 1480 4476
rect 1440 4440 1480 4444
rect 1520 5516 1560 5520
rect 1520 5484 1524 5516
rect 1556 5484 1560 5516
rect 1520 5436 1560 5484
rect 1520 5404 1524 5436
rect 1556 5404 1560 5436
rect 1520 5356 1560 5404
rect 1520 5324 1524 5356
rect 1556 5324 1560 5356
rect 1520 5276 1560 5324
rect 1520 5244 1524 5276
rect 1556 5244 1560 5276
rect 1520 5196 1560 5244
rect 1520 5164 1524 5196
rect 1556 5164 1560 5196
rect 1520 5116 1560 5164
rect 1520 5084 1524 5116
rect 1556 5084 1560 5116
rect 1520 5036 1560 5084
rect 1520 5004 1524 5036
rect 1556 5004 1560 5036
rect 1520 4956 1560 5004
rect 1520 4924 1524 4956
rect 1556 4924 1560 4956
rect 1520 4876 1560 4924
rect 1520 4844 1524 4876
rect 1556 4844 1560 4876
rect 1520 4796 1560 4844
rect 1520 4764 1524 4796
rect 1556 4764 1560 4796
rect 1520 4716 1560 4764
rect 1520 4684 1524 4716
rect 1556 4684 1560 4716
rect 1520 4636 1560 4684
rect 1520 4604 1524 4636
rect 1556 4604 1560 4636
rect 1520 4556 1560 4604
rect 1520 4524 1524 4556
rect 1556 4524 1560 4556
rect 1520 4476 1560 4524
rect 1520 4444 1524 4476
rect 1556 4444 1560 4476
rect 1520 4440 1560 4444
rect 1600 5516 1640 5520
rect 1600 5484 1604 5516
rect 1636 5484 1640 5516
rect 1600 5436 1640 5484
rect 1600 5404 1604 5436
rect 1636 5404 1640 5436
rect 1600 5356 1640 5404
rect 1600 5324 1604 5356
rect 1636 5324 1640 5356
rect 1600 5276 1640 5324
rect 1600 5244 1604 5276
rect 1636 5244 1640 5276
rect 1600 5196 1640 5244
rect 1600 5164 1604 5196
rect 1636 5164 1640 5196
rect 1600 5116 1640 5164
rect 1600 5084 1604 5116
rect 1636 5084 1640 5116
rect 1600 5036 1640 5084
rect 1600 5004 1604 5036
rect 1636 5004 1640 5036
rect 1600 4956 1640 5004
rect 1600 4924 1604 4956
rect 1636 4924 1640 4956
rect 1600 4876 1640 4924
rect 1600 4844 1604 4876
rect 1636 4844 1640 4876
rect 1600 4796 1640 4844
rect 1600 4764 1604 4796
rect 1636 4764 1640 4796
rect 1600 4716 1640 4764
rect 1600 4684 1604 4716
rect 1636 4684 1640 4716
rect 1600 4636 1640 4684
rect 1600 4604 1604 4636
rect 1636 4604 1640 4636
rect 1600 4556 1640 4604
rect 1600 4524 1604 4556
rect 1636 4524 1640 4556
rect 1600 4476 1640 4524
rect 1600 4444 1604 4476
rect 1636 4444 1640 4476
rect 1600 4440 1640 4444
rect 1680 5516 1720 5520
rect 1680 5484 1684 5516
rect 1716 5484 1720 5516
rect 1680 5436 1720 5484
rect 1680 5404 1684 5436
rect 1716 5404 1720 5436
rect 1680 5356 1720 5404
rect 1680 5324 1684 5356
rect 1716 5324 1720 5356
rect 1680 5276 1720 5324
rect 1680 5244 1684 5276
rect 1716 5244 1720 5276
rect 1680 5196 1720 5244
rect 1680 5164 1684 5196
rect 1716 5164 1720 5196
rect 1680 5116 1720 5164
rect 1680 5084 1684 5116
rect 1716 5084 1720 5116
rect 1680 5036 1720 5084
rect 1680 5004 1684 5036
rect 1716 5004 1720 5036
rect 1680 4956 1720 5004
rect 1680 4924 1684 4956
rect 1716 4924 1720 4956
rect 1680 4876 1720 4924
rect 1680 4844 1684 4876
rect 1716 4844 1720 4876
rect 1680 4796 1720 4844
rect 1680 4764 1684 4796
rect 1716 4764 1720 4796
rect 1680 4716 1720 4764
rect 1680 4684 1684 4716
rect 1716 4684 1720 4716
rect 1680 4636 1720 4684
rect 1680 4604 1684 4636
rect 1716 4604 1720 4636
rect 1680 4556 1720 4604
rect 1680 4524 1684 4556
rect 1716 4524 1720 4556
rect 1680 4476 1720 4524
rect 1680 4444 1684 4476
rect 1716 4444 1720 4476
rect 1680 4440 1720 4444
rect 1760 5516 1800 5520
rect 1760 5484 1764 5516
rect 1796 5484 1800 5516
rect 1760 5436 1800 5484
rect 1760 5404 1764 5436
rect 1796 5404 1800 5436
rect 1760 5356 1800 5404
rect 1760 5324 1764 5356
rect 1796 5324 1800 5356
rect 1760 5276 1800 5324
rect 1760 5244 1764 5276
rect 1796 5244 1800 5276
rect 1760 5196 1800 5244
rect 1760 5164 1764 5196
rect 1796 5164 1800 5196
rect 1760 5116 1800 5164
rect 1760 5084 1764 5116
rect 1796 5084 1800 5116
rect 1760 5036 1800 5084
rect 1760 5004 1764 5036
rect 1796 5004 1800 5036
rect 1760 4956 1800 5004
rect 1760 4924 1764 4956
rect 1796 4924 1800 4956
rect 1760 4876 1800 4924
rect 1760 4844 1764 4876
rect 1796 4844 1800 4876
rect 1760 4796 1800 4844
rect 1760 4764 1764 4796
rect 1796 4764 1800 4796
rect 1760 4716 1800 4764
rect 1760 4684 1764 4716
rect 1796 4684 1800 4716
rect 1760 4636 1800 4684
rect 1760 4604 1764 4636
rect 1796 4604 1800 4636
rect 1760 4556 1800 4604
rect 1760 4524 1764 4556
rect 1796 4524 1800 4556
rect 1760 4476 1800 4524
rect 1760 4444 1764 4476
rect 1796 4444 1800 4476
rect 1760 4440 1800 4444
rect 1840 5516 1880 5520
rect 1840 5484 1844 5516
rect 1876 5484 1880 5516
rect 1840 5436 1880 5484
rect 1840 5404 1844 5436
rect 1876 5404 1880 5436
rect 1840 5356 1880 5404
rect 1840 5324 1844 5356
rect 1876 5324 1880 5356
rect 1840 5276 1880 5324
rect 1840 5244 1844 5276
rect 1876 5244 1880 5276
rect 1840 5196 1880 5244
rect 1840 5164 1844 5196
rect 1876 5164 1880 5196
rect 1840 5116 1880 5164
rect 1840 5084 1844 5116
rect 1876 5084 1880 5116
rect 1840 5036 1880 5084
rect 1840 5004 1844 5036
rect 1876 5004 1880 5036
rect 1840 4956 1880 5004
rect 1840 4924 1844 4956
rect 1876 4924 1880 4956
rect 1840 4876 1880 4924
rect 1840 4844 1844 4876
rect 1876 4844 1880 4876
rect 1840 4796 1880 4844
rect 1840 4764 1844 4796
rect 1876 4764 1880 4796
rect 1840 4716 1880 4764
rect 1840 4684 1844 4716
rect 1876 4684 1880 4716
rect 1840 4636 1880 4684
rect 1840 4604 1844 4636
rect 1876 4604 1880 4636
rect 1840 4556 1880 4604
rect 1840 4524 1844 4556
rect 1876 4524 1880 4556
rect 1840 4476 1880 4524
rect 1840 4444 1844 4476
rect 1876 4444 1880 4476
rect 1840 4440 1880 4444
rect 1920 5516 1960 5520
rect 1920 5484 1924 5516
rect 1956 5484 1960 5516
rect 1920 5436 1960 5484
rect 1920 5404 1924 5436
rect 1956 5404 1960 5436
rect 1920 5356 1960 5404
rect 1920 5324 1924 5356
rect 1956 5324 1960 5356
rect 1920 5276 1960 5324
rect 1920 5244 1924 5276
rect 1956 5244 1960 5276
rect 1920 5196 1960 5244
rect 1920 5164 1924 5196
rect 1956 5164 1960 5196
rect 1920 5116 1960 5164
rect 1920 5084 1924 5116
rect 1956 5084 1960 5116
rect 1920 5036 1960 5084
rect 1920 5004 1924 5036
rect 1956 5004 1960 5036
rect 1920 4956 1960 5004
rect 1920 4924 1924 4956
rect 1956 4924 1960 4956
rect 1920 4876 1960 4924
rect 1920 4844 1924 4876
rect 1956 4844 1960 4876
rect 1920 4796 1960 4844
rect 1920 4764 1924 4796
rect 1956 4764 1960 4796
rect 1920 4716 1960 4764
rect 1920 4684 1924 4716
rect 1956 4684 1960 4716
rect 1920 4636 1960 4684
rect 1920 4604 1924 4636
rect 1956 4604 1960 4636
rect 1920 4556 1960 4604
rect 1920 4524 1924 4556
rect 1956 4524 1960 4556
rect 1920 4476 1960 4524
rect 1920 4444 1924 4476
rect 1956 4444 1960 4476
rect 1920 4440 1960 4444
rect 2000 5516 2040 5520
rect 2000 5484 2004 5516
rect 2036 5484 2040 5516
rect 2000 5436 2040 5484
rect 2000 5404 2004 5436
rect 2036 5404 2040 5436
rect 2000 5356 2040 5404
rect 2000 5324 2004 5356
rect 2036 5324 2040 5356
rect 2000 5276 2040 5324
rect 2000 5244 2004 5276
rect 2036 5244 2040 5276
rect 2000 5196 2040 5244
rect 2000 5164 2004 5196
rect 2036 5164 2040 5196
rect 2000 5116 2040 5164
rect 2000 5084 2004 5116
rect 2036 5084 2040 5116
rect 2000 5036 2040 5084
rect 2000 5004 2004 5036
rect 2036 5004 2040 5036
rect 2000 4956 2040 5004
rect 2000 4924 2004 4956
rect 2036 4924 2040 4956
rect 2000 4876 2040 4924
rect 2000 4844 2004 4876
rect 2036 4844 2040 4876
rect 2000 4796 2040 4844
rect 2000 4764 2004 4796
rect 2036 4764 2040 4796
rect 2000 4716 2040 4764
rect 2000 4684 2004 4716
rect 2036 4684 2040 4716
rect 2000 4636 2040 4684
rect 2000 4604 2004 4636
rect 2036 4604 2040 4636
rect 2000 4556 2040 4604
rect 2000 4524 2004 4556
rect 2036 4524 2040 4556
rect 2000 4476 2040 4524
rect 2000 4444 2004 4476
rect 2036 4444 2040 4476
rect 2000 4440 2040 4444
rect 2080 5516 2120 5520
rect 2080 5484 2084 5516
rect 2116 5484 2120 5516
rect 2080 5436 2120 5484
rect 2080 5404 2084 5436
rect 2116 5404 2120 5436
rect 2080 5356 2120 5404
rect 2080 5324 2084 5356
rect 2116 5324 2120 5356
rect 2080 5276 2120 5324
rect 2080 5244 2084 5276
rect 2116 5244 2120 5276
rect 2080 5196 2120 5244
rect 2080 5164 2084 5196
rect 2116 5164 2120 5196
rect 2080 5116 2120 5164
rect 2080 5084 2084 5116
rect 2116 5084 2120 5116
rect 2080 5036 2120 5084
rect 2080 5004 2084 5036
rect 2116 5004 2120 5036
rect 2080 4956 2120 5004
rect 2080 4924 2084 4956
rect 2116 4924 2120 4956
rect 2080 4876 2120 4924
rect 2080 4844 2084 4876
rect 2116 4844 2120 4876
rect 2080 4796 2120 4844
rect 2080 4764 2084 4796
rect 2116 4764 2120 4796
rect 2080 4716 2120 4764
rect 2080 4684 2084 4716
rect 2116 4684 2120 4716
rect 2080 4636 2120 4684
rect 2080 4604 2084 4636
rect 2116 4604 2120 4636
rect 2080 4556 2120 4604
rect 2080 4524 2084 4556
rect 2116 4524 2120 4556
rect 2080 4476 2120 4524
rect 2080 4444 2084 4476
rect 2116 4444 2120 4476
rect 2080 4440 2120 4444
rect 2160 5516 2200 5520
rect 2160 5484 2164 5516
rect 2196 5484 2200 5516
rect 2160 5436 2200 5484
rect 2160 5404 2164 5436
rect 2196 5404 2200 5436
rect 2160 5356 2200 5404
rect 2160 5324 2164 5356
rect 2196 5324 2200 5356
rect 2160 5276 2200 5324
rect 2160 5244 2164 5276
rect 2196 5244 2200 5276
rect 2160 5196 2200 5244
rect 2160 5164 2164 5196
rect 2196 5164 2200 5196
rect 2160 5116 2200 5164
rect 2160 5084 2164 5116
rect 2196 5084 2200 5116
rect 2160 5036 2200 5084
rect 2160 5004 2164 5036
rect 2196 5004 2200 5036
rect 2160 4956 2200 5004
rect 2160 4924 2164 4956
rect 2196 4924 2200 4956
rect 2160 4876 2200 4924
rect 2160 4844 2164 4876
rect 2196 4844 2200 4876
rect 2160 4796 2200 4844
rect 2160 4764 2164 4796
rect 2196 4764 2200 4796
rect 2160 4716 2200 4764
rect 2160 4684 2164 4716
rect 2196 4684 2200 4716
rect 2160 4636 2200 4684
rect 2160 4604 2164 4636
rect 2196 4604 2200 4636
rect 2160 4556 2200 4604
rect 2160 4524 2164 4556
rect 2196 4524 2200 4556
rect 2160 4476 2200 4524
rect 2160 4444 2164 4476
rect 2196 4444 2200 4476
rect 2160 4440 2200 4444
rect 2240 5516 2280 5520
rect 2240 5484 2244 5516
rect 2276 5484 2280 5516
rect 2240 5436 2280 5484
rect 2240 5404 2244 5436
rect 2276 5404 2280 5436
rect 2240 5356 2280 5404
rect 2240 5324 2244 5356
rect 2276 5324 2280 5356
rect 2240 5276 2280 5324
rect 2240 5244 2244 5276
rect 2276 5244 2280 5276
rect 2240 5196 2280 5244
rect 2240 5164 2244 5196
rect 2276 5164 2280 5196
rect 2240 5116 2280 5164
rect 2240 5084 2244 5116
rect 2276 5084 2280 5116
rect 2240 5036 2280 5084
rect 2240 5004 2244 5036
rect 2276 5004 2280 5036
rect 2240 4956 2280 5004
rect 2240 4924 2244 4956
rect 2276 4924 2280 4956
rect 2240 4876 2280 4924
rect 2240 4844 2244 4876
rect 2276 4844 2280 4876
rect 2240 4796 2280 4844
rect 2240 4764 2244 4796
rect 2276 4764 2280 4796
rect 2240 4716 2280 4764
rect 2240 4684 2244 4716
rect 2276 4684 2280 4716
rect 2240 4636 2280 4684
rect 2240 4604 2244 4636
rect 2276 4604 2280 4636
rect 2240 4556 2280 4604
rect 2240 4524 2244 4556
rect 2276 4524 2280 4556
rect 2240 4476 2280 4524
rect 2240 4444 2244 4476
rect 2276 4444 2280 4476
rect 2240 4440 2280 4444
rect 2320 5516 2360 5520
rect 2320 5484 2324 5516
rect 2356 5484 2360 5516
rect 2320 5436 2360 5484
rect 2320 5404 2324 5436
rect 2356 5404 2360 5436
rect 2320 5356 2360 5404
rect 2320 5324 2324 5356
rect 2356 5324 2360 5356
rect 2320 5276 2360 5324
rect 2320 5244 2324 5276
rect 2356 5244 2360 5276
rect 2320 5196 2360 5244
rect 2320 5164 2324 5196
rect 2356 5164 2360 5196
rect 2320 5116 2360 5164
rect 2320 5084 2324 5116
rect 2356 5084 2360 5116
rect 2320 5036 2360 5084
rect 2320 5004 2324 5036
rect 2356 5004 2360 5036
rect 2320 4956 2360 5004
rect 2320 4924 2324 4956
rect 2356 4924 2360 4956
rect 2320 4876 2360 4924
rect 2320 4844 2324 4876
rect 2356 4844 2360 4876
rect 2320 4796 2360 4844
rect 2320 4764 2324 4796
rect 2356 4764 2360 4796
rect 2320 4716 2360 4764
rect 2320 4684 2324 4716
rect 2356 4684 2360 4716
rect 2320 4636 2360 4684
rect 2320 4604 2324 4636
rect 2356 4604 2360 4636
rect 2320 4556 2360 4604
rect 2320 4524 2324 4556
rect 2356 4524 2360 4556
rect 2320 4476 2360 4524
rect 2320 4444 2324 4476
rect 2356 4444 2360 4476
rect 2320 4440 2360 4444
rect 2400 5516 2440 5520
rect 2400 5484 2404 5516
rect 2436 5484 2440 5516
rect 2400 5436 2440 5484
rect 2400 5404 2404 5436
rect 2436 5404 2440 5436
rect 2400 5356 2440 5404
rect 2400 5324 2404 5356
rect 2436 5324 2440 5356
rect 2400 5276 2440 5324
rect 2400 5244 2404 5276
rect 2436 5244 2440 5276
rect 2400 5196 2440 5244
rect 2400 5164 2404 5196
rect 2436 5164 2440 5196
rect 2400 5116 2440 5164
rect 2400 5084 2404 5116
rect 2436 5084 2440 5116
rect 2400 5036 2440 5084
rect 2400 5004 2404 5036
rect 2436 5004 2440 5036
rect 2400 4956 2440 5004
rect 2400 4924 2404 4956
rect 2436 4924 2440 4956
rect 2400 4876 2440 4924
rect 2400 4844 2404 4876
rect 2436 4844 2440 4876
rect 2400 4796 2440 4844
rect 2400 4764 2404 4796
rect 2436 4764 2440 4796
rect 2400 4716 2440 4764
rect 2400 4684 2404 4716
rect 2436 4684 2440 4716
rect 2400 4636 2440 4684
rect 2400 4604 2404 4636
rect 2436 4604 2440 4636
rect 2400 4556 2440 4604
rect 2400 4524 2404 4556
rect 2436 4524 2440 4556
rect 2400 4476 2440 4524
rect 2400 4444 2404 4476
rect 2436 4444 2440 4476
rect 2400 4440 2440 4444
rect 2480 5516 2520 5520
rect 2480 5484 2484 5516
rect 2516 5484 2520 5516
rect 2480 5436 2520 5484
rect 2480 5404 2484 5436
rect 2516 5404 2520 5436
rect 2480 5356 2520 5404
rect 2480 5324 2484 5356
rect 2516 5324 2520 5356
rect 2480 5276 2520 5324
rect 2480 5244 2484 5276
rect 2516 5244 2520 5276
rect 2480 5196 2520 5244
rect 2480 5164 2484 5196
rect 2516 5164 2520 5196
rect 2480 5116 2520 5164
rect 2480 5084 2484 5116
rect 2516 5084 2520 5116
rect 2480 5036 2520 5084
rect 2480 5004 2484 5036
rect 2516 5004 2520 5036
rect 2480 4956 2520 5004
rect 2480 4924 2484 4956
rect 2516 4924 2520 4956
rect 2480 4876 2520 4924
rect 2480 4844 2484 4876
rect 2516 4844 2520 4876
rect 2480 4796 2520 4844
rect 2480 4764 2484 4796
rect 2516 4764 2520 4796
rect 2480 4716 2520 4764
rect 2480 4684 2484 4716
rect 2516 4684 2520 4716
rect 2480 4636 2520 4684
rect 2480 4604 2484 4636
rect 2516 4604 2520 4636
rect 2480 4556 2520 4604
rect 2480 4524 2484 4556
rect 2516 4524 2520 4556
rect 2480 4476 2520 4524
rect 2480 4444 2484 4476
rect 2516 4444 2520 4476
rect 2480 4440 2520 4444
rect 2560 5516 2600 5520
rect 2560 5484 2564 5516
rect 2596 5484 2600 5516
rect 2560 5436 2600 5484
rect 2560 5404 2564 5436
rect 2596 5404 2600 5436
rect 2560 5356 2600 5404
rect 2560 5324 2564 5356
rect 2596 5324 2600 5356
rect 2560 5276 2600 5324
rect 2560 5244 2564 5276
rect 2596 5244 2600 5276
rect 2560 5196 2600 5244
rect 2560 5164 2564 5196
rect 2596 5164 2600 5196
rect 2560 5116 2600 5164
rect 2560 5084 2564 5116
rect 2596 5084 2600 5116
rect 2560 5036 2600 5084
rect 2560 5004 2564 5036
rect 2596 5004 2600 5036
rect 2560 4956 2600 5004
rect 2560 4924 2564 4956
rect 2596 4924 2600 4956
rect 2560 4876 2600 4924
rect 2560 4844 2564 4876
rect 2596 4844 2600 4876
rect 2560 4796 2600 4844
rect 2560 4764 2564 4796
rect 2596 4764 2600 4796
rect 2560 4716 2600 4764
rect 2560 4684 2564 4716
rect 2596 4684 2600 4716
rect 2560 4636 2600 4684
rect 2560 4604 2564 4636
rect 2596 4604 2600 4636
rect 2560 4556 2600 4604
rect 2560 4524 2564 4556
rect 2596 4524 2600 4556
rect 2560 4476 2600 4524
rect 2560 4444 2564 4476
rect 2596 4444 2600 4476
rect 2560 4440 2600 4444
rect 2640 5516 2680 5520
rect 2640 5484 2644 5516
rect 2676 5484 2680 5516
rect 2640 5436 2680 5484
rect 2640 5404 2644 5436
rect 2676 5404 2680 5436
rect 2640 5356 2680 5404
rect 2640 5324 2644 5356
rect 2676 5324 2680 5356
rect 2640 5276 2680 5324
rect 2640 5244 2644 5276
rect 2676 5244 2680 5276
rect 2640 5196 2680 5244
rect 2640 5164 2644 5196
rect 2676 5164 2680 5196
rect 2640 5116 2680 5164
rect 2640 5084 2644 5116
rect 2676 5084 2680 5116
rect 2640 5036 2680 5084
rect 2640 5004 2644 5036
rect 2676 5004 2680 5036
rect 2640 4956 2680 5004
rect 2640 4924 2644 4956
rect 2676 4924 2680 4956
rect 2640 4876 2680 4924
rect 2640 4844 2644 4876
rect 2676 4844 2680 4876
rect 2640 4796 2680 4844
rect 2640 4764 2644 4796
rect 2676 4764 2680 4796
rect 2640 4716 2680 4764
rect 2640 4684 2644 4716
rect 2676 4684 2680 4716
rect 2640 4636 2680 4684
rect 2640 4604 2644 4636
rect 2676 4604 2680 4636
rect 2640 4556 2680 4604
rect 2640 4524 2644 4556
rect 2676 4524 2680 4556
rect 2640 4476 2680 4524
rect 2640 4444 2644 4476
rect 2676 4444 2680 4476
rect 2640 4440 2680 4444
rect 2720 5516 2760 5520
rect 2720 5484 2724 5516
rect 2756 5484 2760 5516
rect 2720 5436 2760 5484
rect 2720 5404 2724 5436
rect 2756 5404 2760 5436
rect 2720 5356 2760 5404
rect 2720 5324 2724 5356
rect 2756 5324 2760 5356
rect 2720 5276 2760 5324
rect 2720 5244 2724 5276
rect 2756 5244 2760 5276
rect 2720 5196 2760 5244
rect 2720 5164 2724 5196
rect 2756 5164 2760 5196
rect 2720 5116 2760 5164
rect 2720 5084 2724 5116
rect 2756 5084 2760 5116
rect 2720 5036 2760 5084
rect 2720 5004 2724 5036
rect 2756 5004 2760 5036
rect 2720 4956 2760 5004
rect 2720 4924 2724 4956
rect 2756 4924 2760 4956
rect 2720 4876 2760 4924
rect 2720 4844 2724 4876
rect 2756 4844 2760 4876
rect 2720 4796 2760 4844
rect 2720 4764 2724 4796
rect 2756 4764 2760 4796
rect 2720 4716 2760 4764
rect 2720 4684 2724 4716
rect 2756 4684 2760 4716
rect 2720 4636 2760 4684
rect 2720 4604 2724 4636
rect 2756 4604 2760 4636
rect 2720 4556 2760 4604
rect 2720 4524 2724 4556
rect 2756 4524 2760 4556
rect 2720 4476 2760 4524
rect 2720 4444 2724 4476
rect 2756 4444 2760 4476
rect 2720 4440 2760 4444
rect 2800 5516 2840 5520
rect 2800 5484 2804 5516
rect 2836 5484 2840 5516
rect 2800 5436 2840 5484
rect 2800 5404 2804 5436
rect 2836 5404 2840 5436
rect 2800 5356 2840 5404
rect 2800 5324 2804 5356
rect 2836 5324 2840 5356
rect 2800 5276 2840 5324
rect 2800 5244 2804 5276
rect 2836 5244 2840 5276
rect 2800 5196 2840 5244
rect 2800 5164 2804 5196
rect 2836 5164 2840 5196
rect 2800 5116 2840 5164
rect 2800 5084 2804 5116
rect 2836 5084 2840 5116
rect 2800 5036 2840 5084
rect 2800 5004 2804 5036
rect 2836 5004 2840 5036
rect 2800 4956 2840 5004
rect 2800 4924 2804 4956
rect 2836 4924 2840 4956
rect 2800 4876 2840 4924
rect 2800 4844 2804 4876
rect 2836 4844 2840 4876
rect 2800 4796 2840 4844
rect 2800 4764 2804 4796
rect 2836 4764 2840 4796
rect 2800 4716 2840 4764
rect 2800 4684 2804 4716
rect 2836 4684 2840 4716
rect 2800 4636 2840 4684
rect 2800 4604 2804 4636
rect 2836 4604 2840 4636
rect 2800 4556 2840 4604
rect 2800 4524 2804 4556
rect 2836 4524 2840 4556
rect 2800 4476 2840 4524
rect 2800 4444 2804 4476
rect 2836 4444 2840 4476
rect 2800 4440 2840 4444
rect 2880 5516 2920 5520
rect 2880 5484 2884 5516
rect 2916 5484 2920 5516
rect 2880 5436 2920 5484
rect 2880 5404 2884 5436
rect 2916 5404 2920 5436
rect 2880 5356 2920 5404
rect 2880 5324 2884 5356
rect 2916 5324 2920 5356
rect 2880 5276 2920 5324
rect 2880 5244 2884 5276
rect 2916 5244 2920 5276
rect 2880 5196 2920 5244
rect 2880 5164 2884 5196
rect 2916 5164 2920 5196
rect 2880 5116 2920 5164
rect 2880 5084 2884 5116
rect 2916 5084 2920 5116
rect 2880 5036 2920 5084
rect 2880 5004 2884 5036
rect 2916 5004 2920 5036
rect 2880 4956 2920 5004
rect 2880 4924 2884 4956
rect 2916 4924 2920 4956
rect 2880 4876 2920 4924
rect 2880 4844 2884 4876
rect 2916 4844 2920 4876
rect 2880 4796 2920 4844
rect 2880 4764 2884 4796
rect 2916 4764 2920 4796
rect 2880 4716 2920 4764
rect 2880 4684 2884 4716
rect 2916 4684 2920 4716
rect 2880 4636 2920 4684
rect 2880 4604 2884 4636
rect 2916 4604 2920 4636
rect 2880 4556 2920 4604
rect 2880 4524 2884 4556
rect 2916 4524 2920 4556
rect 2880 4476 2920 4524
rect 2880 4444 2884 4476
rect 2916 4444 2920 4476
rect 2880 4440 2920 4444
rect 2960 5516 3000 5520
rect 2960 5484 2964 5516
rect 2996 5484 3000 5516
rect 2960 5436 3000 5484
rect 2960 5404 2964 5436
rect 2996 5404 3000 5436
rect 2960 5356 3000 5404
rect 2960 5324 2964 5356
rect 2996 5324 3000 5356
rect 2960 5276 3000 5324
rect 2960 5244 2964 5276
rect 2996 5244 3000 5276
rect 2960 5196 3000 5244
rect 2960 5164 2964 5196
rect 2996 5164 3000 5196
rect 2960 5116 3000 5164
rect 2960 5084 2964 5116
rect 2996 5084 3000 5116
rect 2960 5036 3000 5084
rect 2960 5004 2964 5036
rect 2996 5004 3000 5036
rect 2960 4956 3000 5004
rect 2960 4924 2964 4956
rect 2996 4924 3000 4956
rect 2960 4876 3000 4924
rect 2960 4844 2964 4876
rect 2996 4844 3000 4876
rect 2960 4796 3000 4844
rect 2960 4764 2964 4796
rect 2996 4764 3000 4796
rect 2960 4716 3000 4764
rect 2960 4684 2964 4716
rect 2996 4684 3000 4716
rect 2960 4636 3000 4684
rect 2960 4604 2964 4636
rect 2996 4604 3000 4636
rect 2960 4556 3000 4604
rect 2960 4524 2964 4556
rect 2996 4524 3000 4556
rect 2960 4476 3000 4524
rect 2960 4444 2964 4476
rect 2996 4444 3000 4476
rect 2960 4440 3000 4444
rect 3040 5516 3080 5520
rect 3040 5484 3044 5516
rect 3076 5484 3080 5516
rect 3040 5436 3080 5484
rect 3040 5404 3044 5436
rect 3076 5404 3080 5436
rect 3040 5356 3080 5404
rect 3040 5324 3044 5356
rect 3076 5324 3080 5356
rect 3040 5276 3080 5324
rect 3040 5244 3044 5276
rect 3076 5244 3080 5276
rect 3040 5196 3080 5244
rect 3040 5164 3044 5196
rect 3076 5164 3080 5196
rect 3040 5116 3080 5164
rect 3040 5084 3044 5116
rect 3076 5084 3080 5116
rect 3040 5036 3080 5084
rect 3040 5004 3044 5036
rect 3076 5004 3080 5036
rect 3040 4956 3080 5004
rect 3040 4924 3044 4956
rect 3076 4924 3080 4956
rect 3040 4876 3080 4924
rect 3040 4844 3044 4876
rect 3076 4844 3080 4876
rect 3040 4796 3080 4844
rect 3040 4764 3044 4796
rect 3076 4764 3080 4796
rect 3040 4716 3080 4764
rect 3040 4684 3044 4716
rect 3076 4684 3080 4716
rect 3040 4636 3080 4684
rect 3040 4604 3044 4636
rect 3076 4604 3080 4636
rect 3040 4556 3080 4604
rect 3040 4524 3044 4556
rect 3076 4524 3080 4556
rect 3040 4476 3080 4524
rect 3040 4444 3044 4476
rect 3076 4444 3080 4476
rect 3040 4440 3080 4444
rect 3120 5516 3160 5520
rect 3120 5484 3124 5516
rect 3156 5484 3160 5516
rect 3120 5436 3160 5484
rect 3120 5404 3124 5436
rect 3156 5404 3160 5436
rect 3120 5356 3160 5404
rect 3120 5324 3124 5356
rect 3156 5324 3160 5356
rect 3120 5276 3160 5324
rect 3120 5244 3124 5276
rect 3156 5244 3160 5276
rect 3120 5196 3160 5244
rect 3120 5164 3124 5196
rect 3156 5164 3160 5196
rect 3120 5116 3160 5164
rect 3120 5084 3124 5116
rect 3156 5084 3160 5116
rect 3120 5036 3160 5084
rect 3120 5004 3124 5036
rect 3156 5004 3160 5036
rect 3120 4956 3160 5004
rect 3120 4924 3124 4956
rect 3156 4924 3160 4956
rect 3120 4876 3160 4924
rect 3120 4844 3124 4876
rect 3156 4844 3160 4876
rect 3120 4796 3160 4844
rect 3120 4764 3124 4796
rect 3156 4764 3160 4796
rect 3120 4716 3160 4764
rect 3120 4684 3124 4716
rect 3156 4684 3160 4716
rect 3120 4636 3160 4684
rect 3120 4604 3124 4636
rect 3156 4604 3160 4636
rect 3120 4556 3160 4604
rect 3120 4524 3124 4556
rect 3156 4524 3160 4556
rect 3120 4476 3160 4524
rect 3120 4444 3124 4476
rect 3156 4444 3160 4476
rect 3120 4440 3160 4444
rect 3200 5516 3240 5520
rect 3200 5484 3204 5516
rect 3236 5484 3240 5516
rect 3200 5436 3240 5484
rect 3200 5404 3204 5436
rect 3236 5404 3240 5436
rect 3200 5356 3240 5404
rect 3200 5324 3204 5356
rect 3236 5324 3240 5356
rect 3200 5276 3240 5324
rect 3200 5244 3204 5276
rect 3236 5244 3240 5276
rect 3200 5196 3240 5244
rect 3200 5164 3204 5196
rect 3236 5164 3240 5196
rect 3200 5116 3240 5164
rect 3200 5084 3204 5116
rect 3236 5084 3240 5116
rect 3200 5036 3240 5084
rect 3200 5004 3204 5036
rect 3236 5004 3240 5036
rect 3200 4956 3240 5004
rect 3200 4924 3204 4956
rect 3236 4924 3240 4956
rect 3200 4876 3240 4924
rect 3200 4844 3204 4876
rect 3236 4844 3240 4876
rect 3200 4796 3240 4844
rect 3200 4764 3204 4796
rect 3236 4764 3240 4796
rect 3200 4716 3240 4764
rect 3200 4684 3204 4716
rect 3236 4684 3240 4716
rect 3200 4636 3240 4684
rect 3200 4604 3204 4636
rect 3236 4604 3240 4636
rect 3200 4556 3240 4604
rect 3200 4524 3204 4556
rect 3236 4524 3240 4556
rect 3200 4476 3240 4524
rect 3200 4444 3204 4476
rect 3236 4444 3240 4476
rect 3200 4440 3240 4444
rect 3280 5516 3320 5520
rect 3280 5484 3284 5516
rect 3316 5484 3320 5516
rect 3280 5436 3320 5484
rect 3280 5404 3284 5436
rect 3316 5404 3320 5436
rect 3280 5356 3320 5404
rect 3280 5324 3284 5356
rect 3316 5324 3320 5356
rect 3280 5276 3320 5324
rect 3280 5244 3284 5276
rect 3316 5244 3320 5276
rect 3280 5196 3320 5244
rect 3280 5164 3284 5196
rect 3316 5164 3320 5196
rect 3280 5116 3320 5164
rect 3280 5084 3284 5116
rect 3316 5084 3320 5116
rect 3280 5036 3320 5084
rect 3280 5004 3284 5036
rect 3316 5004 3320 5036
rect 3280 4956 3320 5004
rect 3280 4924 3284 4956
rect 3316 4924 3320 4956
rect 3280 4876 3320 4924
rect 3280 4844 3284 4876
rect 3316 4844 3320 4876
rect 3280 4796 3320 4844
rect 3280 4764 3284 4796
rect 3316 4764 3320 4796
rect 3280 4716 3320 4764
rect 3280 4684 3284 4716
rect 3316 4684 3320 4716
rect 3280 4636 3320 4684
rect 3280 4604 3284 4636
rect 3316 4604 3320 4636
rect 3280 4556 3320 4604
rect 3280 4524 3284 4556
rect 3316 4524 3320 4556
rect 3280 4476 3320 4524
rect 3280 4444 3284 4476
rect 3316 4444 3320 4476
rect 3280 4440 3320 4444
rect 3360 5516 3400 5520
rect 3360 5484 3364 5516
rect 3396 5484 3400 5516
rect 3360 5436 3400 5484
rect 3360 5404 3364 5436
rect 3396 5404 3400 5436
rect 3360 5356 3400 5404
rect 3360 5324 3364 5356
rect 3396 5324 3400 5356
rect 3360 5276 3400 5324
rect 3360 5244 3364 5276
rect 3396 5244 3400 5276
rect 3360 5196 3400 5244
rect 3360 5164 3364 5196
rect 3396 5164 3400 5196
rect 3360 5116 3400 5164
rect 3360 5084 3364 5116
rect 3396 5084 3400 5116
rect 3360 5036 3400 5084
rect 3360 5004 3364 5036
rect 3396 5004 3400 5036
rect 3360 4956 3400 5004
rect 3360 4924 3364 4956
rect 3396 4924 3400 4956
rect 3360 4876 3400 4924
rect 3360 4844 3364 4876
rect 3396 4844 3400 4876
rect 3360 4796 3400 4844
rect 3360 4764 3364 4796
rect 3396 4764 3400 4796
rect 3360 4716 3400 4764
rect 3360 4684 3364 4716
rect 3396 4684 3400 4716
rect 3360 4636 3400 4684
rect 3360 4604 3364 4636
rect 3396 4604 3400 4636
rect 3360 4556 3400 4604
rect 3360 4524 3364 4556
rect 3396 4524 3400 4556
rect 3360 4476 3400 4524
rect 3360 4444 3364 4476
rect 3396 4444 3400 4476
rect 3360 4440 3400 4444
rect 3440 5516 3480 5520
rect 3440 5484 3444 5516
rect 3476 5484 3480 5516
rect 3440 5436 3480 5484
rect 3440 5404 3444 5436
rect 3476 5404 3480 5436
rect 3440 5356 3480 5404
rect 3440 5324 3444 5356
rect 3476 5324 3480 5356
rect 3440 5276 3480 5324
rect 3440 5244 3444 5276
rect 3476 5244 3480 5276
rect 3440 5196 3480 5244
rect 3440 5164 3444 5196
rect 3476 5164 3480 5196
rect 3440 5116 3480 5164
rect 3440 5084 3444 5116
rect 3476 5084 3480 5116
rect 3440 5036 3480 5084
rect 3440 5004 3444 5036
rect 3476 5004 3480 5036
rect 3440 4956 3480 5004
rect 3440 4924 3444 4956
rect 3476 4924 3480 4956
rect 3440 4876 3480 4924
rect 3440 4844 3444 4876
rect 3476 4844 3480 4876
rect 3440 4796 3480 4844
rect 3440 4764 3444 4796
rect 3476 4764 3480 4796
rect 3440 4716 3480 4764
rect 3440 4684 3444 4716
rect 3476 4684 3480 4716
rect 3440 4636 3480 4684
rect 3440 4604 3444 4636
rect 3476 4604 3480 4636
rect 3440 4556 3480 4604
rect 3440 4524 3444 4556
rect 3476 4524 3480 4556
rect 3440 4476 3480 4524
rect 3440 4444 3444 4476
rect 3476 4444 3480 4476
rect 3440 4440 3480 4444
rect 3520 5516 3560 5520
rect 3520 5484 3524 5516
rect 3556 5484 3560 5516
rect 3520 5436 3560 5484
rect 3520 5404 3524 5436
rect 3556 5404 3560 5436
rect 3520 5356 3560 5404
rect 3520 5324 3524 5356
rect 3556 5324 3560 5356
rect 3520 5276 3560 5324
rect 3520 5244 3524 5276
rect 3556 5244 3560 5276
rect 3520 5196 3560 5244
rect 3520 5164 3524 5196
rect 3556 5164 3560 5196
rect 3520 5116 3560 5164
rect 3520 5084 3524 5116
rect 3556 5084 3560 5116
rect 3520 5036 3560 5084
rect 3520 5004 3524 5036
rect 3556 5004 3560 5036
rect 3520 4956 3560 5004
rect 3520 4924 3524 4956
rect 3556 4924 3560 4956
rect 3520 4876 3560 4924
rect 3520 4844 3524 4876
rect 3556 4844 3560 4876
rect 3520 4796 3560 4844
rect 3520 4764 3524 4796
rect 3556 4764 3560 4796
rect 3520 4716 3560 4764
rect 3520 4684 3524 4716
rect 3556 4684 3560 4716
rect 3520 4636 3560 4684
rect 3520 4604 3524 4636
rect 3556 4604 3560 4636
rect 3520 4556 3560 4604
rect 3520 4524 3524 4556
rect 3556 4524 3560 4556
rect 3520 4476 3560 4524
rect 3520 4444 3524 4476
rect 3556 4444 3560 4476
rect 3520 4440 3560 4444
rect 3600 5516 3640 5520
rect 3600 5484 3604 5516
rect 3636 5484 3640 5516
rect 3600 5436 3640 5484
rect 3600 5404 3604 5436
rect 3636 5404 3640 5436
rect 3600 5356 3640 5404
rect 3600 5324 3604 5356
rect 3636 5324 3640 5356
rect 3600 5276 3640 5324
rect 3600 5244 3604 5276
rect 3636 5244 3640 5276
rect 3600 5196 3640 5244
rect 3600 5164 3604 5196
rect 3636 5164 3640 5196
rect 3600 5116 3640 5164
rect 3600 5084 3604 5116
rect 3636 5084 3640 5116
rect 3600 5036 3640 5084
rect 3600 5004 3604 5036
rect 3636 5004 3640 5036
rect 3600 4956 3640 5004
rect 3600 4924 3604 4956
rect 3636 4924 3640 4956
rect 3600 4876 3640 4924
rect 3600 4844 3604 4876
rect 3636 4844 3640 4876
rect 3600 4796 3640 4844
rect 3600 4764 3604 4796
rect 3636 4764 3640 4796
rect 3600 4716 3640 4764
rect 3600 4684 3604 4716
rect 3636 4684 3640 4716
rect 3600 4636 3640 4684
rect 3600 4604 3604 4636
rect 3636 4604 3640 4636
rect 3600 4556 3640 4604
rect 3600 4524 3604 4556
rect 3636 4524 3640 4556
rect 3600 4476 3640 4524
rect 3600 4444 3604 4476
rect 3636 4444 3640 4476
rect 3600 4440 3640 4444
rect 3680 5516 3720 5520
rect 3680 5484 3684 5516
rect 3716 5484 3720 5516
rect 3680 5436 3720 5484
rect 3680 5404 3684 5436
rect 3716 5404 3720 5436
rect 3680 5356 3720 5404
rect 3680 5324 3684 5356
rect 3716 5324 3720 5356
rect 3680 5276 3720 5324
rect 3680 5244 3684 5276
rect 3716 5244 3720 5276
rect 3680 5196 3720 5244
rect 3680 5164 3684 5196
rect 3716 5164 3720 5196
rect 3680 5116 3720 5164
rect 3680 5084 3684 5116
rect 3716 5084 3720 5116
rect 3680 5036 3720 5084
rect 3680 5004 3684 5036
rect 3716 5004 3720 5036
rect 3680 4956 3720 5004
rect 3680 4924 3684 4956
rect 3716 4924 3720 4956
rect 3680 4876 3720 4924
rect 3680 4844 3684 4876
rect 3716 4844 3720 4876
rect 3680 4796 3720 4844
rect 3680 4764 3684 4796
rect 3716 4764 3720 4796
rect 3680 4716 3720 4764
rect 3680 4684 3684 4716
rect 3716 4684 3720 4716
rect 3680 4636 3720 4684
rect 3680 4604 3684 4636
rect 3716 4604 3720 4636
rect 3680 4556 3720 4604
rect 3680 4524 3684 4556
rect 3716 4524 3720 4556
rect 3680 4476 3720 4524
rect 3680 4444 3684 4476
rect 3716 4444 3720 4476
rect 3680 4440 3720 4444
rect 3760 5516 3800 5520
rect 3760 5484 3764 5516
rect 3796 5484 3800 5516
rect 3760 5436 3800 5484
rect 3760 5404 3764 5436
rect 3796 5404 3800 5436
rect 3760 5356 3800 5404
rect 3760 5324 3764 5356
rect 3796 5324 3800 5356
rect 3760 5276 3800 5324
rect 3760 5244 3764 5276
rect 3796 5244 3800 5276
rect 3760 5196 3800 5244
rect 3760 5164 3764 5196
rect 3796 5164 3800 5196
rect 3760 5116 3800 5164
rect 3760 5084 3764 5116
rect 3796 5084 3800 5116
rect 3760 5036 3800 5084
rect 3760 5004 3764 5036
rect 3796 5004 3800 5036
rect 3760 4956 3800 5004
rect 3760 4924 3764 4956
rect 3796 4924 3800 4956
rect 3760 4876 3800 4924
rect 3760 4844 3764 4876
rect 3796 4844 3800 4876
rect 3760 4796 3800 4844
rect 3760 4764 3764 4796
rect 3796 4764 3800 4796
rect 3760 4716 3800 4764
rect 3760 4684 3764 4716
rect 3796 4684 3800 4716
rect 3760 4636 3800 4684
rect 3760 4604 3764 4636
rect 3796 4604 3800 4636
rect 3760 4556 3800 4604
rect 3760 4524 3764 4556
rect 3796 4524 3800 4556
rect 3760 4476 3800 4524
rect 3760 4444 3764 4476
rect 3796 4444 3800 4476
rect 3760 4440 3800 4444
rect 3840 5516 3880 5520
rect 3840 5484 3844 5516
rect 3876 5484 3880 5516
rect 3840 5436 3880 5484
rect 3840 5404 3844 5436
rect 3876 5404 3880 5436
rect 3840 5356 3880 5404
rect 3840 5324 3844 5356
rect 3876 5324 3880 5356
rect 3840 5276 3880 5324
rect 3840 5244 3844 5276
rect 3876 5244 3880 5276
rect 3840 5196 3880 5244
rect 3840 5164 3844 5196
rect 3876 5164 3880 5196
rect 3840 5116 3880 5164
rect 3840 5084 3844 5116
rect 3876 5084 3880 5116
rect 3840 5036 3880 5084
rect 3840 5004 3844 5036
rect 3876 5004 3880 5036
rect 3840 4956 3880 5004
rect 3840 4924 3844 4956
rect 3876 4924 3880 4956
rect 3840 4876 3880 4924
rect 3840 4844 3844 4876
rect 3876 4844 3880 4876
rect 3840 4796 3880 4844
rect 3840 4764 3844 4796
rect 3876 4764 3880 4796
rect 3840 4716 3880 4764
rect 3840 4684 3844 4716
rect 3876 4684 3880 4716
rect 3840 4636 3880 4684
rect 3840 4604 3844 4636
rect 3876 4604 3880 4636
rect 3840 4556 3880 4604
rect 3840 4524 3844 4556
rect 3876 4524 3880 4556
rect 3840 4476 3880 4524
rect 3840 4444 3844 4476
rect 3876 4444 3880 4476
rect 3840 4440 3880 4444
rect 3920 5516 3960 5520
rect 3920 5484 3924 5516
rect 3956 5484 3960 5516
rect 3920 5436 3960 5484
rect 3920 5404 3924 5436
rect 3956 5404 3960 5436
rect 3920 5356 3960 5404
rect 3920 5324 3924 5356
rect 3956 5324 3960 5356
rect 3920 5276 3960 5324
rect 3920 5244 3924 5276
rect 3956 5244 3960 5276
rect 3920 5196 3960 5244
rect 3920 5164 3924 5196
rect 3956 5164 3960 5196
rect 3920 5116 3960 5164
rect 3920 5084 3924 5116
rect 3956 5084 3960 5116
rect 3920 5036 3960 5084
rect 3920 5004 3924 5036
rect 3956 5004 3960 5036
rect 3920 4956 3960 5004
rect 3920 4924 3924 4956
rect 3956 4924 3960 4956
rect 3920 4876 3960 4924
rect 3920 4844 3924 4876
rect 3956 4844 3960 4876
rect 3920 4796 3960 4844
rect 3920 4764 3924 4796
rect 3956 4764 3960 4796
rect 3920 4716 3960 4764
rect 3920 4684 3924 4716
rect 3956 4684 3960 4716
rect 3920 4636 3960 4684
rect 3920 4604 3924 4636
rect 3956 4604 3960 4636
rect 3920 4556 3960 4604
rect 3920 4524 3924 4556
rect 3956 4524 3960 4556
rect 3920 4476 3960 4524
rect 3920 4444 3924 4476
rect 3956 4444 3960 4476
rect 3920 4440 3960 4444
rect 4000 5516 4040 5520
rect 4000 5484 4004 5516
rect 4036 5484 4040 5516
rect 4000 5436 4040 5484
rect 4000 5404 4004 5436
rect 4036 5404 4040 5436
rect 4000 5356 4040 5404
rect 4000 5324 4004 5356
rect 4036 5324 4040 5356
rect 4000 5276 4040 5324
rect 4000 5244 4004 5276
rect 4036 5244 4040 5276
rect 4000 5196 4040 5244
rect 4000 5164 4004 5196
rect 4036 5164 4040 5196
rect 4000 5116 4040 5164
rect 4000 5084 4004 5116
rect 4036 5084 4040 5116
rect 4000 5036 4040 5084
rect 4000 5004 4004 5036
rect 4036 5004 4040 5036
rect 4000 4956 4040 5004
rect 4000 4924 4004 4956
rect 4036 4924 4040 4956
rect 4000 4876 4040 4924
rect 4000 4844 4004 4876
rect 4036 4844 4040 4876
rect 4000 4796 4040 4844
rect 4000 4764 4004 4796
rect 4036 4764 4040 4796
rect 4000 4716 4040 4764
rect 4000 4684 4004 4716
rect 4036 4684 4040 4716
rect 4000 4636 4040 4684
rect 4000 4604 4004 4636
rect 4036 4604 4040 4636
rect 4000 4556 4040 4604
rect 4000 4524 4004 4556
rect 4036 4524 4040 4556
rect 4000 4476 4040 4524
rect 4000 4444 4004 4476
rect 4036 4444 4040 4476
rect 4000 4440 4040 4444
rect 4080 5516 4120 5520
rect 4080 5484 4084 5516
rect 4116 5484 4120 5516
rect 4080 5436 4120 5484
rect 4080 5404 4084 5436
rect 4116 5404 4120 5436
rect 4080 5356 4120 5404
rect 4080 5324 4084 5356
rect 4116 5324 4120 5356
rect 4080 5276 4120 5324
rect 4080 5244 4084 5276
rect 4116 5244 4120 5276
rect 4080 5196 4120 5244
rect 4080 5164 4084 5196
rect 4116 5164 4120 5196
rect 4080 5116 4120 5164
rect 4080 5084 4084 5116
rect 4116 5084 4120 5116
rect 4080 5036 4120 5084
rect 4080 5004 4084 5036
rect 4116 5004 4120 5036
rect 4080 4956 4120 5004
rect 4080 4924 4084 4956
rect 4116 4924 4120 4956
rect 4080 4876 4120 4924
rect 4080 4844 4084 4876
rect 4116 4844 4120 4876
rect 4080 4796 4120 4844
rect 4080 4764 4084 4796
rect 4116 4764 4120 4796
rect 4080 4716 4120 4764
rect 4080 4684 4084 4716
rect 4116 4684 4120 4716
rect 4080 4636 4120 4684
rect 4080 4604 4084 4636
rect 4116 4604 4120 4636
rect 4080 4556 4120 4604
rect 4080 4524 4084 4556
rect 4116 4524 4120 4556
rect 4080 4476 4120 4524
rect 4080 4444 4084 4476
rect 4116 4444 4120 4476
rect 4080 4440 4120 4444
rect 4160 5516 4200 5520
rect 4160 5484 4164 5516
rect 4196 5484 4200 5516
rect 4160 5436 4200 5484
rect 4160 5404 4164 5436
rect 4196 5404 4200 5436
rect 4160 5356 4200 5404
rect 4160 5324 4164 5356
rect 4196 5324 4200 5356
rect 4160 5276 4200 5324
rect 4160 5244 4164 5276
rect 4196 5244 4200 5276
rect 4160 5196 4200 5244
rect 4160 5164 4164 5196
rect 4196 5164 4200 5196
rect 4160 5116 4200 5164
rect 4160 5084 4164 5116
rect 4196 5084 4200 5116
rect 4160 5036 4200 5084
rect 4160 5004 4164 5036
rect 4196 5004 4200 5036
rect 4160 4956 4200 5004
rect 4160 4924 4164 4956
rect 4196 4924 4200 4956
rect 4160 4876 4200 4924
rect 4160 4844 4164 4876
rect 4196 4844 4200 4876
rect 4160 4796 4200 4844
rect 4160 4764 4164 4796
rect 4196 4764 4200 4796
rect 4160 4716 4200 4764
rect 4160 4684 4164 4716
rect 4196 4684 4200 4716
rect 4160 4636 4200 4684
rect 4160 4604 4164 4636
rect 4196 4604 4200 4636
rect 4160 4556 4200 4604
rect 4160 4524 4164 4556
rect 4196 4524 4200 4556
rect 4160 4476 4200 4524
rect 4160 4444 4164 4476
rect 4196 4444 4200 4476
rect 4160 4440 4200 4444
rect 4240 5516 4280 5520
rect 4240 5484 4244 5516
rect 4276 5484 4280 5516
rect 4240 5436 4280 5484
rect 4240 5404 4244 5436
rect 4276 5404 4280 5436
rect 4240 5356 4280 5404
rect 4240 5324 4244 5356
rect 4276 5324 4280 5356
rect 4240 5276 4280 5324
rect 4240 5244 4244 5276
rect 4276 5244 4280 5276
rect 4240 5196 4280 5244
rect 4240 5164 4244 5196
rect 4276 5164 4280 5196
rect 4240 5116 4280 5164
rect 4240 5084 4244 5116
rect 4276 5084 4280 5116
rect 4240 5036 4280 5084
rect 4240 5004 4244 5036
rect 4276 5004 4280 5036
rect 4240 4956 4280 5004
rect 4240 4924 4244 4956
rect 4276 4924 4280 4956
rect 4240 4876 4280 4924
rect 4240 4844 4244 4876
rect 4276 4844 4280 4876
rect 4240 4796 4280 4844
rect 4240 4764 4244 4796
rect 4276 4764 4280 4796
rect 4240 4716 4280 4764
rect 4240 4684 4244 4716
rect 4276 4684 4280 4716
rect 4240 4636 4280 4684
rect 4240 4604 4244 4636
rect 4276 4604 4280 4636
rect 4240 4556 4280 4604
rect 4240 4524 4244 4556
rect 4276 4524 4280 4556
rect 4240 4476 4280 4524
rect 4240 4444 4244 4476
rect 4276 4444 4280 4476
rect 4240 4440 4280 4444
rect 4320 5516 4360 5520
rect 4320 5484 4324 5516
rect 4356 5484 4360 5516
rect 4320 5436 4360 5484
rect 4320 5404 4324 5436
rect 4356 5404 4360 5436
rect 4320 5356 4360 5404
rect 4320 5324 4324 5356
rect 4356 5324 4360 5356
rect 4320 5276 4360 5324
rect 4320 5244 4324 5276
rect 4356 5244 4360 5276
rect 4320 5196 4360 5244
rect 4320 5164 4324 5196
rect 4356 5164 4360 5196
rect 4320 5116 4360 5164
rect 4320 5084 4324 5116
rect 4356 5084 4360 5116
rect 4320 5036 4360 5084
rect 4320 5004 4324 5036
rect 4356 5004 4360 5036
rect 4320 4956 4360 5004
rect 4320 4924 4324 4956
rect 4356 4924 4360 4956
rect 4320 4876 4360 4924
rect 4320 4844 4324 4876
rect 4356 4844 4360 4876
rect 4320 4796 4360 4844
rect 4320 4764 4324 4796
rect 4356 4764 4360 4796
rect 4320 4716 4360 4764
rect 4320 4684 4324 4716
rect 4356 4684 4360 4716
rect 4320 4636 4360 4684
rect 4320 4604 4324 4636
rect 4356 4604 4360 4636
rect 4320 4556 4360 4604
rect 4320 4524 4324 4556
rect 4356 4524 4360 4556
rect 4320 4476 4360 4524
rect 4320 4444 4324 4476
rect 4356 4444 4360 4476
rect 4320 4440 4360 4444
rect 4400 5516 4440 5520
rect 4400 5484 4404 5516
rect 4436 5484 4440 5516
rect 4400 5436 4440 5484
rect 4400 5404 4404 5436
rect 4436 5404 4440 5436
rect 4400 5356 4440 5404
rect 4400 5324 4404 5356
rect 4436 5324 4440 5356
rect 4400 5276 4440 5324
rect 4400 5244 4404 5276
rect 4436 5244 4440 5276
rect 4400 5196 4440 5244
rect 4400 5164 4404 5196
rect 4436 5164 4440 5196
rect 4400 5116 4440 5164
rect 4400 5084 4404 5116
rect 4436 5084 4440 5116
rect 4400 5036 4440 5084
rect 4400 5004 4404 5036
rect 4436 5004 4440 5036
rect 4400 4956 4440 5004
rect 4400 4924 4404 4956
rect 4436 4924 4440 4956
rect 4400 4876 4440 4924
rect 4400 4844 4404 4876
rect 4436 4844 4440 4876
rect 4400 4796 4440 4844
rect 4400 4764 4404 4796
rect 4436 4764 4440 4796
rect 4400 4716 4440 4764
rect 4400 4684 4404 4716
rect 4436 4684 4440 4716
rect 4400 4636 4440 4684
rect 4400 4604 4404 4636
rect 4436 4604 4440 4636
rect 4400 4556 4440 4604
rect 4400 4524 4404 4556
rect 4436 4524 4440 4556
rect 4400 4476 4440 4524
rect 4400 4444 4404 4476
rect 4436 4444 4440 4476
rect 4400 4440 4440 4444
rect 4480 5516 4520 5520
rect 4480 5484 4484 5516
rect 4516 5484 4520 5516
rect 4480 5436 4520 5484
rect 4480 5404 4484 5436
rect 4516 5404 4520 5436
rect 4480 5356 4520 5404
rect 4480 5324 4484 5356
rect 4516 5324 4520 5356
rect 4480 5276 4520 5324
rect 4480 5244 4484 5276
rect 4516 5244 4520 5276
rect 4480 5196 4520 5244
rect 4480 5164 4484 5196
rect 4516 5164 4520 5196
rect 4480 5116 4520 5164
rect 4480 5084 4484 5116
rect 4516 5084 4520 5116
rect 4480 5036 4520 5084
rect 4480 5004 4484 5036
rect 4516 5004 4520 5036
rect 4480 4956 4520 5004
rect 4480 4924 4484 4956
rect 4516 4924 4520 4956
rect 4480 4876 4520 4924
rect 4480 4844 4484 4876
rect 4516 4844 4520 4876
rect 4480 4796 4520 4844
rect 4480 4764 4484 4796
rect 4516 4764 4520 4796
rect 4480 4716 4520 4764
rect 4480 4684 4484 4716
rect 4516 4684 4520 4716
rect 4480 4636 4520 4684
rect 4480 4604 4484 4636
rect 4516 4604 4520 4636
rect 4480 4556 4520 4604
rect 4480 4524 4484 4556
rect 4516 4524 4520 4556
rect 4480 4476 4520 4524
rect 4480 4444 4484 4476
rect 4516 4444 4520 4476
rect 4480 4440 4520 4444
rect 4560 5516 4600 5520
rect 4560 5484 4564 5516
rect 4596 5484 4600 5516
rect 4560 5436 4600 5484
rect 4560 5404 4564 5436
rect 4596 5404 4600 5436
rect 4560 5356 4600 5404
rect 4560 5324 4564 5356
rect 4596 5324 4600 5356
rect 4560 5276 4600 5324
rect 4560 5244 4564 5276
rect 4596 5244 4600 5276
rect 4560 5196 4600 5244
rect 4560 5164 4564 5196
rect 4596 5164 4600 5196
rect 4560 5116 4600 5164
rect 4560 5084 4564 5116
rect 4596 5084 4600 5116
rect 4560 5036 4600 5084
rect 4560 5004 4564 5036
rect 4596 5004 4600 5036
rect 4560 4956 4600 5004
rect 4560 4924 4564 4956
rect 4596 4924 4600 4956
rect 4560 4876 4600 4924
rect 4560 4844 4564 4876
rect 4596 4844 4600 4876
rect 4560 4796 4600 4844
rect 4560 4764 4564 4796
rect 4596 4764 4600 4796
rect 4560 4716 4600 4764
rect 4560 4684 4564 4716
rect 4596 4684 4600 4716
rect 4560 4636 4600 4684
rect 4560 4604 4564 4636
rect 4596 4604 4600 4636
rect 4560 4556 4600 4604
rect 4560 4524 4564 4556
rect 4596 4524 4600 4556
rect 4560 4476 4600 4524
rect 4560 4444 4564 4476
rect 4596 4444 4600 4476
rect 4560 4440 4600 4444
rect 4640 5516 4680 5520
rect 4640 5484 4644 5516
rect 4676 5484 4680 5516
rect 4640 5436 4680 5484
rect 4640 5404 4644 5436
rect 4676 5404 4680 5436
rect 4640 5356 4680 5404
rect 4640 5324 4644 5356
rect 4676 5324 4680 5356
rect 4640 5276 4680 5324
rect 4640 5244 4644 5276
rect 4676 5244 4680 5276
rect 4640 5196 4680 5244
rect 4640 5164 4644 5196
rect 4676 5164 4680 5196
rect 4640 5116 4680 5164
rect 4640 5084 4644 5116
rect 4676 5084 4680 5116
rect 4640 5036 4680 5084
rect 4640 5004 4644 5036
rect 4676 5004 4680 5036
rect 4640 4956 4680 5004
rect 4640 4924 4644 4956
rect 4676 4924 4680 4956
rect 4640 4876 4680 4924
rect 4640 4844 4644 4876
rect 4676 4844 4680 4876
rect 4640 4796 4680 4844
rect 4640 4764 4644 4796
rect 4676 4764 4680 4796
rect 4640 4716 4680 4764
rect 4640 4684 4644 4716
rect 4676 4684 4680 4716
rect 4640 4636 4680 4684
rect 4640 4604 4644 4636
rect 4676 4604 4680 4636
rect 4640 4556 4680 4604
rect 4640 4524 4644 4556
rect 4676 4524 4680 4556
rect 4640 4476 4680 4524
rect 4640 4444 4644 4476
rect 4676 4444 4680 4476
rect 4640 4440 4680 4444
rect 4720 5516 4760 5520
rect 4720 5484 4724 5516
rect 4756 5484 4760 5516
rect 4720 5436 4760 5484
rect 4720 5404 4724 5436
rect 4756 5404 4760 5436
rect 4720 5356 4760 5404
rect 4720 5324 4724 5356
rect 4756 5324 4760 5356
rect 4720 5276 4760 5324
rect 4720 5244 4724 5276
rect 4756 5244 4760 5276
rect 4720 5196 4760 5244
rect 4720 5164 4724 5196
rect 4756 5164 4760 5196
rect 4720 5116 4760 5164
rect 4720 5084 4724 5116
rect 4756 5084 4760 5116
rect 4720 5036 4760 5084
rect 4720 5004 4724 5036
rect 4756 5004 4760 5036
rect 4720 4956 4760 5004
rect 4720 4924 4724 4956
rect 4756 4924 4760 4956
rect 4720 4876 4760 4924
rect 4720 4844 4724 4876
rect 4756 4844 4760 4876
rect 4720 4796 4760 4844
rect 4720 4764 4724 4796
rect 4756 4764 4760 4796
rect 4720 4716 4760 4764
rect 4720 4684 4724 4716
rect 4756 4684 4760 4716
rect 4720 4636 4760 4684
rect 4720 4604 4724 4636
rect 4756 4604 4760 4636
rect 4720 4556 4760 4604
rect 4720 4524 4724 4556
rect 4756 4524 4760 4556
rect 4720 4476 4760 4524
rect 4720 4444 4724 4476
rect 4756 4444 4760 4476
rect 4720 4440 4760 4444
rect 4800 5516 4840 5520
rect 4800 5484 4804 5516
rect 4836 5484 4840 5516
rect 4800 5436 4840 5484
rect 4800 5404 4804 5436
rect 4836 5404 4840 5436
rect 4800 5356 4840 5404
rect 4800 5324 4804 5356
rect 4836 5324 4840 5356
rect 4800 5276 4840 5324
rect 4800 5244 4804 5276
rect 4836 5244 4840 5276
rect 4800 5196 4840 5244
rect 4800 5164 4804 5196
rect 4836 5164 4840 5196
rect 4800 5116 4840 5164
rect 4800 5084 4804 5116
rect 4836 5084 4840 5116
rect 4800 5036 4840 5084
rect 4800 5004 4804 5036
rect 4836 5004 4840 5036
rect 4800 4956 4840 5004
rect 4800 4924 4804 4956
rect 4836 4924 4840 4956
rect 4800 4876 4840 4924
rect 4800 4844 4804 4876
rect 4836 4844 4840 4876
rect 4800 4796 4840 4844
rect 4800 4764 4804 4796
rect 4836 4764 4840 4796
rect 4800 4716 4840 4764
rect 4800 4684 4804 4716
rect 4836 4684 4840 4716
rect 4800 4636 4840 4684
rect 4800 4604 4804 4636
rect 4836 4604 4840 4636
rect 4800 4556 4840 4604
rect 4800 4524 4804 4556
rect 4836 4524 4840 4556
rect 4800 4476 4840 4524
rect 4800 4444 4804 4476
rect 4836 4444 4840 4476
rect 4800 4440 4840 4444
rect 4880 5516 4920 5564
rect 4880 5484 4884 5516
rect 4916 5484 4920 5516
rect 4880 5436 4920 5484
rect 4880 5404 4884 5436
rect 4916 5404 4920 5436
rect 4880 5356 4920 5404
rect 4880 5324 4884 5356
rect 4916 5324 4920 5356
rect 4880 5276 4920 5324
rect 4880 5244 4884 5276
rect 4916 5244 4920 5276
rect 4880 5196 4920 5244
rect 4880 5164 4884 5196
rect 4916 5164 4920 5196
rect 4880 5116 4920 5164
rect 4880 5084 4884 5116
rect 4916 5084 4920 5116
rect 4880 5036 4920 5084
rect 4880 5004 4884 5036
rect 4916 5004 4920 5036
rect 4880 4956 4920 5004
rect 4880 4924 4884 4956
rect 4916 4924 4920 4956
rect 4880 4876 4920 4924
rect 4880 4844 4884 4876
rect 4916 4844 4920 4876
rect 4880 4796 4920 4844
rect 4880 4764 4884 4796
rect 4916 4764 4920 4796
rect 4880 4716 4920 4764
rect 4880 4684 4884 4716
rect 4916 4684 4920 4716
rect 4880 4636 4920 4684
rect 4880 4604 4884 4636
rect 4916 4604 4920 4636
rect 4880 4556 4920 4604
rect 4880 4524 4884 4556
rect 4916 4524 4920 4556
rect 4880 4476 4920 4524
rect 4880 4444 4884 4476
rect 4916 4444 4920 4476
rect -880 4364 -876 4396
rect -844 4364 -840 4396
rect -880 4316 -840 4364
rect -880 4284 -876 4316
rect -844 4284 -840 4316
rect -880 4236 -840 4284
rect -880 4204 -876 4236
rect -844 4204 -840 4236
rect -880 4156 -840 4204
rect -880 4124 -876 4156
rect -844 4124 -840 4156
rect -880 4076 -840 4124
rect -880 4044 -876 4076
rect -844 4044 -840 4076
rect -880 3996 -840 4044
rect -880 3964 -876 3996
rect -844 3964 -840 3996
rect -880 3916 -840 3964
rect -880 3884 -876 3916
rect -844 3884 -840 3916
rect -880 3836 -840 3884
rect -880 3804 -876 3836
rect -844 3804 -840 3836
rect -880 3756 -840 3804
rect -880 3724 -876 3756
rect -844 3724 -840 3756
rect -880 3676 -840 3724
rect -880 3644 -876 3676
rect -844 3644 -840 3676
rect -880 3596 -840 3644
rect -800 4396 -760 4400
rect -800 4364 -796 4396
rect -764 4364 -760 4396
rect -800 4316 -760 4364
rect -800 4284 -796 4316
rect -764 4284 -760 4316
rect -800 4236 -760 4284
rect -800 4204 -796 4236
rect -764 4204 -760 4236
rect -800 4156 -760 4204
rect -800 4124 -796 4156
rect -764 4124 -760 4156
rect -800 4076 -760 4124
rect -800 4044 -796 4076
rect -764 4044 -760 4076
rect -800 3996 -760 4044
rect -800 3964 -796 3996
rect -764 3964 -760 3996
rect -800 3916 -760 3964
rect -800 3884 -796 3916
rect -764 3884 -760 3916
rect -800 3836 -760 3884
rect -800 3804 -796 3836
rect -764 3804 -760 3836
rect -800 3756 -760 3804
rect -800 3724 -796 3756
rect -764 3724 -760 3756
rect -800 3676 -760 3724
rect -800 3644 -796 3676
rect -764 3644 -760 3676
rect -800 3640 -760 3644
rect -720 4396 -680 4400
rect -720 4364 -716 4396
rect -684 4364 -680 4396
rect -720 4316 -680 4364
rect -720 4284 -716 4316
rect -684 4284 -680 4316
rect -720 4236 -680 4284
rect -720 4204 -716 4236
rect -684 4204 -680 4236
rect -720 4156 -680 4204
rect -720 4124 -716 4156
rect -684 4124 -680 4156
rect -720 4076 -680 4124
rect -720 4044 -716 4076
rect -684 4044 -680 4076
rect -720 3996 -680 4044
rect -720 3964 -716 3996
rect -684 3964 -680 3996
rect -720 3916 -680 3964
rect -720 3884 -716 3916
rect -684 3884 -680 3916
rect -720 3836 -680 3884
rect -720 3804 -716 3836
rect -684 3804 -680 3836
rect -720 3756 -680 3804
rect -720 3724 -716 3756
rect -684 3724 -680 3756
rect -720 3676 -680 3724
rect -720 3644 -716 3676
rect -684 3644 -680 3676
rect -720 3640 -680 3644
rect -640 4396 -600 4400
rect -640 4364 -636 4396
rect -604 4364 -600 4396
rect -640 4316 -600 4364
rect -640 4284 -636 4316
rect -604 4284 -600 4316
rect -640 4236 -600 4284
rect -640 4204 -636 4236
rect -604 4204 -600 4236
rect -640 4156 -600 4204
rect -640 4124 -636 4156
rect -604 4124 -600 4156
rect -640 4076 -600 4124
rect -640 4044 -636 4076
rect -604 4044 -600 4076
rect -640 3996 -600 4044
rect -640 3964 -636 3996
rect -604 3964 -600 3996
rect -640 3916 -600 3964
rect -640 3884 -636 3916
rect -604 3884 -600 3916
rect -640 3836 -600 3884
rect -640 3804 -636 3836
rect -604 3804 -600 3836
rect -640 3756 -600 3804
rect -640 3724 -636 3756
rect -604 3724 -600 3756
rect -640 3676 -600 3724
rect -640 3644 -636 3676
rect -604 3644 -600 3676
rect -640 3640 -600 3644
rect -560 4396 -520 4400
rect -560 4364 -556 4396
rect -524 4364 -520 4396
rect -560 4316 -520 4364
rect -560 4284 -556 4316
rect -524 4284 -520 4316
rect -560 4236 -520 4284
rect -560 4204 -556 4236
rect -524 4204 -520 4236
rect -560 4156 -520 4204
rect -560 4124 -556 4156
rect -524 4124 -520 4156
rect -560 4076 -520 4124
rect -560 4044 -556 4076
rect -524 4044 -520 4076
rect -560 3996 -520 4044
rect -560 3964 -556 3996
rect -524 3964 -520 3996
rect -560 3916 -520 3964
rect -560 3884 -556 3916
rect -524 3884 -520 3916
rect -560 3836 -520 3884
rect -560 3804 -556 3836
rect -524 3804 -520 3836
rect -560 3756 -520 3804
rect -560 3724 -556 3756
rect -524 3724 -520 3756
rect -560 3676 -520 3724
rect -560 3644 -556 3676
rect -524 3644 -520 3676
rect -560 3640 -520 3644
rect -480 4396 -440 4400
rect -480 4364 -476 4396
rect -444 4364 -440 4396
rect -480 4316 -440 4364
rect -480 4284 -476 4316
rect -444 4284 -440 4316
rect -480 4236 -440 4284
rect -480 4204 -476 4236
rect -444 4204 -440 4236
rect -480 4156 -440 4204
rect -480 4124 -476 4156
rect -444 4124 -440 4156
rect -480 4076 -440 4124
rect -480 4044 -476 4076
rect -444 4044 -440 4076
rect -480 3996 -440 4044
rect -480 3964 -476 3996
rect -444 3964 -440 3996
rect -480 3916 -440 3964
rect -480 3884 -476 3916
rect -444 3884 -440 3916
rect -480 3836 -440 3884
rect -480 3804 -476 3836
rect -444 3804 -440 3836
rect -480 3756 -440 3804
rect -480 3724 -476 3756
rect -444 3724 -440 3756
rect -480 3676 -440 3724
rect -480 3644 -476 3676
rect -444 3644 -440 3676
rect -480 3640 -440 3644
rect -400 4396 -360 4400
rect -400 4364 -396 4396
rect -364 4364 -360 4396
rect -400 4316 -360 4364
rect -400 4284 -396 4316
rect -364 4284 -360 4316
rect -400 4236 -360 4284
rect -400 4204 -396 4236
rect -364 4204 -360 4236
rect -400 4156 -360 4204
rect -400 4124 -396 4156
rect -364 4124 -360 4156
rect -400 4076 -360 4124
rect -400 4044 -396 4076
rect -364 4044 -360 4076
rect -400 3996 -360 4044
rect -400 3964 -396 3996
rect -364 3964 -360 3996
rect -400 3916 -360 3964
rect -400 3884 -396 3916
rect -364 3884 -360 3916
rect -400 3836 -360 3884
rect -400 3804 -396 3836
rect -364 3804 -360 3836
rect -400 3756 -360 3804
rect -400 3724 -396 3756
rect -364 3724 -360 3756
rect -400 3676 -360 3724
rect -400 3644 -396 3676
rect -364 3644 -360 3676
rect -400 3640 -360 3644
rect -320 4396 -280 4400
rect -320 4364 -316 4396
rect -284 4364 -280 4396
rect -320 4316 -280 4364
rect -320 4284 -316 4316
rect -284 4284 -280 4316
rect -320 4236 -280 4284
rect -320 4204 -316 4236
rect -284 4204 -280 4236
rect -320 4156 -280 4204
rect -320 4124 -316 4156
rect -284 4124 -280 4156
rect -320 4076 -280 4124
rect -320 4044 -316 4076
rect -284 4044 -280 4076
rect -320 3996 -280 4044
rect -320 3964 -316 3996
rect -284 3964 -280 3996
rect -320 3916 -280 3964
rect -320 3884 -316 3916
rect -284 3884 -280 3916
rect -320 3836 -280 3884
rect -320 3804 -316 3836
rect -284 3804 -280 3836
rect -320 3756 -280 3804
rect -320 3724 -316 3756
rect -284 3724 -280 3756
rect -320 3676 -280 3724
rect -320 3644 -316 3676
rect -284 3644 -280 3676
rect -320 3640 -280 3644
rect -240 4396 -200 4400
rect -240 4364 -236 4396
rect -204 4364 -200 4396
rect -240 4316 -200 4364
rect -240 4284 -236 4316
rect -204 4284 -200 4316
rect -240 4236 -200 4284
rect -240 4204 -236 4236
rect -204 4204 -200 4236
rect -240 4156 -200 4204
rect -240 4124 -236 4156
rect -204 4124 -200 4156
rect -240 4076 -200 4124
rect -240 4044 -236 4076
rect -204 4044 -200 4076
rect -240 3996 -200 4044
rect -240 3964 -236 3996
rect -204 3964 -200 3996
rect -240 3916 -200 3964
rect -240 3884 -236 3916
rect -204 3884 -200 3916
rect -240 3836 -200 3884
rect -240 3804 -236 3836
rect -204 3804 -200 3836
rect -240 3756 -200 3804
rect -240 3724 -236 3756
rect -204 3724 -200 3756
rect -240 3676 -200 3724
rect -240 3644 -236 3676
rect -204 3644 -200 3676
rect -240 3640 -200 3644
rect -160 4396 -120 4400
rect -160 4364 -156 4396
rect -124 4364 -120 4396
rect -160 4316 -120 4364
rect -160 4284 -156 4316
rect -124 4284 -120 4316
rect -160 4236 -120 4284
rect -160 4204 -156 4236
rect -124 4204 -120 4236
rect -160 4156 -120 4204
rect -160 4124 -156 4156
rect -124 4124 -120 4156
rect -160 4076 -120 4124
rect -160 4044 -156 4076
rect -124 4044 -120 4076
rect -160 3996 -120 4044
rect -160 3964 -156 3996
rect -124 3964 -120 3996
rect -160 3916 -120 3964
rect -160 3884 -156 3916
rect -124 3884 -120 3916
rect -160 3836 -120 3884
rect -160 3804 -156 3836
rect -124 3804 -120 3836
rect -160 3756 -120 3804
rect -160 3724 -156 3756
rect -124 3724 -120 3756
rect -160 3676 -120 3724
rect -160 3644 -156 3676
rect -124 3644 -120 3676
rect -160 3640 -120 3644
rect -80 4396 -40 4400
rect -80 4364 -76 4396
rect -44 4364 -40 4396
rect -80 4316 -40 4364
rect -80 4284 -76 4316
rect -44 4284 -40 4316
rect -80 4236 -40 4284
rect -80 4204 -76 4236
rect -44 4204 -40 4236
rect -80 4156 -40 4204
rect -80 4124 -76 4156
rect -44 4124 -40 4156
rect -80 4076 -40 4124
rect -80 4044 -76 4076
rect -44 4044 -40 4076
rect -80 3996 -40 4044
rect -80 3964 -76 3996
rect -44 3964 -40 3996
rect -80 3916 -40 3964
rect -80 3884 -76 3916
rect -44 3884 -40 3916
rect -80 3836 -40 3884
rect -80 3804 -76 3836
rect -44 3804 -40 3836
rect -80 3756 -40 3804
rect -80 3724 -76 3756
rect -44 3724 -40 3756
rect -80 3676 -40 3724
rect -80 3644 -76 3676
rect -44 3644 -40 3676
rect -80 3640 -40 3644
rect 0 4396 40 4400
rect 0 4364 4 4396
rect 36 4364 40 4396
rect 0 4316 40 4364
rect 0 4284 4 4316
rect 36 4284 40 4316
rect 0 4236 40 4284
rect 0 4204 4 4236
rect 36 4204 40 4236
rect 0 4156 40 4204
rect 0 4124 4 4156
rect 36 4124 40 4156
rect 0 4076 40 4124
rect 0 4044 4 4076
rect 36 4044 40 4076
rect 0 3996 40 4044
rect 0 3964 4 3996
rect 36 3964 40 3996
rect 0 3916 40 3964
rect 0 3884 4 3916
rect 36 3884 40 3916
rect 0 3836 40 3884
rect 0 3804 4 3836
rect 36 3804 40 3836
rect 0 3756 40 3804
rect 0 3724 4 3756
rect 36 3724 40 3756
rect 0 3676 40 3724
rect 0 3644 4 3676
rect 36 3644 40 3676
rect 0 3640 40 3644
rect 80 4396 120 4400
rect 80 4364 84 4396
rect 116 4364 120 4396
rect 80 4316 120 4364
rect 80 4284 84 4316
rect 116 4284 120 4316
rect 80 4236 120 4284
rect 80 4204 84 4236
rect 116 4204 120 4236
rect 80 4156 120 4204
rect 80 4124 84 4156
rect 116 4124 120 4156
rect 80 4076 120 4124
rect 80 4044 84 4076
rect 116 4044 120 4076
rect 80 3996 120 4044
rect 80 3964 84 3996
rect 116 3964 120 3996
rect 80 3916 120 3964
rect 80 3884 84 3916
rect 116 3884 120 3916
rect 80 3836 120 3884
rect 80 3804 84 3836
rect 116 3804 120 3836
rect 80 3756 120 3804
rect 80 3724 84 3756
rect 116 3724 120 3756
rect 80 3676 120 3724
rect 80 3644 84 3676
rect 116 3644 120 3676
rect 80 3640 120 3644
rect 160 4396 200 4400
rect 160 4364 164 4396
rect 196 4364 200 4396
rect 160 4316 200 4364
rect 160 4284 164 4316
rect 196 4284 200 4316
rect 160 4236 200 4284
rect 160 4204 164 4236
rect 196 4204 200 4236
rect 160 4156 200 4204
rect 160 4124 164 4156
rect 196 4124 200 4156
rect 160 4076 200 4124
rect 160 4044 164 4076
rect 196 4044 200 4076
rect 160 3996 200 4044
rect 160 3964 164 3996
rect 196 3964 200 3996
rect 160 3916 200 3964
rect 160 3884 164 3916
rect 196 3884 200 3916
rect 160 3836 200 3884
rect 160 3804 164 3836
rect 196 3804 200 3836
rect 160 3756 200 3804
rect 160 3724 164 3756
rect 196 3724 200 3756
rect 160 3676 200 3724
rect 160 3644 164 3676
rect 196 3644 200 3676
rect 160 3640 200 3644
rect 240 4396 280 4400
rect 240 4364 244 4396
rect 276 4364 280 4396
rect 240 4316 280 4364
rect 240 4284 244 4316
rect 276 4284 280 4316
rect 240 4236 280 4284
rect 240 4204 244 4236
rect 276 4204 280 4236
rect 240 4156 280 4204
rect 240 4124 244 4156
rect 276 4124 280 4156
rect 240 4076 280 4124
rect 240 4044 244 4076
rect 276 4044 280 4076
rect 240 3996 280 4044
rect 240 3964 244 3996
rect 276 3964 280 3996
rect 240 3916 280 3964
rect 240 3884 244 3916
rect 276 3884 280 3916
rect 240 3836 280 3884
rect 240 3804 244 3836
rect 276 3804 280 3836
rect 240 3756 280 3804
rect 240 3724 244 3756
rect 276 3724 280 3756
rect 240 3676 280 3724
rect 240 3644 244 3676
rect 276 3644 280 3676
rect 240 3640 280 3644
rect 320 4396 360 4400
rect 320 4364 324 4396
rect 356 4364 360 4396
rect 320 4316 360 4364
rect 320 4284 324 4316
rect 356 4284 360 4316
rect 320 4236 360 4284
rect 320 4204 324 4236
rect 356 4204 360 4236
rect 320 4156 360 4204
rect 320 4124 324 4156
rect 356 4124 360 4156
rect 320 4076 360 4124
rect 320 4044 324 4076
rect 356 4044 360 4076
rect 320 3996 360 4044
rect 320 3964 324 3996
rect 356 3964 360 3996
rect 320 3916 360 3964
rect 320 3884 324 3916
rect 356 3884 360 3916
rect 320 3836 360 3884
rect 320 3804 324 3836
rect 356 3804 360 3836
rect 320 3756 360 3804
rect 320 3724 324 3756
rect 356 3724 360 3756
rect 320 3676 360 3724
rect 320 3644 324 3676
rect 356 3644 360 3676
rect 320 3640 360 3644
rect 400 4396 440 4400
rect 400 4364 404 4396
rect 436 4364 440 4396
rect 400 4316 440 4364
rect 400 4284 404 4316
rect 436 4284 440 4316
rect 400 4236 440 4284
rect 400 4204 404 4236
rect 436 4204 440 4236
rect 400 4156 440 4204
rect 400 4124 404 4156
rect 436 4124 440 4156
rect 400 4076 440 4124
rect 400 4044 404 4076
rect 436 4044 440 4076
rect 400 3996 440 4044
rect 400 3964 404 3996
rect 436 3964 440 3996
rect 400 3916 440 3964
rect 400 3884 404 3916
rect 436 3884 440 3916
rect 400 3836 440 3884
rect 400 3804 404 3836
rect 436 3804 440 3836
rect 400 3756 440 3804
rect 400 3724 404 3756
rect 436 3724 440 3756
rect 400 3676 440 3724
rect 400 3644 404 3676
rect 436 3644 440 3676
rect 400 3640 440 3644
rect 480 4396 520 4400
rect 480 4364 484 4396
rect 516 4364 520 4396
rect 480 4316 520 4364
rect 480 4284 484 4316
rect 516 4284 520 4316
rect 480 4236 520 4284
rect 480 4204 484 4236
rect 516 4204 520 4236
rect 480 4156 520 4204
rect 480 4124 484 4156
rect 516 4124 520 4156
rect 480 4076 520 4124
rect 480 4044 484 4076
rect 516 4044 520 4076
rect 480 3996 520 4044
rect 480 3964 484 3996
rect 516 3964 520 3996
rect 480 3916 520 3964
rect 480 3884 484 3916
rect 516 3884 520 3916
rect 480 3836 520 3884
rect 480 3804 484 3836
rect 516 3804 520 3836
rect 480 3756 520 3804
rect 480 3724 484 3756
rect 516 3724 520 3756
rect 480 3676 520 3724
rect 480 3644 484 3676
rect 516 3644 520 3676
rect 480 3640 520 3644
rect 560 4396 600 4400
rect 560 4364 564 4396
rect 596 4364 600 4396
rect 560 4316 600 4364
rect 560 4284 564 4316
rect 596 4284 600 4316
rect 560 4236 600 4284
rect 560 4204 564 4236
rect 596 4204 600 4236
rect 560 4156 600 4204
rect 560 4124 564 4156
rect 596 4124 600 4156
rect 560 4076 600 4124
rect 560 4044 564 4076
rect 596 4044 600 4076
rect 560 3996 600 4044
rect 560 3964 564 3996
rect 596 3964 600 3996
rect 560 3916 600 3964
rect 560 3884 564 3916
rect 596 3884 600 3916
rect 560 3836 600 3884
rect 560 3804 564 3836
rect 596 3804 600 3836
rect 560 3756 600 3804
rect 560 3724 564 3756
rect 596 3724 600 3756
rect 560 3676 600 3724
rect 560 3644 564 3676
rect 596 3644 600 3676
rect 560 3640 600 3644
rect 640 4396 680 4400
rect 640 4364 644 4396
rect 676 4364 680 4396
rect 640 4316 680 4364
rect 640 4284 644 4316
rect 676 4284 680 4316
rect 640 4236 680 4284
rect 640 4204 644 4236
rect 676 4204 680 4236
rect 640 4156 680 4204
rect 640 4124 644 4156
rect 676 4124 680 4156
rect 640 4076 680 4124
rect 640 4044 644 4076
rect 676 4044 680 4076
rect 640 3996 680 4044
rect 640 3964 644 3996
rect 676 3964 680 3996
rect 640 3916 680 3964
rect 640 3884 644 3916
rect 676 3884 680 3916
rect 640 3836 680 3884
rect 640 3804 644 3836
rect 676 3804 680 3836
rect 640 3756 680 3804
rect 640 3724 644 3756
rect 676 3724 680 3756
rect 640 3676 680 3724
rect 640 3644 644 3676
rect 676 3644 680 3676
rect 640 3640 680 3644
rect 720 4396 760 4400
rect 720 4364 724 4396
rect 756 4364 760 4396
rect 720 4316 760 4364
rect 720 4284 724 4316
rect 756 4284 760 4316
rect 720 4236 760 4284
rect 720 4204 724 4236
rect 756 4204 760 4236
rect 720 4156 760 4204
rect 720 4124 724 4156
rect 756 4124 760 4156
rect 720 4076 760 4124
rect 720 4044 724 4076
rect 756 4044 760 4076
rect 720 3996 760 4044
rect 720 3964 724 3996
rect 756 3964 760 3996
rect 720 3916 760 3964
rect 720 3884 724 3916
rect 756 3884 760 3916
rect 720 3836 760 3884
rect 720 3804 724 3836
rect 756 3804 760 3836
rect 720 3756 760 3804
rect 720 3724 724 3756
rect 756 3724 760 3756
rect 720 3676 760 3724
rect 720 3644 724 3676
rect 756 3644 760 3676
rect 720 3640 760 3644
rect 800 4396 840 4400
rect 800 4364 804 4396
rect 836 4364 840 4396
rect 800 4316 840 4364
rect 800 4284 804 4316
rect 836 4284 840 4316
rect 800 4236 840 4284
rect 800 4204 804 4236
rect 836 4204 840 4236
rect 800 4156 840 4204
rect 800 4124 804 4156
rect 836 4124 840 4156
rect 800 4076 840 4124
rect 800 4044 804 4076
rect 836 4044 840 4076
rect 800 3996 840 4044
rect 800 3964 804 3996
rect 836 3964 840 3996
rect 800 3916 840 3964
rect 800 3884 804 3916
rect 836 3884 840 3916
rect 800 3836 840 3884
rect 800 3804 804 3836
rect 836 3804 840 3836
rect 800 3756 840 3804
rect 800 3724 804 3756
rect 836 3724 840 3756
rect 800 3676 840 3724
rect 800 3644 804 3676
rect 836 3644 840 3676
rect 800 3640 840 3644
rect 880 4396 920 4400
rect 880 4364 884 4396
rect 916 4364 920 4396
rect 880 4316 920 4364
rect 880 4284 884 4316
rect 916 4284 920 4316
rect 880 4236 920 4284
rect 880 4204 884 4236
rect 916 4204 920 4236
rect 880 4156 920 4204
rect 880 4124 884 4156
rect 916 4124 920 4156
rect 880 4076 920 4124
rect 880 4044 884 4076
rect 916 4044 920 4076
rect 880 3996 920 4044
rect 880 3964 884 3996
rect 916 3964 920 3996
rect 880 3916 920 3964
rect 880 3884 884 3916
rect 916 3884 920 3916
rect 880 3836 920 3884
rect 880 3804 884 3836
rect 916 3804 920 3836
rect 880 3756 920 3804
rect 880 3724 884 3756
rect 916 3724 920 3756
rect 880 3676 920 3724
rect 880 3644 884 3676
rect 916 3644 920 3676
rect 880 3640 920 3644
rect 960 4396 1000 4400
rect 960 4364 964 4396
rect 996 4364 1000 4396
rect 960 4316 1000 4364
rect 960 4284 964 4316
rect 996 4284 1000 4316
rect 960 4236 1000 4284
rect 960 4204 964 4236
rect 996 4204 1000 4236
rect 960 4156 1000 4204
rect 960 4124 964 4156
rect 996 4124 1000 4156
rect 960 4076 1000 4124
rect 960 4044 964 4076
rect 996 4044 1000 4076
rect 960 3996 1000 4044
rect 960 3964 964 3996
rect 996 3964 1000 3996
rect 960 3916 1000 3964
rect 960 3884 964 3916
rect 996 3884 1000 3916
rect 960 3836 1000 3884
rect 960 3804 964 3836
rect 996 3804 1000 3836
rect 960 3756 1000 3804
rect 960 3724 964 3756
rect 996 3724 1000 3756
rect 960 3676 1000 3724
rect 960 3644 964 3676
rect 996 3644 1000 3676
rect 960 3640 1000 3644
rect 1040 4396 1080 4400
rect 1040 4364 1044 4396
rect 1076 4364 1080 4396
rect 1040 4316 1080 4364
rect 1040 4284 1044 4316
rect 1076 4284 1080 4316
rect 1040 4236 1080 4284
rect 1040 4204 1044 4236
rect 1076 4204 1080 4236
rect 1040 4156 1080 4204
rect 1040 4124 1044 4156
rect 1076 4124 1080 4156
rect 1040 4076 1080 4124
rect 1040 4044 1044 4076
rect 1076 4044 1080 4076
rect 1040 3996 1080 4044
rect 1040 3964 1044 3996
rect 1076 3964 1080 3996
rect 1040 3916 1080 3964
rect 1040 3884 1044 3916
rect 1076 3884 1080 3916
rect 1040 3836 1080 3884
rect 1040 3804 1044 3836
rect 1076 3804 1080 3836
rect 1040 3756 1080 3804
rect 1040 3724 1044 3756
rect 1076 3724 1080 3756
rect 1040 3676 1080 3724
rect 1040 3644 1044 3676
rect 1076 3644 1080 3676
rect 1040 3640 1080 3644
rect 1120 4396 1160 4400
rect 1120 4364 1124 4396
rect 1156 4364 1160 4396
rect 1120 4316 1160 4364
rect 1120 4284 1124 4316
rect 1156 4284 1160 4316
rect 1120 4236 1160 4284
rect 1120 4204 1124 4236
rect 1156 4204 1160 4236
rect 1120 4156 1160 4204
rect 1120 4124 1124 4156
rect 1156 4124 1160 4156
rect 1120 4076 1160 4124
rect 1120 4044 1124 4076
rect 1156 4044 1160 4076
rect 1120 3996 1160 4044
rect 1120 3964 1124 3996
rect 1156 3964 1160 3996
rect 1120 3916 1160 3964
rect 1120 3884 1124 3916
rect 1156 3884 1160 3916
rect 1120 3836 1160 3884
rect 1120 3804 1124 3836
rect 1156 3804 1160 3836
rect 1120 3756 1160 3804
rect 1120 3724 1124 3756
rect 1156 3724 1160 3756
rect 1120 3676 1160 3724
rect 1120 3644 1124 3676
rect 1156 3644 1160 3676
rect 1120 3640 1160 3644
rect 1200 4396 1240 4400
rect 1200 4364 1204 4396
rect 1236 4364 1240 4396
rect 1200 4316 1240 4364
rect 1200 4284 1204 4316
rect 1236 4284 1240 4316
rect 1200 4236 1240 4284
rect 1200 4204 1204 4236
rect 1236 4204 1240 4236
rect 1200 4156 1240 4204
rect 1200 4124 1204 4156
rect 1236 4124 1240 4156
rect 1200 4076 1240 4124
rect 1200 4044 1204 4076
rect 1236 4044 1240 4076
rect 1200 3996 1240 4044
rect 1200 3964 1204 3996
rect 1236 3964 1240 3996
rect 1200 3916 1240 3964
rect 1200 3884 1204 3916
rect 1236 3884 1240 3916
rect 1200 3836 1240 3884
rect 1200 3804 1204 3836
rect 1236 3804 1240 3836
rect 1200 3756 1240 3804
rect 1200 3724 1204 3756
rect 1236 3724 1240 3756
rect 1200 3676 1240 3724
rect 1200 3644 1204 3676
rect 1236 3644 1240 3676
rect 1200 3640 1240 3644
rect 1280 4396 1320 4400
rect 1280 4364 1284 4396
rect 1316 4364 1320 4396
rect 1280 4316 1320 4364
rect 1280 4284 1284 4316
rect 1316 4284 1320 4316
rect 1280 4236 1320 4284
rect 1280 4204 1284 4236
rect 1316 4204 1320 4236
rect 1280 4156 1320 4204
rect 1280 4124 1284 4156
rect 1316 4124 1320 4156
rect 1280 4076 1320 4124
rect 1280 4044 1284 4076
rect 1316 4044 1320 4076
rect 1280 3996 1320 4044
rect 1280 3964 1284 3996
rect 1316 3964 1320 3996
rect 1280 3916 1320 3964
rect 1280 3884 1284 3916
rect 1316 3884 1320 3916
rect 1280 3836 1320 3884
rect 1280 3804 1284 3836
rect 1316 3804 1320 3836
rect 1280 3756 1320 3804
rect 1280 3724 1284 3756
rect 1316 3724 1320 3756
rect 1280 3676 1320 3724
rect 1280 3644 1284 3676
rect 1316 3644 1320 3676
rect 1280 3640 1320 3644
rect 1360 4396 1400 4400
rect 1360 4364 1364 4396
rect 1396 4364 1400 4396
rect 1360 4316 1400 4364
rect 1360 4284 1364 4316
rect 1396 4284 1400 4316
rect 1360 4236 1400 4284
rect 1360 4204 1364 4236
rect 1396 4204 1400 4236
rect 1360 4156 1400 4204
rect 1360 4124 1364 4156
rect 1396 4124 1400 4156
rect 1360 4076 1400 4124
rect 1360 4044 1364 4076
rect 1396 4044 1400 4076
rect 1360 3996 1400 4044
rect 1360 3964 1364 3996
rect 1396 3964 1400 3996
rect 1360 3916 1400 3964
rect 1360 3884 1364 3916
rect 1396 3884 1400 3916
rect 1360 3836 1400 3884
rect 1360 3804 1364 3836
rect 1396 3804 1400 3836
rect 1360 3756 1400 3804
rect 1360 3724 1364 3756
rect 1396 3724 1400 3756
rect 1360 3676 1400 3724
rect 1360 3644 1364 3676
rect 1396 3644 1400 3676
rect 1360 3640 1400 3644
rect 1440 4396 1480 4400
rect 1440 4364 1444 4396
rect 1476 4364 1480 4396
rect 1440 4316 1480 4364
rect 1440 4284 1444 4316
rect 1476 4284 1480 4316
rect 1440 4236 1480 4284
rect 1440 4204 1444 4236
rect 1476 4204 1480 4236
rect 1440 4156 1480 4204
rect 1440 4124 1444 4156
rect 1476 4124 1480 4156
rect 1440 4076 1480 4124
rect 1440 4044 1444 4076
rect 1476 4044 1480 4076
rect 1440 3996 1480 4044
rect 1440 3964 1444 3996
rect 1476 3964 1480 3996
rect 1440 3916 1480 3964
rect 1440 3884 1444 3916
rect 1476 3884 1480 3916
rect 1440 3836 1480 3884
rect 1440 3804 1444 3836
rect 1476 3804 1480 3836
rect 1440 3756 1480 3804
rect 1440 3724 1444 3756
rect 1476 3724 1480 3756
rect 1440 3676 1480 3724
rect 1440 3644 1444 3676
rect 1476 3644 1480 3676
rect 1440 3640 1480 3644
rect 1520 4396 1560 4400
rect 1520 4364 1524 4396
rect 1556 4364 1560 4396
rect 1520 4316 1560 4364
rect 1520 4284 1524 4316
rect 1556 4284 1560 4316
rect 1520 4236 1560 4284
rect 1520 4204 1524 4236
rect 1556 4204 1560 4236
rect 1520 4156 1560 4204
rect 1520 4124 1524 4156
rect 1556 4124 1560 4156
rect 1520 4076 1560 4124
rect 1520 4044 1524 4076
rect 1556 4044 1560 4076
rect 1520 3996 1560 4044
rect 1520 3964 1524 3996
rect 1556 3964 1560 3996
rect 1520 3916 1560 3964
rect 1520 3884 1524 3916
rect 1556 3884 1560 3916
rect 1520 3836 1560 3884
rect 1520 3804 1524 3836
rect 1556 3804 1560 3836
rect 1520 3756 1560 3804
rect 1520 3724 1524 3756
rect 1556 3724 1560 3756
rect 1520 3676 1560 3724
rect 1520 3644 1524 3676
rect 1556 3644 1560 3676
rect 1520 3640 1560 3644
rect 1600 4396 1640 4400
rect 1600 4364 1604 4396
rect 1636 4364 1640 4396
rect 1600 4316 1640 4364
rect 1600 4284 1604 4316
rect 1636 4284 1640 4316
rect 1600 4236 1640 4284
rect 1600 4204 1604 4236
rect 1636 4204 1640 4236
rect 1600 4156 1640 4204
rect 1600 4124 1604 4156
rect 1636 4124 1640 4156
rect 1600 4076 1640 4124
rect 1600 4044 1604 4076
rect 1636 4044 1640 4076
rect 1600 3996 1640 4044
rect 1600 3964 1604 3996
rect 1636 3964 1640 3996
rect 1600 3916 1640 3964
rect 1600 3884 1604 3916
rect 1636 3884 1640 3916
rect 1600 3836 1640 3884
rect 1600 3804 1604 3836
rect 1636 3804 1640 3836
rect 1600 3756 1640 3804
rect 1600 3724 1604 3756
rect 1636 3724 1640 3756
rect 1600 3676 1640 3724
rect 1600 3644 1604 3676
rect 1636 3644 1640 3676
rect 1600 3640 1640 3644
rect 1680 4396 1720 4400
rect 1680 4364 1684 4396
rect 1716 4364 1720 4396
rect 1680 4316 1720 4364
rect 1680 4284 1684 4316
rect 1716 4284 1720 4316
rect 1680 4236 1720 4284
rect 1680 4204 1684 4236
rect 1716 4204 1720 4236
rect 1680 4156 1720 4204
rect 1680 4124 1684 4156
rect 1716 4124 1720 4156
rect 1680 4076 1720 4124
rect 1680 4044 1684 4076
rect 1716 4044 1720 4076
rect 1680 3996 1720 4044
rect 1680 3964 1684 3996
rect 1716 3964 1720 3996
rect 1680 3916 1720 3964
rect 1680 3884 1684 3916
rect 1716 3884 1720 3916
rect 1680 3836 1720 3884
rect 1680 3804 1684 3836
rect 1716 3804 1720 3836
rect 1680 3756 1720 3804
rect 1680 3724 1684 3756
rect 1716 3724 1720 3756
rect 1680 3676 1720 3724
rect 1680 3644 1684 3676
rect 1716 3644 1720 3676
rect 1680 3640 1720 3644
rect 1760 4396 1800 4400
rect 1760 4364 1764 4396
rect 1796 4364 1800 4396
rect 1760 4316 1800 4364
rect 1760 4284 1764 4316
rect 1796 4284 1800 4316
rect 1760 4236 1800 4284
rect 1760 4204 1764 4236
rect 1796 4204 1800 4236
rect 1760 4156 1800 4204
rect 1760 4124 1764 4156
rect 1796 4124 1800 4156
rect 1760 4076 1800 4124
rect 1760 4044 1764 4076
rect 1796 4044 1800 4076
rect 1760 3996 1800 4044
rect 1760 3964 1764 3996
rect 1796 3964 1800 3996
rect 1760 3916 1800 3964
rect 1760 3884 1764 3916
rect 1796 3884 1800 3916
rect 1760 3836 1800 3884
rect 1760 3804 1764 3836
rect 1796 3804 1800 3836
rect 1760 3756 1800 3804
rect 1760 3724 1764 3756
rect 1796 3724 1800 3756
rect 1760 3676 1800 3724
rect 1760 3644 1764 3676
rect 1796 3644 1800 3676
rect 1760 3640 1800 3644
rect 1840 4396 1880 4400
rect 1840 4364 1844 4396
rect 1876 4364 1880 4396
rect 1840 4316 1880 4364
rect 1840 4284 1844 4316
rect 1876 4284 1880 4316
rect 1840 4236 1880 4284
rect 1840 4204 1844 4236
rect 1876 4204 1880 4236
rect 1840 4156 1880 4204
rect 1840 4124 1844 4156
rect 1876 4124 1880 4156
rect 1840 4076 1880 4124
rect 1840 4044 1844 4076
rect 1876 4044 1880 4076
rect 1840 3996 1880 4044
rect 1840 3964 1844 3996
rect 1876 3964 1880 3996
rect 1840 3916 1880 3964
rect 1840 3884 1844 3916
rect 1876 3884 1880 3916
rect 1840 3836 1880 3884
rect 1840 3804 1844 3836
rect 1876 3804 1880 3836
rect 1840 3756 1880 3804
rect 1840 3724 1844 3756
rect 1876 3724 1880 3756
rect 1840 3676 1880 3724
rect 1840 3644 1844 3676
rect 1876 3644 1880 3676
rect 1840 3640 1880 3644
rect 1920 4396 1960 4400
rect 1920 4364 1924 4396
rect 1956 4364 1960 4396
rect 1920 4316 1960 4364
rect 1920 4284 1924 4316
rect 1956 4284 1960 4316
rect 1920 4236 1960 4284
rect 1920 4204 1924 4236
rect 1956 4204 1960 4236
rect 1920 4156 1960 4204
rect 1920 4124 1924 4156
rect 1956 4124 1960 4156
rect 1920 4076 1960 4124
rect 1920 4044 1924 4076
rect 1956 4044 1960 4076
rect 1920 3996 1960 4044
rect 1920 3964 1924 3996
rect 1956 3964 1960 3996
rect 1920 3916 1960 3964
rect 1920 3884 1924 3916
rect 1956 3884 1960 3916
rect 1920 3836 1960 3884
rect 1920 3804 1924 3836
rect 1956 3804 1960 3836
rect 1920 3756 1960 3804
rect 1920 3724 1924 3756
rect 1956 3724 1960 3756
rect 1920 3676 1960 3724
rect 1920 3644 1924 3676
rect 1956 3644 1960 3676
rect 1920 3640 1960 3644
rect 2000 4396 2040 4400
rect 2000 4364 2004 4396
rect 2036 4364 2040 4396
rect 2000 4316 2040 4364
rect 2000 4284 2004 4316
rect 2036 4284 2040 4316
rect 2000 4236 2040 4284
rect 2000 4204 2004 4236
rect 2036 4204 2040 4236
rect 2000 4156 2040 4204
rect 2000 4124 2004 4156
rect 2036 4124 2040 4156
rect 2000 4076 2040 4124
rect 2000 4044 2004 4076
rect 2036 4044 2040 4076
rect 2000 3996 2040 4044
rect 2000 3964 2004 3996
rect 2036 3964 2040 3996
rect 2000 3916 2040 3964
rect 2000 3884 2004 3916
rect 2036 3884 2040 3916
rect 2000 3836 2040 3884
rect 2000 3804 2004 3836
rect 2036 3804 2040 3836
rect 2000 3756 2040 3804
rect 2000 3724 2004 3756
rect 2036 3724 2040 3756
rect 2000 3676 2040 3724
rect 2000 3644 2004 3676
rect 2036 3644 2040 3676
rect 2000 3640 2040 3644
rect 2080 4396 2120 4400
rect 2080 4364 2084 4396
rect 2116 4364 2120 4396
rect 2080 4316 2120 4364
rect 2080 4284 2084 4316
rect 2116 4284 2120 4316
rect 2080 4236 2120 4284
rect 2080 4204 2084 4236
rect 2116 4204 2120 4236
rect 2080 4156 2120 4204
rect 2080 4124 2084 4156
rect 2116 4124 2120 4156
rect 2080 4076 2120 4124
rect 2080 4044 2084 4076
rect 2116 4044 2120 4076
rect 2080 3996 2120 4044
rect 2080 3964 2084 3996
rect 2116 3964 2120 3996
rect 2080 3916 2120 3964
rect 2080 3884 2084 3916
rect 2116 3884 2120 3916
rect 2080 3836 2120 3884
rect 2080 3804 2084 3836
rect 2116 3804 2120 3836
rect 2080 3756 2120 3804
rect 2080 3724 2084 3756
rect 2116 3724 2120 3756
rect 2080 3676 2120 3724
rect 2080 3644 2084 3676
rect 2116 3644 2120 3676
rect 2080 3640 2120 3644
rect 2160 4396 2200 4400
rect 2160 4364 2164 4396
rect 2196 4364 2200 4396
rect 2160 4316 2200 4364
rect 2160 4284 2164 4316
rect 2196 4284 2200 4316
rect 2160 4236 2200 4284
rect 2160 4204 2164 4236
rect 2196 4204 2200 4236
rect 2160 4156 2200 4204
rect 2160 4124 2164 4156
rect 2196 4124 2200 4156
rect 2160 4076 2200 4124
rect 2160 4044 2164 4076
rect 2196 4044 2200 4076
rect 2160 3996 2200 4044
rect 2160 3964 2164 3996
rect 2196 3964 2200 3996
rect 2160 3916 2200 3964
rect 2160 3884 2164 3916
rect 2196 3884 2200 3916
rect 2160 3836 2200 3884
rect 2160 3804 2164 3836
rect 2196 3804 2200 3836
rect 2160 3756 2200 3804
rect 2160 3724 2164 3756
rect 2196 3724 2200 3756
rect 2160 3676 2200 3724
rect 2160 3644 2164 3676
rect 2196 3644 2200 3676
rect 2160 3640 2200 3644
rect 2240 4396 2280 4400
rect 2240 4364 2244 4396
rect 2276 4364 2280 4396
rect 2240 4316 2280 4364
rect 2240 4284 2244 4316
rect 2276 4284 2280 4316
rect 2240 4236 2280 4284
rect 2240 4204 2244 4236
rect 2276 4204 2280 4236
rect 2240 4156 2280 4204
rect 2240 4124 2244 4156
rect 2276 4124 2280 4156
rect 2240 4076 2280 4124
rect 2240 4044 2244 4076
rect 2276 4044 2280 4076
rect 2240 3996 2280 4044
rect 2240 3964 2244 3996
rect 2276 3964 2280 3996
rect 2240 3916 2280 3964
rect 2240 3884 2244 3916
rect 2276 3884 2280 3916
rect 2240 3836 2280 3884
rect 2240 3804 2244 3836
rect 2276 3804 2280 3836
rect 2240 3756 2280 3804
rect 2240 3724 2244 3756
rect 2276 3724 2280 3756
rect 2240 3676 2280 3724
rect 2240 3644 2244 3676
rect 2276 3644 2280 3676
rect 2240 3640 2280 3644
rect 2320 4396 2360 4400
rect 2320 4364 2324 4396
rect 2356 4364 2360 4396
rect 2320 4316 2360 4364
rect 2320 4284 2324 4316
rect 2356 4284 2360 4316
rect 2320 4236 2360 4284
rect 2320 4204 2324 4236
rect 2356 4204 2360 4236
rect 2320 4156 2360 4204
rect 2320 4124 2324 4156
rect 2356 4124 2360 4156
rect 2320 4076 2360 4124
rect 2320 4044 2324 4076
rect 2356 4044 2360 4076
rect 2320 3996 2360 4044
rect 2320 3964 2324 3996
rect 2356 3964 2360 3996
rect 2320 3916 2360 3964
rect 2320 3884 2324 3916
rect 2356 3884 2360 3916
rect 2320 3836 2360 3884
rect 2320 3804 2324 3836
rect 2356 3804 2360 3836
rect 2320 3756 2360 3804
rect 2320 3724 2324 3756
rect 2356 3724 2360 3756
rect 2320 3676 2360 3724
rect 2320 3644 2324 3676
rect 2356 3644 2360 3676
rect 2320 3640 2360 3644
rect 2400 4396 2440 4400
rect 2400 4364 2404 4396
rect 2436 4364 2440 4396
rect 2400 4316 2440 4364
rect 2400 4284 2404 4316
rect 2436 4284 2440 4316
rect 2400 4236 2440 4284
rect 2400 4204 2404 4236
rect 2436 4204 2440 4236
rect 2400 4156 2440 4204
rect 2400 4124 2404 4156
rect 2436 4124 2440 4156
rect 2400 4076 2440 4124
rect 2400 4044 2404 4076
rect 2436 4044 2440 4076
rect 2400 3996 2440 4044
rect 2400 3964 2404 3996
rect 2436 3964 2440 3996
rect 2400 3916 2440 3964
rect 2400 3884 2404 3916
rect 2436 3884 2440 3916
rect 2400 3836 2440 3884
rect 2400 3804 2404 3836
rect 2436 3804 2440 3836
rect 2400 3756 2440 3804
rect 2400 3724 2404 3756
rect 2436 3724 2440 3756
rect 2400 3676 2440 3724
rect 2400 3644 2404 3676
rect 2436 3644 2440 3676
rect 2400 3640 2440 3644
rect 2480 4396 2520 4400
rect 2480 4364 2484 4396
rect 2516 4364 2520 4396
rect 2480 4316 2520 4364
rect 2480 4284 2484 4316
rect 2516 4284 2520 4316
rect 2480 4236 2520 4284
rect 2480 4204 2484 4236
rect 2516 4204 2520 4236
rect 2480 4156 2520 4204
rect 2480 4124 2484 4156
rect 2516 4124 2520 4156
rect 2480 4076 2520 4124
rect 2480 4044 2484 4076
rect 2516 4044 2520 4076
rect 2480 3996 2520 4044
rect 2480 3964 2484 3996
rect 2516 3964 2520 3996
rect 2480 3916 2520 3964
rect 2480 3884 2484 3916
rect 2516 3884 2520 3916
rect 2480 3836 2520 3884
rect 2480 3804 2484 3836
rect 2516 3804 2520 3836
rect 2480 3756 2520 3804
rect 2480 3724 2484 3756
rect 2516 3724 2520 3756
rect 2480 3676 2520 3724
rect 2480 3644 2484 3676
rect 2516 3644 2520 3676
rect 2480 3640 2520 3644
rect 2560 4396 2600 4400
rect 2560 4364 2564 4396
rect 2596 4364 2600 4396
rect 2560 4316 2600 4364
rect 2560 4284 2564 4316
rect 2596 4284 2600 4316
rect 2560 4236 2600 4284
rect 2560 4204 2564 4236
rect 2596 4204 2600 4236
rect 2560 4156 2600 4204
rect 2560 4124 2564 4156
rect 2596 4124 2600 4156
rect 2560 4076 2600 4124
rect 2560 4044 2564 4076
rect 2596 4044 2600 4076
rect 2560 3996 2600 4044
rect 2560 3964 2564 3996
rect 2596 3964 2600 3996
rect 2560 3916 2600 3964
rect 2560 3884 2564 3916
rect 2596 3884 2600 3916
rect 2560 3836 2600 3884
rect 2560 3804 2564 3836
rect 2596 3804 2600 3836
rect 2560 3756 2600 3804
rect 2560 3724 2564 3756
rect 2596 3724 2600 3756
rect 2560 3676 2600 3724
rect 2560 3644 2564 3676
rect 2596 3644 2600 3676
rect 2560 3640 2600 3644
rect 2640 4396 2680 4400
rect 2640 4364 2644 4396
rect 2676 4364 2680 4396
rect 2640 4316 2680 4364
rect 2640 4284 2644 4316
rect 2676 4284 2680 4316
rect 2640 4236 2680 4284
rect 2640 4204 2644 4236
rect 2676 4204 2680 4236
rect 2640 4156 2680 4204
rect 2640 4124 2644 4156
rect 2676 4124 2680 4156
rect 2640 4076 2680 4124
rect 2640 4044 2644 4076
rect 2676 4044 2680 4076
rect 2640 3996 2680 4044
rect 2640 3964 2644 3996
rect 2676 3964 2680 3996
rect 2640 3916 2680 3964
rect 2640 3884 2644 3916
rect 2676 3884 2680 3916
rect 2640 3836 2680 3884
rect 2640 3804 2644 3836
rect 2676 3804 2680 3836
rect 2640 3756 2680 3804
rect 2640 3724 2644 3756
rect 2676 3724 2680 3756
rect 2640 3676 2680 3724
rect 2640 3644 2644 3676
rect 2676 3644 2680 3676
rect 2640 3640 2680 3644
rect 2720 4396 2760 4400
rect 2720 4364 2724 4396
rect 2756 4364 2760 4396
rect 2720 4316 2760 4364
rect 2720 4284 2724 4316
rect 2756 4284 2760 4316
rect 2720 4236 2760 4284
rect 2720 4204 2724 4236
rect 2756 4204 2760 4236
rect 2720 4156 2760 4204
rect 2720 4124 2724 4156
rect 2756 4124 2760 4156
rect 2720 4076 2760 4124
rect 2720 4044 2724 4076
rect 2756 4044 2760 4076
rect 2720 3996 2760 4044
rect 2720 3964 2724 3996
rect 2756 3964 2760 3996
rect 2720 3916 2760 3964
rect 2720 3884 2724 3916
rect 2756 3884 2760 3916
rect 2720 3836 2760 3884
rect 2720 3804 2724 3836
rect 2756 3804 2760 3836
rect 2720 3756 2760 3804
rect 2720 3724 2724 3756
rect 2756 3724 2760 3756
rect 2720 3676 2760 3724
rect 2720 3644 2724 3676
rect 2756 3644 2760 3676
rect 2720 3640 2760 3644
rect 2800 4396 2840 4400
rect 2800 4364 2804 4396
rect 2836 4364 2840 4396
rect 2800 4316 2840 4364
rect 2800 4284 2804 4316
rect 2836 4284 2840 4316
rect 2800 4236 2840 4284
rect 2800 4204 2804 4236
rect 2836 4204 2840 4236
rect 2800 4156 2840 4204
rect 2800 4124 2804 4156
rect 2836 4124 2840 4156
rect 2800 4076 2840 4124
rect 2800 4044 2804 4076
rect 2836 4044 2840 4076
rect 2800 3996 2840 4044
rect 2800 3964 2804 3996
rect 2836 3964 2840 3996
rect 2800 3916 2840 3964
rect 2800 3884 2804 3916
rect 2836 3884 2840 3916
rect 2800 3836 2840 3884
rect 2800 3804 2804 3836
rect 2836 3804 2840 3836
rect 2800 3756 2840 3804
rect 2800 3724 2804 3756
rect 2836 3724 2840 3756
rect 2800 3676 2840 3724
rect 2800 3644 2804 3676
rect 2836 3644 2840 3676
rect 2800 3640 2840 3644
rect 2880 4396 2920 4400
rect 2880 4364 2884 4396
rect 2916 4364 2920 4396
rect 2880 4316 2920 4364
rect 2880 4284 2884 4316
rect 2916 4284 2920 4316
rect 2880 4236 2920 4284
rect 2880 4204 2884 4236
rect 2916 4204 2920 4236
rect 2880 4156 2920 4204
rect 2880 4124 2884 4156
rect 2916 4124 2920 4156
rect 2880 4076 2920 4124
rect 2880 4044 2884 4076
rect 2916 4044 2920 4076
rect 2880 3996 2920 4044
rect 2880 3964 2884 3996
rect 2916 3964 2920 3996
rect 2880 3916 2920 3964
rect 2880 3884 2884 3916
rect 2916 3884 2920 3916
rect 2880 3836 2920 3884
rect 2880 3804 2884 3836
rect 2916 3804 2920 3836
rect 2880 3756 2920 3804
rect 2880 3724 2884 3756
rect 2916 3724 2920 3756
rect 2880 3676 2920 3724
rect 2880 3644 2884 3676
rect 2916 3644 2920 3676
rect 2880 3640 2920 3644
rect 2960 4396 3000 4400
rect 2960 4364 2964 4396
rect 2996 4364 3000 4396
rect 2960 4316 3000 4364
rect 2960 4284 2964 4316
rect 2996 4284 3000 4316
rect 2960 4236 3000 4284
rect 2960 4204 2964 4236
rect 2996 4204 3000 4236
rect 2960 4156 3000 4204
rect 2960 4124 2964 4156
rect 2996 4124 3000 4156
rect 2960 4076 3000 4124
rect 2960 4044 2964 4076
rect 2996 4044 3000 4076
rect 2960 3996 3000 4044
rect 2960 3964 2964 3996
rect 2996 3964 3000 3996
rect 2960 3916 3000 3964
rect 2960 3884 2964 3916
rect 2996 3884 3000 3916
rect 2960 3836 3000 3884
rect 2960 3804 2964 3836
rect 2996 3804 3000 3836
rect 2960 3756 3000 3804
rect 2960 3724 2964 3756
rect 2996 3724 3000 3756
rect 2960 3676 3000 3724
rect 2960 3644 2964 3676
rect 2996 3644 3000 3676
rect 2960 3640 3000 3644
rect 3040 4396 3080 4400
rect 3040 4364 3044 4396
rect 3076 4364 3080 4396
rect 3040 4316 3080 4364
rect 3040 4284 3044 4316
rect 3076 4284 3080 4316
rect 3040 4236 3080 4284
rect 3040 4204 3044 4236
rect 3076 4204 3080 4236
rect 3040 4156 3080 4204
rect 3040 4124 3044 4156
rect 3076 4124 3080 4156
rect 3040 4076 3080 4124
rect 3040 4044 3044 4076
rect 3076 4044 3080 4076
rect 3040 3996 3080 4044
rect 3040 3964 3044 3996
rect 3076 3964 3080 3996
rect 3040 3916 3080 3964
rect 3040 3884 3044 3916
rect 3076 3884 3080 3916
rect 3040 3836 3080 3884
rect 3040 3804 3044 3836
rect 3076 3804 3080 3836
rect 3040 3756 3080 3804
rect 3040 3724 3044 3756
rect 3076 3724 3080 3756
rect 3040 3676 3080 3724
rect 3040 3644 3044 3676
rect 3076 3644 3080 3676
rect 3040 3640 3080 3644
rect 3120 4396 3160 4400
rect 3120 4364 3124 4396
rect 3156 4364 3160 4396
rect 3120 4316 3160 4364
rect 3120 4284 3124 4316
rect 3156 4284 3160 4316
rect 3120 4236 3160 4284
rect 3120 4204 3124 4236
rect 3156 4204 3160 4236
rect 3120 4156 3160 4204
rect 3120 4124 3124 4156
rect 3156 4124 3160 4156
rect 3120 4076 3160 4124
rect 3120 4044 3124 4076
rect 3156 4044 3160 4076
rect 3120 3996 3160 4044
rect 3120 3964 3124 3996
rect 3156 3964 3160 3996
rect 3120 3916 3160 3964
rect 3120 3884 3124 3916
rect 3156 3884 3160 3916
rect 3120 3836 3160 3884
rect 3120 3804 3124 3836
rect 3156 3804 3160 3836
rect 3120 3756 3160 3804
rect 3120 3724 3124 3756
rect 3156 3724 3160 3756
rect 3120 3676 3160 3724
rect 3120 3644 3124 3676
rect 3156 3644 3160 3676
rect 3120 3640 3160 3644
rect 3200 4396 3240 4400
rect 3200 4364 3204 4396
rect 3236 4364 3240 4396
rect 3200 4316 3240 4364
rect 3200 4284 3204 4316
rect 3236 4284 3240 4316
rect 3200 4236 3240 4284
rect 3200 4204 3204 4236
rect 3236 4204 3240 4236
rect 3200 4156 3240 4204
rect 3200 4124 3204 4156
rect 3236 4124 3240 4156
rect 3200 4076 3240 4124
rect 3200 4044 3204 4076
rect 3236 4044 3240 4076
rect 3200 3996 3240 4044
rect 3200 3964 3204 3996
rect 3236 3964 3240 3996
rect 3200 3916 3240 3964
rect 3200 3884 3204 3916
rect 3236 3884 3240 3916
rect 3200 3836 3240 3884
rect 3200 3804 3204 3836
rect 3236 3804 3240 3836
rect 3200 3756 3240 3804
rect 3200 3724 3204 3756
rect 3236 3724 3240 3756
rect 3200 3676 3240 3724
rect 3200 3644 3204 3676
rect 3236 3644 3240 3676
rect 3200 3640 3240 3644
rect 3280 4396 3320 4400
rect 3280 4364 3284 4396
rect 3316 4364 3320 4396
rect 3280 4316 3320 4364
rect 3280 4284 3284 4316
rect 3316 4284 3320 4316
rect 3280 4236 3320 4284
rect 3280 4204 3284 4236
rect 3316 4204 3320 4236
rect 3280 4156 3320 4204
rect 3280 4124 3284 4156
rect 3316 4124 3320 4156
rect 3280 4076 3320 4124
rect 3280 4044 3284 4076
rect 3316 4044 3320 4076
rect 3280 3996 3320 4044
rect 3280 3964 3284 3996
rect 3316 3964 3320 3996
rect 3280 3916 3320 3964
rect 3280 3884 3284 3916
rect 3316 3884 3320 3916
rect 3280 3836 3320 3884
rect 3280 3804 3284 3836
rect 3316 3804 3320 3836
rect 3280 3756 3320 3804
rect 3280 3724 3284 3756
rect 3316 3724 3320 3756
rect 3280 3676 3320 3724
rect 3280 3644 3284 3676
rect 3316 3644 3320 3676
rect 3280 3640 3320 3644
rect 3360 4396 3400 4400
rect 3360 4364 3364 4396
rect 3396 4364 3400 4396
rect 3360 4316 3400 4364
rect 3360 4284 3364 4316
rect 3396 4284 3400 4316
rect 3360 4236 3400 4284
rect 3360 4204 3364 4236
rect 3396 4204 3400 4236
rect 3360 4156 3400 4204
rect 3360 4124 3364 4156
rect 3396 4124 3400 4156
rect 3360 4076 3400 4124
rect 3360 4044 3364 4076
rect 3396 4044 3400 4076
rect 3360 3996 3400 4044
rect 3360 3964 3364 3996
rect 3396 3964 3400 3996
rect 3360 3916 3400 3964
rect 3360 3884 3364 3916
rect 3396 3884 3400 3916
rect 3360 3836 3400 3884
rect 3360 3804 3364 3836
rect 3396 3804 3400 3836
rect 3360 3756 3400 3804
rect 3360 3724 3364 3756
rect 3396 3724 3400 3756
rect 3360 3676 3400 3724
rect 3360 3644 3364 3676
rect 3396 3644 3400 3676
rect 3360 3640 3400 3644
rect 3440 4396 3480 4400
rect 3440 4364 3444 4396
rect 3476 4364 3480 4396
rect 3440 4316 3480 4364
rect 3440 4284 3444 4316
rect 3476 4284 3480 4316
rect 3440 4236 3480 4284
rect 3440 4204 3444 4236
rect 3476 4204 3480 4236
rect 3440 4156 3480 4204
rect 3440 4124 3444 4156
rect 3476 4124 3480 4156
rect 3440 4076 3480 4124
rect 3440 4044 3444 4076
rect 3476 4044 3480 4076
rect 3440 3996 3480 4044
rect 3440 3964 3444 3996
rect 3476 3964 3480 3996
rect 3440 3916 3480 3964
rect 3440 3884 3444 3916
rect 3476 3884 3480 3916
rect 3440 3836 3480 3884
rect 3440 3804 3444 3836
rect 3476 3804 3480 3836
rect 3440 3756 3480 3804
rect 3440 3724 3444 3756
rect 3476 3724 3480 3756
rect 3440 3676 3480 3724
rect 3440 3644 3444 3676
rect 3476 3644 3480 3676
rect 3440 3640 3480 3644
rect 3520 4396 3560 4400
rect 3520 4364 3524 4396
rect 3556 4364 3560 4396
rect 3520 4316 3560 4364
rect 3520 4284 3524 4316
rect 3556 4284 3560 4316
rect 3520 4236 3560 4284
rect 3520 4204 3524 4236
rect 3556 4204 3560 4236
rect 3520 4156 3560 4204
rect 3520 4124 3524 4156
rect 3556 4124 3560 4156
rect 3520 4076 3560 4124
rect 3520 4044 3524 4076
rect 3556 4044 3560 4076
rect 3520 3996 3560 4044
rect 3520 3964 3524 3996
rect 3556 3964 3560 3996
rect 3520 3916 3560 3964
rect 3520 3884 3524 3916
rect 3556 3884 3560 3916
rect 3520 3836 3560 3884
rect 3520 3804 3524 3836
rect 3556 3804 3560 3836
rect 3520 3756 3560 3804
rect 3520 3724 3524 3756
rect 3556 3724 3560 3756
rect 3520 3676 3560 3724
rect 3520 3644 3524 3676
rect 3556 3644 3560 3676
rect 3520 3640 3560 3644
rect 3600 4396 3640 4400
rect 3600 4364 3604 4396
rect 3636 4364 3640 4396
rect 3600 4316 3640 4364
rect 3600 4284 3604 4316
rect 3636 4284 3640 4316
rect 3600 4236 3640 4284
rect 3600 4204 3604 4236
rect 3636 4204 3640 4236
rect 3600 4156 3640 4204
rect 3600 4124 3604 4156
rect 3636 4124 3640 4156
rect 3600 4076 3640 4124
rect 3600 4044 3604 4076
rect 3636 4044 3640 4076
rect 3600 3996 3640 4044
rect 3600 3964 3604 3996
rect 3636 3964 3640 3996
rect 3600 3916 3640 3964
rect 3600 3884 3604 3916
rect 3636 3884 3640 3916
rect 3600 3836 3640 3884
rect 3600 3804 3604 3836
rect 3636 3804 3640 3836
rect 3600 3756 3640 3804
rect 3600 3724 3604 3756
rect 3636 3724 3640 3756
rect 3600 3676 3640 3724
rect 3600 3644 3604 3676
rect 3636 3644 3640 3676
rect 3600 3640 3640 3644
rect 3680 4396 3720 4400
rect 3680 4364 3684 4396
rect 3716 4364 3720 4396
rect 3680 4316 3720 4364
rect 3680 4284 3684 4316
rect 3716 4284 3720 4316
rect 3680 4236 3720 4284
rect 3680 4204 3684 4236
rect 3716 4204 3720 4236
rect 3680 4156 3720 4204
rect 3680 4124 3684 4156
rect 3716 4124 3720 4156
rect 3680 4076 3720 4124
rect 3680 4044 3684 4076
rect 3716 4044 3720 4076
rect 3680 3996 3720 4044
rect 3680 3964 3684 3996
rect 3716 3964 3720 3996
rect 3680 3916 3720 3964
rect 3680 3884 3684 3916
rect 3716 3884 3720 3916
rect 3680 3836 3720 3884
rect 3680 3804 3684 3836
rect 3716 3804 3720 3836
rect 3680 3756 3720 3804
rect 3680 3724 3684 3756
rect 3716 3724 3720 3756
rect 3680 3676 3720 3724
rect 3680 3644 3684 3676
rect 3716 3644 3720 3676
rect 3680 3640 3720 3644
rect 3760 4396 3800 4400
rect 3760 4364 3764 4396
rect 3796 4364 3800 4396
rect 3760 4316 3800 4364
rect 3760 4284 3764 4316
rect 3796 4284 3800 4316
rect 3760 4236 3800 4284
rect 3760 4204 3764 4236
rect 3796 4204 3800 4236
rect 3760 4156 3800 4204
rect 3760 4124 3764 4156
rect 3796 4124 3800 4156
rect 3760 4076 3800 4124
rect 3760 4044 3764 4076
rect 3796 4044 3800 4076
rect 3760 3996 3800 4044
rect 3760 3964 3764 3996
rect 3796 3964 3800 3996
rect 3760 3916 3800 3964
rect 3760 3884 3764 3916
rect 3796 3884 3800 3916
rect 3760 3836 3800 3884
rect 3760 3804 3764 3836
rect 3796 3804 3800 3836
rect 3760 3756 3800 3804
rect 3760 3724 3764 3756
rect 3796 3724 3800 3756
rect 3760 3676 3800 3724
rect 3760 3644 3764 3676
rect 3796 3644 3800 3676
rect 3760 3640 3800 3644
rect 3840 4396 3880 4400
rect 3840 4364 3844 4396
rect 3876 4364 3880 4396
rect 3840 4316 3880 4364
rect 3840 4284 3844 4316
rect 3876 4284 3880 4316
rect 3840 4236 3880 4284
rect 3840 4204 3844 4236
rect 3876 4204 3880 4236
rect 3840 4156 3880 4204
rect 3840 4124 3844 4156
rect 3876 4124 3880 4156
rect 3840 4076 3880 4124
rect 3840 4044 3844 4076
rect 3876 4044 3880 4076
rect 3840 3996 3880 4044
rect 3840 3964 3844 3996
rect 3876 3964 3880 3996
rect 3840 3916 3880 3964
rect 3840 3884 3844 3916
rect 3876 3884 3880 3916
rect 3840 3836 3880 3884
rect 3840 3804 3844 3836
rect 3876 3804 3880 3836
rect 3840 3756 3880 3804
rect 3840 3724 3844 3756
rect 3876 3724 3880 3756
rect 3840 3676 3880 3724
rect 3840 3644 3844 3676
rect 3876 3644 3880 3676
rect 3840 3640 3880 3644
rect 3920 4396 3960 4400
rect 3920 4364 3924 4396
rect 3956 4364 3960 4396
rect 3920 4316 3960 4364
rect 3920 4284 3924 4316
rect 3956 4284 3960 4316
rect 3920 4236 3960 4284
rect 3920 4204 3924 4236
rect 3956 4204 3960 4236
rect 3920 4156 3960 4204
rect 3920 4124 3924 4156
rect 3956 4124 3960 4156
rect 3920 4076 3960 4124
rect 3920 4044 3924 4076
rect 3956 4044 3960 4076
rect 3920 3996 3960 4044
rect 3920 3964 3924 3996
rect 3956 3964 3960 3996
rect 3920 3916 3960 3964
rect 3920 3884 3924 3916
rect 3956 3884 3960 3916
rect 3920 3836 3960 3884
rect 3920 3804 3924 3836
rect 3956 3804 3960 3836
rect 3920 3756 3960 3804
rect 3920 3724 3924 3756
rect 3956 3724 3960 3756
rect 3920 3676 3960 3724
rect 3920 3644 3924 3676
rect 3956 3644 3960 3676
rect 3920 3640 3960 3644
rect 4000 4396 4040 4400
rect 4000 4364 4004 4396
rect 4036 4364 4040 4396
rect 4000 4316 4040 4364
rect 4000 4284 4004 4316
rect 4036 4284 4040 4316
rect 4000 4236 4040 4284
rect 4000 4204 4004 4236
rect 4036 4204 4040 4236
rect 4000 4156 4040 4204
rect 4000 4124 4004 4156
rect 4036 4124 4040 4156
rect 4000 4076 4040 4124
rect 4000 4044 4004 4076
rect 4036 4044 4040 4076
rect 4000 3996 4040 4044
rect 4000 3964 4004 3996
rect 4036 3964 4040 3996
rect 4000 3916 4040 3964
rect 4000 3884 4004 3916
rect 4036 3884 4040 3916
rect 4000 3836 4040 3884
rect 4000 3804 4004 3836
rect 4036 3804 4040 3836
rect 4000 3756 4040 3804
rect 4000 3724 4004 3756
rect 4036 3724 4040 3756
rect 4000 3676 4040 3724
rect 4000 3644 4004 3676
rect 4036 3644 4040 3676
rect 4000 3640 4040 3644
rect 4080 4396 4120 4400
rect 4080 4364 4084 4396
rect 4116 4364 4120 4396
rect 4080 4316 4120 4364
rect 4080 4284 4084 4316
rect 4116 4284 4120 4316
rect 4080 4236 4120 4284
rect 4080 4204 4084 4236
rect 4116 4204 4120 4236
rect 4080 4156 4120 4204
rect 4080 4124 4084 4156
rect 4116 4124 4120 4156
rect 4080 4076 4120 4124
rect 4080 4044 4084 4076
rect 4116 4044 4120 4076
rect 4080 3996 4120 4044
rect 4080 3964 4084 3996
rect 4116 3964 4120 3996
rect 4080 3916 4120 3964
rect 4080 3884 4084 3916
rect 4116 3884 4120 3916
rect 4080 3836 4120 3884
rect 4080 3804 4084 3836
rect 4116 3804 4120 3836
rect 4080 3756 4120 3804
rect 4080 3724 4084 3756
rect 4116 3724 4120 3756
rect 4080 3676 4120 3724
rect 4080 3644 4084 3676
rect 4116 3644 4120 3676
rect 4080 3640 4120 3644
rect 4160 4396 4200 4400
rect 4160 4364 4164 4396
rect 4196 4364 4200 4396
rect 4160 4316 4200 4364
rect 4160 4284 4164 4316
rect 4196 4284 4200 4316
rect 4160 4236 4200 4284
rect 4160 4204 4164 4236
rect 4196 4204 4200 4236
rect 4160 4156 4200 4204
rect 4160 4124 4164 4156
rect 4196 4124 4200 4156
rect 4160 4076 4200 4124
rect 4160 4044 4164 4076
rect 4196 4044 4200 4076
rect 4160 3996 4200 4044
rect 4160 3964 4164 3996
rect 4196 3964 4200 3996
rect 4160 3916 4200 3964
rect 4160 3884 4164 3916
rect 4196 3884 4200 3916
rect 4160 3836 4200 3884
rect 4160 3804 4164 3836
rect 4196 3804 4200 3836
rect 4160 3756 4200 3804
rect 4160 3724 4164 3756
rect 4196 3724 4200 3756
rect 4160 3676 4200 3724
rect 4160 3644 4164 3676
rect 4196 3644 4200 3676
rect 4160 3640 4200 3644
rect 4240 4396 4280 4400
rect 4240 4364 4244 4396
rect 4276 4364 4280 4396
rect 4240 4316 4280 4364
rect 4240 4284 4244 4316
rect 4276 4284 4280 4316
rect 4240 4236 4280 4284
rect 4240 4204 4244 4236
rect 4276 4204 4280 4236
rect 4240 4156 4280 4204
rect 4240 4124 4244 4156
rect 4276 4124 4280 4156
rect 4240 4076 4280 4124
rect 4240 4044 4244 4076
rect 4276 4044 4280 4076
rect 4240 3996 4280 4044
rect 4240 3964 4244 3996
rect 4276 3964 4280 3996
rect 4240 3916 4280 3964
rect 4240 3884 4244 3916
rect 4276 3884 4280 3916
rect 4240 3836 4280 3884
rect 4240 3804 4244 3836
rect 4276 3804 4280 3836
rect 4240 3756 4280 3804
rect 4240 3724 4244 3756
rect 4276 3724 4280 3756
rect 4240 3676 4280 3724
rect 4240 3644 4244 3676
rect 4276 3644 4280 3676
rect 4240 3640 4280 3644
rect 4320 4396 4360 4400
rect 4320 4364 4324 4396
rect 4356 4364 4360 4396
rect 4320 4316 4360 4364
rect 4320 4284 4324 4316
rect 4356 4284 4360 4316
rect 4320 4236 4360 4284
rect 4320 4204 4324 4236
rect 4356 4204 4360 4236
rect 4320 4156 4360 4204
rect 4320 4124 4324 4156
rect 4356 4124 4360 4156
rect 4320 4076 4360 4124
rect 4320 4044 4324 4076
rect 4356 4044 4360 4076
rect 4320 3996 4360 4044
rect 4320 3964 4324 3996
rect 4356 3964 4360 3996
rect 4320 3916 4360 3964
rect 4320 3884 4324 3916
rect 4356 3884 4360 3916
rect 4320 3836 4360 3884
rect 4320 3804 4324 3836
rect 4356 3804 4360 3836
rect 4320 3756 4360 3804
rect 4320 3724 4324 3756
rect 4356 3724 4360 3756
rect 4320 3676 4360 3724
rect 4320 3644 4324 3676
rect 4356 3644 4360 3676
rect 4320 3640 4360 3644
rect 4400 4396 4440 4400
rect 4400 4364 4404 4396
rect 4436 4364 4440 4396
rect 4400 4316 4440 4364
rect 4400 4284 4404 4316
rect 4436 4284 4440 4316
rect 4400 4236 4440 4284
rect 4400 4204 4404 4236
rect 4436 4204 4440 4236
rect 4400 4156 4440 4204
rect 4400 4124 4404 4156
rect 4436 4124 4440 4156
rect 4400 4076 4440 4124
rect 4400 4044 4404 4076
rect 4436 4044 4440 4076
rect 4400 3996 4440 4044
rect 4400 3964 4404 3996
rect 4436 3964 4440 3996
rect 4400 3916 4440 3964
rect 4400 3884 4404 3916
rect 4436 3884 4440 3916
rect 4400 3836 4440 3884
rect 4400 3804 4404 3836
rect 4436 3804 4440 3836
rect 4400 3756 4440 3804
rect 4400 3724 4404 3756
rect 4436 3724 4440 3756
rect 4400 3676 4440 3724
rect 4400 3644 4404 3676
rect 4436 3644 4440 3676
rect 4400 3640 4440 3644
rect 4480 4396 4520 4400
rect 4480 4364 4484 4396
rect 4516 4364 4520 4396
rect 4480 4316 4520 4364
rect 4480 4284 4484 4316
rect 4516 4284 4520 4316
rect 4480 4236 4520 4284
rect 4480 4204 4484 4236
rect 4516 4204 4520 4236
rect 4480 4156 4520 4204
rect 4480 4124 4484 4156
rect 4516 4124 4520 4156
rect 4480 4076 4520 4124
rect 4480 4044 4484 4076
rect 4516 4044 4520 4076
rect 4480 3996 4520 4044
rect 4480 3964 4484 3996
rect 4516 3964 4520 3996
rect 4480 3916 4520 3964
rect 4480 3884 4484 3916
rect 4516 3884 4520 3916
rect 4480 3836 4520 3884
rect 4480 3804 4484 3836
rect 4516 3804 4520 3836
rect 4480 3756 4520 3804
rect 4480 3724 4484 3756
rect 4516 3724 4520 3756
rect 4480 3676 4520 3724
rect 4480 3644 4484 3676
rect 4516 3644 4520 3676
rect 4480 3640 4520 3644
rect 4560 4396 4600 4400
rect 4560 4364 4564 4396
rect 4596 4364 4600 4396
rect 4560 4316 4600 4364
rect 4560 4284 4564 4316
rect 4596 4284 4600 4316
rect 4560 4236 4600 4284
rect 4560 4204 4564 4236
rect 4596 4204 4600 4236
rect 4560 4156 4600 4204
rect 4560 4124 4564 4156
rect 4596 4124 4600 4156
rect 4560 4076 4600 4124
rect 4560 4044 4564 4076
rect 4596 4044 4600 4076
rect 4560 3996 4600 4044
rect 4560 3964 4564 3996
rect 4596 3964 4600 3996
rect 4560 3916 4600 3964
rect 4560 3884 4564 3916
rect 4596 3884 4600 3916
rect 4560 3836 4600 3884
rect 4560 3804 4564 3836
rect 4596 3804 4600 3836
rect 4560 3756 4600 3804
rect 4560 3724 4564 3756
rect 4596 3724 4600 3756
rect 4560 3676 4600 3724
rect 4560 3644 4564 3676
rect 4596 3644 4600 3676
rect 4560 3640 4600 3644
rect 4640 4396 4680 4400
rect 4640 4364 4644 4396
rect 4676 4364 4680 4396
rect 4640 4316 4680 4364
rect 4640 4284 4644 4316
rect 4676 4284 4680 4316
rect 4640 4236 4680 4284
rect 4640 4204 4644 4236
rect 4676 4204 4680 4236
rect 4640 4156 4680 4204
rect 4640 4124 4644 4156
rect 4676 4124 4680 4156
rect 4640 4076 4680 4124
rect 4640 4044 4644 4076
rect 4676 4044 4680 4076
rect 4640 3996 4680 4044
rect 4640 3964 4644 3996
rect 4676 3964 4680 3996
rect 4640 3916 4680 3964
rect 4640 3884 4644 3916
rect 4676 3884 4680 3916
rect 4640 3836 4680 3884
rect 4640 3804 4644 3836
rect 4676 3804 4680 3836
rect 4640 3756 4680 3804
rect 4640 3724 4644 3756
rect 4676 3724 4680 3756
rect 4640 3676 4680 3724
rect 4640 3644 4644 3676
rect 4676 3644 4680 3676
rect 4640 3640 4680 3644
rect 4720 4396 4760 4400
rect 4720 4364 4724 4396
rect 4756 4364 4760 4396
rect 4720 4316 4760 4364
rect 4720 4284 4724 4316
rect 4756 4284 4760 4316
rect 4720 4236 4760 4284
rect 4720 4204 4724 4236
rect 4756 4204 4760 4236
rect 4720 4156 4760 4204
rect 4720 4124 4724 4156
rect 4756 4124 4760 4156
rect 4720 4076 4760 4124
rect 4720 4044 4724 4076
rect 4756 4044 4760 4076
rect 4720 3996 4760 4044
rect 4720 3964 4724 3996
rect 4756 3964 4760 3996
rect 4720 3916 4760 3964
rect 4720 3884 4724 3916
rect 4756 3884 4760 3916
rect 4720 3836 4760 3884
rect 4720 3804 4724 3836
rect 4756 3804 4760 3836
rect 4720 3756 4760 3804
rect 4720 3724 4724 3756
rect 4756 3724 4760 3756
rect 4720 3676 4760 3724
rect 4720 3644 4724 3676
rect 4756 3644 4760 3676
rect 4720 3640 4760 3644
rect 4800 4396 4840 4400
rect 4800 4364 4804 4396
rect 4836 4364 4840 4396
rect 4800 4316 4840 4364
rect 4800 4284 4804 4316
rect 4836 4284 4840 4316
rect 4800 4236 4840 4284
rect 4800 4204 4804 4236
rect 4836 4204 4840 4236
rect 4800 4156 4840 4204
rect 4800 4124 4804 4156
rect 4836 4124 4840 4156
rect 4800 4076 4840 4124
rect 4800 4044 4804 4076
rect 4836 4044 4840 4076
rect 4800 3996 4840 4044
rect 4800 3964 4804 3996
rect 4836 3964 4840 3996
rect 4800 3916 4840 3964
rect 4800 3884 4804 3916
rect 4836 3884 4840 3916
rect 4800 3836 4840 3884
rect 4800 3804 4804 3836
rect 4836 3804 4840 3836
rect 4800 3756 4840 3804
rect 4800 3724 4804 3756
rect 4836 3724 4840 3756
rect 4800 3676 4840 3724
rect 4800 3644 4804 3676
rect 4836 3644 4840 3676
rect 4800 3640 4840 3644
rect 4880 4396 4920 4444
rect 4880 4364 4884 4396
rect 4916 4364 4920 4396
rect 4880 4316 4920 4364
rect 4880 4284 4884 4316
rect 4916 4284 4920 4316
rect 4880 4236 4920 4284
rect 4880 4204 4884 4236
rect 4916 4204 4920 4236
rect 4880 4156 4920 4204
rect 4880 4124 4884 4156
rect 4916 4124 4920 4156
rect 4880 4076 4920 4124
rect 4880 4044 4884 4076
rect 4916 4044 4920 4076
rect 4880 3996 4920 4044
rect 4880 3964 4884 3996
rect 4916 3964 4920 3996
rect 4880 3916 4920 3964
rect 4880 3884 4884 3916
rect 4916 3884 4920 3916
rect 4880 3836 4920 3884
rect 4880 3804 4884 3836
rect 4916 3804 4920 3836
rect 4880 3756 4920 3804
rect 4880 3724 4884 3756
rect 4916 3724 4920 3756
rect 4880 3676 4920 3724
rect 4880 3644 4884 3676
rect 4916 3644 4920 3676
rect -880 3564 -876 3596
rect -844 3564 -840 3596
rect -880 3516 -840 3564
rect -880 3484 -876 3516
rect -844 3484 -840 3516
rect -880 3436 -840 3484
rect -880 3404 -876 3436
rect -844 3404 -840 3436
rect -880 3356 -840 3404
rect -880 3324 -876 3356
rect -844 3324 -840 3356
rect -880 3276 -840 3324
rect -880 3244 -876 3276
rect -844 3244 -840 3276
rect -880 3196 -840 3244
rect -880 3164 -876 3196
rect -844 3164 -840 3196
rect -880 3116 -840 3164
rect -880 3084 -876 3116
rect -844 3084 -840 3116
rect -880 3036 -840 3084
rect -880 3004 -876 3036
rect -844 3004 -840 3036
rect -880 2956 -840 3004
rect -880 2924 -876 2956
rect -844 2924 -840 2956
rect -880 2876 -840 2924
rect -880 2844 -876 2876
rect -844 2844 -840 2876
rect -880 2796 -840 2844
rect -880 2764 -876 2796
rect -844 2764 -840 2796
rect -880 2716 -840 2764
rect -880 2684 -876 2716
rect -844 2684 -840 2716
rect -880 2636 -840 2684
rect -880 2604 -876 2636
rect -844 2604 -840 2636
rect -880 2556 -840 2604
rect -880 2524 -876 2556
rect -844 2524 -840 2556
rect -880 2476 -840 2524
rect -800 3596 -760 3600
rect -800 3564 -796 3596
rect -764 3564 -760 3596
rect -800 3516 -760 3564
rect -800 3484 -796 3516
rect -764 3484 -760 3516
rect -800 3436 -760 3484
rect -800 3404 -796 3436
rect -764 3404 -760 3436
rect -800 3356 -760 3404
rect -800 3324 -796 3356
rect -764 3324 -760 3356
rect -800 3276 -760 3324
rect -800 3244 -796 3276
rect -764 3244 -760 3276
rect -800 3196 -760 3244
rect -800 3164 -796 3196
rect -764 3164 -760 3196
rect -800 3116 -760 3164
rect -800 3084 -796 3116
rect -764 3084 -760 3116
rect -800 3036 -760 3084
rect -800 3004 -796 3036
rect -764 3004 -760 3036
rect -800 2956 -760 3004
rect -800 2924 -796 2956
rect -764 2924 -760 2956
rect -800 2876 -760 2924
rect -800 2844 -796 2876
rect -764 2844 -760 2876
rect -800 2796 -760 2844
rect -800 2764 -796 2796
rect -764 2764 -760 2796
rect -800 2716 -760 2764
rect -800 2684 -796 2716
rect -764 2684 -760 2716
rect -800 2636 -760 2684
rect -800 2604 -796 2636
rect -764 2604 -760 2636
rect -800 2556 -760 2604
rect -800 2524 -796 2556
rect -764 2524 -760 2556
rect -800 2520 -760 2524
rect -720 3596 -680 3600
rect -720 3564 -716 3596
rect -684 3564 -680 3596
rect -720 3516 -680 3564
rect -720 3484 -716 3516
rect -684 3484 -680 3516
rect -720 3436 -680 3484
rect -720 3404 -716 3436
rect -684 3404 -680 3436
rect -720 3356 -680 3404
rect -720 3324 -716 3356
rect -684 3324 -680 3356
rect -720 3276 -680 3324
rect -720 3244 -716 3276
rect -684 3244 -680 3276
rect -720 3196 -680 3244
rect -720 3164 -716 3196
rect -684 3164 -680 3196
rect -720 3116 -680 3164
rect -720 3084 -716 3116
rect -684 3084 -680 3116
rect -720 3036 -680 3084
rect -720 3004 -716 3036
rect -684 3004 -680 3036
rect -720 2956 -680 3004
rect -720 2924 -716 2956
rect -684 2924 -680 2956
rect -720 2876 -680 2924
rect -720 2844 -716 2876
rect -684 2844 -680 2876
rect -720 2796 -680 2844
rect -720 2764 -716 2796
rect -684 2764 -680 2796
rect -720 2716 -680 2764
rect -720 2684 -716 2716
rect -684 2684 -680 2716
rect -720 2636 -680 2684
rect -720 2604 -716 2636
rect -684 2604 -680 2636
rect -720 2556 -680 2604
rect -720 2524 -716 2556
rect -684 2524 -680 2556
rect -720 2520 -680 2524
rect -640 3596 -600 3600
rect -640 3564 -636 3596
rect -604 3564 -600 3596
rect -640 3516 -600 3564
rect -640 3484 -636 3516
rect -604 3484 -600 3516
rect -640 3436 -600 3484
rect -640 3404 -636 3436
rect -604 3404 -600 3436
rect -640 3356 -600 3404
rect -640 3324 -636 3356
rect -604 3324 -600 3356
rect -640 3276 -600 3324
rect -640 3244 -636 3276
rect -604 3244 -600 3276
rect -640 3196 -600 3244
rect -640 3164 -636 3196
rect -604 3164 -600 3196
rect -640 3116 -600 3164
rect -640 3084 -636 3116
rect -604 3084 -600 3116
rect -640 3036 -600 3084
rect -640 3004 -636 3036
rect -604 3004 -600 3036
rect -640 2956 -600 3004
rect -640 2924 -636 2956
rect -604 2924 -600 2956
rect -640 2876 -600 2924
rect -640 2844 -636 2876
rect -604 2844 -600 2876
rect -640 2796 -600 2844
rect -640 2764 -636 2796
rect -604 2764 -600 2796
rect -640 2716 -600 2764
rect -640 2684 -636 2716
rect -604 2684 -600 2716
rect -640 2636 -600 2684
rect -640 2604 -636 2636
rect -604 2604 -600 2636
rect -640 2556 -600 2604
rect -640 2524 -636 2556
rect -604 2524 -600 2556
rect -640 2520 -600 2524
rect -560 3596 -520 3600
rect -560 3564 -556 3596
rect -524 3564 -520 3596
rect -560 3516 -520 3564
rect -560 3484 -556 3516
rect -524 3484 -520 3516
rect -560 3436 -520 3484
rect -560 3404 -556 3436
rect -524 3404 -520 3436
rect -560 3356 -520 3404
rect -560 3324 -556 3356
rect -524 3324 -520 3356
rect -560 3276 -520 3324
rect -560 3244 -556 3276
rect -524 3244 -520 3276
rect -560 3196 -520 3244
rect -560 3164 -556 3196
rect -524 3164 -520 3196
rect -560 3116 -520 3164
rect -560 3084 -556 3116
rect -524 3084 -520 3116
rect -560 3036 -520 3084
rect -560 3004 -556 3036
rect -524 3004 -520 3036
rect -560 2956 -520 3004
rect -560 2924 -556 2956
rect -524 2924 -520 2956
rect -560 2876 -520 2924
rect -560 2844 -556 2876
rect -524 2844 -520 2876
rect -560 2796 -520 2844
rect -560 2764 -556 2796
rect -524 2764 -520 2796
rect -560 2716 -520 2764
rect -560 2684 -556 2716
rect -524 2684 -520 2716
rect -560 2636 -520 2684
rect -560 2604 -556 2636
rect -524 2604 -520 2636
rect -560 2556 -520 2604
rect -560 2524 -556 2556
rect -524 2524 -520 2556
rect -560 2520 -520 2524
rect -480 3596 -440 3600
rect -480 3564 -476 3596
rect -444 3564 -440 3596
rect -480 3516 -440 3564
rect -480 3484 -476 3516
rect -444 3484 -440 3516
rect -480 3436 -440 3484
rect -480 3404 -476 3436
rect -444 3404 -440 3436
rect -480 3356 -440 3404
rect -480 3324 -476 3356
rect -444 3324 -440 3356
rect -480 3276 -440 3324
rect -480 3244 -476 3276
rect -444 3244 -440 3276
rect -480 3196 -440 3244
rect -480 3164 -476 3196
rect -444 3164 -440 3196
rect -480 3116 -440 3164
rect -480 3084 -476 3116
rect -444 3084 -440 3116
rect -480 3036 -440 3084
rect -480 3004 -476 3036
rect -444 3004 -440 3036
rect -480 2956 -440 3004
rect -480 2924 -476 2956
rect -444 2924 -440 2956
rect -480 2876 -440 2924
rect -480 2844 -476 2876
rect -444 2844 -440 2876
rect -480 2796 -440 2844
rect -480 2764 -476 2796
rect -444 2764 -440 2796
rect -480 2716 -440 2764
rect -480 2684 -476 2716
rect -444 2684 -440 2716
rect -480 2636 -440 2684
rect -480 2604 -476 2636
rect -444 2604 -440 2636
rect -480 2556 -440 2604
rect -480 2524 -476 2556
rect -444 2524 -440 2556
rect -480 2520 -440 2524
rect -400 3596 -360 3600
rect -400 3564 -396 3596
rect -364 3564 -360 3596
rect -400 3516 -360 3564
rect -400 3484 -396 3516
rect -364 3484 -360 3516
rect -400 3436 -360 3484
rect -400 3404 -396 3436
rect -364 3404 -360 3436
rect -400 3356 -360 3404
rect -400 3324 -396 3356
rect -364 3324 -360 3356
rect -400 3276 -360 3324
rect -400 3244 -396 3276
rect -364 3244 -360 3276
rect -400 3196 -360 3244
rect -400 3164 -396 3196
rect -364 3164 -360 3196
rect -400 3116 -360 3164
rect -400 3084 -396 3116
rect -364 3084 -360 3116
rect -400 3036 -360 3084
rect -400 3004 -396 3036
rect -364 3004 -360 3036
rect -400 2956 -360 3004
rect -400 2924 -396 2956
rect -364 2924 -360 2956
rect -400 2876 -360 2924
rect -400 2844 -396 2876
rect -364 2844 -360 2876
rect -400 2796 -360 2844
rect -400 2764 -396 2796
rect -364 2764 -360 2796
rect -400 2716 -360 2764
rect -400 2684 -396 2716
rect -364 2684 -360 2716
rect -400 2636 -360 2684
rect -400 2604 -396 2636
rect -364 2604 -360 2636
rect -400 2556 -360 2604
rect -400 2524 -396 2556
rect -364 2524 -360 2556
rect -400 2520 -360 2524
rect -320 3596 -280 3600
rect -320 3564 -316 3596
rect -284 3564 -280 3596
rect -320 3516 -280 3564
rect -320 3484 -316 3516
rect -284 3484 -280 3516
rect -320 3436 -280 3484
rect -320 3404 -316 3436
rect -284 3404 -280 3436
rect -320 3356 -280 3404
rect -320 3324 -316 3356
rect -284 3324 -280 3356
rect -320 3276 -280 3324
rect -320 3244 -316 3276
rect -284 3244 -280 3276
rect -320 3196 -280 3244
rect -320 3164 -316 3196
rect -284 3164 -280 3196
rect -320 3116 -280 3164
rect -320 3084 -316 3116
rect -284 3084 -280 3116
rect -320 3036 -280 3084
rect -320 3004 -316 3036
rect -284 3004 -280 3036
rect -320 2956 -280 3004
rect -320 2924 -316 2956
rect -284 2924 -280 2956
rect -320 2876 -280 2924
rect -320 2844 -316 2876
rect -284 2844 -280 2876
rect -320 2796 -280 2844
rect -320 2764 -316 2796
rect -284 2764 -280 2796
rect -320 2716 -280 2764
rect -320 2684 -316 2716
rect -284 2684 -280 2716
rect -320 2636 -280 2684
rect -320 2604 -316 2636
rect -284 2604 -280 2636
rect -320 2556 -280 2604
rect -320 2524 -316 2556
rect -284 2524 -280 2556
rect -320 2520 -280 2524
rect -240 3596 -200 3600
rect -240 3564 -236 3596
rect -204 3564 -200 3596
rect -240 3516 -200 3564
rect -240 3484 -236 3516
rect -204 3484 -200 3516
rect -240 3436 -200 3484
rect -240 3404 -236 3436
rect -204 3404 -200 3436
rect -240 3356 -200 3404
rect -240 3324 -236 3356
rect -204 3324 -200 3356
rect -240 3276 -200 3324
rect -240 3244 -236 3276
rect -204 3244 -200 3276
rect -240 3196 -200 3244
rect -240 3164 -236 3196
rect -204 3164 -200 3196
rect -240 3116 -200 3164
rect -240 3084 -236 3116
rect -204 3084 -200 3116
rect -240 3036 -200 3084
rect -240 3004 -236 3036
rect -204 3004 -200 3036
rect -240 2956 -200 3004
rect -240 2924 -236 2956
rect -204 2924 -200 2956
rect -240 2876 -200 2924
rect -240 2844 -236 2876
rect -204 2844 -200 2876
rect -240 2796 -200 2844
rect -240 2764 -236 2796
rect -204 2764 -200 2796
rect -240 2716 -200 2764
rect -240 2684 -236 2716
rect -204 2684 -200 2716
rect -240 2636 -200 2684
rect -240 2604 -236 2636
rect -204 2604 -200 2636
rect -240 2556 -200 2604
rect -240 2524 -236 2556
rect -204 2524 -200 2556
rect -240 2520 -200 2524
rect -160 3596 -120 3600
rect -160 3564 -156 3596
rect -124 3564 -120 3596
rect -160 3516 -120 3564
rect -160 3484 -156 3516
rect -124 3484 -120 3516
rect -160 3436 -120 3484
rect -160 3404 -156 3436
rect -124 3404 -120 3436
rect -160 3356 -120 3404
rect -160 3324 -156 3356
rect -124 3324 -120 3356
rect -160 3276 -120 3324
rect -160 3244 -156 3276
rect -124 3244 -120 3276
rect -160 3196 -120 3244
rect -160 3164 -156 3196
rect -124 3164 -120 3196
rect -160 3116 -120 3164
rect -160 3084 -156 3116
rect -124 3084 -120 3116
rect -160 3036 -120 3084
rect -160 3004 -156 3036
rect -124 3004 -120 3036
rect -160 2956 -120 3004
rect -160 2924 -156 2956
rect -124 2924 -120 2956
rect -160 2876 -120 2924
rect -160 2844 -156 2876
rect -124 2844 -120 2876
rect -160 2796 -120 2844
rect -160 2764 -156 2796
rect -124 2764 -120 2796
rect -160 2716 -120 2764
rect -160 2684 -156 2716
rect -124 2684 -120 2716
rect -160 2636 -120 2684
rect -160 2604 -156 2636
rect -124 2604 -120 2636
rect -160 2556 -120 2604
rect -160 2524 -156 2556
rect -124 2524 -120 2556
rect -160 2520 -120 2524
rect -80 3596 -40 3600
rect -80 3564 -76 3596
rect -44 3564 -40 3596
rect -80 3516 -40 3564
rect -80 3484 -76 3516
rect -44 3484 -40 3516
rect -80 3436 -40 3484
rect -80 3404 -76 3436
rect -44 3404 -40 3436
rect -80 3356 -40 3404
rect -80 3324 -76 3356
rect -44 3324 -40 3356
rect -80 3276 -40 3324
rect -80 3244 -76 3276
rect -44 3244 -40 3276
rect -80 3196 -40 3244
rect -80 3164 -76 3196
rect -44 3164 -40 3196
rect -80 3116 -40 3164
rect -80 3084 -76 3116
rect -44 3084 -40 3116
rect -80 3036 -40 3084
rect -80 3004 -76 3036
rect -44 3004 -40 3036
rect -80 2956 -40 3004
rect -80 2924 -76 2956
rect -44 2924 -40 2956
rect -80 2876 -40 2924
rect -80 2844 -76 2876
rect -44 2844 -40 2876
rect -80 2796 -40 2844
rect -80 2764 -76 2796
rect -44 2764 -40 2796
rect -80 2716 -40 2764
rect -80 2684 -76 2716
rect -44 2684 -40 2716
rect -80 2636 -40 2684
rect -80 2604 -76 2636
rect -44 2604 -40 2636
rect -80 2556 -40 2604
rect -80 2524 -76 2556
rect -44 2524 -40 2556
rect -80 2520 -40 2524
rect 0 3596 40 3600
rect 0 3564 4 3596
rect 36 3564 40 3596
rect 0 3516 40 3564
rect 0 3484 4 3516
rect 36 3484 40 3516
rect 0 3436 40 3484
rect 0 3404 4 3436
rect 36 3404 40 3436
rect 0 3356 40 3404
rect 0 3324 4 3356
rect 36 3324 40 3356
rect 0 3276 40 3324
rect 0 3244 4 3276
rect 36 3244 40 3276
rect 0 3196 40 3244
rect 0 3164 4 3196
rect 36 3164 40 3196
rect 0 3116 40 3164
rect 0 3084 4 3116
rect 36 3084 40 3116
rect 0 3036 40 3084
rect 0 3004 4 3036
rect 36 3004 40 3036
rect 0 2956 40 3004
rect 0 2924 4 2956
rect 36 2924 40 2956
rect 0 2876 40 2924
rect 0 2844 4 2876
rect 36 2844 40 2876
rect 0 2796 40 2844
rect 0 2764 4 2796
rect 36 2764 40 2796
rect 0 2716 40 2764
rect 0 2684 4 2716
rect 36 2684 40 2716
rect 0 2636 40 2684
rect 0 2604 4 2636
rect 36 2604 40 2636
rect 0 2556 40 2604
rect 0 2524 4 2556
rect 36 2524 40 2556
rect 0 2520 40 2524
rect 80 3596 120 3600
rect 80 3564 84 3596
rect 116 3564 120 3596
rect 80 3516 120 3564
rect 80 3484 84 3516
rect 116 3484 120 3516
rect 80 3436 120 3484
rect 80 3404 84 3436
rect 116 3404 120 3436
rect 80 3356 120 3404
rect 80 3324 84 3356
rect 116 3324 120 3356
rect 80 3276 120 3324
rect 80 3244 84 3276
rect 116 3244 120 3276
rect 80 3196 120 3244
rect 80 3164 84 3196
rect 116 3164 120 3196
rect 80 3116 120 3164
rect 80 3084 84 3116
rect 116 3084 120 3116
rect 80 3036 120 3084
rect 80 3004 84 3036
rect 116 3004 120 3036
rect 80 2956 120 3004
rect 80 2924 84 2956
rect 116 2924 120 2956
rect 80 2876 120 2924
rect 80 2844 84 2876
rect 116 2844 120 2876
rect 80 2796 120 2844
rect 80 2764 84 2796
rect 116 2764 120 2796
rect 80 2716 120 2764
rect 80 2684 84 2716
rect 116 2684 120 2716
rect 80 2636 120 2684
rect 80 2604 84 2636
rect 116 2604 120 2636
rect 80 2556 120 2604
rect 80 2524 84 2556
rect 116 2524 120 2556
rect 80 2520 120 2524
rect 160 3596 200 3600
rect 160 3564 164 3596
rect 196 3564 200 3596
rect 160 3516 200 3564
rect 160 3484 164 3516
rect 196 3484 200 3516
rect 160 3436 200 3484
rect 160 3404 164 3436
rect 196 3404 200 3436
rect 160 3356 200 3404
rect 160 3324 164 3356
rect 196 3324 200 3356
rect 160 3276 200 3324
rect 160 3244 164 3276
rect 196 3244 200 3276
rect 160 3196 200 3244
rect 160 3164 164 3196
rect 196 3164 200 3196
rect 160 3116 200 3164
rect 160 3084 164 3116
rect 196 3084 200 3116
rect 160 3036 200 3084
rect 160 3004 164 3036
rect 196 3004 200 3036
rect 160 2956 200 3004
rect 160 2924 164 2956
rect 196 2924 200 2956
rect 160 2876 200 2924
rect 160 2844 164 2876
rect 196 2844 200 2876
rect 160 2796 200 2844
rect 160 2764 164 2796
rect 196 2764 200 2796
rect 160 2716 200 2764
rect 160 2684 164 2716
rect 196 2684 200 2716
rect 160 2636 200 2684
rect 160 2604 164 2636
rect 196 2604 200 2636
rect 160 2556 200 2604
rect 160 2524 164 2556
rect 196 2524 200 2556
rect 160 2520 200 2524
rect 240 3596 280 3600
rect 240 3564 244 3596
rect 276 3564 280 3596
rect 240 3516 280 3564
rect 240 3484 244 3516
rect 276 3484 280 3516
rect 240 3436 280 3484
rect 240 3404 244 3436
rect 276 3404 280 3436
rect 240 3356 280 3404
rect 240 3324 244 3356
rect 276 3324 280 3356
rect 240 3276 280 3324
rect 240 3244 244 3276
rect 276 3244 280 3276
rect 240 3196 280 3244
rect 240 3164 244 3196
rect 276 3164 280 3196
rect 240 3116 280 3164
rect 240 3084 244 3116
rect 276 3084 280 3116
rect 240 3036 280 3084
rect 240 3004 244 3036
rect 276 3004 280 3036
rect 240 2956 280 3004
rect 240 2924 244 2956
rect 276 2924 280 2956
rect 240 2876 280 2924
rect 240 2844 244 2876
rect 276 2844 280 2876
rect 240 2796 280 2844
rect 240 2764 244 2796
rect 276 2764 280 2796
rect 240 2716 280 2764
rect 240 2684 244 2716
rect 276 2684 280 2716
rect 240 2636 280 2684
rect 240 2604 244 2636
rect 276 2604 280 2636
rect 240 2556 280 2604
rect 240 2524 244 2556
rect 276 2524 280 2556
rect 240 2520 280 2524
rect 320 3596 360 3600
rect 320 3564 324 3596
rect 356 3564 360 3596
rect 320 3516 360 3564
rect 320 3484 324 3516
rect 356 3484 360 3516
rect 320 3436 360 3484
rect 320 3404 324 3436
rect 356 3404 360 3436
rect 320 3356 360 3404
rect 320 3324 324 3356
rect 356 3324 360 3356
rect 320 3276 360 3324
rect 320 3244 324 3276
rect 356 3244 360 3276
rect 320 3196 360 3244
rect 320 3164 324 3196
rect 356 3164 360 3196
rect 320 3116 360 3164
rect 320 3084 324 3116
rect 356 3084 360 3116
rect 320 3036 360 3084
rect 320 3004 324 3036
rect 356 3004 360 3036
rect 320 2956 360 3004
rect 320 2924 324 2956
rect 356 2924 360 2956
rect 320 2876 360 2924
rect 320 2844 324 2876
rect 356 2844 360 2876
rect 320 2796 360 2844
rect 320 2764 324 2796
rect 356 2764 360 2796
rect 320 2716 360 2764
rect 320 2684 324 2716
rect 356 2684 360 2716
rect 320 2636 360 2684
rect 320 2604 324 2636
rect 356 2604 360 2636
rect 320 2556 360 2604
rect 320 2524 324 2556
rect 356 2524 360 2556
rect 320 2520 360 2524
rect 400 3596 440 3600
rect 400 3564 404 3596
rect 436 3564 440 3596
rect 400 3516 440 3564
rect 400 3484 404 3516
rect 436 3484 440 3516
rect 400 3436 440 3484
rect 400 3404 404 3436
rect 436 3404 440 3436
rect 400 3356 440 3404
rect 400 3324 404 3356
rect 436 3324 440 3356
rect 400 3276 440 3324
rect 400 3244 404 3276
rect 436 3244 440 3276
rect 400 3196 440 3244
rect 400 3164 404 3196
rect 436 3164 440 3196
rect 400 3116 440 3164
rect 400 3084 404 3116
rect 436 3084 440 3116
rect 400 3036 440 3084
rect 400 3004 404 3036
rect 436 3004 440 3036
rect 400 2956 440 3004
rect 400 2924 404 2956
rect 436 2924 440 2956
rect 400 2876 440 2924
rect 400 2844 404 2876
rect 436 2844 440 2876
rect 400 2796 440 2844
rect 400 2764 404 2796
rect 436 2764 440 2796
rect 400 2716 440 2764
rect 400 2684 404 2716
rect 436 2684 440 2716
rect 400 2636 440 2684
rect 400 2604 404 2636
rect 436 2604 440 2636
rect 400 2556 440 2604
rect 400 2524 404 2556
rect 436 2524 440 2556
rect 400 2520 440 2524
rect 480 3596 520 3600
rect 480 3564 484 3596
rect 516 3564 520 3596
rect 480 3516 520 3564
rect 480 3484 484 3516
rect 516 3484 520 3516
rect 480 3436 520 3484
rect 480 3404 484 3436
rect 516 3404 520 3436
rect 480 3356 520 3404
rect 480 3324 484 3356
rect 516 3324 520 3356
rect 480 3276 520 3324
rect 480 3244 484 3276
rect 516 3244 520 3276
rect 480 3196 520 3244
rect 480 3164 484 3196
rect 516 3164 520 3196
rect 480 3116 520 3164
rect 480 3084 484 3116
rect 516 3084 520 3116
rect 480 3036 520 3084
rect 480 3004 484 3036
rect 516 3004 520 3036
rect 480 2956 520 3004
rect 480 2924 484 2956
rect 516 2924 520 2956
rect 480 2876 520 2924
rect 480 2844 484 2876
rect 516 2844 520 2876
rect 480 2796 520 2844
rect 480 2764 484 2796
rect 516 2764 520 2796
rect 480 2716 520 2764
rect 480 2684 484 2716
rect 516 2684 520 2716
rect 480 2636 520 2684
rect 480 2604 484 2636
rect 516 2604 520 2636
rect 480 2556 520 2604
rect 480 2524 484 2556
rect 516 2524 520 2556
rect 480 2520 520 2524
rect 560 3596 600 3600
rect 560 3564 564 3596
rect 596 3564 600 3596
rect 560 3516 600 3564
rect 560 3484 564 3516
rect 596 3484 600 3516
rect 560 3436 600 3484
rect 560 3404 564 3436
rect 596 3404 600 3436
rect 560 3356 600 3404
rect 560 3324 564 3356
rect 596 3324 600 3356
rect 560 3276 600 3324
rect 560 3244 564 3276
rect 596 3244 600 3276
rect 560 3196 600 3244
rect 560 3164 564 3196
rect 596 3164 600 3196
rect 560 3116 600 3164
rect 560 3084 564 3116
rect 596 3084 600 3116
rect 560 3036 600 3084
rect 560 3004 564 3036
rect 596 3004 600 3036
rect 560 2956 600 3004
rect 560 2924 564 2956
rect 596 2924 600 2956
rect 560 2876 600 2924
rect 560 2844 564 2876
rect 596 2844 600 2876
rect 560 2796 600 2844
rect 560 2764 564 2796
rect 596 2764 600 2796
rect 560 2716 600 2764
rect 560 2684 564 2716
rect 596 2684 600 2716
rect 560 2636 600 2684
rect 560 2604 564 2636
rect 596 2604 600 2636
rect 560 2556 600 2604
rect 560 2524 564 2556
rect 596 2524 600 2556
rect 560 2520 600 2524
rect 640 3596 680 3600
rect 640 3564 644 3596
rect 676 3564 680 3596
rect 640 3516 680 3564
rect 640 3484 644 3516
rect 676 3484 680 3516
rect 640 3436 680 3484
rect 640 3404 644 3436
rect 676 3404 680 3436
rect 640 3356 680 3404
rect 640 3324 644 3356
rect 676 3324 680 3356
rect 640 3276 680 3324
rect 640 3244 644 3276
rect 676 3244 680 3276
rect 640 3196 680 3244
rect 640 3164 644 3196
rect 676 3164 680 3196
rect 640 3116 680 3164
rect 640 3084 644 3116
rect 676 3084 680 3116
rect 640 3036 680 3084
rect 640 3004 644 3036
rect 676 3004 680 3036
rect 640 2956 680 3004
rect 640 2924 644 2956
rect 676 2924 680 2956
rect 640 2876 680 2924
rect 640 2844 644 2876
rect 676 2844 680 2876
rect 640 2796 680 2844
rect 640 2764 644 2796
rect 676 2764 680 2796
rect 640 2716 680 2764
rect 640 2684 644 2716
rect 676 2684 680 2716
rect 640 2636 680 2684
rect 640 2604 644 2636
rect 676 2604 680 2636
rect 640 2556 680 2604
rect 640 2524 644 2556
rect 676 2524 680 2556
rect 640 2520 680 2524
rect 720 3596 760 3600
rect 720 3564 724 3596
rect 756 3564 760 3596
rect 720 3516 760 3564
rect 720 3484 724 3516
rect 756 3484 760 3516
rect 720 3436 760 3484
rect 720 3404 724 3436
rect 756 3404 760 3436
rect 720 3356 760 3404
rect 720 3324 724 3356
rect 756 3324 760 3356
rect 720 3276 760 3324
rect 720 3244 724 3276
rect 756 3244 760 3276
rect 720 3196 760 3244
rect 720 3164 724 3196
rect 756 3164 760 3196
rect 720 3116 760 3164
rect 720 3084 724 3116
rect 756 3084 760 3116
rect 720 3036 760 3084
rect 720 3004 724 3036
rect 756 3004 760 3036
rect 720 2956 760 3004
rect 720 2924 724 2956
rect 756 2924 760 2956
rect 720 2876 760 2924
rect 720 2844 724 2876
rect 756 2844 760 2876
rect 720 2796 760 2844
rect 720 2764 724 2796
rect 756 2764 760 2796
rect 720 2716 760 2764
rect 720 2684 724 2716
rect 756 2684 760 2716
rect 720 2636 760 2684
rect 720 2604 724 2636
rect 756 2604 760 2636
rect 720 2556 760 2604
rect 720 2524 724 2556
rect 756 2524 760 2556
rect 720 2520 760 2524
rect 800 3596 840 3600
rect 800 3564 804 3596
rect 836 3564 840 3596
rect 800 3516 840 3564
rect 800 3484 804 3516
rect 836 3484 840 3516
rect 800 3436 840 3484
rect 800 3404 804 3436
rect 836 3404 840 3436
rect 800 3356 840 3404
rect 800 3324 804 3356
rect 836 3324 840 3356
rect 800 3276 840 3324
rect 800 3244 804 3276
rect 836 3244 840 3276
rect 800 3196 840 3244
rect 800 3164 804 3196
rect 836 3164 840 3196
rect 800 3116 840 3164
rect 800 3084 804 3116
rect 836 3084 840 3116
rect 800 3036 840 3084
rect 800 3004 804 3036
rect 836 3004 840 3036
rect 800 2956 840 3004
rect 800 2924 804 2956
rect 836 2924 840 2956
rect 800 2876 840 2924
rect 800 2844 804 2876
rect 836 2844 840 2876
rect 800 2796 840 2844
rect 800 2764 804 2796
rect 836 2764 840 2796
rect 800 2716 840 2764
rect 800 2684 804 2716
rect 836 2684 840 2716
rect 800 2636 840 2684
rect 800 2604 804 2636
rect 836 2604 840 2636
rect 800 2556 840 2604
rect 800 2524 804 2556
rect 836 2524 840 2556
rect 800 2520 840 2524
rect 880 3596 920 3600
rect 880 3564 884 3596
rect 916 3564 920 3596
rect 880 3516 920 3564
rect 880 3484 884 3516
rect 916 3484 920 3516
rect 880 3436 920 3484
rect 880 3404 884 3436
rect 916 3404 920 3436
rect 880 3356 920 3404
rect 880 3324 884 3356
rect 916 3324 920 3356
rect 880 3276 920 3324
rect 880 3244 884 3276
rect 916 3244 920 3276
rect 880 3196 920 3244
rect 880 3164 884 3196
rect 916 3164 920 3196
rect 880 3116 920 3164
rect 880 3084 884 3116
rect 916 3084 920 3116
rect 880 3036 920 3084
rect 880 3004 884 3036
rect 916 3004 920 3036
rect 880 2956 920 3004
rect 880 2924 884 2956
rect 916 2924 920 2956
rect 880 2876 920 2924
rect 880 2844 884 2876
rect 916 2844 920 2876
rect 880 2796 920 2844
rect 880 2764 884 2796
rect 916 2764 920 2796
rect 880 2716 920 2764
rect 880 2684 884 2716
rect 916 2684 920 2716
rect 880 2636 920 2684
rect 880 2604 884 2636
rect 916 2604 920 2636
rect 880 2556 920 2604
rect 880 2524 884 2556
rect 916 2524 920 2556
rect 880 2520 920 2524
rect 960 3596 1000 3600
rect 960 3564 964 3596
rect 996 3564 1000 3596
rect 960 3516 1000 3564
rect 960 3484 964 3516
rect 996 3484 1000 3516
rect 960 3436 1000 3484
rect 960 3404 964 3436
rect 996 3404 1000 3436
rect 960 3356 1000 3404
rect 960 3324 964 3356
rect 996 3324 1000 3356
rect 960 3276 1000 3324
rect 960 3244 964 3276
rect 996 3244 1000 3276
rect 960 3196 1000 3244
rect 960 3164 964 3196
rect 996 3164 1000 3196
rect 960 3116 1000 3164
rect 960 3084 964 3116
rect 996 3084 1000 3116
rect 960 3036 1000 3084
rect 960 3004 964 3036
rect 996 3004 1000 3036
rect 960 2956 1000 3004
rect 960 2924 964 2956
rect 996 2924 1000 2956
rect 960 2876 1000 2924
rect 960 2844 964 2876
rect 996 2844 1000 2876
rect 960 2796 1000 2844
rect 960 2764 964 2796
rect 996 2764 1000 2796
rect 960 2716 1000 2764
rect 960 2684 964 2716
rect 996 2684 1000 2716
rect 960 2636 1000 2684
rect 960 2604 964 2636
rect 996 2604 1000 2636
rect 960 2556 1000 2604
rect 960 2524 964 2556
rect 996 2524 1000 2556
rect 960 2520 1000 2524
rect 1040 3596 1080 3600
rect 1040 3564 1044 3596
rect 1076 3564 1080 3596
rect 1040 3516 1080 3564
rect 1040 3484 1044 3516
rect 1076 3484 1080 3516
rect 1040 3436 1080 3484
rect 1040 3404 1044 3436
rect 1076 3404 1080 3436
rect 1040 3356 1080 3404
rect 1040 3324 1044 3356
rect 1076 3324 1080 3356
rect 1040 3276 1080 3324
rect 1040 3244 1044 3276
rect 1076 3244 1080 3276
rect 1040 3196 1080 3244
rect 1040 3164 1044 3196
rect 1076 3164 1080 3196
rect 1040 3116 1080 3164
rect 1040 3084 1044 3116
rect 1076 3084 1080 3116
rect 1040 3036 1080 3084
rect 1040 3004 1044 3036
rect 1076 3004 1080 3036
rect 1040 2956 1080 3004
rect 1040 2924 1044 2956
rect 1076 2924 1080 2956
rect 1040 2876 1080 2924
rect 1040 2844 1044 2876
rect 1076 2844 1080 2876
rect 1040 2796 1080 2844
rect 1040 2764 1044 2796
rect 1076 2764 1080 2796
rect 1040 2716 1080 2764
rect 1040 2684 1044 2716
rect 1076 2684 1080 2716
rect 1040 2636 1080 2684
rect 1040 2604 1044 2636
rect 1076 2604 1080 2636
rect 1040 2556 1080 2604
rect 1040 2524 1044 2556
rect 1076 2524 1080 2556
rect 1040 2520 1080 2524
rect 1120 3596 1160 3600
rect 1120 3564 1124 3596
rect 1156 3564 1160 3596
rect 1120 3516 1160 3564
rect 1120 3484 1124 3516
rect 1156 3484 1160 3516
rect 1120 3436 1160 3484
rect 1120 3404 1124 3436
rect 1156 3404 1160 3436
rect 1120 3356 1160 3404
rect 1120 3324 1124 3356
rect 1156 3324 1160 3356
rect 1120 3276 1160 3324
rect 1120 3244 1124 3276
rect 1156 3244 1160 3276
rect 1120 3196 1160 3244
rect 1120 3164 1124 3196
rect 1156 3164 1160 3196
rect 1120 3116 1160 3164
rect 1120 3084 1124 3116
rect 1156 3084 1160 3116
rect 1120 3036 1160 3084
rect 1120 3004 1124 3036
rect 1156 3004 1160 3036
rect 1120 2956 1160 3004
rect 1120 2924 1124 2956
rect 1156 2924 1160 2956
rect 1120 2876 1160 2924
rect 1120 2844 1124 2876
rect 1156 2844 1160 2876
rect 1120 2796 1160 2844
rect 1120 2764 1124 2796
rect 1156 2764 1160 2796
rect 1120 2716 1160 2764
rect 1120 2684 1124 2716
rect 1156 2684 1160 2716
rect 1120 2636 1160 2684
rect 1120 2604 1124 2636
rect 1156 2604 1160 2636
rect 1120 2556 1160 2604
rect 1120 2524 1124 2556
rect 1156 2524 1160 2556
rect 1120 2520 1160 2524
rect 1200 3596 1240 3600
rect 1200 3564 1204 3596
rect 1236 3564 1240 3596
rect 1200 3516 1240 3564
rect 1200 3484 1204 3516
rect 1236 3484 1240 3516
rect 1200 3436 1240 3484
rect 1200 3404 1204 3436
rect 1236 3404 1240 3436
rect 1200 3356 1240 3404
rect 1200 3324 1204 3356
rect 1236 3324 1240 3356
rect 1200 3276 1240 3324
rect 1200 3244 1204 3276
rect 1236 3244 1240 3276
rect 1200 3196 1240 3244
rect 1200 3164 1204 3196
rect 1236 3164 1240 3196
rect 1200 3116 1240 3164
rect 1200 3084 1204 3116
rect 1236 3084 1240 3116
rect 1200 3036 1240 3084
rect 1200 3004 1204 3036
rect 1236 3004 1240 3036
rect 1200 2956 1240 3004
rect 1200 2924 1204 2956
rect 1236 2924 1240 2956
rect 1200 2876 1240 2924
rect 1200 2844 1204 2876
rect 1236 2844 1240 2876
rect 1200 2796 1240 2844
rect 1200 2764 1204 2796
rect 1236 2764 1240 2796
rect 1200 2716 1240 2764
rect 1200 2684 1204 2716
rect 1236 2684 1240 2716
rect 1200 2636 1240 2684
rect 1200 2604 1204 2636
rect 1236 2604 1240 2636
rect 1200 2556 1240 2604
rect 1200 2524 1204 2556
rect 1236 2524 1240 2556
rect 1200 2520 1240 2524
rect 1280 3596 1320 3600
rect 1280 3564 1284 3596
rect 1316 3564 1320 3596
rect 1280 3516 1320 3564
rect 1280 3484 1284 3516
rect 1316 3484 1320 3516
rect 1280 3436 1320 3484
rect 1280 3404 1284 3436
rect 1316 3404 1320 3436
rect 1280 3356 1320 3404
rect 1280 3324 1284 3356
rect 1316 3324 1320 3356
rect 1280 3276 1320 3324
rect 1280 3244 1284 3276
rect 1316 3244 1320 3276
rect 1280 3196 1320 3244
rect 1280 3164 1284 3196
rect 1316 3164 1320 3196
rect 1280 3116 1320 3164
rect 1280 3084 1284 3116
rect 1316 3084 1320 3116
rect 1280 3036 1320 3084
rect 1280 3004 1284 3036
rect 1316 3004 1320 3036
rect 1280 2956 1320 3004
rect 1280 2924 1284 2956
rect 1316 2924 1320 2956
rect 1280 2876 1320 2924
rect 1280 2844 1284 2876
rect 1316 2844 1320 2876
rect 1280 2796 1320 2844
rect 1280 2764 1284 2796
rect 1316 2764 1320 2796
rect 1280 2716 1320 2764
rect 1280 2684 1284 2716
rect 1316 2684 1320 2716
rect 1280 2636 1320 2684
rect 1280 2604 1284 2636
rect 1316 2604 1320 2636
rect 1280 2556 1320 2604
rect 1280 2524 1284 2556
rect 1316 2524 1320 2556
rect 1280 2520 1320 2524
rect 1360 3596 1400 3600
rect 1360 3564 1364 3596
rect 1396 3564 1400 3596
rect 1360 3516 1400 3564
rect 1360 3484 1364 3516
rect 1396 3484 1400 3516
rect 1360 3436 1400 3484
rect 1360 3404 1364 3436
rect 1396 3404 1400 3436
rect 1360 3356 1400 3404
rect 1360 3324 1364 3356
rect 1396 3324 1400 3356
rect 1360 3276 1400 3324
rect 1360 3244 1364 3276
rect 1396 3244 1400 3276
rect 1360 3196 1400 3244
rect 1360 3164 1364 3196
rect 1396 3164 1400 3196
rect 1360 3116 1400 3164
rect 1360 3084 1364 3116
rect 1396 3084 1400 3116
rect 1360 3036 1400 3084
rect 1360 3004 1364 3036
rect 1396 3004 1400 3036
rect 1360 2956 1400 3004
rect 1360 2924 1364 2956
rect 1396 2924 1400 2956
rect 1360 2876 1400 2924
rect 1360 2844 1364 2876
rect 1396 2844 1400 2876
rect 1360 2796 1400 2844
rect 1360 2764 1364 2796
rect 1396 2764 1400 2796
rect 1360 2716 1400 2764
rect 1360 2684 1364 2716
rect 1396 2684 1400 2716
rect 1360 2636 1400 2684
rect 1360 2604 1364 2636
rect 1396 2604 1400 2636
rect 1360 2556 1400 2604
rect 1360 2524 1364 2556
rect 1396 2524 1400 2556
rect 1360 2520 1400 2524
rect 1440 3596 1480 3600
rect 1440 3564 1444 3596
rect 1476 3564 1480 3596
rect 1440 3516 1480 3564
rect 1440 3484 1444 3516
rect 1476 3484 1480 3516
rect 1440 3436 1480 3484
rect 1440 3404 1444 3436
rect 1476 3404 1480 3436
rect 1440 3356 1480 3404
rect 1440 3324 1444 3356
rect 1476 3324 1480 3356
rect 1440 3276 1480 3324
rect 1440 3244 1444 3276
rect 1476 3244 1480 3276
rect 1440 3196 1480 3244
rect 1440 3164 1444 3196
rect 1476 3164 1480 3196
rect 1440 3116 1480 3164
rect 1440 3084 1444 3116
rect 1476 3084 1480 3116
rect 1440 3036 1480 3084
rect 1440 3004 1444 3036
rect 1476 3004 1480 3036
rect 1440 2956 1480 3004
rect 1440 2924 1444 2956
rect 1476 2924 1480 2956
rect 1440 2876 1480 2924
rect 1440 2844 1444 2876
rect 1476 2844 1480 2876
rect 1440 2796 1480 2844
rect 1440 2764 1444 2796
rect 1476 2764 1480 2796
rect 1440 2716 1480 2764
rect 1440 2684 1444 2716
rect 1476 2684 1480 2716
rect 1440 2636 1480 2684
rect 1440 2604 1444 2636
rect 1476 2604 1480 2636
rect 1440 2556 1480 2604
rect 1440 2524 1444 2556
rect 1476 2524 1480 2556
rect 1440 2520 1480 2524
rect 1520 3596 1560 3600
rect 1520 3564 1524 3596
rect 1556 3564 1560 3596
rect 1520 3516 1560 3564
rect 1520 3484 1524 3516
rect 1556 3484 1560 3516
rect 1520 3436 1560 3484
rect 1520 3404 1524 3436
rect 1556 3404 1560 3436
rect 1520 3356 1560 3404
rect 1520 3324 1524 3356
rect 1556 3324 1560 3356
rect 1520 3276 1560 3324
rect 1520 3244 1524 3276
rect 1556 3244 1560 3276
rect 1520 3196 1560 3244
rect 1520 3164 1524 3196
rect 1556 3164 1560 3196
rect 1520 3116 1560 3164
rect 1520 3084 1524 3116
rect 1556 3084 1560 3116
rect 1520 3036 1560 3084
rect 1520 3004 1524 3036
rect 1556 3004 1560 3036
rect 1520 2956 1560 3004
rect 1520 2924 1524 2956
rect 1556 2924 1560 2956
rect 1520 2876 1560 2924
rect 1520 2844 1524 2876
rect 1556 2844 1560 2876
rect 1520 2796 1560 2844
rect 1520 2764 1524 2796
rect 1556 2764 1560 2796
rect 1520 2716 1560 2764
rect 1520 2684 1524 2716
rect 1556 2684 1560 2716
rect 1520 2636 1560 2684
rect 1520 2604 1524 2636
rect 1556 2604 1560 2636
rect 1520 2556 1560 2604
rect 1520 2524 1524 2556
rect 1556 2524 1560 2556
rect 1520 2520 1560 2524
rect 1600 3596 1640 3600
rect 1600 3564 1604 3596
rect 1636 3564 1640 3596
rect 1600 3516 1640 3564
rect 1600 3484 1604 3516
rect 1636 3484 1640 3516
rect 1600 3436 1640 3484
rect 1600 3404 1604 3436
rect 1636 3404 1640 3436
rect 1600 3356 1640 3404
rect 1600 3324 1604 3356
rect 1636 3324 1640 3356
rect 1600 3276 1640 3324
rect 1600 3244 1604 3276
rect 1636 3244 1640 3276
rect 1600 3196 1640 3244
rect 1600 3164 1604 3196
rect 1636 3164 1640 3196
rect 1600 3116 1640 3164
rect 1600 3084 1604 3116
rect 1636 3084 1640 3116
rect 1600 3036 1640 3084
rect 1600 3004 1604 3036
rect 1636 3004 1640 3036
rect 1600 2956 1640 3004
rect 1600 2924 1604 2956
rect 1636 2924 1640 2956
rect 1600 2876 1640 2924
rect 1600 2844 1604 2876
rect 1636 2844 1640 2876
rect 1600 2796 1640 2844
rect 1600 2764 1604 2796
rect 1636 2764 1640 2796
rect 1600 2716 1640 2764
rect 1600 2684 1604 2716
rect 1636 2684 1640 2716
rect 1600 2636 1640 2684
rect 1600 2604 1604 2636
rect 1636 2604 1640 2636
rect 1600 2556 1640 2604
rect 1600 2524 1604 2556
rect 1636 2524 1640 2556
rect 1600 2520 1640 2524
rect 1680 3596 1720 3600
rect 1680 3564 1684 3596
rect 1716 3564 1720 3596
rect 1680 3516 1720 3564
rect 1680 3484 1684 3516
rect 1716 3484 1720 3516
rect 1680 3436 1720 3484
rect 1680 3404 1684 3436
rect 1716 3404 1720 3436
rect 1680 3356 1720 3404
rect 1680 3324 1684 3356
rect 1716 3324 1720 3356
rect 1680 3276 1720 3324
rect 1680 3244 1684 3276
rect 1716 3244 1720 3276
rect 1680 3196 1720 3244
rect 1680 3164 1684 3196
rect 1716 3164 1720 3196
rect 1680 3116 1720 3164
rect 1680 3084 1684 3116
rect 1716 3084 1720 3116
rect 1680 3036 1720 3084
rect 1680 3004 1684 3036
rect 1716 3004 1720 3036
rect 1680 2956 1720 3004
rect 1680 2924 1684 2956
rect 1716 2924 1720 2956
rect 1680 2876 1720 2924
rect 1680 2844 1684 2876
rect 1716 2844 1720 2876
rect 1680 2796 1720 2844
rect 1680 2764 1684 2796
rect 1716 2764 1720 2796
rect 1680 2716 1720 2764
rect 1680 2684 1684 2716
rect 1716 2684 1720 2716
rect 1680 2636 1720 2684
rect 1680 2604 1684 2636
rect 1716 2604 1720 2636
rect 1680 2556 1720 2604
rect 1680 2524 1684 2556
rect 1716 2524 1720 2556
rect 1680 2520 1720 2524
rect 1760 3596 1800 3600
rect 1760 3564 1764 3596
rect 1796 3564 1800 3596
rect 1760 3516 1800 3564
rect 1760 3484 1764 3516
rect 1796 3484 1800 3516
rect 1760 3436 1800 3484
rect 1760 3404 1764 3436
rect 1796 3404 1800 3436
rect 1760 3356 1800 3404
rect 1760 3324 1764 3356
rect 1796 3324 1800 3356
rect 1760 3276 1800 3324
rect 1760 3244 1764 3276
rect 1796 3244 1800 3276
rect 1760 3196 1800 3244
rect 1760 3164 1764 3196
rect 1796 3164 1800 3196
rect 1760 3116 1800 3164
rect 1760 3084 1764 3116
rect 1796 3084 1800 3116
rect 1760 3036 1800 3084
rect 1760 3004 1764 3036
rect 1796 3004 1800 3036
rect 1760 2956 1800 3004
rect 1760 2924 1764 2956
rect 1796 2924 1800 2956
rect 1760 2876 1800 2924
rect 1760 2844 1764 2876
rect 1796 2844 1800 2876
rect 1760 2796 1800 2844
rect 1760 2764 1764 2796
rect 1796 2764 1800 2796
rect 1760 2716 1800 2764
rect 1760 2684 1764 2716
rect 1796 2684 1800 2716
rect 1760 2636 1800 2684
rect 1760 2604 1764 2636
rect 1796 2604 1800 2636
rect 1760 2556 1800 2604
rect 1760 2524 1764 2556
rect 1796 2524 1800 2556
rect 1760 2520 1800 2524
rect 1840 3596 1880 3600
rect 1840 3564 1844 3596
rect 1876 3564 1880 3596
rect 1840 3516 1880 3564
rect 1840 3484 1844 3516
rect 1876 3484 1880 3516
rect 1840 3436 1880 3484
rect 1840 3404 1844 3436
rect 1876 3404 1880 3436
rect 1840 3356 1880 3404
rect 1840 3324 1844 3356
rect 1876 3324 1880 3356
rect 1840 3276 1880 3324
rect 1840 3244 1844 3276
rect 1876 3244 1880 3276
rect 1840 3196 1880 3244
rect 1840 3164 1844 3196
rect 1876 3164 1880 3196
rect 1840 3116 1880 3164
rect 1840 3084 1844 3116
rect 1876 3084 1880 3116
rect 1840 3036 1880 3084
rect 1840 3004 1844 3036
rect 1876 3004 1880 3036
rect 1840 2956 1880 3004
rect 1840 2924 1844 2956
rect 1876 2924 1880 2956
rect 1840 2876 1880 2924
rect 1840 2844 1844 2876
rect 1876 2844 1880 2876
rect 1840 2796 1880 2844
rect 1840 2764 1844 2796
rect 1876 2764 1880 2796
rect 1840 2716 1880 2764
rect 1840 2684 1844 2716
rect 1876 2684 1880 2716
rect 1840 2636 1880 2684
rect 1840 2604 1844 2636
rect 1876 2604 1880 2636
rect 1840 2556 1880 2604
rect 1840 2524 1844 2556
rect 1876 2524 1880 2556
rect 1840 2520 1880 2524
rect 1920 3596 1960 3600
rect 1920 3564 1924 3596
rect 1956 3564 1960 3596
rect 1920 3516 1960 3564
rect 1920 3484 1924 3516
rect 1956 3484 1960 3516
rect 1920 3436 1960 3484
rect 1920 3404 1924 3436
rect 1956 3404 1960 3436
rect 1920 3356 1960 3404
rect 1920 3324 1924 3356
rect 1956 3324 1960 3356
rect 1920 3276 1960 3324
rect 1920 3244 1924 3276
rect 1956 3244 1960 3276
rect 1920 3196 1960 3244
rect 1920 3164 1924 3196
rect 1956 3164 1960 3196
rect 1920 3116 1960 3164
rect 1920 3084 1924 3116
rect 1956 3084 1960 3116
rect 1920 3036 1960 3084
rect 1920 3004 1924 3036
rect 1956 3004 1960 3036
rect 1920 2956 1960 3004
rect 1920 2924 1924 2956
rect 1956 2924 1960 2956
rect 1920 2876 1960 2924
rect 1920 2844 1924 2876
rect 1956 2844 1960 2876
rect 1920 2796 1960 2844
rect 1920 2764 1924 2796
rect 1956 2764 1960 2796
rect 1920 2716 1960 2764
rect 1920 2684 1924 2716
rect 1956 2684 1960 2716
rect 1920 2636 1960 2684
rect 1920 2604 1924 2636
rect 1956 2604 1960 2636
rect 1920 2556 1960 2604
rect 1920 2524 1924 2556
rect 1956 2524 1960 2556
rect 1920 2520 1960 2524
rect 2000 3596 2040 3600
rect 2000 3564 2004 3596
rect 2036 3564 2040 3596
rect 2000 3516 2040 3564
rect 2000 3484 2004 3516
rect 2036 3484 2040 3516
rect 2000 3436 2040 3484
rect 2000 3404 2004 3436
rect 2036 3404 2040 3436
rect 2000 3356 2040 3404
rect 2000 3324 2004 3356
rect 2036 3324 2040 3356
rect 2000 3276 2040 3324
rect 2000 3244 2004 3276
rect 2036 3244 2040 3276
rect 2000 3196 2040 3244
rect 2000 3164 2004 3196
rect 2036 3164 2040 3196
rect 2000 3116 2040 3164
rect 2000 3084 2004 3116
rect 2036 3084 2040 3116
rect 2000 3036 2040 3084
rect 2000 3004 2004 3036
rect 2036 3004 2040 3036
rect 2000 2956 2040 3004
rect 2000 2924 2004 2956
rect 2036 2924 2040 2956
rect 2000 2876 2040 2924
rect 2000 2844 2004 2876
rect 2036 2844 2040 2876
rect 2000 2796 2040 2844
rect 2000 2764 2004 2796
rect 2036 2764 2040 2796
rect 2000 2716 2040 2764
rect 2000 2684 2004 2716
rect 2036 2684 2040 2716
rect 2000 2636 2040 2684
rect 2000 2604 2004 2636
rect 2036 2604 2040 2636
rect 2000 2556 2040 2604
rect 2000 2524 2004 2556
rect 2036 2524 2040 2556
rect 2000 2520 2040 2524
rect 2080 3596 2120 3600
rect 2080 3564 2084 3596
rect 2116 3564 2120 3596
rect 2080 3516 2120 3564
rect 2080 3484 2084 3516
rect 2116 3484 2120 3516
rect 2080 3436 2120 3484
rect 2080 3404 2084 3436
rect 2116 3404 2120 3436
rect 2080 3356 2120 3404
rect 2080 3324 2084 3356
rect 2116 3324 2120 3356
rect 2080 3276 2120 3324
rect 2080 3244 2084 3276
rect 2116 3244 2120 3276
rect 2080 3196 2120 3244
rect 2080 3164 2084 3196
rect 2116 3164 2120 3196
rect 2080 3116 2120 3164
rect 2080 3084 2084 3116
rect 2116 3084 2120 3116
rect 2080 3036 2120 3084
rect 2080 3004 2084 3036
rect 2116 3004 2120 3036
rect 2080 2956 2120 3004
rect 2080 2924 2084 2956
rect 2116 2924 2120 2956
rect 2080 2876 2120 2924
rect 2080 2844 2084 2876
rect 2116 2844 2120 2876
rect 2080 2796 2120 2844
rect 2080 2764 2084 2796
rect 2116 2764 2120 2796
rect 2080 2716 2120 2764
rect 2080 2684 2084 2716
rect 2116 2684 2120 2716
rect 2080 2636 2120 2684
rect 2080 2604 2084 2636
rect 2116 2604 2120 2636
rect 2080 2556 2120 2604
rect 2080 2524 2084 2556
rect 2116 2524 2120 2556
rect 2080 2520 2120 2524
rect 2160 3596 2200 3600
rect 2160 3564 2164 3596
rect 2196 3564 2200 3596
rect 2160 3516 2200 3564
rect 2160 3484 2164 3516
rect 2196 3484 2200 3516
rect 2160 3436 2200 3484
rect 2160 3404 2164 3436
rect 2196 3404 2200 3436
rect 2160 3356 2200 3404
rect 2160 3324 2164 3356
rect 2196 3324 2200 3356
rect 2160 3276 2200 3324
rect 2160 3244 2164 3276
rect 2196 3244 2200 3276
rect 2160 3196 2200 3244
rect 2160 3164 2164 3196
rect 2196 3164 2200 3196
rect 2160 3116 2200 3164
rect 2160 3084 2164 3116
rect 2196 3084 2200 3116
rect 2160 3036 2200 3084
rect 2160 3004 2164 3036
rect 2196 3004 2200 3036
rect 2160 2956 2200 3004
rect 2160 2924 2164 2956
rect 2196 2924 2200 2956
rect 2160 2876 2200 2924
rect 2160 2844 2164 2876
rect 2196 2844 2200 2876
rect 2160 2796 2200 2844
rect 2160 2764 2164 2796
rect 2196 2764 2200 2796
rect 2160 2716 2200 2764
rect 2160 2684 2164 2716
rect 2196 2684 2200 2716
rect 2160 2636 2200 2684
rect 2160 2604 2164 2636
rect 2196 2604 2200 2636
rect 2160 2556 2200 2604
rect 2160 2524 2164 2556
rect 2196 2524 2200 2556
rect 2160 2520 2200 2524
rect 2240 3596 2280 3600
rect 2240 3564 2244 3596
rect 2276 3564 2280 3596
rect 2240 3516 2280 3564
rect 2240 3484 2244 3516
rect 2276 3484 2280 3516
rect 2240 3436 2280 3484
rect 2240 3404 2244 3436
rect 2276 3404 2280 3436
rect 2240 3356 2280 3404
rect 2240 3324 2244 3356
rect 2276 3324 2280 3356
rect 2240 3276 2280 3324
rect 2240 3244 2244 3276
rect 2276 3244 2280 3276
rect 2240 3196 2280 3244
rect 2240 3164 2244 3196
rect 2276 3164 2280 3196
rect 2240 3116 2280 3164
rect 2240 3084 2244 3116
rect 2276 3084 2280 3116
rect 2240 3036 2280 3084
rect 2240 3004 2244 3036
rect 2276 3004 2280 3036
rect 2240 2956 2280 3004
rect 2240 2924 2244 2956
rect 2276 2924 2280 2956
rect 2240 2876 2280 2924
rect 2240 2844 2244 2876
rect 2276 2844 2280 2876
rect 2240 2796 2280 2844
rect 2240 2764 2244 2796
rect 2276 2764 2280 2796
rect 2240 2716 2280 2764
rect 2240 2684 2244 2716
rect 2276 2684 2280 2716
rect 2240 2636 2280 2684
rect 2240 2604 2244 2636
rect 2276 2604 2280 2636
rect 2240 2556 2280 2604
rect 2240 2524 2244 2556
rect 2276 2524 2280 2556
rect 2240 2520 2280 2524
rect 2320 3596 2360 3600
rect 2320 3564 2324 3596
rect 2356 3564 2360 3596
rect 2320 3516 2360 3564
rect 2320 3484 2324 3516
rect 2356 3484 2360 3516
rect 2320 3436 2360 3484
rect 2320 3404 2324 3436
rect 2356 3404 2360 3436
rect 2320 3356 2360 3404
rect 2320 3324 2324 3356
rect 2356 3324 2360 3356
rect 2320 3276 2360 3324
rect 2320 3244 2324 3276
rect 2356 3244 2360 3276
rect 2320 3196 2360 3244
rect 2320 3164 2324 3196
rect 2356 3164 2360 3196
rect 2320 3116 2360 3164
rect 2320 3084 2324 3116
rect 2356 3084 2360 3116
rect 2320 3036 2360 3084
rect 2320 3004 2324 3036
rect 2356 3004 2360 3036
rect 2320 2956 2360 3004
rect 2320 2924 2324 2956
rect 2356 2924 2360 2956
rect 2320 2876 2360 2924
rect 2320 2844 2324 2876
rect 2356 2844 2360 2876
rect 2320 2796 2360 2844
rect 2320 2764 2324 2796
rect 2356 2764 2360 2796
rect 2320 2716 2360 2764
rect 2320 2684 2324 2716
rect 2356 2684 2360 2716
rect 2320 2636 2360 2684
rect 2320 2604 2324 2636
rect 2356 2604 2360 2636
rect 2320 2556 2360 2604
rect 2320 2524 2324 2556
rect 2356 2524 2360 2556
rect 2320 2520 2360 2524
rect 2400 3596 2440 3600
rect 2400 3564 2404 3596
rect 2436 3564 2440 3596
rect 2400 3516 2440 3564
rect 2400 3484 2404 3516
rect 2436 3484 2440 3516
rect 2400 3436 2440 3484
rect 2400 3404 2404 3436
rect 2436 3404 2440 3436
rect 2400 3356 2440 3404
rect 2400 3324 2404 3356
rect 2436 3324 2440 3356
rect 2400 3276 2440 3324
rect 2400 3244 2404 3276
rect 2436 3244 2440 3276
rect 2400 3196 2440 3244
rect 2400 3164 2404 3196
rect 2436 3164 2440 3196
rect 2400 3116 2440 3164
rect 2400 3084 2404 3116
rect 2436 3084 2440 3116
rect 2400 3036 2440 3084
rect 2400 3004 2404 3036
rect 2436 3004 2440 3036
rect 2400 2956 2440 3004
rect 2400 2924 2404 2956
rect 2436 2924 2440 2956
rect 2400 2876 2440 2924
rect 2400 2844 2404 2876
rect 2436 2844 2440 2876
rect 2400 2796 2440 2844
rect 2400 2764 2404 2796
rect 2436 2764 2440 2796
rect 2400 2716 2440 2764
rect 2400 2684 2404 2716
rect 2436 2684 2440 2716
rect 2400 2636 2440 2684
rect 2400 2604 2404 2636
rect 2436 2604 2440 2636
rect 2400 2556 2440 2604
rect 2400 2524 2404 2556
rect 2436 2524 2440 2556
rect 2400 2520 2440 2524
rect 2480 3596 2520 3600
rect 2480 3564 2484 3596
rect 2516 3564 2520 3596
rect 2480 3516 2520 3564
rect 2480 3484 2484 3516
rect 2516 3484 2520 3516
rect 2480 3436 2520 3484
rect 2480 3404 2484 3436
rect 2516 3404 2520 3436
rect 2480 3356 2520 3404
rect 2480 3324 2484 3356
rect 2516 3324 2520 3356
rect 2480 3276 2520 3324
rect 2480 3244 2484 3276
rect 2516 3244 2520 3276
rect 2480 3196 2520 3244
rect 2480 3164 2484 3196
rect 2516 3164 2520 3196
rect 2480 3116 2520 3164
rect 2480 3084 2484 3116
rect 2516 3084 2520 3116
rect 2480 3036 2520 3084
rect 2480 3004 2484 3036
rect 2516 3004 2520 3036
rect 2480 2956 2520 3004
rect 2480 2924 2484 2956
rect 2516 2924 2520 2956
rect 2480 2876 2520 2924
rect 2480 2844 2484 2876
rect 2516 2844 2520 2876
rect 2480 2796 2520 2844
rect 2480 2764 2484 2796
rect 2516 2764 2520 2796
rect 2480 2716 2520 2764
rect 2480 2684 2484 2716
rect 2516 2684 2520 2716
rect 2480 2636 2520 2684
rect 2480 2604 2484 2636
rect 2516 2604 2520 2636
rect 2480 2556 2520 2604
rect 2480 2524 2484 2556
rect 2516 2524 2520 2556
rect 2480 2520 2520 2524
rect 2560 3596 2600 3600
rect 2560 3564 2564 3596
rect 2596 3564 2600 3596
rect 2560 3516 2600 3564
rect 2560 3484 2564 3516
rect 2596 3484 2600 3516
rect 2560 3436 2600 3484
rect 2560 3404 2564 3436
rect 2596 3404 2600 3436
rect 2560 3356 2600 3404
rect 2560 3324 2564 3356
rect 2596 3324 2600 3356
rect 2560 3276 2600 3324
rect 2560 3244 2564 3276
rect 2596 3244 2600 3276
rect 2560 3196 2600 3244
rect 2560 3164 2564 3196
rect 2596 3164 2600 3196
rect 2560 3116 2600 3164
rect 2560 3084 2564 3116
rect 2596 3084 2600 3116
rect 2560 3036 2600 3084
rect 2560 3004 2564 3036
rect 2596 3004 2600 3036
rect 2560 2956 2600 3004
rect 2560 2924 2564 2956
rect 2596 2924 2600 2956
rect 2560 2876 2600 2924
rect 2560 2844 2564 2876
rect 2596 2844 2600 2876
rect 2560 2796 2600 2844
rect 2560 2764 2564 2796
rect 2596 2764 2600 2796
rect 2560 2716 2600 2764
rect 2560 2684 2564 2716
rect 2596 2684 2600 2716
rect 2560 2636 2600 2684
rect 2560 2604 2564 2636
rect 2596 2604 2600 2636
rect 2560 2556 2600 2604
rect 2560 2524 2564 2556
rect 2596 2524 2600 2556
rect 2560 2520 2600 2524
rect 2640 3596 2680 3600
rect 2640 3564 2644 3596
rect 2676 3564 2680 3596
rect 2640 3516 2680 3564
rect 2640 3484 2644 3516
rect 2676 3484 2680 3516
rect 2640 3436 2680 3484
rect 2640 3404 2644 3436
rect 2676 3404 2680 3436
rect 2640 3356 2680 3404
rect 2640 3324 2644 3356
rect 2676 3324 2680 3356
rect 2640 3276 2680 3324
rect 2640 3244 2644 3276
rect 2676 3244 2680 3276
rect 2640 3196 2680 3244
rect 2640 3164 2644 3196
rect 2676 3164 2680 3196
rect 2640 3116 2680 3164
rect 2640 3084 2644 3116
rect 2676 3084 2680 3116
rect 2640 3036 2680 3084
rect 2640 3004 2644 3036
rect 2676 3004 2680 3036
rect 2640 2956 2680 3004
rect 2640 2924 2644 2956
rect 2676 2924 2680 2956
rect 2640 2876 2680 2924
rect 2640 2844 2644 2876
rect 2676 2844 2680 2876
rect 2640 2796 2680 2844
rect 2640 2764 2644 2796
rect 2676 2764 2680 2796
rect 2640 2716 2680 2764
rect 2640 2684 2644 2716
rect 2676 2684 2680 2716
rect 2640 2636 2680 2684
rect 2640 2604 2644 2636
rect 2676 2604 2680 2636
rect 2640 2556 2680 2604
rect 2640 2524 2644 2556
rect 2676 2524 2680 2556
rect 2640 2520 2680 2524
rect 2720 3596 2760 3600
rect 2720 3564 2724 3596
rect 2756 3564 2760 3596
rect 2720 3516 2760 3564
rect 2720 3484 2724 3516
rect 2756 3484 2760 3516
rect 2720 3436 2760 3484
rect 2720 3404 2724 3436
rect 2756 3404 2760 3436
rect 2720 3356 2760 3404
rect 2720 3324 2724 3356
rect 2756 3324 2760 3356
rect 2720 3276 2760 3324
rect 2720 3244 2724 3276
rect 2756 3244 2760 3276
rect 2720 3196 2760 3244
rect 2720 3164 2724 3196
rect 2756 3164 2760 3196
rect 2720 3116 2760 3164
rect 2720 3084 2724 3116
rect 2756 3084 2760 3116
rect 2720 3036 2760 3084
rect 2720 3004 2724 3036
rect 2756 3004 2760 3036
rect 2720 2956 2760 3004
rect 2720 2924 2724 2956
rect 2756 2924 2760 2956
rect 2720 2876 2760 2924
rect 2720 2844 2724 2876
rect 2756 2844 2760 2876
rect 2720 2796 2760 2844
rect 2720 2764 2724 2796
rect 2756 2764 2760 2796
rect 2720 2716 2760 2764
rect 2720 2684 2724 2716
rect 2756 2684 2760 2716
rect 2720 2636 2760 2684
rect 2720 2604 2724 2636
rect 2756 2604 2760 2636
rect 2720 2556 2760 2604
rect 2720 2524 2724 2556
rect 2756 2524 2760 2556
rect 2720 2520 2760 2524
rect 2800 3596 2840 3600
rect 2800 3564 2804 3596
rect 2836 3564 2840 3596
rect 2800 3516 2840 3564
rect 2800 3484 2804 3516
rect 2836 3484 2840 3516
rect 2800 3436 2840 3484
rect 2800 3404 2804 3436
rect 2836 3404 2840 3436
rect 2800 3356 2840 3404
rect 2800 3324 2804 3356
rect 2836 3324 2840 3356
rect 2800 3276 2840 3324
rect 2800 3244 2804 3276
rect 2836 3244 2840 3276
rect 2800 3196 2840 3244
rect 2800 3164 2804 3196
rect 2836 3164 2840 3196
rect 2800 3116 2840 3164
rect 2800 3084 2804 3116
rect 2836 3084 2840 3116
rect 2800 3036 2840 3084
rect 2800 3004 2804 3036
rect 2836 3004 2840 3036
rect 2800 2956 2840 3004
rect 2800 2924 2804 2956
rect 2836 2924 2840 2956
rect 2800 2876 2840 2924
rect 2800 2844 2804 2876
rect 2836 2844 2840 2876
rect 2800 2796 2840 2844
rect 2800 2764 2804 2796
rect 2836 2764 2840 2796
rect 2800 2716 2840 2764
rect 2800 2684 2804 2716
rect 2836 2684 2840 2716
rect 2800 2636 2840 2684
rect 2800 2604 2804 2636
rect 2836 2604 2840 2636
rect 2800 2556 2840 2604
rect 2800 2524 2804 2556
rect 2836 2524 2840 2556
rect 2800 2520 2840 2524
rect 2880 3596 2920 3600
rect 2880 3564 2884 3596
rect 2916 3564 2920 3596
rect 2880 3516 2920 3564
rect 2880 3484 2884 3516
rect 2916 3484 2920 3516
rect 2880 3436 2920 3484
rect 2880 3404 2884 3436
rect 2916 3404 2920 3436
rect 2880 3356 2920 3404
rect 2880 3324 2884 3356
rect 2916 3324 2920 3356
rect 2880 3276 2920 3324
rect 2880 3244 2884 3276
rect 2916 3244 2920 3276
rect 2880 3196 2920 3244
rect 2880 3164 2884 3196
rect 2916 3164 2920 3196
rect 2880 3116 2920 3164
rect 2880 3084 2884 3116
rect 2916 3084 2920 3116
rect 2880 3036 2920 3084
rect 2880 3004 2884 3036
rect 2916 3004 2920 3036
rect 2880 2956 2920 3004
rect 2880 2924 2884 2956
rect 2916 2924 2920 2956
rect 2880 2876 2920 2924
rect 2880 2844 2884 2876
rect 2916 2844 2920 2876
rect 2880 2796 2920 2844
rect 2880 2764 2884 2796
rect 2916 2764 2920 2796
rect 2880 2716 2920 2764
rect 2880 2684 2884 2716
rect 2916 2684 2920 2716
rect 2880 2636 2920 2684
rect 2880 2604 2884 2636
rect 2916 2604 2920 2636
rect 2880 2556 2920 2604
rect 2880 2524 2884 2556
rect 2916 2524 2920 2556
rect 2880 2520 2920 2524
rect 2960 3596 3000 3600
rect 2960 3564 2964 3596
rect 2996 3564 3000 3596
rect 2960 3516 3000 3564
rect 2960 3484 2964 3516
rect 2996 3484 3000 3516
rect 2960 3436 3000 3484
rect 2960 3404 2964 3436
rect 2996 3404 3000 3436
rect 2960 3356 3000 3404
rect 2960 3324 2964 3356
rect 2996 3324 3000 3356
rect 2960 3276 3000 3324
rect 2960 3244 2964 3276
rect 2996 3244 3000 3276
rect 2960 3196 3000 3244
rect 2960 3164 2964 3196
rect 2996 3164 3000 3196
rect 2960 3116 3000 3164
rect 2960 3084 2964 3116
rect 2996 3084 3000 3116
rect 2960 3036 3000 3084
rect 2960 3004 2964 3036
rect 2996 3004 3000 3036
rect 2960 2956 3000 3004
rect 2960 2924 2964 2956
rect 2996 2924 3000 2956
rect 2960 2876 3000 2924
rect 2960 2844 2964 2876
rect 2996 2844 3000 2876
rect 2960 2796 3000 2844
rect 2960 2764 2964 2796
rect 2996 2764 3000 2796
rect 2960 2716 3000 2764
rect 2960 2684 2964 2716
rect 2996 2684 3000 2716
rect 2960 2636 3000 2684
rect 2960 2604 2964 2636
rect 2996 2604 3000 2636
rect 2960 2556 3000 2604
rect 2960 2524 2964 2556
rect 2996 2524 3000 2556
rect 2960 2520 3000 2524
rect 3040 3596 3080 3600
rect 3040 3564 3044 3596
rect 3076 3564 3080 3596
rect 3040 3516 3080 3564
rect 3040 3484 3044 3516
rect 3076 3484 3080 3516
rect 3040 3436 3080 3484
rect 3040 3404 3044 3436
rect 3076 3404 3080 3436
rect 3040 3356 3080 3404
rect 3040 3324 3044 3356
rect 3076 3324 3080 3356
rect 3040 3276 3080 3324
rect 3040 3244 3044 3276
rect 3076 3244 3080 3276
rect 3040 3196 3080 3244
rect 3040 3164 3044 3196
rect 3076 3164 3080 3196
rect 3040 3116 3080 3164
rect 3040 3084 3044 3116
rect 3076 3084 3080 3116
rect 3040 3036 3080 3084
rect 3040 3004 3044 3036
rect 3076 3004 3080 3036
rect 3040 2956 3080 3004
rect 3040 2924 3044 2956
rect 3076 2924 3080 2956
rect 3040 2876 3080 2924
rect 3040 2844 3044 2876
rect 3076 2844 3080 2876
rect 3040 2796 3080 2844
rect 3040 2764 3044 2796
rect 3076 2764 3080 2796
rect 3040 2716 3080 2764
rect 3040 2684 3044 2716
rect 3076 2684 3080 2716
rect 3040 2636 3080 2684
rect 3040 2604 3044 2636
rect 3076 2604 3080 2636
rect 3040 2556 3080 2604
rect 3040 2524 3044 2556
rect 3076 2524 3080 2556
rect 3040 2520 3080 2524
rect 3120 3596 3160 3600
rect 3120 3564 3124 3596
rect 3156 3564 3160 3596
rect 3120 3516 3160 3564
rect 3120 3484 3124 3516
rect 3156 3484 3160 3516
rect 3120 3436 3160 3484
rect 3120 3404 3124 3436
rect 3156 3404 3160 3436
rect 3120 3356 3160 3404
rect 3120 3324 3124 3356
rect 3156 3324 3160 3356
rect 3120 3276 3160 3324
rect 3120 3244 3124 3276
rect 3156 3244 3160 3276
rect 3120 3196 3160 3244
rect 3120 3164 3124 3196
rect 3156 3164 3160 3196
rect 3120 3116 3160 3164
rect 3120 3084 3124 3116
rect 3156 3084 3160 3116
rect 3120 3036 3160 3084
rect 3120 3004 3124 3036
rect 3156 3004 3160 3036
rect 3120 2956 3160 3004
rect 3120 2924 3124 2956
rect 3156 2924 3160 2956
rect 3120 2876 3160 2924
rect 3120 2844 3124 2876
rect 3156 2844 3160 2876
rect 3120 2796 3160 2844
rect 3120 2764 3124 2796
rect 3156 2764 3160 2796
rect 3120 2716 3160 2764
rect 3120 2684 3124 2716
rect 3156 2684 3160 2716
rect 3120 2636 3160 2684
rect 3120 2604 3124 2636
rect 3156 2604 3160 2636
rect 3120 2556 3160 2604
rect 3120 2524 3124 2556
rect 3156 2524 3160 2556
rect 3120 2520 3160 2524
rect 3200 3596 3240 3600
rect 3200 3564 3204 3596
rect 3236 3564 3240 3596
rect 3200 3516 3240 3564
rect 3200 3484 3204 3516
rect 3236 3484 3240 3516
rect 3200 3436 3240 3484
rect 3200 3404 3204 3436
rect 3236 3404 3240 3436
rect 3200 3356 3240 3404
rect 3200 3324 3204 3356
rect 3236 3324 3240 3356
rect 3200 3276 3240 3324
rect 3200 3244 3204 3276
rect 3236 3244 3240 3276
rect 3200 3196 3240 3244
rect 3200 3164 3204 3196
rect 3236 3164 3240 3196
rect 3200 3116 3240 3164
rect 3200 3084 3204 3116
rect 3236 3084 3240 3116
rect 3200 3036 3240 3084
rect 3200 3004 3204 3036
rect 3236 3004 3240 3036
rect 3200 2956 3240 3004
rect 3200 2924 3204 2956
rect 3236 2924 3240 2956
rect 3200 2876 3240 2924
rect 3200 2844 3204 2876
rect 3236 2844 3240 2876
rect 3200 2796 3240 2844
rect 3200 2764 3204 2796
rect 3236 2764 3240 2796
rect 3200 2716 3240 2764
rect 3200 2684 3204 2716
rect 3236 2684 3240 2716
rect 3200 2636 3240 2684
rect 3200 2604 3204 2636
rect 3236 2604 3240 2636
rect 3200 2556 3240 2604
rect 3200 2524 3204 2556
rect 3236 2524 3240 2556
rect 3200 2520 3240 2524
rect 3280 3596 3320 3600
rect 3280 3564 3284 3596
rect 3316 3564 3320 3596
rect 3280 3516 3320 3564
rect 3280 3484 3284 3516
rect 3316 3484 3320 3516
rect 3280 3436 3320 3484
rect 3280 3404 3284 3436
rect 3316 3404 3320 3436
rect 3280 3356 3320 3404
rect 3280 3324 3284 3356
rect 3316 3324 3320 3356
rect 3280 3276 3320 3324
rect 3280 3244 3284 3276
rect 3316 3244 3320 3276
rect 3280 3196 3320 3244
rect 3280 3164 3284 3196
rect 3316 3164 3320 3196
rect 3280 3116 3320 3164
rect 3280 3084 3284 3116
rect 3316 3084 3320 3116
rect 3280 3036 3320 3084
rect 3280 3004 3284 3036
rect 3316 3004 3320 3036
rect 3280 2956 3320 3004
rect 3280 2924 3284 2956
rect 3316 2924 3320 2956
rect 3280 2876 3320 2924
rect 3280 2844 3284 2876
rect 3316 2844 3320 2876
rect 3280 2796 3320 2844
rect 3280 2764 3284 2796
rect 3316 2764 3320 2796
rect 3280 2716 3320 2764
rect 3280 2684 3284 2716
rect 3316 2684 3320 2716
rect 3280 2636 3320 2684
rect 3280 2604 3284 2636
rect 3316 2604 3320 2636
rect 3280 2556 3320 2604
rect 3280 2524 3284 2556
rect 3316 2524 3320 2556
rect 3280 2520 3320 2524
rect 3360 3596 3400 3600
rect 3360 3564 3364 3596
rect 3396 3564 3400 3596
rect 3360 3516 3400 3564
rect 3360 3484 3364 3516
rect 3396 3484 3400 3516
rect 3360 3436 3400 3484
rect 3360 3404 3364 3436
rect 3396 3404 3400 3436
rect 3360 3356 3400 3404
rect 3360 3324 3364 3356
rect 3396 3324 3400 3356
rect 3360 3276 3400 3324
rect 3360 3244 3364 3276
rect 3396 3244 3400 3276
rect 3360 3196 3400 3244
rect 3360 3164 3364 3196
rect 3396 3164 3400 3196
rect 3360 3116 3400 3164
rect 3360 3084 3364 3116
rect 3396 3084 3400 3116
rect 3360 3036 3400 3084
rect 3360 3004 3364 3036
rect 3396 3004 3400 3036
rect 3360 2956 3400 3004
rect 3360 2924 3364 2956
rect 3396 2924 3400 2956
rect 3360 2876 3400 2924
rect 3360 2844 3364 2876
rect 3396 2844 3400 2876
rect 3360 2796 3400 2844
rect 3360 2764 3364 2796
rect 3396 2764 3400 2796
rect 3360 2716 3400 2764
rect 3360 2684 3364 2716
rect 3396 2684 3400 2716
rect 3360 2636 3400 2684
rect 3360 2604 3364 2636
rect 3396 2604 3400 2636
rect 3360 2556 3400 2604
rect 3360 2524 3364 2556
rect 3396 2524 3400 2556
rect 3360 2520 3400 2524
rect 3440 3596 3480 3600
rect 3440 3564 3444 3596
rect 3476 3564 3480 3596
rect 3440 3516 3480 3564
rect 3440 3484 3444 3516
rect 3476 3484 3480 3516
rect 3440 3436 3480 3484
rect 3440 3404 3444 3436
rect 3476 3404 3480 3436
rect 3440 3356 3480 3404
rect 3440 3324 3444 3356
rect 3476 3324 3480 3356
rect 3440 3276 3480 3324
rect 3440 3244 3444 3276
rect 3476 3244 3480 3276
rect 3440 3196 3480 3244
rect 3440 3164 3444 3196
rect 3476 3164 3480 3196
rect 3440 3116 3480 3164
rect 3440 3084 3444 3116
rect 3476 3084 3480 3116
rect 3440 3036 3480 3084
rect 3440 3004 3444 3036
rect 3476 3004 3480 3036
rect 3440 2956 3480 3004
rect 3440 2924 3444 2956
rect 3476 2924 3480 2956
rect 3440 2876 3480 2924
rect 3440 2844 3444 2876
rect 3476 2844 3480 2876
rect 3440 2796 3480 2844
rect 3440 2764 3444 2796
rect 3476 2764 3480 2796
rect 3440 2716 3480 2764
rect 3440 2684 3444 2716
rect 3476 2684 3480 2716
rect 3440 2636 3480 2684
rect 3440 2604 3444 2636
rect 3476 2604 3480 2636
rect 3440 2556 3480 2604
rect 3440 2524 3444 2556
rect 3476 2524 3480 2556
rect 3440 2520 3480 2524
rect 3520 3596 3560 3600
rect 3520 3564 3524 3596
rect 3556 3564 3560 3596
rect 3520 3516 3560 3564
rect 3520 3484 3524 3516
rect 3556 3484 3560 3516
rect 3520 3436 3560 3484
rect 3520 3404 3524 3436
rect 3556 3404 3560 3436
rect 3520 3356 3560 3404
rect 3520 3324 3524 3356
rect 3556 3324 3560 3356
rect 3520 3276 3560 3324
rect 3520 3244 3524 3276
rect 3556 3244 3560 3276
rect 3520 3196 3560 3244
rect 3520 3164 3524 3196
rect 3556 3164 3560 3196
rect 3520 3116 3560 3164
rect 3520 3084 3524 3116
rect 3556 3084 3560 3116
rect 3520 3036 3560 3084
rect 3520 3004 3524 3036
rect 3556 3004 3560 3036
rect 3520 2956 3560 3004
rect 3520 2924 3524 2956
rect 3556 2924 3560 2956
rect 3520 2876 3560 2924
rect 3520 2844 3524 2876
rect 3556 2844 3560 2876
rect 3520 2796 3560 2844
rect 3520 2764 3524 2796
rect 3556 2764 3560 2796
rect 3520 2716 3560 2764
rect 3520 2684 3524 2716
rect 3556 2684 3560 2716
rect 3520 2636 3560 2684
rect 3520 2604 3524 2636
rect 3556 2604 3560 2636
rect 3520 2556 3560 2604
rect 3520 2524 3524 2556
rect 3556 2524 3560 2556
rect 3520 2520 3560 2524
rect 3600 3596 3640 3600
rect 3600 3564 3604 3596
rect 3636 3564 3640 3596
rect 3600 3516 3640 3564
rect 3600 3484 3604 3516
rect 3636 3484 3640 3516
rect 3600 3436 3640 3484
rect 3600 3404 3604 3436
rect 3636 3404 3640 3436
rect 3600 3356 3640 3404
rect 3600 3324 3604 3356
rect 3636 3324 3640 3356
rect 3600 3276 3640 3324
rect 3600 3244 3604 3276
rect 3636 3244 3640 3276
rect 3600 3196 3640 3244
rect 3600 3164 3604 3196
rect 3636 3164 3640 3196
rect 3600 3116 3640 3164
rect 3600 3084 3604 3116
rect 3636 3084 3640 3116
rect 3600 3036 3640 3084
rect 3600 3004 3604 3036
rect 3636 3004 3640 3036
rect 3600 2956 3640 3004
rect 3600 2924 3604 2956
rect 3636 2924 3640 2956
rect 3600 2876 3640 2924
rect 3600 2844 3604 2876
rect 3636 2844 3640 2876
rect 3600 2796 3640 2844
rect 3600 2764 3604 2796
rect 3636 2764 3640 2796
rect 3600 2716 3640 2764
rect 3600 2684 3604 2716
rect 3636 2684 3640 2716
rect 3600 2636 3640 2684
rect 3600 2604 3604 2636
rect 3636 2604 3640 2636
rect 3600 2556 3640 2604
rect 3600 2524 3604 2556
rect 3636 2524 3640 2556
rect 3600 2520 3640 2524
rect 3680 3596 3720 3600
rect 3680 3564 3684 3596
rect 3716 3564 3720 3596
rect 3680 3516 3720 3564
rect 3680 3484 3684 3516
rect 3716 3484 3720 3516
rect 3680 3436 3720 3484
rect 3680 3404 3684 3436
rect 3716 3404 3720 3436
rect 3680 3356 3720 3404
rect 3680 3324 3684 3356
rect 3716 3324 3720 3356
rect 3680 3276 3720 3324
rect 3680 3244 3684 3276
rect 3716 3244 3720 3276
rect 3680 3196 3720 3244
rect 3680 3164 3684 3196
rect 3716 3164 3720 3196
rect 3680 3116 3720 3164
rect 3680 3084 3684 3116
rect 3716 3084 3720 3116
rect 3680 3036 3720 3084
rect 3680 3004 3684 3036
rect 3716 3004 3720 3036
rect 3680 2956 3720 3004
rect 3680 2924 3684 2956
rect 3716 2924 3720 2956
rect 3680 2876 3720 2924
rect 3680 2844 3684 2876
rect 3716 2844 3720 2876
rect 3680 2796 3720 2844
rect 3680 2764 3684 2796
rect 3716 2764 3720 2796
rect 3680 2716 3720 2764
rect 3680 2684 3684 2716
rect 3716 2684 3720 2716
rect 3680 2636 3720 2684
rect 3680 2604 3684 2636
rect 3716 2604 3720 2636
rect 3680 2556 3720 2604
rect 3680 2524 3684 2556
rect 3716 2524 3720 2556
rect 3680 2520 3720 2524
rect 3760 3596 3800 3600
rect 3760 3564 3764 3596
rect 3796 3564 3800 3596
rect 3760 3516 3800 3564
rect 3760 3484 3764 3516
rect 3796 3484 3800 3516
rect 3760 3436 3800 3484
rect 3760 3404 3764 3436
rect 3796 3404 3800 3436
rect 3760 3356 3800 3404
rect 3760 3324 3764 3356
rect 3796 3324 3800 3356
rect 3760 3276 3800 3324
rect 3760 3244 3764 3276
rect 3796 3244 3800 3276
rect 3760 3196 3800 3244
rect 3760 3164 3764 3196
rect 3796 3164 3800 3196
rect 3760 3116 3800 3164
rect 3760 3084 3764 3116
rect 3796 3084 3800 3116
rect 3760 3036 3800 3084
rect 3760 3004 3764 3036
rect 3796 3004 3800 3036
rect 3760 2956 3800 3004
rect 3760 2924 3764 2956
rect 3796 2924 3800 2956
rect 3760 2876 3800 2924
rect 3760 2844 3764 2876
rect 3796 2844 3800 2876
rect 3760 2796 3800 2844
rect 3760 2764 3764 2796
rect 3796 2764 3800 2796
rect 3760 2716 3800 2764
rect 3760 2684 3764 2716
rect 3796 2684 3800 2716
rect 3760 2636 3800 2684
rect 3760 2604 3764 2636
rect 3796 2604 3800 2636
rect 3760 2556 3800 2604
rect 3760 2524 3764 2556
rect 3796 2524 3800 2556
rect 3760 2520 3800 2524
rect 3840 3596 3880 3600
rect 3840 3564 3844 3596
rect 3876 3564 3880 3596
rect 3840 3516 3880 3564
rect 3840 3484 3844 3516
rect 3876 3484 3880 3516
rect 3840 3436 3880 3484
rect 3840 3404 3844 3436
rect 3876 3404 3880 3436
rect 3840 3356 3880 3404
rect 3840 3324 3844 3356
rect 3876 3324 3880 3356
rect 3840 3276 3880 3324
rect 3840 3244 3844 3276
rect 3876 3244 3880 3276
rect 3840 3196 3880 3244
rect 3840 3164 3844 3196
rect 3876 3164 3880 3196
rect 3840 3116 3880 3164
rect 3840 3084 3844 3116
rect 3876 3084 3880 3116
rect 3840 3036 3880 3084
rect 3840 3004 3844 3036
rect 3876 3004 3880 3036
rect 3840 2956 3880 3004
rect 3840 2924 3844 2956
rect 3876 2924 3880 2956
rect 3840 2876 3880 2924
rect 3840 2844 3844 2876
rect 3876 2844 3880 2876
rect 3840 2796 3880 2844
rect 3840 2764 3844 2796
rect 3876 2764 3880 2796
rect 3840 2716 3880 2764
rect 3840 2684 3844 2716
rect 3876 2684 3880 2716
rect 3840 2636 3880 2684
rect 3840 2604 3844 2636
rect 3876 2604 3880 2636
rect 3840 2556 3880 2604
rect 3840 2524 3844 2556
rect 3876 2524 3880 2556
rect 3840 2520 3880 2524
rect 3920 3596 3960 3600
rect 3920 3564 3924 3596
rect 3956 3564 3960 3596
rect 3920 3516 3960 3564
rect 3920 3484 3924 3516
rect 3956 3484 3960 3516
rect 3920 3436 3960 3484
rect 3920 3404 3924 3436
rect 3956 3404 3960 3436
rect 3920 3356 3960 3404
rect 3920 3324 3924 3356
rect 3956 3324 3960 3356
rect 3920 3276 3960 3324
rect 3920 3244 3924 3276
rect 3956 3244 3960 3276
rect 3920 3196 3960 3244
rect 3920 3164 3924 3196
rect 3956 3164 3960 3196
rect 3920 3116 3960 3164
rect 3920 3084 3924 3116
rect 3956 3084 3960 3116
rect 3920 3036 3960 3084
rect 3920 3004 3924 3036
rect 3956 3004 3960 3036
rect 3920 2956 3960 3004
rect 3920 2924 3924 2956
rect 3956 2924 3960 2956
rect 3920 2876 3960 2924
rect 3920 2844 3924 2876
rect 3956 2844 3960 2876
rect 3920 2796 3960 2844
rect 3920 2764 3924 2796
rect 3956 2764 3960 2796
rect 3920 2716 3960 2764
rect 3920 2684 3924 2716
rect 3956 2684 3960 2716
rect 3920 2636 3960 2684
rect 3920 2604 3924 2636
rect 3956 2604 3960 2636
rect 3920 2556 3960 2604
rect 3920 2524 3924 2556
rect 3956 2524 3960 2556
rect 3920 2520 3960 2524
rect 4000 3596 4040 3600
rect 4000 3564 4004 3596
rect 4036 3564 4040 3596
rect 4000 3516 4040 3564
rect 4000 3484 4004 3516
rect 4036 3484 4040 3516
rect 4000 3436 4040 3484
rect 4000 3404 4004 3436
rect 4036 3404 4040 3436
rect 4000 3356 4040 3404
rect 4000 3324 4004 3356
rect 4036 3324 4040 3356
rect 4000 3276 4040 3324
rect 4000 3244 4004 3276
rect 4036 3244 4040 3276
rect 4000 3196 4040 3244
rect 4000 3164 4004 3196
rect 4036 3164 4040 3196
rect 4000 3116 4040 3164
rect 4000 3084 4004 3116
rect 4036 3084 4040 3116
rect 4000 3036 4040 3084
rect 4000 3004 4004 3036
rect 4036 3004 4040 3036
rect 4000 2956 4040 3004
rect 4000 2924 4004 2956
rect 4036 2924 4040 2956
rect 4000 2876 4040 2924
rect 4000 2844 4004 2876
rect 4036 2844 4040 2876
rect 4000 2796 4040 2844
rect 4000 2764 4004 2796
rect 4036 2764 4040 2796
rect 4000 2716 4040 2764
rect 4000 2684 4004 2716
rect 4036 2684 4040 2716
rect 4000 2636 4040 2684
rect 4000 2604 4004 2636
rect 4036 2604 4040 2636
rect 4000 2556 4040 2604
rect 4000 2524 4004 2556
rect 4036 2524 4040 2556
rect 4000 2520 4040 2524
rect 4080 3596 4120 3600
rect 4080 3564 4084 3596
rect 4116 3564 4120 3596
rect 4080 3516 4120 3564
rect 4080 3484 4084 3516
rect 4116 3484 4120 3516
rect 4080 3436 4120 3484
rect 4080 3404 4084 3436
rect 4116 3404 4120 3436
rect 4080 3356 4120 3404
rect 4080 3324 4084 3356
rect 4116 3324 4120 3356
rect 4080 3276 4120 3324
rect 4080 3244 4084 3276
rect 4116 3244 4120 3276
rect 4080 3196 4120 3244
rect 4080 3164 4084 3196
rect 4116 3164 4120 3196
rect 4080 3116 4120 3164
rect 4080 3084 4084 3116
rect 4116 3084 4120 3116
rect 4080 3036 4120 3084
rect 4080 3004 4084 3036
rect 4116 3004 4120 3036
rect 4080 2956 4120 3004
rect 4080 2924 4084 2956
rect 4116 2924 4120 2956
rect 4080 2876 4120 2924
rect 4080 2844 4084 2876
rect 4116 2844 4120 2876
rect 4080 2796 4120 2844
rect 4080 2764 4084 2796
rect 4116 2764 4120 2796
rect 4080 2716 4120 2764
rect 4080 2684 4084 2716
rect 4116 2684 4120 2716
rect 4080 2636 4120 2684
rect 4080 2604 4084 2636
rect 4116 2604 4120 2636
rect 4080 2556 4120 2604
rect 4080 2524 4084 2556
rect 4116 2524 4120 2556
rect 4080 2520 4120 2524
rect 4160 3596 4200 3600
rect 4160 3564 4164 3596
rect 4196 3564 4200 3596
rect 4160 3516 4200 3564
rect 4160 3484 4164 3516
rect 4196 3484 4200 3516
rect 4160 3436 4200 3484
rect 4160 3404 4164 3436
rect 4196 3404 4200 3436
rect 4160 3356 4200 3404
rect 4160 3324 4164 3356
rect 4196 3324 4200 3356
rect 4160 3276 4200 3324
rect 4160 3244 4164 3276
rect 4196 3244 4200 3276
rect 4160 3196 4200 3244
rect 4160 3164 4164 3196
rect 4196 3164 4200 3196
rect 4160 3116 4200 3164
rect 4160 3084 4164 3116
rect 4196 3084 4200 3116
rect 4160 3036 4200 3084
rect 4160 3004 4164 3036
rect 4196 3004 4200 3036
rect 4160 2956 4200 3004
rect 4160 2924 4164 2956
rect 4196 2924 4200 2956
rect 4160 2876 4200 2924
rect 4160 2844 4164 2876
rect 4196 2844 4200 2876
rect 4160 2796 4200 2844
rect 4160 2764 4164 2796
rect 4196 2764 4200 2796
rect 4160 2716 4200 2764
rect 4160 2684 4164 2716
rect 4196 2684 4200 2716
rect 4160 2636 4200 2684
rect 4160 2604 4164 2636
rect 4196 2604 4200 2636
rect 4160 2556 4200 2604
rect 4160 2524 4164 2556
rect 4196 2524 4200 2556
rect 4160 2520 4200 2524
rect 4240 3596 4280 3600
rect 4240 3564 4244 3596
rect 4276 3564 4280 3596
rect 4240 3516 4280 3564
rect 4240 3484 4244 3516
rect 4276 3484 4280 3516
rect 4240 3436 4280 3484
rect 4240 3404 4244 3436
rect 4276 3404 4280 3436
rect 4240 3356 4280 3404
rect 4240 3324 4244 3356
rect 4276 3324 4280 3356
rect 4240 3276 4280 3324
rect 4240 3244 4244 3276
rect 4276 3244 4280 3276
rect 4240 3196 4280 3244
rect 4240 3164 4244 3196
rect 4276 3164 4280 3196
rect 4240 3116 4280 3164
rect 4240 3084 4244 3116
rect 4276 3084 4280 3116
rect 4240 3036 4280 3084
rect 4240 3004 4244 3036
rect 4276 3004 4280 3036
rect 4240 2956 4280 3004
rect 4240 2924 4244 2956
rect 4276 2924 4280 2956
rect 4240 2876 4280 2924
rect 4240 2844 4244 2876
rect 4276 2844 4280 2876
rect 4240 2796 4280 2844
rect 4240 2764 4244 2796
rect 4276 2764 4280 2796
rect 4240 2716 4280 2764
rect 4240 2684 4244 2716
rect 4276 2684 4280 2716
rect 4240 2636 4280 2684
rect 4240 2604 4244 2636
rect 4276 2604 4280 2636
rect 4240 2556 4280 2604
rect 4240 2524 4244 2556
rect 4276 2524 4280 2556
rect 4240 2520 4280 2524
rect 4320 3596 4360 3600
rect 4320 3564 4324 3596
rect 4356 3564 4360 3596
rect 4320 3516 4360 3564
rect 4320 3484 4324 3516
rect 4356 3484 4360 3516
rect 4320 3436 4360 3484
rect 4320 3404 4324 3436
rect 4356 3404 4360 3436
rect 4320 3356 4360 3404
rect 4320 3324 4324 3356
rect 4356 3324 4360 3356
rect 4320 3276 4360 3324
rect 4320 3244 4324 3276
rect 4356 3244 4360 3276
rect 4320 3196 4360 3244
rect 4320 3164 4324 3196
rect 4356 3164 4360 3196
rect 4320 3116 4360 3164
rect 4320 3084 4324 3116
rect 4356 3084 4360 3116
rect 4320 3036 4360 3084
rect 4320 3004 4324 3036
rect 4356 3004 4360 3036
rect 4320 2956 4360 3004
rect 4320 2924 4324 2956
rect 4356 2924 4360 2956
rect 4320 2876 4360 2924
rect 4320 2844 4324 2876
rect 4356 2844 4360 2876
rect 4320 2796 4360 2844
rect 4320 2764 4324 2796
rect 4356 2764 4360 2796
rect 4320 2716 4360 2764
rect 4320 2684 4324 2716
rect 4356 2684 4360 2716
rect 4320 2636 4360 2684
rect 4320 2604 4324 2636
rect 4356 2604 4360 2636
rect 4320 2556 4360 2604
rect 4320 2524 4324 2556
rect 4356 2524 4360 2556
rect 4320 2520 4360 2524
rect 4400 3596 4440 3600
rect 4400 3564 4404 3596
rect 4436 3564 4440 3596
rect 4400 3516 4440 3564
rect 4400 3484 4404 3516
rect 4436 3484 4440 3516
rect 4400 3436 4440 3484
rect 4400 3404 4404 3436
rect 4436 3404 4440 3436
rect 4400 3356 4440 3404
rect 4400 3324 4404 3356
rect 4436 3324 4440 3356
rect 4400 3276 4440 3324
rect 4400 3244 4404 3276
rect 4436 3244 4440 3276
rect 4400 3196 4440 3244
rect 4400 3164 4404 3196
rect 4436 3164 4440 3196
rect 4400 3116 4440 3164
rect 4400 3084 4404 3116
rect 4436 3084 4440 3116
rect 4400 3036 4440 3084
rect 4400 3004 4404 3036
rect 4436 3004 4440 3036
rect 4400 2956 4440 3004
rect 4400 2924 4404 2956
rect 4436 2924 4440 2956
rect 4400 2876 4440 2924
rect 4400 2844 4404 2876
rect 4436 2844 4440 2876
rect 4400 2796 4440 2844
rect 4400 2764 4404 2796
rect 4436 2764 4440 2796
rect 4400 2716 4440 2764
rect 4400 2684 4404 2716
rect 4436 2684 4440 2716
rect 4400 2636 4440 2684
rect 4400 2604 4404 2636
rect 4436 2604 4440 2636
rect 4400 2556 4440 2604
rect 4400 2524 4404 2556
rect 4436 2524 4440 2556
rect 4400 2520 4440 2524
rect 4480 3596 4520 3600
rect 4480 3564 4484 3596
rect 4516 3564 4520 3596
rect 4480 3516 4520 3564
rect 4480 3484 4484 3516
rect 4516 3484 4520 3516
rect 4480 3436 4520 3484
rect 4480 3404 4484 3436
rect 4516 3404 4520 3436
rect 4480 3356 4520 3404
rect 4480 3324 4484 3356
rect 4516 3324 4520 3356
rect 4480 3276 4520 3324
rect 4480 3244 4484 3276
rect 4516 3244 4520 3276
rect 4480 3196 4520 3244
rect 4480 3164 4484 3196
rect 4516 3164 4520 3196
rect 4480 3116 4520 3164
rect 4480 3084 4484 3116
rect 4516 3084 4520 3116
rect 4480 3036 4520 3084
rect 4480 3004 4484 3036
rect 4516 3004 4520 3036
rect 4480 2956 4520 3004
rect 4480 2924 4484 2956
rect 4516 2924 4520 2956
rect 4480 2876 4520 2924
rect 4480 2844 4484 2876
rect 4516 2844 4520 2876
rect 4480 2796 4520 2844
rect 4480 2764 4484 2796
rect 4516 2764 4520 2796
rect 4480 2716 4520 2764
rect 4480 2684 4484 2716
rect 4516 2684 4520 2716
rect 4480 2636 4520 2684
rect 4480 2604 4484 2636
rect 4516 2604 4520 2636
rect 4480 2556 4520 2604
rect 4480 2524 4484 2556
rect 4516 2524 4520 2556
rect 4480 2520 4520 2524
rect 4560 3596 4600 3600
rect 4560 3564 4564 3596
rect 4596 3564 4600 3596
rect 4560 3516 4600 3564
rect 4560 3484 4564 3516
rect 4596 3484 4600 3516
rect 4560 3436 4600 3484
rect 4560 3404 4564 3436
rect 4596 3404 4600 3436
rect 4560 3356 4600 3404
rect 4560 3324 4564 3356
rect 4596 3324 4600 3356
rect 4560 3276 4600 3324
rect 4560 3244 4564 3276
rect 4596 3244 4600 3276
rect 4560 3196 4600 3244
rect 4560 3164 4564 3196
rect 4596 3164 4600 3196
rect 4560 3116 4600 3164
rect 4560 3084 4564 3116
rect 4596 3084 4600 3116
rect 4560 3036 4600 3084
rect 4560 3004 4564 3036
rect 4596 3004 4600 3036
rect 4560 2956 4600 3004
rect 4560 2924 4564 2956
rect 4596 2924 4600 2956
rect 4560 2876 4600 2924
rect 4560 2844 4564 2876
rect 4596 2844 4600 2876
rect 4560 2796 4600 2844
rect 4560 2764 4564 2796
rect 4596 2764 4600 2796
rect 4560 2716 4600 2764
rect 4560 2684 4564 2716
rect 4596 2684 4600 2716
rect 4560 2636 4600 2684
rect 4560 2604 4564 2636
rect 4596 2604 4600 2636
rect 4560 2556 4600 2604
rect 4560 2524 4564 2556
rect 4596 2524 4600 2556
rect 4560 2520 4600 2524
rect 4640 3596 4680 3600
rect 4640 3564 4644 3596
rect 4676 3564 4680 3596
rect 4640 3516 4680 3564
rect 4640 3484 4644 3516
rect 4676 3484 4680 3516
rect 4640 3436 4680 3484
rect 4640 3404 4644 3436
rect 4676 3404 4680 3436
rect 4640 3356 4680 3404
rect 4640 3324 4644 3356
rect 4676 3324 4680 3356
rect 4640 3276 4680 3324
rect 4640 3244 4644 3276
rect 4676 3244 4680 3276
rect 4640 3196 4680 3244
rect 4640 3164 4644 3196
rect 4676 3164 4680 3196
rect 4640 3116 4680 3164
rect 4640 3084 4644 3116
rect 4676 3084 4680 3116
rect 4640 3036 4680 3084
rect 4640 3004 4644 3036
rect 4676 3004 4680 3036
rect 4640 2956 4680 3004
rect 4640 2924 4644 2956
rect 4676 2924 4680 2956
rect 4640 2876 4680 2924
rect 4640 2844 4644 2876
rect 4676 2844 4680 2876
rect 4640 2796 4680 2844
rect 4640 2764 4644 2796
rect 4676 2764 4680 2796
rect 4640 2716 4680 2764
rect 4640 2684 4644 2716
rect 4676 2684 4680 2716
rect 4640 2636 4680 2684
rect 4640 2604 4644 2636
rect 4676 2604 4680 2636
rect 4640 2556 4680 2604
rect 4640 2524 4644 2556
rect 4676 2524 4680 2556
rect 4640 2520 4680 2524
rect 4720 3596 4760 3600
rect 4720 3564 4724 3596
rect 4756 3564 4760 3596
rect 4720 3516 4760 3564
rect 4720 3484 4724 3516
rect 4756 3484 4760 3516
rect 4720 3436 4760 3484
rect 4720 3404 4724 3436
rect 4756 3404 4760 3436
rect 4720 3356 4760 3404
rect 4720 3324 4724 3356
rect 4756 3324 4760 3356
rect 4720 3276 4760 3324
rect 4720 3244 4724 3276
rect 4756 3244 4760 3276
rect 4720 3196 4760 3244
rect 4720 3164 4724 3196
rect 4756 3164 4760 3196
rect 4720 3116 4760 3164
rect 4720 3084 4724 3116
rect 4756 3084 4760 3116
rect 4720 3036 4760 3084
rect 4720 3004 4724 3036
rect 4756 3004 4760 3036
rect 4720 2956 4760 3004
rect 4720 2924 4724 2956
rect 4756 2924 4760 2956
rect 4720 2876 4760 2924
rect 4720 2844 4724 2876
rect 4756 2844 4760 2876
rect 4720 2796 4760 2844
rect 4720 2764 4724 2796
rect 4756 2764 4760 2796
rect 4720 2716 4760 2764
rect 4720 2684 4724 2716
rect 4756 2684 4760 2716
rect 4720 2636 4760 2684
rect 4720 2604 4724 2636
rect 4756 2604 4760 2636
rect 4720 2556 4760 2604
rect 4720 2524 4724 2556
rect 4756 2524 4760 2556
rect 4720 2520 4760 2524
rect 4800 3596 4840 3600
rect 4800 3564 4804 3596
rect 4836 3564 4840 3596
rect 4800 3516 4840 3564
rect 4800 3484 4804 3516
rect 4836 3484 4840 3516
rect 4800 3436 4840 3484
rect 4800 3404 4804 3436
rect 4836 3404 4840 3436
rect 4800 3356 4840 3404
rect 4800 3324 4804 3356
rect 4836 3324 4840 3356
rect 4800 3276 4840 3324
rect 4800 3244 4804 3276
rect 4836 3244 4840 3276
rect 4800 3196 4840 3244
rect 4800 3164 4804 3196
rect 4836 3164 4840 3196
rect 4800 3116 4840 3164
rect 4800 3084 4804 3116
rect 4836 3084 4840 3116
rect 4800 3036 4840 3084
rect 4800 3004 4804 3036
rect 4836 3004 4840 3036
rect 4800 2956 4840 3004
rect 4800 2924 4804 2956
rect 4836 2924 4840 2956
rect 4800 2876 4840 2924
rect 4800 2844 4804 2876
rect 4836 2844 4840 2876
rect 4800 2796 4840 2844
rect 4800 2764 4804 2796
rect 4836 2764 4840 2796
rect 4800 2716 4840 2764
rect 4800 2684 4804 2716
rect 4836 2684 4840 2716
rect 4800 2636 4840 2684
rect 4800 2604 4804 2636
rect 4836 2604 4840 2636
rect 4800 2556 4840 2604
rect 4800 2524 4804 2556
rect 4836 2524 4840 2556
rect 4800 2520 4840 2524
rect 4880 3596 4920 3644
rect 4880 3564 4884 3596
rect 4916 3564 4920 3596
rect 4880 3516 4920 3564
rect 4880 3484 4884 3516
rect 4916 3484 4920 3516
rect 4880 3436 4920 3484
rect 4880 3404 4884 3436
rect 4916 3404 4920 3436
rect 4880 3356 4920 3404
rect 4880 3324 4884 3356
rect 4916 3324 4920 3356
rect 4880 3276 4920 3324
rect 4880 3244 4884 3276
rect 4916 3244 4920 3276
rect 4880 3196 4920 3244
rect 4880 3164 4884 3196
rect 4916 3164 4920 3196
rect 4880 3116 4920 3164
rect 4880 3084 4884 3116
rect 4916 3084 4920 3116
rect 4880 3036 4920 3084
rect 4880 3004 4884 3036
rect 4916 3004 4920 3036
rect 4880 2956 4920 3004
rect 4880 2924 4884 2956
rect 4916 2924 4920 2956
rect 4880 2876 4920 2924
rect 4880 2844 4884 2876
rect 4916 2844 4920 2876
rect 4880 2796 4920 2844
rect 4880 2764 4884 2796
rect 4916 2764 4920 2796
rect 4880 2716 4920 2764
rect 4880 2684 4884 2716
rect 4916 2684 4920 2716
rect 4880 2636 4920 2684
rect 4880 2604 4884 2636
rect 4916 2604 4920 2636
rect 4880 2556 4920 2604
rect 4880 2524 4884 2556
rect 4916 2524 4920 2556
rect -880 2444 -876 2476
rect -844 2444 -840 2476
rect -880 2396 -840 2444
rect -880 2364 -876 2396
rect -844 2364 -840 2396
rect -880 2316 -840 2364
rect -880 2284 -876 2316
rect -844 2284 -840 2316
rect -880 2236 -840 2284
rect -880 2204 -876 2236
rect -844 2204 -840 2236
rect -880 2156 -840 2204
rect -880 2124 -876 2156
rect -844 2124 -840 2156
rect -880 2076 -840 2124
rect -880 2044 -876 2076
rect -844 2044 -840 2076
rect -880 1996 -840 2044
rect -880 1964 -876 1996
rect -844 1964 -840 1996
rect -880 1916 -840 1964
rect -880 1884 -876 1916
rect -844 1884 -840 1916
rect -880 1836 -840 1884
rect -880 1804 -876 1836
rect -844 1804 -840 1836
rect -880 1756 -840 1804
rect -880 1724 -876 1756
rect -844 1724 -840 1756
rect -880 1676 -840 1724
rect -800 2476 -760 2480
rect -800 2444 -796 2476
rect -764 2444 -760 2476
rect -800 2396 -760 2444
rect -800 2364 -796 2396
rect -764 2364 -760 2396
rect -800 2316 -760 2364
rect -800 2284 -796 2316
rect -764 2284 -760 2316
rect -800 2236 -760 2284
rect -800 2204 -796 2236
rect -764 2204 -760 2236
rect -800 2156 -760 2204
rect -800 2124 -796 2156
rect -764 2124 -760 2156
rect -800 2076 -760 2124
rect -800 2044 -796 2076
rect -764 2044 -760 2076
rect -800 1996 -760 2044
rect -800 1964 -796 1996
rect -764 1964 -760 1996
rect -800 1916 -760 1964
rect -800 1884 -796 1916
rect -764 1884 -760 1916
rect -800 1836 -760 1884
rect -800 1804 -796 1836
rect -764 1804 -760 1836
rect -800 1756 -760 1804
rect -800 1724 -796 1756
rect -764 1724 -760 1756
rect -800 1720 -760 1724
rect -720 2476 -680 2480
rect -720 2444 -716 2476
rect -684 2444 -680 2476
rect -720 2396 -680 2444
rect -720 2364 -716 2396
rect -684 2364 -680 2396
rect -720 2316 -680 2364
rect -720 2284 -716 2316
rect -684 2284 -680 2316
rect -720 2236 -680 2284
rect -720 2204 -716 2236
rect -684 2204 -680 2236
rect -720 2156 -680 2204
rect -720 2124 -716 2156
rect -684 2124 -680 2156
rect -720 2076 -680 2124
rect -720 2044 -716 2076
rect -684 2044 -680 2076
rect -720 1996 -680 2044
rect -720 1964 -716 1996
rect -684 1964 -680 1996
rect -720 1916 -680 1964
rect -720 1884 -716 1916
rect -684 1884 -680 1916
rect -720 1836 -680 1884
rect -720 1804 -716 1836
rect -684 1804 -680 1836
rect -720 1756 -680 1804
rect -720 1724 -716 1756
rect -684 1724 -680 1756
rect -720 1720 -680 1724
rect -640 2476 -600 2480
rect -640 2444 -636 2476
rect -604 2444 -600 2476
rect -640 2396 -600 2444
rect -640 2364 -636 2396
rect -604 2364 -600 2396
rect -640 2316 -600 2364
rect -640 2284 -636 2316
rect -604 2284 -600 2316
rect -640 2236 -600 2284
rect -640 2204 -636 2236
rect -604 2204 -600 2236
rect -640 2156 -600 2204
rect -640 2124 -636 2156
rect -604 2124 -600 2156
rect -640 2076 -600 2124
rect -640 2044 -636 2076
rect -604 2044 -600 2076
rect -640 1996 -600 2044
rect -640 1964 -636 1996
rect -604 1964 -600 1996
rect -640 1916 -600 1964
rect -640 1884 -636 1916
rect -604 1884 -600 1916
rect -640 1836 -600 1884
rect -640 1804 -636 1836
rect -604 1804 -600 1836
rect -640 1756 -600 1804
rect -640 1724 -636 1756
rect -604 1724 -600 1756
rect -640 1720 -600 1724
rect -560 2476 -520 2480
rect -560 2444 -556 2476
rect -524 2444 -520 2476
rect -560 2396 -520 2444
rect -560 2364 -556 2396
rect -524 2364 -520 2396
rect -560 2316 -520 2364
rect -560 2284 -556 2316
rect -524 2284 -520 2316
rect -560 2236 -520 2284
rect -560 2204 -556 2236
rect -524 2204 -520 2236
rect -560 2156 -520 2204
rect -560 2124 -556 2156
rect -524 2124 -520 2156
rect -560 2076 -520 2124
rect -560 2044 -556 2076
rect -524 2044 -520 2076
rect -560 1996 -520 2044
rect -560 1964 -556 1996
rect -524 1964 -520 1996
rect -560 1916 -520 1964
rect -560 1884 -556 1916
rect -524 1884 -520 1916
rect -560 1836 -520 1884
rect -560 1804 -556 1836
rect -524 1804 -520 1836
rect -560 1756 -520 1804
rect -560 1724 -556 1756
rect -524 1724 -520 1756
rect -560 1720 -520 1724
rect -480 2476 -440 2480
rect -480 2444 -476 2476
rect -444 2444 -440 2476
rect -480 2396 -440 2444
rect -480 2364 -476 2396
rect -444 2364 -440 2396
rect -480 2316 -440 2364
rect -480 2284 -476 2316
rect -444 2284 -440 2316
rect -480 2236 -440 2284
rect -480 2204 -476 2236
rect -444 2204 -440 2236
rect -480 2156 -440 2204
rect -480 2124 -476 2156
rect -444 2124 -440 2156
rect -480 2076 -440 2124
rect -480 2044 -476 2076
rect -444 2044 -440 2076
rect -480 1996 -440 2044
rect -480 1964 -476 1996
rect -444 1964 -440 1996
rect -480 1916 -440 1964
rect -480 1884 -476 1916
rect -444 1884 -440 1916
rect -480 1836 -440 1884
rect -480 1804 -476 1836
rect -444 1804 -440 1836
rect -480 1756 -440 1804
rect -480 1724 -476 1756
rect -444 1724 -440 1756
rect -480 1720 -440 1724
rect -400 2476 -360 2480
rect -400 2444 -396 2476
rect -364 2444 -360 2476
rect -400 2396 -360 2444
rect -400 2364 -396 2396
rect -364 2364 -360 2396
rect -400 2316 -360 2364
rect -400 2284 -396 2316
rect -364 2284 -360 2316
rect -400 2236 -360 2284
rect -400 2204 -396 2236
rect -364 2204 -360 2236
rect -400 2156 -360 2204
rect -400 2124 -396 2156
rect -364 2124 -360 2156
rect -400 2076 -360 2124
rect -400 2044 -396 2076
rect -364 2044 -360 2076
rect -400 1996 -360 2044
rect -400 1964 -396 1996
rect -364 1964 -360 1996
rect -400 1916 -360 1964
rect -400 1884 -396 1916
rect -364 1884 -360 1916
rect -400 1836 -360 1884
rect -400 1804 -396 1836
rect -364 1804 -360 1836
rect -400 1756 -360 1804
rect -400 1724 -396 1756
rect -364 1724 -360 1756
rect -400 1720 -360 1724
rect -320 2476 -280 2480
rect -320 2444 -316 2476
rect -284 2444 -280 2476
rect -320 2396 -280 2444
rect -320 2364 -316 2396
rect -284 2364 -280 2396
rect -320 2316 -280 2364
rect -320 2284 -316 2316
rect -284 2284 -280 2316
rect -320 2236 -280 2284
rect -320 2204 -316 2236
rect -284 2204 -280 2236
rect -320 2156 -280 2204
rect -320 2124 -316 2156
rect -284 2124 -280 2156
rect -320 2076 -280 2124
rect -320 2044 -316 2076
rect -284 2044 -280 2076
rect -320 1996 -280 2044
rect -320 1964 -316 1996
rect -284 1964 -280 1996
rect -320 1916 -280 1964
rect -320 1884 -316 1916
rect -284 1884 -280 1916
rect -320 1836 -280 1884
rect -320 1804 -316 1836
rect -284 1804 -280 1836
rect -320 1756 -280 1804
rect -320 1724 -316 1756
rect -284 1724 -280 1756
rect -320 1720 -280 1724
rect -240 2476 -200 2480
rect -240 2444 -236 2476
rect -204 2444 -200 2476
rect -240 2396 -200 2444
rect -240 2364 -236 2396
rect -204 2364 -200 2396
rect -240 2316 -200 2364
rect -240 2284 -236 2316
rect -204 2284 -200 2316
rect -240 2236 -200 2284
rect -240 2204 -236 2236
rect -204 2204 -200 2236
rect -240 2156 -200 2204
rect -240 2124 -236 2156
rect -204 2124 -200 2156
rect -240 2076 -200 2124
rect -240 2044 -236 2076
rect -204 2044 -200 2076
rect -240 1996 -200 2044
rect -240 1964 -236 1996
rect -204 1964 -200 1996
rect -240 1916 -200 1964
rect -240 1884 -236 1916
rect -204 1884 -200 1916
rect -240 1836 -200 1884
rect -240 1804 -236 1836
rect -204 1804 -200 1836
rect -240 1756 -200 1804
rect -240 1724 -236 1756
rect -204 1724 -200 1756
rect -240 1720 -200 1724
rect -160 2476 -120 2480
rect -160 2444 -156 2476
rect -124 2444 -120 2476
rect -160 2396 -120 2444
rect -160 2364 -156 2396
rect -124 2364 -120 2396
rect -160 2316 -120 2364
rect -160 2284 -156 2316
rect -124 2284 -120 2316
rect -160 2236 -120 2284
rect -160 2204 -156 2236
rect -124 2204 -120 2236
rect -160 2156 -120 2204
rect -160 2124 -156 2156
rect -124 2124 -120 2156
rect -160 2076 -120 2124
rect -160 2044 -156 2076
rect -124 2044 -120 2076
rect -160 1996 -120 2044
rect -160 1964 -156 1996
rect -124 1964 -120 1996
rect -160 1916 -120 1964
rect -160 1884 -156 1916
rect -124 1884 -120 1916
rect -160 1836 -120 1884
rect -160 1804 -156 1836
rect -124 1804 -120 1836
rect -160 1756 -120 1804
rect -160 1724 -156 1756
rect -124 1724 -120 1756
rect -160 1720 -120 1724
rect -80 2476 -40 2480
rect -80 2444 -76 2476
rect -44 2444 -40 2476
rect -80 2396 -40 2444
rect -80 2364 -76 2396
rect -44 2364 -40 2396
rect -80 2316 -40 2364
rect -80 2284 -76 2316
rect -44 2284 -40 2316
rect -80 2236 -40 2284
rect -80 2204 -76 2236
rect -44 2204 -40 2236
rect -80 2156 -40 2204
rect -80 2124 -76 2156
rect -44 2124 -40 2156
rect -80 2076 -40 2124
rect -80 2044 -76 2076
rect -44 2044 -40 2076
rect -80 1996 -40 2044
rect -80 1964 -76 1996
rect -44 1964 -40 1996
rect -80 1916 -40 1964
rect -80 1884 -76 1916
rect -44 1884 -40 1916
rect -80 1836 -40 1884
rect -80 1804 -76 1836
rect -44 1804 -40 1836
rect -80 1756 -40 1804
rect -80 1724 -76 1756
rect -44 1724 -40 1756
rect -80 1720 -40 1724
rect 0 2476 40 2480
rect 0 2444 4 2476
rect 36 2444 40 2476
rect 0 2396 40 2444
rect 0 2364 4 2396
rect 36 2364 40 2396
rect 0 2316 40 2364
rect 0 2284 4 2316
rect 36 2284 40 2316
rect 0 2236 40 2284
rect 0 2204 4 2236
rect 36 2204 40 2236
rect 0 2156 40 2204
rect 0 2124 4 2156
rect 36 2124 40 2156
rect 0 2076 40 2124
rect 0 2044 4 2076
rect 36 2044 40 2076
rect 0 1996 40 2044
rect 0 1964 4 1996
rect 36 1964 40 1996
rect 0 1916 40 1964
rect 0 1884 4 1916
rect 36 1884 40 1916
rect 0 1836 40 1884
rect 0 1804 4 1836
rect 36 1804 40 1836
rect 0 1756 40 1804
rect 0 1724 4 1756
rect 36 1724 40 1756
rect 0 1720 40 1724
rect 80 2476 120 2480
rect 80 2444 84 2476
rect 116 2444 120 2476
rect 80 2396 120 2444
rect 80 2364 84 2396
rect 116 2364 120 2396
rect 80 2316 120 2364
rect 80 2284 84 2316
rect 116 2284 120 2316
rect 80 2236 120 2284
rect 80 2204 84 2236
rect 116 2204 120 2236
rect 80 2156 120 2204
rect 80 2124 84 2156
rect 116 2124 120 2156
rect 80 2076 120 2124
rect 80 2044 84 2076
rect 116 2044 120 2076
rect 80 1996 120 2044
rect 80 1964 84 1996
rect 116 1964 120 1996
rect 80 1916 120 1964
rect 80 1884 84 1916
rect 116 1884 120 1916
rect 80 1836 120 1884
rect 80 1804 84 1836
rect 116 1804 120 1836
rect 80 1756 120 1804
rect 80 1724 84 1756
rect 116 1724 120 1756
rect 80 1720 120 1724
rect 160 2476 200 2480
rect 160 2444 164 2476
rect 196 2444 200 2476
rect 160 2396 200 2444
rect 160 2364 164 2396
rect 196 2364 200 2396
rect 160 2316 200 2364
rect 160 2284 164 2316
rect 196 2284 200 2316
rect 160 2236 200 2284
rect 160 2204 164 2236
rect 196 2204 200 2236
rect 160 2156 200 2204
rect 160 2124 164 2156
rect 196 2124 200 2156
rect 160 2076 200 2124
rect 160 2044 164 2076
rect 196 2044 200 2076
rect 160 1996 200 2044
rect 160 1964 164 1996
rect 196 1964 200 1996
rect 160 1916 200 1964
rect 160 1884 164 1916
rect 196 1884 200 1916
rect 160 1836 200 1884
rect 160 1804 164 1836
rect 196 1804 200 1836
rect 160 1756 200 1804
rect 160 1724 164 1756
rect 196 1724 200 1756
rect 160 1720 200 1724
rect 240 2476 280 2480
rect 240 2444 244 2476
rect 276 2444 280 2476
rect 240 2396 280 2444
rect 240 2364 244 2396
rect 276 2364 280 2396
rect 240 2316 280 2364
rect 240 2284 244 2316
rect 276 2284 280 2316
rect 240 2236 280 2284
rect 240 2204 244 2236
rect 276 2204 280 2236
rect 240 2156 280 2204
rect 240 2124 244 2156
rect 276 2124 280 2156
rect 240 2076 280 2124
rect 240 2044 244 2076
rect 276 2044 280 2076
rect 240 1996 280 2044
rect 240 1964 244 1996
rect 276 1964 280 1996
rect 240 1916 280 1964
rect 240 1884 244 1916
rect 276 1884 280 1916
rect 240 1836 280 1884
rect 240 1804 244 1836
rect 276 1804 280 1836
rect 240 1756 280 1804
rect 240 1724 244 1756
rect 276 1724 280 1756
rect 240 1720 280 1724
rect 320 2476 360 2480
rect 320 2444 324 2476
rect 356 2444 360 2476
rect 320 2396 360 2444
rect 320 2364 324 2396
rect 356 2364 360 2396
rect 320 2316 360 2364
rect 320 2284 324 2316
rect 356 2284 360 2316
rect 320 2236 360 2284
rect 320 2204 324 2236
rect 356 2204 360 2236
rect 320 2156 360 2204
rect 320 2124 324 2156
rect 356 2124 360 2156
rect 320 2076 360 2124
rect 320 2044 324 2076
rect 356 2044 360 2076
rect 320 1996 360 2044
rect 320 1964 324 1996
rect 356 1964 360 1996
rect 320 1916 360 1964
rect 320 1884 324 1916
rect 356 1884 360 1916
rect 320 1836 360 1884
rect 320 1804 324 1836
rect 356 1804 360 1836
rect 320 1756 360 1804
rect 320 1724 324 1756
rect 356 1724 360 1756
rect 320 1720 360 1724
rect 400 2476 440 2480
rect 400 2444 404 2476
rect 436 2444 440 2476
rect 400 2396 440 2444
rect 400 2364 404 2396
rect 436 2364 440 2396
rect 400 2316 440 2364
rect 400 2284 404 2316
rect 436 2284 440 2316
rect 400 2236 440 2284
rect 400 2204 404 2236
rect 436 2204 440 2236
rect 400 2156 440 2204
rect 400 2124 404 2156
rect 436 2124 440 2156
rect 400 2076 440 2124
rect 400 2044 404 2076
rect 436 2044 440 2076
rect 400 1996 440 2044
rect 400 1964 404 1996
rect 436 1964 440 1996
rect 400 1916 440 1964
rect 400 1884 404 1916
rect 436 1884 440 1916
rect 400 1836 440 1884
rect 400 1804 404 1836
rect 436 1804 440 1836
rect 400 1756 440 1804
rect 400 1724 404 1756
rect 436 1724 440 1756
rect 400 1720 440 1724
rect 480 2476 520 2480
rect 480 2444 484 2476
rect 516 2444 520 2476
rect 480 2396 520 2444
rect 480 2364 484 2396
rect 516 2364 520 2396
rect 480 2316 520 2364
rect 480 2284 484 2316
rect 516 2284 520 2316
rect 480 2236 520 2284
rect 480 2204 484 2236
rect 516 2204 520 2236
rect 480 2156 520 2204
rect 480 2124 484 2156
rect 516 2124 520 2156
rect 480 2076 520 2124
rect 480 2044 484 2076
rect 516 2044 520 2076
rect 480 1996 520 2044
rect 480 1964 484 1996
rect 516 1964 520 1996
rect 480 1916 520 1964
rect 480 1884 484 1916
rect 516 1884 520 1916
rect 480 1836 520 1884
rect 480 1804 484 1836
rect 516 1804 520 1836
rect 480 1756 520 1804
rect 480 1724 484 1756
rect 516 1724 520 1756
rect 480 1720 520 1724
rect 560 2476 600 2480
rect 560 2444 564 2476
rect 596 2444 600 2476
rect 560 2396 600 2444
rect 560 2364 564 2396
rect 596 2364 600 2396
rect 560 2316 600 2364
rect 560 2284 564 2316
rect 596 2284 600 2316
rect 560 2236 600 2284
rect 560 2204 564 2236
rect 596 2204 600 2236
rect 560 2156 600 2204
rect 560 2124 564 2156
rect 596 2124 600 2156
rect 560 2076 600 2124
rect 560 2044 564 2076
rect 596 2044 600 2076
rect 560 1996 600 2044
rect 560 1964 564 1996
rect 596 1964 600 1996
rect 560 1916 600 1964
rect 560 1884 564 1916
rect 596 1884 600 1916
rect 560 1836 600 1884
rect 560 1804 564 1836
rect 596 1804 600 1836
rect 560 1756 600 1804
rect 560 1724 564 1756
rect 596 1724 600 1756
rect 560 1720 600 1724
rect 640 2476 680 2480
rect 640 2444 644 2476
rect 676 2444 680 2476
rect 640 2396 680 2444
rect 640 2364 644 2396
rect 676 2364 680 2396
rect 640 2316 680 2364
rect 640 2284 644 2316
rect 676 2284 680 2316
rect 640 2236 680 2284
rect 640 2204 644 2236
rect 676 2204 680 2236
rect 640 2156 680 2204
rect 640 2124 644 2156
rect 676 2124 680 2156
rect 640 2076 680 2124
rect 640 2044 644 2076
rect 676 2044 680 2076
rect 640 1996 680 2044
rect 640 1964 644 1996
rect 676 1964 680 1996
rect 640 1916 680 1964
rect 640 1884 644 1916
rect 676 1884 680 1916
rect 640 1836 680 1884
rect 640 1804 644 1836
rect 676 1804 680 1836
rect 640 1756 680 1804
rect 640 1724 644 1756
rect 676 1724 680 1756
rect 640 1720 680 1724
rect 720 2476 760 2480
rect 720 2444 724 2476
rect 756 2444 760 2476
rect 720 2396 760 2444
rect 720 2364 724 2396
rect 756 2364 760 2396
rect 720 2316 760 2364
rect 720 2284 724 2316
rect 756 2284 760 2316
rect 720 2236 760 2284
rect 720 2204 724 2236
rect 756 2204 760 2236
rect 720 2156 760 2204
rect 720 2124 724 2156
rect 756 2124 760 2156
rect 720 2076 760 2124
rect 720 2044 724 2076
rect 756 2044 760 2076
rect 720 1996 760 2044
rect 720 1964 724 1996
rect 756 1964 760 1996
rect 720 1916 760 1964
rect 720 1884 724 1916
rect 756 1884 760 1916
rect 720 1836 760 1884
rect 720 1804 724 1836
rect 756 1804 760 1836
rect 720 1756 760 1804
rect 720 1724 724 1756
rect 756 1724 760 1756
rect 720 1720 760 1724
rect 800 2476 840 2480
rect 800 2444 804 2476
rect 836 2444 840 2476
rect 800 2396 840 2444
rect 800 2364 804 2396
rect 836 2364 840 2396
rect 800 2316 840 2364
rect 800 2284 804 2316
rect 836 2284 840 2316
rect 800 2236 840 2284
rect 800 2204 804 2236
rect 836 2204 840 2236
rect 800 2156 840 2204
rect 800 2124 804 2156
rect 836 2124 840 2156
rect 800 2076 840 2124
rect 800 2044 804 2076
rect 836 2044 840 2076
rect 800 1996 840 2044
rect 800 1964 804 1996
rect 836 1964 840 1996
rect 800 1916 840 1964
rect 800 1884 804 1916
rect 836 1884 840 1916
rect 800 1836 840 1884
rect 800 1804 804 1836
rect 836 1804 840 1836
rect 800 1756 840 1804
rect 800 1724 804 1756
rect 836 1724 840 1756
rect 800 1720 840 1724
rect 880 2476 920 2480
rect 880 2444 884 2476
rect 916 2444 920 2476
rect 880 2396 920 2444
rect 880 2364 884 2396
rect 916 2364 920 2396
rect 880 2316 920 2364
rect 880 2284 884 2316
rect 916 2284 920 2316
rect 880 2236 920 2284
rect 880 2204 884 2236
rect 916 2204 920 2236
rect 880 2156 920 2204
rect 880 2124 884 2156
rect 916 2124 920 2156
rect 880 2076 920 2124
rect 880 2044 884 2076
rect 916 2044 920 2076
rect 880 1996 920 2044
rect 880 1964 884 1996
rect 916 1964 920 1996
rect 880 1916 920 1964
rect 880 1884 884 1916
rect 916 1884 920 1916
rect 880 1836 920 1884
rect 880 1804 884 1836
rect 916 1804 920 1836
rect 880 1756 920 1804
rect 880 1724 884 1756
rect 916 1724 920 1756
rect 880 1720 920 1724
rect 960 2476 1000 2480
rect 960 2444 964 2476
rect 996 2444 1000 2476
rect 960 2396 1000 2444
rect 960 2364 964 2396
rect 996 2364 1000 2396
rect 960 2316 1000 2364
rect 960 2284 964 2316
rect 996 2284 1000 2316
rect 960 2236 1000 2284
rect 960 2204 964 2236
rect 996 2204 1000 2236
rect 960 2156 1000 2204
rect 960 2124 964 2156
rect 996 2124 1000 2156
rect 960 2076 1000 2124
rect 960 2044 964 2076
rect 996 2044 1000 2076
rect 960 1996 1000 2044
rect 960 1964 964 1996
rect 996 1964 1000 1996
rect 960 1916 1000 1964
rect 960 1884 964 1916
rect 996 1884 1000 1916
rect 960 1836 1000 1884
rect 960 1804 964 1836
rect 996 1804 1000 1836
rect 960 1756 1000 1804
rect 960 1724 964 1756
rect 996 1724 1000 1756
rect 960 1720 1000 1724
rect 1040 2476 1080 2480
rect 1040 2444 1044 2476
rect 1076 2444 1080 2476
rect 1040 2396 1080 2444
rect 1040 2364 1044 2396
rect 1076 2364 1080 2396
rect 1040 2316 1080 2364
rect 1040 2284 1044 2316
rect 1076 2284 1080 2316
rect 1040 2236 1080 2284
rect 1040 2204 1044 2236
rect 1076 2204 1080 2236
rect 1040 2156 1080 2204
rect 1040 2124 1044 2156
rect 1076 2124 1080 2156
rect 1040 2076 1080 2124
rect 1040 2044 1044 2076
rect 1076 2044 1080 2076
rect 1040 1996 1080 2044
rect 1040 1964 1044 1996
rect 1076 1964 1080 1996
rect 1040 1916 1080 1964
rect 1040 1884 1044 1916
rect 1076 1884 1080 1916
rect 1040 1836 1080 1884
rect 1040 1804 1044 1836
rect 1076 1804 1080 1836
rect 1040 1756 1080 1804
rect 1040 1724 1044 1756
rect 1076 1724 1080 1756
rect 1040 1720 1080 1724
rect 1120 2476 1160 2480
rect 1120 2444 1124 2476
rect 1156 2444 1160 2476
rect 1120 2396 1160 2444
rect 1120 2364 1124 2396
rect 1156 2364 1160 2396
rect 1120 2316 1160 2364
rect 1120 2284 1124 2316
rect 1156 2284 1160 2316
rect 1120 2236 1160 2284
rect 1120 2204 1124 2236
rect 1156 2204 1160 2236
rect 1120 2156 1160 2204
rect 1120 2124 1124 2156
rect 1156 2124 1160 2156
rect 1120 2076 1160 2124
rect 1120 2044 1124 2076
rect 1156 2044 1160 2076
rect 1120 1996 1160 2044
rect 1120 1964 1124 1996
rect 1156 1964 1160 1996
rect 1120 1916 1160 1964
rect 1120 1884 1124 1916
rect 1156 1884 1160 1916
rect 1120 1836 1160 1884
rect 1120 1804 1124 1836
rect 1156 1804 1160 1836
rect 1120 1756 1160 1804
rect 1120 1724 1124 1756
rect 1156 1724 1160 1756
rect 1120 1720 1160 1724
rect 1200 2476 1240 2480
rect 1200 2444 1204 2476
rect 1236 2444 1240 2476
rect 1200 2396 1240 2444
rect 1200 2364 1204 2396
rect 1236 2364 1240 2396
rect 1200 2316 1240 2364
rect 1200 2284 1204 2316
rect 1236 2284 1240 2316
rect 1200 2236 1240 2284
rect 1200 2204 1204 2236
rect 1236 2204 1240 2236
rect 1200 2156 1240 2204
rect 1200 2124 1204 2156
rect 1236 2124 1240 2156
rect 1200 2076 1240 2124
rect 1200 2044 1204 2076
rect 1236 2044 1240 2076
rect 1200 1996 1240 2044
rect 1200 1964 1204 1996
rect 1236 1964 1240 1996
rect 1200 1916 1240 1964
rect 1200 1884 1204 1916
rect 1236 1884 1240 1916
rect 1200 1836 1240 1884
rect 1200 1804 1204 1836
rect 1236 1804 1240 1836
rect 1200 1756 1240 1804
rect 1200 1724 1204 1756
rect 1236 1724 1240 1756
rect 1200 1720 1240 1724
rect 1280 2476 1320 2480
rect 1280 2444 1284 2476
rect 1316 2444 1320 2476
rect 1280 2396 1320 2444
rect 1280 2364 1284 2396
rect 1316 2364 1320 2396
rect 1280 2316 1320 2364
rect 1280 2284 1284 2316
rect 1316 2284 1320 2316
rect 1280 2236 1320 2284
rect 1280 2204 1284 2236
rect 1316 2204 1320 2236
rect 1280 2156 1320 2204
rect 1280 2124 1284 2156
rect 1316 2124 1320 2156
rect 1280 2076 1320 2124
rect 1280 2044 1284 2076
rect 1316 2044 1320 2076
rect 1280 1996 1320 2044
rect 1280 1964 1284 1996
rect 1316 1964 1320 1996
rect 1280 1916 1320 1964
rect 1280 1884 1284 1916
rect 1316 1884 1320 1916
rect 1280 1836 1320 1884
rect 1280 1804 1284 1836
rect 1316 1804 1320 1836
rect 1280 1756 1320 1804
rect 1280 1724 1284 1756
rect 1316 1724 1320 1756
rect 1280 1720 1320 1724
rect 1360 2476 1400 2480
rect 1360 2444 1364 2476
rect 1396 2444 1400 2476
rect 1360 2396 1400 2444
rect 1360 2364 1364 2396
rect 1396 2364 1400 2396
rect 1360 2316 1400 2364
rect 1360 2284 1364 2316
rect 1396 2284 1400 2316
rect 1360 2236 1400 2284
rect 1360 2204 1364 2236
rect 1396 2204 1400 2236
rect 1360 2156 1400 2204
rect 1360 2124 1364 2156
rect 1396 2124 1400 2156
rect 1360 2076 1400 2124
rect 1360 2044 1364 2076
rect 1396 2044 1400 2076
rect 1360 1996 1400 2044
rect 1360 1964 1364 1996
rect 1396 1964 1400 1996
rect 1360 1916 1400 1964
rect 1360 1884 1364 1916
rect 1396 1884 1400 1916
rect 1360 1836 1400 1884
rect 1360 1804 1364 1836
rect 1396 1804 1400 1836
rect 1360 1756 1400 1804
rect 1360 1724 1364 1756
rect 1396 1724 1400 1756
rect 1360 1720 1400 1724
rect 1440 2476 1480 2480
rect 1440 2444 1444 2476
rect 1476 2444 1480 2476
rect 1440 2396 1480 2444
rect 1440 2364 1444 2396
rect 1476 2364 1480 2396
rect 1440 2316 1480 2364
rect 1440 2284 1444 2316
rect 1476 2284 1480 2316
rect 1440 2236 1480 2284
rect 1440 2204 1444 2236
rect 1476 2204 1480 2236
rect 1440 2156 1480 2204
rect 1440 2124 1444 2156
rect 1476 2124 1480 2156
rect 1440 2076 1480 2124
rect 1440 2044 1444 2076
rect 1476 2044 1480 2076
rect 1440 1996 1480 2044
rect 1440 1964 1444 1996
rect 1476 1964 1480 1996
rect 1440 1916 1480 1964
rect 1440 1884 1444 1916
rect 1476 1884 1480 1916
rect 1440 1836 1480 1884
rect 1440 1804 1444 1836
rect 1476 1804 1480 1836
rect 1440 1756 1480 1804
rect 1440 1724 1444 1756
rect 1476 1724 1480 1756
rect 1440 1720 1480 1724
rect 1520 2476 1560 2480
rect 1520 2444 1524 2476
rect 1556 2444 1560 2476
rect 1520 2396 1560 2444
rect 1520 2364 1524 2396
rect 1556 2364 1560 2396
rect 1520 2316 1560 2364
rect 1520 2284 1524 2316
rect 1556 2284 1560 2316
rect 1520 2236 1560 2284
rect 1520 2204 1524 2236
rect 1556 2204 1560 2236
rect 1520 2156 1560 2204
rect 1520 2124 1524 2156
rect 1556 2124 1560 2156
rect 1520 2076 1560 2124
rect 1520 2044 1524 2076
rect 1556 2044 1560 2076
rect 1520 1996 1560 2044
rect 1520 1964 1524 1996
rect 1556 1964 1560 1996
rect 1520 1916 1560 1964
rect 1520 1884 1524 1916
rect 1556 1884 1560 1916
rect 1520 1836 1560 1884
rect 1520 1804 1524 1836
rect 1556 1804 1560 1836
rect 1520 1756 1560 1804
rect 1520 1724 1524 1756
rect 1556 1724 1560 1756
rect 1520 1720 1560 1724
rect 1600 2476 1640 2480
rect 1600 2444 1604 2476
rect 1636 2444 1640 2476
rect 1600 2396 1640 2444
rect 1600 2364 1604 2396
rect 1636 2364 1640 2396
rect 1600 2316 1640 2364
rect 1600 2284 1604 2316
rect 1636 2284 1640 2316
rect 1600 2236 1640 2284
rect 1600 2204 1604 2236
rect 1636 2204 1640 2236
rect 1600 2156 1640 2204
rect 1600 2124 1604 2156
rect 1636 2124 1640 2156
rect 1600 2076 1640 2124
rect 1600 2044 1604 2076
rect 1636 2044 1640 2076
rect 1600 1996 1640 2044
rect 1600 1964 1604 1996
rect 1636 1964 1640 1996
rect 1600 1916 1640 1964
rect 1600 1884 1604 1916
rect 1636 1884 1640 1916
rect 1600 1836 1640 1884
rect 1600 1804 1604 1836
rect 1636 1804 1640 1836
rect 1600 1756 1640 1804
rect 1600 1724 1604 1756
rect 1636 1724 1640 1756
rect 1600 1720 1640 1724
rect 1680 2476 1720 2480
rect 1680 2444 1684 2476
rect 1716 2444 1720 2476
rect 1680 2396 1720 2444
rect 1680 2364 1684 2396
rect 1716 2364 1720 2396
rect 1680 2316 1720 2364
rect 1680 2284 1684 2316
rect 1716 2284 1720 2316
rect 1680 2236 1720 2284
rect 1680 2204 1684 2236
rect 1716 2204 1720 2236
rect 1680 2156 1720 2204
rect 1680 2124 1684 2156
rect 1716 2124 1720 2156
rect 1680 2076 1720 2124
rect 1680 2044 1684 2076
rect 1716 2044 1720 2076
rect 1680 1996 1720 2044
rect 1680 1964 1684 1996
rect 1716 1964 1720 1996
rect 1680 1916 1720 1964
rect 1680 1884 1684 1916
rect 1716 1884 1720 1916
rect 1680 1836 1720 1884
rect 1680 1804 1684 1836
rect 1716 1804 1720 1836
rect 1680 1756 1720 1804
rect 1680 1724 1684 1756
rect 1716 1724 1720 1756
rect 1680 1720 1720 1724
rect 1760 2476 1800 2480
rect 1760 2444 1764 2476
rect 1796 2444 1800 2476
rect 1760 2396 1800 2444
rect 1760 2364 1764 2396
rect 1796 2364 1800 2396
rect 1760 2316 1800 2364
rect 1760 2284 1764 2316
rect 1796 2284 1800 2316
rect 1760 2236 1800 2284
rect 1760 2204 1764 2236
rect 1796 2204 1800 2236
rect 1760 2156 1800 2204
rect 1760 2124 1764 2156
rect 1796 2124 1800 2156
rect 1760 2076 1800 2124
rect 1760 2044 1764 2076
rect 1796 2044 1800 2076
rect 1760 1996 1800 2044
rect 1760 1964 1764 1996
rect 1796 1964 1800 1996
rect 1760 1916 1800 1964
rect 1760 1884 1764 1916
rect 1796 1884 1800 1916
rect 1760 1836 1800 1884
rect 1760 1804 1764 1836
rect 1796 1804 1800 1836
rect 1760 1756 1800 1804
rect 1760 1724 1764 1756
rect 1796 1724 1800 1756
rect 1760 1720 1800 1724
rect 1840 2476 1880 2480
rect 1840 2444 1844 2476
rect 1876 2444 1880 2476
rect 1840 2396 1880 2444
rect 1840 2364 1844 2396
rect 1876 2364 1880 2396
rect 1840 2316 1880 2364
rect 1840 2284 1844 2316
rect 1876 2284 1880 2316
rect 1840 2236 1880 2284
rect 1840 2204 1844 2236
rect 1876 2204 1880 2236
rect 1840 2156 1880 2204
rect 1840 2124 1844 2156
rect 1876 2124 1880 2156
rect 1840 2076 1880 2124
rect 1840 2044 1844 2076
rect 1876 2044 1880 2076
rect 1840 1996 1880 2044
rect 1840 1964 1844 1996
rect 1876 1964 1880 1996
rect 1840 1916 1880 1964
rect 1840 1884 1844 1916
rect 1876 1884 1880 1916
rect 1840 1836 1880 1884
rect 1840 1804 1844 1836
rect 1876 1804 1880 1836
rect 1840 1756 1880 1804
rect 1840 1724 1844 1756
rect 1876 1724 1880 1756
rect 1840 1720 1880 1724
rect 1920 2476 1960 2480
rect 1920 2444 1924 2476
rect 1956 2444 1960 2476
rect 1920 2396 1960 2444
rect 1920 2364 1924 2396
rect 1956 2364 1960 2396
rect 1920 2316 1960 2364
rect 1920 2284 1924 2316
rect 1956 2284 1960 2316
rect 1920 2236 1960 2284
rect 1920 2204 1924 2236
rect 1956 2204 1960 2236
rect 1920 2156 1960 2204
rect 1920 2124 1924 2156
rect 1956 2124 1960 2156
rect 1920 2076 1960 2124
rect 1920 2044 1924 2076
rect 1956 2044 1960 2076
rect 1920 1996 1960 2044
rect 1920 1964 1924 1996
rect 1956 1964 1960 1996
rect 1920 1916 1960 1964
rect 1920 1884 1924 1916
rect 1956 1884 1960 1916
rect 1920 1836 1960 1884
rect 1920 1804 1924 1836
rect 1956 1804 1960 1836
rect 1920 1756 1960 1804
rect 1920 1724 1924 1756
rect 1956 1724 1960 1756
rect 1920 1720 1960 1724
rect 2000 2476 2040 2480
rect 2000 2444 2004 2476
rect 2036 2444 2040 2476
rect 2000 2396 2040 2444
rect 2000 2364 2004 2396
rect 2036 2364 2040 2396
rect 2000 2316 2040 2364
rect 2000 2284 2004 2316
rect 2036 2284 2040 2316
rect 2000 2236 2040 2284
rect 2000 2204 2004 2236
rect 2036 2204 2040 2236
rect 2000 2156 2040 2204
rect 2000 2124 2004 2156
rect 2036 2124 2040 2156
rect 2000 2076 2040 2124
rect 2000 2044 2004 2076
rect 2036 2044 2040 2076
rect 2000 1996 2040 2044
rect 2000 1964 2004 1996
rect 2036 1964 2040 1996
rect 2000 1916 2040 1964
rect 2000 1884 2004 1916
rect 2036 1884 2040 1916
rect 2000 1836 2040 1884
rect 2000 1804 2004 1836
rect 2036 1804 2040 1836
rect 2000 1756 2040 1804
rect 2000 1724 2004 1756
rect 2036 1724 2040 1756
rect 2000 1720 2040 1724
rect 2080 2476 2120 2480
rect 2080 2444 2084 2476
rect 2116 2444 2120 2476
rect 2080 2396 2120 2444
rect 2080 2364 2084 2396
rect 2116 2364 2120 2396
rect 2080 2316 2120 2364
rect 2080 2284 2084 2316
rect 2116 2284 2120 2316
rect 2080 2236 2120 2284
rect 2080 2204 2084 2236
rect 2116 2204 2120 2236
rect 2080 2156 2120 2204
rect 2080 2124 2084 2156
rect 2116 2124 2120 2156
rect 2080 2076 2120 2124
rect 2080 2044 2084 2076
rect 2116 2044 2120 2076
rect 2080 1996 2120 2044
rect 2080 1964 2084 1996
rect 2116 1964 2120 1996
rect 2080 1916 2120 1964
rect 2080 1884 2084 1916
rect 2116 1884 2120 1916
rect 2080 1836 2120 1884
rect 2080 1804 2084 1836
rect 2116 1804 2120 1836
rect 2080 1756 2120 1804
rect 2080 1724 2084 1756
rect 2116 1724 2120 1756
rect 2080 1720 2120 1724
rect 2160 2476 2200 2480
rect 2160 2444 2164 2476
rect 2196 2444 2200 2476
rect 2160 2396 2200 2444
rect 2160 2364 2164 2396
rect 2196 2364 2200 2396
rect 2160 2316 2200 2364
rect 2160 2284 2164 2316
rect 2196 2284 2200 2316
rect 2160 2236 2200 2284
rect 2160 2204 2164 2236
rect 2196 2204 2200 2236
rect 2160 2156 2200 2204
rect 2160 2124 2164 2156
rect 2196 2124 2200 2156
rect 2160 2076 2200 2124
rect 2160 2044 2164 2076
rect 2196 2044 2200 2076
rect 2160 1996 2200 2044
rect 2160 1964 2164 1996
rect 2196 1964 2200 1996
rect 2160 1916 2200 1964
rect 2160 1884 2164 1916
rect 2196 1884 2200 1916
rect 2160 1836 2200 1884
rect 2160 1804 2164 1836
rect 2196 1804 2200 1836
rect 2160 1756 2200 1804
rect 2160 1724 2164 1756
rect 2196 1724 2200 1756
rect 2160 1720 2200 1724
rect 2240 2476 2280 2480
rect 2240 2444 2244 2476
rect 2276 2444 2280 2476
rect 2240 2396 2280 2444
rect 2240 2364 2244 2396
rect 2276 2364 2280 2396
rect 2240 2316 2280 2364
rect 2240 2284 2244 2316
rect 2276 2284 2280 2316
rect 2240 2236 2280 2284
rect 2240 2204 2244 2236
rect 2276 2204 2280 2236
rect 2240 2156 2280 2204
rect 2240 2124 2244 2156
rect 2276 2124 2280 2156
rect 2240 2076 2280 2124
rect 2240 2044 2244 2076
rect 2276 2044 2280 2076
rect 2240 1996 2280 2044
rect 2240 1964 2244 1996
rect 2276 1964 2280 1996
rect 2240 1916 2280 1964
rect 2240 1884 2244 1916
rect 2276 1884 2280 1916
rect 2240 1836 2280 1884
rect 2240 1804 2244 1836
rect 2276 1804 2280 1836
rect 2240 1756 2280 1804
rect 2240 1724 2244 1756
rect 2276 1724 2280 1756
rect 2240 1720 2280 1724
rect 2320 2476 2360 2480
rect 2320 2444 2324 2476
rect 2356 2444 2360 2476
rect 2320 2396 2360 2444
rect 2320 2364 2324 2396
rect 2356 2364 2360 2396
rect 2320 2316 2360 2364
rect 2320 2284 2324 2316
rect 2356 2284 2360 2316
rect 2320 2236 2360 2284
rect 2320 2204 2324 2236
rect 2356 2204 2360 2236
rect 2320 2156 2360 2204
rect 2320 2124 2324 2156
rect 2356 2124 2360 2156
rect 2320 2076 2360 2124
rect 2320 2044 2324 2076
rect 2356 2044 2360 2076
rect 2320 1996 2360 2044
rect 2320 1964 2324 1996
rect 2356 1964 2360 1996
rect 2320 1916 2360 1964
rect 2320 1884 2324 1916
rect 2356 1884 2360 1916
rect 2320 1836 2360 1884
rect 2320 1804 2324 1836
rect 2356 1804 2360 1836
rect 2320 1756 2360 1804
rect 2320 1724 2324 1756
rect 2356 1724 2360 1756
rect 2320 1720 2360 1724
rect 2400 2476 2440 2480
rect 2400 2444 2404 2476
rect 2436 2444 2440 2476
rect 2400 2396 2440 2444
rect 2400 2364 2404 2396
rect 2436 2364 2440 2396
rect 2400 2316 2440 2364
rect 2400 2284 2404 2316
rect 2436 2284 2440 2316
rect 2400 2236 2440 2284
rect 2400 2204 2404 2236
rect 2436 2204 2440 2236
rect 2400 2156 2440 2204
rect 2400 2124 2404 2156
rect 2436 2124 2440 2156
rect 2400 2076 2440 2124
rect 2400 2044 2404 2076
rect 2436 2044 2440 2076
rect 2400 1996 2440 2044
rect 2400 1964 2404 1996
rect 2436 1964 2440 1996
rect 2400 1916 2440 1964
rect 2400 1884 2404 1916
rect 2436 1884 2440 1916
rect 2400 1836 2440 1884
rect 2400 1804 2404 1836
rect 2436 1804 2440 1836
rect 2400 1756 2440 1804
rect 2400 1724 2404 1756
rect 2436 1724 2440 1756
rect 2400 1720 2440 1724
rect 2480 2476 2520 2480
rect 2480 2444 2484 2476
rect 2516 2444 2520 2476
rect 2480 2396 2520 2444
rect 2480 2364 2484 2396
rect 2516 2364 2520 2396
rect 2480 2316 2520 2364
rect 2480 2284 2484 2316
rect 2516 2284 2520 2316
rect 2480 2236 2520 2284
rect 2480 2204 2484 2236
rect 2516 2204 2520 2236
rect 2480 2156 2520 2204
rect 2480 2124 2484 2156
rect 2516 2124 2520 2156
rect 2480 2076 2520 2124
rect 2480 2044 2484 2076
rect 2516 2044 2520 2076
rect 2480 1996 2520 2044
rect 2480 1964 2484 1996
rect 2516 1964 2520 1996
rect 2480 1916 2520 1964
rect 2480 1884 2484 1916
rect 2516 1884 2520 1916
rect 2480 1836 2520 1884
rect 2480 1804 2484 1836
rect 2516 1804 2520 1836
rect 2480 1756 2520 1804
rect 2480 1724 2484 1756
rect 2516 1724 2520 1756
rect 2480 1720 2520 1724
rect 2560 2476 2600 2480
rect 2560 2444 2564 2476
rect 2596 2444 2600 2476
rect 2560 2396 2600 2444
rect 2560 2364 2564 2396
rect 2596 2364 2600 2396
rect 2560 2316 2600 2364
rect 2560 2284 2564 2316
rect 2596 2284 2600 2316
rect 2560 2236 2600 2284
rect 2560 2204 2564 2236
rect 2596 2204 2600 2236
rect 2560 2156 2600 2204
rect 2560 2124 2564 2156
rect 2596 2124 2600 2156
rect 2560 2076 2600 2124
rect 2560 2044 2564 2076
rect 2596 2044 2600 2076
rect 2560 1996 2600 2044
rect 2560 1964 2564 1996
rect 2596 1964 2600 1996
rect 2560 1916 2600 1964
rect 2560 1884 2564 1916
rect 2596 1884 2600 1916
rect 2560 1836 2600 1884
rect 2560 1804 2564 1836
rect 2596 1804 2600 1836
rect 2560 1756 2600 1804
rect 2560 1724 2564 1756
rect 2596 1724 2600 1756
rect 2560 1720 2600 1724
rect 2640 2476 2680 2480
rect 2640 2444 2644 2476
rect 2676 2444 2680 2476
rect 2640 2396 2680 2444
rect 2640 2364 2644 2396
rect 2676 2364 2680 2396
rect 2640 2316 2680 2364
rect 2640 2284 2644 2316
rect 2676 2284 2680 2316
rect 2640 2236 2680 2284
rect 2640 2204 2644 2236
rect 2676 2204 2680 2236
rect 2640 2156 2680 2204
rect 2640 2124 2644 2156
rect 2676 2124 2680 2156
rect 2640 2076 2680 2124
rect 2640 2044 2644 2076
rect 2676 2044 2680 2076
rect 2640 1996 2680 2044
rect 2640 1964 2644 1996
rect 2676 1964 2680 1996
rect 2640 1916 2680 1964
rect 2640 1884 2644 1916
rect 2676 1884 2680 1916
rect 2640 1836 2680 1884
rect 2640 1804 2644 1836
rect 2676 1804 2680 1836
rect 2640 1756 2680 1804
rect 2640 1724 2644 1756
rect 2676 1724 2680 1756
rect 2640 1720 2680 1724
rect 2720 2476 2760 2480
rect 2720 2444 2724 2476
rect 2756 2444 2760 2476
rect 2720 2396 2760 2444
rect 2720 2364 2724 2396
rect 2756 2364 2760 2396
rect 2720 2316 2760 2364
rect 2720 2284 2724 2316
rect 2756 2284 2760 2316
rect 2720 2236 2760 2284
rect 2720 2204 2724 2236
rect 2756 2204 2760 2236
rect 2720 2156 2760 2204
rect 2720 2124 2724 2156
rect 2756 2124 2760 2156
rect 2720 2076 2760 2124
rect 2720 2044 2724 2076
rect 2756 2044 2760 2076
rect 2720 1996 2760 2044
rect 2720 1964 2724 1996
rect 2756 1964 2760 1996
rect 2720 1916 2760 1964
rect 2720 1884 2724 1916
rect 2756 1884 2760 1916
rect 2720 1836 2760 1884
rect 2720 1804 2724 1836
rect 2756 1804 2760 1836
rect 2720 1756 2760 1804
rect 2720 1724 2724 1756
rect 2756 1724 2760 1756
rect 2720 1720 2760 1724
rect 2800 2476 2840 2480
rect 2800 2444 2804 2476
rect 2836 2444 2840 2476
rect 2800 2396 2840 2444
rect 2800 2364 2804 2396
rect 2836 2364 2840 2396
rect 2800 2316 2840 2364
rect 2800 2284 2804 2316
rect 2836 2284 2840 2316
rect 2800 2236 2840 2284
rect 2800 2204 2804 2236
rect 2836 2204 2840 2236
rect 2800 2156 2840 2204
rect 2800 2124 2804 2156
rect 2836 2124 2840 2156
rect 2800 2076 2840 2124
rect 2800 2044 2804 2076
rect 2836 2044 2840 2076
rect 2800 1996 2840 2044
rect 2800 1964 2804 1996
rect 2836 1964 2840 1996
rect 2800 1916 2840 1964
rect 2800 1884 2804 1916
rect 2836 1884 2840 1916
rect 2800 1836 2840 1884
rect 2800 1804 2804 1836
rect 2836 1804 2840 1836
rect 2800 1756 2840 1804
rect 2800 1724 2804 1756
rect 2836 1724 2840 1756
rect 2800 1720 2840 1724
rect 2880 2476 2920 2480
rect 2880 2444 2884 2476
rect 2916 2444 2920 2476
rect 2880 2396 2920 2444
rect 2880 2364 2884 2396
rect 2916 2364 2920 2396
rect 2880 2316 2920 2364
rect 2880 2284 2884 2316
rect 2916 2284 2920 2316
rect 2880 2236 2920 2284
rect 2880 2204 2884 2236
rect 2916 2204 2920 2236
rect 2880 2156 2920 2204
rect 2880 2124 2884 2156
rect 2916 2124 2920 2156
rect 2880 2076 2920 2124
rect 2880 2044 2884 2076
rect 2916 2044 2920 2076
rect 2880 1996 2920 2044
rect 2880 1964 2884 1996
rect 2916 1964 2920 1996
rect 2880 1916 2920 1964
rect 2880 1884 2884 1916
rect 2916 1884 2920 1916
rect 2880 1836 2920 1884
rect 2880 1804 2884 1836
rect 2916 1804 2920 1836
rect 2880 1756 2920 1804
rect 2880 1724 2884 1756
rect 2916 1724 2920 1756
rect 2880 1720 2920 1724
rect 2960 2476 3000 2480
rect 2960 2444 2964 2476
rect 2996 2444 3000 2476
rect 2960 2396 3000 2444
rect 2960 2364 2964 2396
rect 2996 2364 3000 2396
rect 2960 2316 3000 2364
rect 2960 2284 2964 2316
rect 2996 2284 3000 2316
rect 2960 2236 3000 2284
rect 2960 2204 2964 2236
rect 2996 2204 3000 2236
rect 2960 2156 3000 2204
rect 2960 2124 2964 2156
rect 2996 2124 3000 2156
rect 2960 2076 3000 2124
rect 2960 2044 2964 2076
rect 2996 2044 3000 2076
rect 2960 1996 3000 2044
rect 2960 1964 2964 1996
rect 2996 1964 3000 1996
rect 2960 1916 3000 1964
rect 2960 1884 2964 1916
rect 2996 1884 3000 1916
rect 2960 1836 3000 1884
rect 2960 1804 2964 1836
rect 2996 1804 3000 1836
rect 2960 1756 3000 1804
rect 2960 1724 2964 1756
rect 2996 1724 3000 1756
rect 2960 1720 3000 1724
rect 3040 2476 3080 2480
rect 3040 2444 3044 2476
rect 3076 2444 3080 2476
rect 3040 2396 3080 2444
rect 3040 2364 3044 2396
rect 3076 2364 3080 2396
rect 3040 2316 3080 2364
rect 3040 2284 3044 2316
rect 3076 2284 3080 2316
rect 3040 2236 3080 2284
rect 3040 2204 3044 2236
rect 3076 2204 3080 2236
rect 3040 2156 3080 2204
rect 3040 2124 3044 2156
rect 3076 2124 3080 2156
rect 3040 2076 3080 2124
rect 3040 2044 3044 2076
rect 3076 2044 3080 2076
rect 3040 1996 3080 2044
rect 3040 1964 3044 1996
rect 3076 1964 3080 1996
rect 3040 1916 3080 1964
rect 3040 1884 3044 1916
rect 3076 1884 3080 1916
rect 3040 1836 3080 1884
rect 3040 1804 3044 1836
rect 3076 1804 3080 1836
rect 3040 1756 3080 1804
rect 3040 1724 3044 1756
rect 3076 1724 3080 1756
rect 3040 1720 3080 1724
rect 3120 2476 3160 2480
rect 3120 2444 3124 2476
rect 3156 2444 3160 2476
rect 3120 2396 3160 2444
rect 3120 2364 3124 2396
rect 3156 2364 3160 2396
rect 3120 2316 3160 2364
rect 3120 2284 3124 2316
rect 3156 2284 3160 2316
rect 3120 2236 3160 2284
rect 3120 2204 3124 2236
rect 3156 2204 3160 2236
rect 3120 2156 3160 2204
rect 3120 2124 3124 2156
rect 3156 2124 3160 2156
rect 3120 2076 3160 2124
rect 3120 2044 3124 2076
rect 3156 2044 3160 2076
rect 3120 1996 3160 2044
rect 3120 1964 3124 1996
rect 3156 1964 3160 1996
rect 3120 1916 3160 1964
rect 3120 1884 3124 1916
rect 3156 1884 3160 1916
rect 3120 1836 3160 1884
rect 3120 1804 3124 1836
rect 3156 1804 3160 1836
rect 3120 1756 3160 1804
rect 3120 1724 3124 1756
rect 3156 1724 3160 1756
rect 3120 1720 3160 1724
rect 3200 2476 3240 2480
rect 3200 2444 3204 2476
rect 3236 2444 3240 2476
rect 3200 2396 3240 2444
rect 3200 2364 3204 2396
rect 3236 2364 3240 2396
rect 3200 2316 3240 2364
rect 3200 2284 3204 2316
rect 3236 2284 3240 2316
rect 3200 2236 3240 2284
rect 3200 2204 3204 2236
rect 3236 2204 3240 2236
rect 3200 2156 3240 2204
rect 3200 2124 3204 2156
rect 3236 2124 3240 2156
rect 3200 2076 3240 2124
rect 3200 2044 3204 2076
rect 3236 2044 3240 2076
rect 3200 1996 3240 2044
rect 3200 1964 3204 1996
rect 3236 1964 3240 1996
rect 3200 1916 3240 1964
rect 3200 1884 3204 1916
rect 3236 1884 3240 1916
rect 3200 1836 3240 1884
rect 3200 1804 3204 1836
rect 3236 1804 3240 1836
rect 3200 1756 3240 1804
rect 3200 1724 3204 1756
rect 3236 1724 3240 1756
rect 3200 1720 3240 1724
rect 3280 2476 3320 2480
rect 3280 2444 3284 2476
rect 3316 2444 3320 2476
rect 3280 2396 3320 2444
rect 3280 2364 3284 2396
rect 3316 2364 3320 2396
rect 3280 2316 3320 2364
rect 3280 2284 3284 2316
rect 3316 2284 3320 2316
rect 3280 2236 3320 2284
rect 3280 2204 3284 2236
rect 3316 2204 3320 2236
rect 3280 2156 3320 2204
rect 3280 2124 3284 2156
rect 3316 2124 3320 2156
rect 3280 2076 3320 2124
rect 3280 2044 3284 2076
rect 3316 2044 3320 2076
rect 3280 1996 3320 2044
rect 3280 1964 3284 1996
rect 3316 1964 3320 1996
rect 3280 1916 3320 1964
rect 3280 1884 3284 1916
rect 3316 1884 3320 1916
rect 3280 1836 3320 1884
rect 3280 1804 3284 1836
rect 3316 1804 3320 1836
rect 3280 1756 3320 1804
rect 3280 1724 3284 1756
rect 3316 1724 3320 1756
rect 3280 1720 3320 1724
rect 3360 2476 3400 2480
rect 3360 2444 3364 2476
rect 3396 2444 3400 2476
rect 3360 2396 3400 2444
rect 3360 2364 3364 2396
rect 3396 2364 3400 2396
rect 3360 2316 3400 2364
rect 3360 2284 3364 2316
rect 3396 2284 3400 2316
rect 3360 2236 3400 2284
rect 3360 2204 3364 2236
rect 3396 2204 3400 2236
rect 3360 2156 3400 2204
rect 3360 2124 3364 2156
rect 3396 2124 3400 2156
rect 3360 2076 3400 2124
rect 3360 2044 3364 2076
rect 3396 2044 3400 2076
rect 3360 1996 3400 2044
rect 3360 1964 3364 1996
rect 3396 1964 3400 1996
rect 3360 1916 3400 1964
rect 3360 1884 3364 1916
rect 3396 1884 3400 1916
rect 3360 1836 3400 1884
rect 3360 1804 3364 1836
rect 3396 1804 3400 1836
rect 3360 1756 3400 1804
rect 3360 1724 3364 1756
rect 3396 1724 3400 1756
rect 3360 1720 3400 1724
rect 3440 2476 3480 2480
rect 3440 2444 3444 2476
rect 3476 2444 3480 2476
rect 3440 2396 3480 2444
rect 3440 2364 3444 2396
rect 3476 2364 3480 2396
rect 3440 2316 3480 2364
rect 3440 2284 3444 2316
rect 3476 2284 3480 2316
rect 3440 2236 3480 2284
rect 3440 2204 3444 2236
rect 3476 2204 3480 2236
rect 3440 2156 3480 2204
rect 3440 2124 3444 2156
rect 3476 2124 3480 2156
rect 3440 2076 3480 2124
rect 3440 2044 3444 2076
rect 3476 2044 3480 2076
rect 3440 1996 3480 2044
rect 3440 1964 3444 1996
rect 3476 1964 3480 1996
rect 3440 1916 3480 1964
rect 3440 1884 3444 1916
rect 3476 1884 3480 1916
rect 3440 1836 3480 1884
rect 3440 1804 3444 1836
rect 3476 1804 3480 1836
rect 3440 1756 3480 1804
rect 3440 1724 3444 1756
rect 3476 1724 3480 1756
rect 3440 1720 3480 1724
rect 3520 2476 3560 2480
rect 3520 2444 3524 2476
rect 3556 2444 3560 2476
rect 3520 2396 3560 2444
rect 3520 2364 3524 2396
rect 3556 2364 3560 2396
rect 3520 2316 3560 2364
rect 3520 2284 3524 2316
rect 3556 2284 3560 2316
rect 3520 2236 3560 2284
rect 3520 2204 3524 2236
rect 3556 2204 3560 2236
rect 3520 2156 3560 2204
rect 3520 2124 3524 2156
rect 3556 2124 3560 2156
rect 3520 2076 3560 2124
rect 3520 2044 3524 2076
rect 3556 2044 3560 2076
rect 3520 1996 3560 2044
rect 3520 1964 3524 1996
rect 3556 1964 3560 1996
rect 3520 1916 3560 1964
rect 3520 1884 3524 1916
rect 3556 1884 3560 1916
rect 3520 1836 3560 1884
rect 3520 1804 3524 1836
rect 3556 1804 3560 1836
rect 3520 1756 3560 1804
rect 3520 1724 3524 1756
rect 3556 1724 3560 1756
rect 3520 1720 3560 1724
rect 3600 2476 3640 2480
rect 3600 2444 3604 2476
rect 3636 2444 3640 2476
rect 3600 2396 3640 2444
rect 3600 2364 3604 2396
rect 3636 2364 3640 2396
rect 3600 2316 3640 2364
rect 3600 2284 3604 2316
rect 3636 2284 3640 2316
rect 3600 2236 3640 2284
rect 3600 2204 3604 2236
rect 3636 2204 3640 2236
rect 3600 2156 3640 2204
rect 3600 2124 3604 2156
rect 3636 2124 3640 2156
rect 3600 2076 3640 2124
rect 3600 2044 3604 2076
rect 3636 2044 3640 2076
rect 3600 1996 3640 2044
rect 3600 1964 3604 1996
rect 3636 1964 3640 1996
rect 3600 1916 3640 1964
rect 3600 1884 3604 1916
rect 3636 1884 3640 1916
rect 3600 1836 3640 1884
rect 3600 1804 3604 1836
rect 3636 1804 3640 1836
rect 3600 1756 3640 1804
rect 3600 1724 3604 1756
rect 3636 1724 3640 1756
rect 3600 1720 3640 1724
rect 3680 2476 3720 2480
rect 3680 2444 3684 2476
rect 3716 2444 3720 2476
rect 3680 2396 3720 2444
rect 3680 2364 3684 2396
rect 3716 2364 3720 2396
rect 3680 2316 3720 2364
rect 3680 2284 3684 2316
rect 3716 2284 3720 2316
rect 3680 2236 3720 2284
rect 3680 2204 3684 2236
rect 3716 2204 3720 2236
rect 3680 2156 3720 2204
rect 3680 2124 3684 2156
rect 3716 2124 3720 2156
rect 3680 2076 3720 2124
rect 3680 2044 3684 2076
rect 3716 2044 3720 2076
rect 3680 1996 3720 2044
rect 3680 1964 3684 1996
rect 3716 1964 3720 1996
rect 3680 1916 3720 1964
rect 3680 1884 3684 1916
rect 3716 1884 3720 1916
rect 3680 1836 3720 1884
rect 3680 1804 3684 1836
rect 3716 1804 3720 1836
rect 3680 1756 3720 1804
rect 3680 1724 3684 1756
rect 3716 1724 3720 1756
rect 3680 1720 3720 1724
rect 3760 2476 3800 2480
rect 3760 2444 3764 2476
rect 3796 2444 3800 2476
rect 3760 2396 3800 2444
rect 3760 2364 3764 2396
rect 3796 2364 3800 2396
rect 3760 2316 3800 2364
rect 3760 2284 3764 2316
rect 3796 2284 3800 2316
rect 3760 2236 3800 2284
rect 3760 2204 3764 2236
rect 3796 2204 3800 2236
rect 3760 2156 3800 2204
rect 3760 2124 3764 2156
rect 3796 2124 3800 2156
rect 3760 2076 3800 2124
rect 3760 2044 3764 2076
rect 3796 2044 3800 2076
rect 3760 1996 3800 2044
rect 3760 1964 3764 1996
rect 3796 1964 3800 1996
rect 3760 1916 3800 1964
rect 3760 1884 3764 1916
rect 3796 1884 3800 1916
rect 3760 1836 3800 1884
rect 3760 1804 3764 1836
rect 3796 1804 3800 1836
rect 3760 1756 3800 1804
rect 3760 1724 3764 1756
rect 3796 1724 3800 1756
rect 3760 1720 3800 1724
rect 3840 2476 3880 2480
rect 3840 2444 3844 2476
rect 3876 2444 3880 2476
rect 3840 2396 3880 2444
rect 3840 2364 3844 2396
rect 3876 2364 3880 2396
rect 3840 2316 3880 2364
rect 3840 2284 3844 2316
rect 3876 2284 3880 2316
rect 3840 2236 3880 2284
rect 3840 2204 3844 2236
rect 3876 2204 3880 2236
rect 3840 2156 3880 2204
rect 3840 2124 3844 2156
rect 3876 2124 3880 2156
rect 3840 2076 3880 2124
rect 3840 2044 3844 2076
rect 3876 2044 3880 2076
rect 3840 1996 3880 2044
rect 3840 1964 3844 1996
rect 3876 1964 3880 1996
rect 3840 1916 3880 1964
rect 3840 1884 3844 1916
rect 3876 1884 3880 1916
rect 3840 1836 3880 1884
rect 3840 1804 3844 1836
rect 3876 1804 3880 1836
rect 3840 1756 3880 1804
rect 3840 1724 3844 1756
rect 3876 1724 3880 1756
rect 3840 1720 3880 1724
rect 3920 2476 3960 2480
rect 3920 2444 3924 2476
rect 3956 2444 3960 2476
rect 3920 2396 3960 2444
rect 3920 2364 3924 2396
rect 3956 2364 3960 2396
rect 3920 2316 3960 2364
rect 3920 2284 3924 2316
rect 3956 2284 3960 2316
rect 3920 2236 3960 2284
rect 3920 2204 3924 2236
rect 3956 2204 3960 2236
rect 3920 2156 3960 2204
rect 3920 2124 3924 2156
rect 3956 2124 3960 2156
rect 3920 2076 3960 2124
rect 3920 2044 3924 2076
rect 3956 2044 3960 2076
rect 3920 1996 3960 2044
rect 3920 1964 3924 1996
rect 3956 1964 3960 1996
rect 3920 1916 3960 1964
rect 3920 1884 3924 1916
rect 3956 1884 3960 1916
rect 3920 1836 3960 1884
rect 3920 1804 3924 1836
rect 3956 1804 3960 1836
rect 3920 1756 3960 1804
rect 3920 1724 3924 1756
rect 3956 1724 3960 1756
rect 3920 1720 3960 1724
rect 4000 2476 4040 2480
rect 4000 2444 4004 2476
rect 4036 2444 4040 2476
rect 4000 2396 4040 2444
rect 4000 2364 4004 2396
rect 4036 2364 4040 2396
rect 4000 2316 4040 2364
rect 4000 2284 4004 2316
rect 4036 2284 4040 2316
rect 4000 2236 4040 2284
rect 4000 2204 4004 2236
rect 4036 2204 4040 2236
rect 4000 2156 4040 2204
rect 4000 2124 4004 2156
rect 4036 2124 4040 2156
rect 4000 2076 4040 2124
rect 4000 2044 4004 2076
rect 4036 2044 4040 2076
rect 4000 1996 4040 2044
rect 4000 1964 4004 1996
rect 4036 1964 4040 1996
rect 4000 1916 4040 1964
rect 4000 1884 4004 1916
rect 4036 1884 4040 1916
rect 4000 1836 4040 1884
rect 4000 1804 4004 1836
rect 4036 1804 4040 1836
rect 4000 1756 4040 1804
rect 4000 1724 4004 1756
rect 4036 1724 4040 1756
rect 4000 1720 4040 1724
rect 4080 2476 4120 2480
rect 4080 2444 4084 2476
rect 4116 2444 4120 2476
rect 4080 2396 4120 2444
rect 4080 2364 4084 2396
rect 4116 2364 4120 2396
rect 4080 2316 4120 2364
rect 4080 2284 4084 2316
rect 4116 2284 4120 2316
rect 4080 2236 4120 2284
rect 4080 2204 4084 2236
rect 4116 2204 4120 2236
rect 4080 2156 4120 2204
rect 4080 2124 4084 2156
rect 4116 2124 4120 2156
rect 4080 2076 4120 2124
rect 4080 2044 4084 2076
rect 4116 2044 4120 2076
rect 4080 1996 4120 2044
rect 4080 1964 4084 1996
rect 4116 1964 4120 1996
rect 4080 1916 4120 1964
rect 4080 1884 4084 1916
rect 4116 1884 4120 1916
rect 4080 1836 4120 1884
rect 4080 1804 4084 1836
rect 4116 1804 4120 1836
rect 4080 1756 4120 1804
rect 4080 1724 4084 1756
rect 4116 1724 4120 1756
rect 4080 1720 4120 1724
rect 4160 2476 4200 2480
rect 4160 2444 4164 2476
rect 4196 2444 4200 2476
rect 4160 2396 4200 2444
rect 4160 2364 4164 2396
rect 4196 2364 4200 2396
rect 4160 2316 4200 2364
rect 4160 2284 4164 2316
rect 4196 2284 4200 2316
rect 4160 2236 4200 2284
rect 4160 2204 4164 2236
rect 4196 2204 4200 2236
rect 4160 2156 4200 2204
rect 4160 2124 4164 2156
rect 4196 2124 4200 2156
rect 4160 2076 4200 2124
rect 4160 2044 4164 2076
rect 4196 2044 4200 2076
rect 4160 1996 4200 2044
rect 4160 1964 4164 1996
rect 4196 1964 4200 1996
rect 4160 1916 4200 1964
rect 4160 1884 4164 1916
rect 4196 1884 4200 1916
rect 4160 1836 4200 1884
rect 4160 1804 4164 1836
rect 4196 1804 4200 1836
rect 4160 1756 4200 1804
rect 4160 1724 4164 1756
rect 4196 1724 4200 1756
rect 4160 1720 4200 1724
rect 4240 2476 4280 2480
rect 4240 2444 4244 2476
rect 4276 2444 4280 2476
rect 4240 2396 4280 2444
rect 4240 2364 4244 2396
rect 4276 2364 4280 2396
rect 4240 2316 4280 2364
rect 4240 2284 4244 2316
rect 4276 2284 4280 2316
rect 4240 2236 4280 2284
rect 4240 2204 4244 2236
rect 4276 2204 4280 2236
rect 4240 2156 4280 2204
rect 4240 2124 4244 2156
rect 4276 2124 4280 2156
rect 4240 2076 4280 2124
rect 4240 2044 4244 2076
rect 4276 2044 4280 2076
rect 4240 1996 4280 2044
rect 4240 1964 4244 1996
rect 4276 1964 4280 1996
rect 4240 1916 4280 1964
rect 4240 1884 4244 1916
rect 4276 1884 4280 1916
rect 4240 1836 4280 1884
rect 4240 1804 4244 1836
rect 4276 1804 4280 1836
rect 4240 1756 4280 1804
rect 4240 1724 4244 1756
rect 4276 1724 4280 1756
rect 4240 1720 4280 1724
rect 4320 2476 4360 2480
rect 4320 2444 4324 2476
rect 4356 2444 4360 2476
rect 4320 2396 4360 2444
rect 4320 2364 4324 2396
rect 4356 2364 4360 2396
rect 4320 2316 4360 2364
rect 4320 2284 4324 2316
rect 4356 2284 4360 2316
rect 4320 2236 4360 2284
rect 4320 2204 4324 2236
rect 4356 2204 4360 2236
rect 4320 2156 4360 2204
rect 4320 2124 4324 2156
rect 4356 2124 4360 2156
rect 4320 2076 4360 2124
rect 4320 2044 4324 2076
rect 4356 2044 4360 2076
rect 4320 1996 4360 2044
rect 4320 1964 4324 1996
rect 4356 1964 4360 1996
rect 4320 1916 4360 1964
rect 4320 1884 4324 1916
rect 4356 1884 4360 1916
rect 4320 1836 4360 1884
rect 4320 1804 4324 1836
rect 4356 1804 4360 1836
rect 4320 1756 4360 1804
rect 4320 1724 4324 1756
rect 4356 1724 4360 1756
rect 4320 1720 4360 1724
rect 4400 2476 4440 2480
rect 4400 2444 4404 2476
rect 4436 2444 4440 2476
rect 4400 2396 4440 2444
rect 4400 2364 4404 2396
rect 4436 2364 4440 2396
rect 4400 2316 4440 2364
rect 4400 2284 4404 2316
rect 4436 2284 4440 2316
rect 4400 2236 4440 2284
rect 4400 2204 4404 2236
rect 4436 2204 4440 2236
rect 4400 2156 4440 2204
rect 4400 2124 4404 2156
rect 4436 2124 4440 2156
rect 4400 2076 4440 2124
rect 4400 2044 4404 2076
rect 4436 2044 4440 2076
rect 4400 1996 4440 2044
rect 4400 1964 4404 1996
rect 4436 1964 4440 1996
rect 4400 1916 4440 1964
rect 4400 1884 4404 1916
rect 4436 1884 4440 1916
rect 4400 1836 4440 1884
rect 4400 1804 4404 1836
rect 4436 1804 4440 1836
rect 4400 1756 4440 1804
rect 4400 1724 4404 1756
rect 4436 1724 4440 1756
rect 4400 1720 4440 1724
rect 4480 2476 4520 2480
rect 4480 2444 4484 2476
rect 4516 2444 4520 2476
rect 4480 2396 4520 2444
rect 4480 2364 4484 2396
rect 4516 2364 4520 2396
rect 4480 2316 4520 2364
rect 4480 2284 4484 2316
rect 4516 2284 4520 2316
rect 4480 2236 4520 2284
rect 4480 2204 4484 2236
rect 4516 2204 4520 2236
rect 4480 2156 4520 2204
rect 4480 2124 4484 2156
rect 4516 2124 4520 2156
rect 4480 2076 4520 2124
rect 4480 2044 4484 2076
rect 4516 2044 4520 2076
rect 4480 1996 4520 2044
rect 4480 1964 4484 1996
rect 4516 1964 4520 1996
rect 4480 1916 4520 1964
rect 4480 1884 4484 1916
rect 4516 1884 4520 1916
rect 4480 1836 4520 1884
rect 4480 1804 4484 1836
rect 4516 1804 4520 1836
rect 4480 1756 4520 1804
rect 4480 1724 4484 1756
rect 4516 1724 4520 1756
rect 4480 1720 4520 1724
rect 4560 2476 4600 2480
rect 4560 2444 4564 2476
rect 4596 2444 4600 2476
rect 4560 2396 4600 2444
rect 4560 2364 4564 2396
rect 4596 2364 4600 2396
rect 4560 2316 4600 2364
rect 4560 2284 4564 2316
rect 4596 2284 4600 2316
rect 4560 2236 4600 2284
rect 4560 2204 4564 2236
rect 4596 2204 4600 2236
rect 4560 2156 4600 2204
rect 4560 2124 4564 2156
rect 4596 2124 4600 2156
rect 4560 2076 4600 2124
rect 4560 2044 4564 2076
rect 4596 2044 4600 2076
rect 4560 1996 4600 2044
rect 4560 1964 4564 1996
rect 4596 1964 4600 1996
rect 4560 1916 4600 1964
rect 4560 1884 4564 1916
rect 4596 1884 4600 1916
rect 4560 1836 4600 1884
rect 4560 1804 4564 1836
rect 4596 1804 4600 1836
rect 4560 1756 4600 1804
rect 4560 1724 4564 1756
rect 4596 1724 4600 1756
rect 4560 1720 4600 1724
rect 4640 2476 4680 2480
rect 4640 2444 4644 2476
rect 4676 2444 4680 2476
rect 4640 2396 4680 2444
rect 4640 2364 4644 2396
rect 4676 2364 4680 2396
rect 4640 2316 4680 2364
rect 4640 2284 4644 2316
rect 4676 2284 4680 2316
rect 4640 2236 4680 2284
rect 4640 2204 4644 2236
rect 4676 2204 4680 2236
rect 4640 2156 4680 2204
rect 4640 2124 4644 2156
rect 4676 2124 4680 2156
rect 4640 2076 4680 2124
rect 4640 2044 4644 2076
rect 4676 2044 4680 2076
rect 4640 1996 4680 2044
rect 4640 1964 4644 1996
rect 4676 1964 4680 1996
rect 4640 1916 4680 1964
rect 4640 1884 4644 1916
rect 4676 1884 4680 1916
rect 4640 1836 4680 1884
rect 4640 1804 4644 1836
rect 4676 1804 4680 1836
rect 4640 1756 4680 1804
rect 4640 1724 4644 1756
rect 4676 1724 4680 1756
rect 4640 1720 4680 1724
rect 4720 2476 4760 2480
rect 4720 2444 4724 2476
rect 4756 2444 4760 2476
rect 4720 2396 4760 2444
rect 4720 2364 4724 2396
rect 4756 2364 4760 2396
rect 4720 2316 4760 2364
rect 4720 2284 4724 2316
rect 4756 2284 4760 2316
rect 4720 2236 4760 2284
rect 4720 2204 4724 2236
rect 4756 2204 4760 2236
rect 4720 2156 4760 2204
rect 4720 2124 4724 2156
rect 4756 2124 4760 2156
rect 4720 2076 4760 2124
rect 4720 2044 4724 2076
rect 4756 2044 4760 2076
rect 4720 1996 4760 2044
rect 4720 1964 4724 1996
rect 4756 1964 4760 1996
rect 4720 1916 4760 1964
rect 4720 1884 4724 1916
rect 4756 1884 4760 1916
rect 4720 1836 4760 1884
rect 4720 1804 4724 1836
rect 4756 1804 4760 1836
rect 4720 1756 4760 1804
rect 4720 1724 4724 1756
rect 4756 1724 4760 1756
rect 4720 1720 4760 1724
rect 4800 2476 4840 2480
rect 4800 2444 4804 2476
rect 4836 2444 4840 2476
rect 4800 2396 4840 2444
rect 4800 2364 4804 2396
rect 4836 2364 4840 2396
rect 4800 2316 4840 2364
rect 4800 2284 4804 2316
rect 4836 2284 4840 2316
rect 4800 2236 4840 2284
rect 4800 2204 4804 2236
rect 4836 2204 4840 2236
rect 4800 2156 4840 2204
rect 4800 2124 4804 2156
rect 4836 2124 4840 2156
rect 4800 2076 4840 2124
rect 4800 2044 4804 2076
rect 4836 2044 4840 2076
rect 4800 1996 4840 2044
rect 4800 1964 4804 1996
rect 4836 1964 4840 1996
rect 4800 1916 4840 1964
rect 4800 1884 4804 1916
rect 4836 1884 4840 1916
rect 4800 1836 4840 1884
rect 4800 1804 4804 1836
rect 4836 1804 4840 1836
rect 4800 1756 4840 1804
rect 4800 1724 4804 1756
rect 4836 1724 4840 1756
rect 4800 1720 4840 1724
rect 4880 2476 4920 2524
rect 4880 2444 4884 2476
rect 4916 2444 4920 2476
rect 4880 2396 4920 2444
rect 4880 2364 4884 2396
rect 4916 2364 4920 2396
rect 4880 2316 4920 2364
rect 4880 2284 4884 2316
rect 4916 2284 4920 2316
rect 4880 2236 4920 2284
rect 4880 2204 4884 2236
rect 4916 2204 4920 2236
rect 4880 2156 4920 2204
rect 4880 2124 4884 2156
rect 4916 2124 4920 2156
rect 4880 2076 4920 2124
rect 4880 2044 4884 2076
rect 4916 2044 4920 2076
rect 4880 1996 4920 2044
rect 4880 1964 4884 1996
rect 4916 1964 4920 1996
rect 4880 1916 4920 1964
rect 4880 1884 4884 1916
rect 4916 1884 4920 1916
rect 4880 1836 4920 1884
rect 4880 1804 4884 1836
rect 4916 1804 4920 1836
rect 4880 1756 4920 1804
rect 4880 1724 4884 1756
rect 4916 1724 4920 1756
rect -880 1644 -876 1676
rect -844 1644 -840 1676
rect -880 1596 -840 1644
rect -880 1564 -876 1596
rect -844 1564 -840 1596
rect -880 1516 -840 1564
rect -880 1484 -876 1516
rect -844 1484 -840 1516
rect -880 1436 -840 1484
rect -880 1404 -876 1436
rect -844 1404 -840 1436
rect -880 1356 -840 1404
rect -880 1324 -876 1356
rect -844 1324 -840 1356
rect -880 1276 -840 1324
rect -880 1244 -876 1276
rect -844 1244 -840 1276
rect -880 1196 -840 1244
rect -880 1164 -876 1196
rect -844 1164 -840 1196
rect -880 1116 -840 1164
rect -880 1084 -876 1116
rect -844 1084 -840 1116
rect -880 1036 -840 1084
rect -880 1004 -876 1036
rect -844 1004 -840 1036
rect -880 956 -840 1004
rect -880 924 -876 956
rect -844 924 -840 956
rect -880 876 -840 924
rect -800 1676 -760 1680
rect -800 1644 -796 1676
rect -764 1644 -760 1676
rect -800 1596 -760 1644
rect -800 1564 -796 1596
rect -764 1564 -760 1596
rect -800 1516 -760 1564
rect -800 1484 -796 1516
rect -764 1484 -760 1516
rect -800 1436 -760 1484
rect -800 1404 -796 1436
rect -764 1404 -760 1436
rect -800 1356 -760 1404
rect -800 1324 -796 1356
rect -764 1324 -760 1356
rect -800 1276 -760 1324
rect -800 1244 -796 1276
rect -764 1244 -760 1276
rect -800 1196 -760 1244
rect -800 1164 -796 1196
rect -764 1164 -760 1196
rect -800 1116 -760 1164
rect -800 1084 -796 1116
rect -764 1084 -760 1116
rect -800 1036 -760 1084
rect -800 1004 -796 1036
rect -764 1004 -760 1036
rect -800 956 -760 1004
rect -800 924 -796 956
rect -764 924 -760 956
rect -800 920 -760 924
rect -720 1676 -680 1680
rect -720 1644 -716 1676
rect -684 1644 -680 1676
rect -720 1596 -680 1644
rect -720 1564 -716 1596
rect -684 1564 -680 1596
rect -720 1516 -680 1564
rect -720 1484 -716 1516
rect -684 1484 -680 1516
rect -720 1436 -680 1484
rect -720 1404 -716 1436
rect -684 1404 -680 1436
rect -720 1356 -680 1404
rect -720 1324 -716 1356
rect -684 1324 -680 1356
rect -720 1276 -680 1324
rect -720 1244 -716 1276
rect -684 1244 -680 1276
rect -720 1196 -680 1244
rect -720 1164 -716 1196
rect -684 1164 -680 1196
rect -720 1116 -680 1164
rect -720 1084 -716 1116
rect -684 1084 -680 1116
rect -720 1036 -680 1084
rect -720 1004 -716 1036
rect -684 1004 -680 1036
rect -720 956 -680 1004
rect -720 924 -716 956
rect -684 924 -680 956
rect -720 920 -680 924
rect -640 1676 -600 1680
rect -640 1644 -636 1676
rect -604 1644 -600 1676
rect -640 1596 -600 1644
rect -640 1564 -636 1596
rect -604 1564 -600 1596
rect -640 1516 -600 1564
rect -640 1484 -636 1516
rect -604 1484 -600 1516
rect -640 1436 -600 1484
rect -640 1404 -636 1436
rect -604 1404 -600 1436
rect -640 1356 -600 1404
rect -640 1324 -636 1356
rect -604 1324 -600 1356
rect -640 1276 -600 1324
rect -640 1244 -636 1276
rect -604 1244 -600 1276
rect -640 1196 -600 1244
rect -640 1164 -636 1196
rect -604 1164 -600 1196
rect -640 1116 -600 1164
rect -640 1084 -636 1116
rect -604 1084 -600 1116
rect -640 1036 -600 1084
rect -640 1004 -636 1036
rect -604 1004 -600 1036
rect -640 956 -600 1004
rect -640 924 -636 956
rect -604 924 -600 956
rect -640 920 -600 924
rect -560 1676 -520 1680
rect -560 1644 -556 1676
rect -524 1644 -520 1676
rect -560 1596 -520 1644
rect -560 1564 -556 1596
rect -524 1564 -520 1596
rect -560 1516 -520 1564
rect -560 1484 -556 1516
rect -524 1484 -520 1516
rect -560 1436 -520 1484
rect -560 1404 -556 1436
rect -524 1404 -520 1436
rect -560 1356 -520 1404
rect -560 1324 -556 1356
rect -524 1324 -520 1356
rect -560 1276 -520 1324
rect -560 1244 -556 1276
rect -524 1244 -520 1276
rect -560 1196 -520 1244
rect -560 1164 -556 1196
rect -524 1164 -520 1196
rect -560 1116 -520 1164
rect -560 1084 -556 1116
rect -524 1084 -520 1116
rect -560 1036 -520 1084
rect -560 1004 -556 1036
rect -524 1004 -520 1036
rect -560 956 -520 1004
rect -560 924 -556 956
rect -524 924 -520 956
rect -560 920 -520 924
rect -480 1676 -440 1680
rect -480 1644 -476 1676
rect -444 1644 -440 1676
rect -480 1596 -440 1644
rect -480 1564 -476 1596
rect -444 1564 -440 1596
rect -480 1516 -440 1564
rect -480 1484 -476 1516
rect -444 1484 -440 1516
rect -480 1436 -440 1484
rect -480 1404 -476 1436
rect -444 1404 -440 1436
rect -480 1356 -440 1404
rect -480 1324 -476 1356
rect -444 1324 -440 1356
rect -480 1276 -440 1324
rect -480 1244 -476 1276
rect -444 1244 -440 1276
rect -480 1196 -440 1244
rect -480 1164 -476 1196
rect -444 1164 -440 1196
rect -480 1116 -440 1164
rect -480 1084 -476 1116
rect -444 1084 -440 1116
rect -480 1036 -440 1084
rect -480 1004 -476 1036
rect -444 1004 -440 1036
rect -480 956 -440 1004
rect -480 924 -476 956
rect -444 924 -440 956
rect -480 920 -440 924
rect -400 1676 -360 1680
rect -400 1644 -396 1676
rect -364 1644 -360 1676
rect -400 1596 -360 1644
rect -400 1564 -396 1596
rect -364 1564 -360 1596
rect -400 1516 -360 1564
rect -400 1484 -396 1516
rect -364 1484 -360 1516
rect -400 1436 -360 1484
rect -400 1404 -396 1436
rect -364 1404 -360 1436
rect -400 1356 -360 1404
rect -400 1324 -396 1356
rect -364 1324 -360 1356
rect -400 1276 -360 1324
rect -400 1244 -396 1276
rect -364 1244 -360 1276
rect -400 1196 -360 1244
rect -400 1164 -396 1196
rect -364 1164 -360 1196
rect -400 1116 -360 1164
rect -400 1084 -396 1116
rect -364 1084 -360 1116
rect -400 1036 -360 1084
rect -400 1004 -396 1036
rect -364 1004 -360 1036
rect -400 956 -360 1004
rect -400 924 -396 956
rect -364 924 -360 956
rect -400 920 -360 924
rect -320 1676 -280 1680
rect -320 1644 -316 1676
rect -284 1644 -280 1676
rect -320 1596 -280 1644
rect -320 1564 -316 1596
rect -284 1564 -280 1596
rect -320 1516 -280 1564
rect -320 1484 -316 1516
rect -284 1484 -280 1516
rect -320 1436 -280 1484
rect -320 1404 -316 1436
rect -284 1404 -280 1436
rect -320 1356 -280 1404
rect -320 1324 -316 1356
rect -284 1324 -280 1356
rect -320 1276 -280 1324
rect -320 1244 -316 1276
rect -284 1244 -280 1276
rect -320 1196 -280 1244
rect -320 1164 -316 1196
rect -284 1164 -280 1196
rect -320 1116 -280 1164
rect -320 1084 -316 1116
rect -284 1084 -280 1116
rect -320 1036 -280 1084
rect -320 1004 -316 1036
rect -284 1004 -280 1036
rect -320 956 -280 1004
rect -320 924 -316 956
rect -284 924 -280 956
rect -320 920 -280 924
rect -240 1676 -200 1680
rect -240 1644 -236 1676
rect -204 1644 -200 1676
rect -240 1596 -200 1644
rect -240 1564 -236 1596
rect -204 1564 -200 1596
rect -240 1516 -200 1564
rect -240 1484 -236 1516
rect -204 1484 -200 1516
rect -240 1436 -200 1484
rect -240 1404 -236 1436
rect -204 1404 -200 1436
rect -240 1356 -200 1404
rect -240 1324 -236 1356
rect -204 1324 -200 1356
rect -240 1276 -200 1324
rect -240 1244 -236 1276
rect -204 1244 -200 1276
rect -240 1196 -200 1244
rect -240 1164 -236 1196
rect -204 1164 -200 1196
rect -240 1116 -200 1164
rect -240 1084 -236 1116
rect -204 1084 -200 1116
rect -240 1036 -200 1084
rect -240 1004 -236 1036
rect -204 1004 -200 1036
rect -240 956 -200 1004
rect -240 924 -236 956
rect -204 924 -200 956
rect -240 920 -200 924
rect -160 1676 -120 1680
rect -160 1644 -156 1676
rect -124 1644 -120 1676
rect -160 1596 -120 1644
rect -160 1564 -156 1596
rect -124 1564 -120 1596
rect -160 1516 -120 1564
rect -160 1484 -156 1516
rect -124 1484 -120 1516
rect -160 1436 -120 1484
rect -160 1404 -156 1436
rect -124 1404 -120 1436
rect -160 1356 -120 1404
rect -160 1324 -156 1356
rect -124 1324 -120 1356
rect -160 1276 -120 1324
rect -160 1244 -156 1276
rect -124 1244 -120 1276
rect -160 1196 -120 1244
rect -160 1164 -156 1196
rect -124 1164 -120 1196
rect -160 1116 -120 1164
rect -160 1084 -156 1116
rect -124 1084 -120 1116
rect -160 1036 -120 1084
rect -160 1004 -156 1036
rect -124 1004 -120 1036
rect -160 956 -120 1004
rect -160 924 -156 956
rect -124 924 -120 956
rect -160 920 -120 924
rect -80 1676 -40 1680
rect -80 1644 -76 1676
rect -44 1644 -40 1676
rect -80 1596 -40 1644
rect -80 1564 -76 1596
rect -44 1564 -40 1596
rect -80 1516 -40 1564
rect -80 1484 -76 1516
rect -44 1484 -40 1516
rect -80 1436 -40 1484
rect -80 1404 -76 1436
rect -44 1404 -40 1436
rect -80 1356 -40 1404
rect -80 1324 -76 1356
rect -44 1324 -40 1356
rect -80 1276 -40 1324
rect -80 1244 -76 1276
rect -44 1244 -40 1276
rect -80 1196 -40 1244
rect -80 1164 -76 1196
rect -44 1164 -40 1196
rect -80 1116 -40 1164
rect -80 1084 -76 1116
rect -44 1084 -40 1116
rect -80 1036 -40 1084
rect -80 1004 -76 1036
rect -44 1004 -40 1036
rect -80 956 -40 1004
rect -80 924 -76 956
rect -44 924 -40 956
rect -80 920 -40 924
rect 0 1676 40 1680
rect 0 1644 4 1676
rect 36 1644 40 1676
rect 0 1596 40 1644
rect 0 1564 4 1596
rect 36 1564 40 1596
rect 0 1516 40 1564
rect 0 1484 4 1516
rect 36 1484 40 1516
rect 0 1436 40 1484
rect 0 1404 4 1436
rect 36 1404 40 1436
rect 0 1356 40 1404
rect 0 1324 4 1356
rect 36 1324 40 1356
rect 0 1276 40 1324
rect 0 1244 4 1276
rect 36 1244 40 1276
rect 0 1196 40 1244
rect 0 1164 4 1196
rect 36 1164 40 1196
rect 0 1116 40 1164
rect 0 1084 4 1116
rect 36 1084 40 1116
rect 0 1036 40 1084
rect 0 1004 4 1036
rect 36 1004 40 1036
rect 0 956 40 1004
rect 0 924 4 956
rect 36 924 40 956
rect 0 920 40 924
rect 80 1676 120 1680
rect 80 1644 84 1676
rect 116 1644 120 1676
rect 80 1596 120 1644
rect 80 1564 84 1596
rect 116 1564 120 1596
rect 80 1516 120 1564
rect 80 1484 84 1516
rect 116 1484 120 1516
rect 80 1436 120 1484
rect 80 1404 84 1436
rect 116 1404 120 1436
rect 80 1356 120 1404
rect 80 1324 84 1356
rect 116 1324 120 1356
rect 80 1276 120 1324
rect 80 1244 84 1276
rect 116 1244 120 1276
rect 80 1196 120 1244
rect 80 1164 84 1196
rect 116 1164 120 1196
rect 80 1116 120 1164
rect 80 1084 84 1116
rect 116 1084 120 1116
rect 80 1036 120 1084
rect 80 1004 84 1036
rect 116 1004 120 1036
rect 80 956 120 1004
rect 80 924 84 956
rect 116 924 120 956
rect 80 920 120 924
rect 160 1676 200 1680
rect 160 1644 164 1676
rect 196 1644 200 1676
rect 160 1596 200 1644
rect 160 1564 164 1596
rect 196 1564 200 1596
rect 160 1516 200 1564
rect 160 1484 164 1516
rect 196 1484 200 1516
rect 160 1436 200 1484
rect 160 1404 164 1436
rect 196 1404 200 1436
rect 160 1356 200 1404
rect 160 1324 164 1356
rect 196 1324 200 1356
rect 160 1276 200 1324
rect 160 1244 164 1276
rect 196 1244 200 1276
rect 160 1196 200 1244
rect 160 1164 164 1196
rect 196 1164 200 1196
rect 160 1116 200 1164
rect 160 1084 164 1116
rect 196 1084 200 1116
rect 160 1036 200 1084
rect 160 1004 164 1036
rect 196 1004 200 1036
rect 160 956 200 1004
rect 160 924 164 956
rect 196 924 200 956
rect 160 920 200 924
rect 240 1676 280 1680
rect 240 1644 244 1676
rect 276 1644 280 1676
rect 240 1596 280 1644
rect 240 1564 244 1596
rect 276 1564 280 1596
rect 240 1516 280 1564
rect 240 1484 244 1516
rect 276 1484 280 1516
rect 240 1436 280 1484
rect 240 1404 244 1436
rect 276 1404 280 1436
rect 240 1356 280 1404
rect 240 1324 244 1356
rect 276 1324 280 1356
rect 240 1276 280 1324
rect 240 1244 244 1276
rect 276 1244 280 1276
rect 240 1196 280 1244
rect 240 1164 244 1196
rect 276 1164 280 1196
rect 240 1116 280 1164
rect 240 1084 244 1116
rect 276 1084 280 1116
rect 240 1036 280 1084
rect 240 1004 244 1036
rect 276 1004 280 1036
rect 240 956 280 1004
rect 240 924 244 956
rect 276 924 280 956
rect 240 920 280 924
rect 320 1676 360 1680
rect 320 1644 324 1676
rect 356 1644 360 1676
rect 320 1596 360 1644
rect 320 1564 324 1596
rect 356 1564 360 1596
rect 320 1516 360 1564
rect 320 1484 324 1516
rect 356 1484 360 1516
rect 320 1436 360 1484
rect 320 1404 324 1436
rect 356 1404 360 1436
rect 320 1356 360 1404
rect 320 1324 324 1356
rect 356 1324 360 1356
rect 320 1276 360 1324
rect 320 1244 324 1276
rect 356 1244 360 1276
rect 320 1196 360 1244
rect 320 1164 324 1196
rect 356 1164 360 1196
rect 320 1116 360 1164
rect 320 1084 324 1116
rect 356 1084 360 1116
rect 320 1036 360 1084
rect 320 1004 324 1036
rect 356 1004 360 1036
rect 320 956 360 1004
rect 320 924 324 956
rect 356 924 360 956
rect 320 920 360 924
rect 400 1676 440 1680
rect 400 1644 404 1676
rect 436 1644 440 1676
rect 400 1596 440 1644
rect 400 1564 404 1596
rect 436 1564 440 1596
rect 400 1516 440 1564
rect 400 1484 404 1516
rect 436 1484 440 1516
rect 400 1436 440 1484
rect 400 1404 404 1436
rect 436 1404 440 1436
rect 400 1356 440 1404
rect 400 1324 404 1356
rect 436 1324 440 1356
rect 400 1276 440 1324
rect 400 1244 404 1276
rect 436 1244 440 1276
rect 400 1196 440 1244
rect 400 1164 404 1196
rect 436 1164 440 1196
rect 400 1116 440 1164
rect 400 1084 404 1116
rect 436 1084 440 1116
rect 400 1036 440 1084
rect 400 1004 404 1036
rect 436 1004 440 1036
rect 400 956 440 1004
rect 400 924 404 956
rect 436 924 440 956
rect 400 920 440 924
rect 480 1676 520 1680
rect 480 1644 484 1676
rect 516 1644 520 1676
rect 480 1596 520 1644
rect 480 1564 484 1596
rect 516 1564 520 1596
rect 480 1516 520 1564
rect 480 1484 484 1516
rect 516 1484 520 1516
rect 480 1436 520 1484
rect 480 1404 484 1436
rect 516 1404 520 1436
rect 480 1356 520 1404
rect 480 1324 484 1356
rect 516 1324 520 1356
rect 480 1276 520 1324
rect 480 1244 484 1276
rect 516 1244 520 1276
rect 480 1196 520 1244
rect 480 1164 484 1196
rect 516 1164 520 1196
rect 480 1116 520 1164
rect 480 1084 484 1116
rect 516 1084 520 1116
rect 480 1036 520 1084
rect 480 1004 484 1036
rect 516 1004 520 1036
rect 480 956 520 1004
rect 480 924 484 956
rect 516 924 520 956
rect 480 920 520 924
rect 560 1676 600 1680
rect 560 1644 564 1676
rect 596 1644 600 1676
rect 560 1596 600 1644
rect 560 1564 564 1596
rect 596 1564 600 1596
rect 560 1516 600 1564
rect 560 1484 564 1516
rect 596 1484 600 1516
rect 560 1436 600 1484
rect 560 1404 564 1436
rect 596 1404 600 1436
rect 560 1356 600 1404
rect 560 1324 564 1356
rect 596 1324 600 1356
rect 560 1276 600 1324
rect 560 1244 564 1276
rect 596 1244 600 1276
rect 560 1196 600 1244
rect 560 1164 564 1196
rect 596 1164 600 1196
rect 560 1116 600 1164
rect 560 1084 564 1116
rect 596 1084 600 1116
rect 560 1036 600 1084
rect 560 1004 564 1036
rect 596 1004 600 1036
rect 560 956 600 1004
rect 560 924 564 956
rect 596 924 600 956
rect 560 920 600 924
rect 640 1676 680 1680
rect 640 1644 644 1676
rect 676 1644 680 1676
rect 640 1596 680 1644
rect 640 1564 644 1596
rect 676 1564 680 1596
rect 640 1516 680 1564
rect 640 1484 644 1516
rect 676 1484 680 1516
rect 640 1436 680 1484
rect 640 1404 644 1436
rect 676 1404 680 1436
rect 640 1356 680 1404
rect 640 1324 644 1356
rect 676 1324 680 1356
rect 640 1276 680 1324
rect 640 1244 644 1276
rect 676 1244 680 1276
rect 640 1196 680 1244
rect 640 1164 644 1196
rect 676 1164 680 1196
rect 640 1116 680 1164
rect 640 1084 644 1116
rect 676 1084 680 1116
rect 640 1036 680 1084
rect 640 1004 644 1036
rect 676 1004 680 1036
rect 640 956 680 1004
rect 640 924 644 956
rect 676 924 680 956
rect 640 920 680 924
rect 720 1676 760 1680
rect 720 1644 724 1676
rect 756 1644 760 1676
rect 720 1596 760 1644
rect 720 1564 724 1596
rect 756 1564 760 1596
rect 720 1516 760 1564
rect 720 1484 724 1516
rect 756 1484 760 1516
rect 720 1436 760 1484
rect 720 1404 724 1436
rect 756 1404 760 1436
rect 720 1356 760 1404
rect 720 1324 724 1356
rect 756 1324 760 1356
rect 720 1276 760 1324
rect 720 1244 724 1276
rect 756 1244 760 1276
rect 720 1196 760 1244
rect 720 1164 724 1196
rect 756 1164 760 1196
rect 720 1116 760 1164
rect 720 1084 724 1116
rect 756 1084 760 1116
rect 720 1036 760 1084
rect 720 1004 724 1036
rect 756 1004 760 1036
rect 720 956 760 1004
rect 720 924 724 956
rect 756 924 760 956
rect 720 920 760 924
rect 800 1676 840 1680
rect 800 1644 804 1676
rect 836 1644 840 1676
rect 800 1596 840 1644
rect 800 1564 804 1596
rect 836 1564 840 1596
rect 800 1516 840 1564
rect 800 1484 804 1516
rect 836 1484 840 1516
rect 800 1436 840 1484
rect 800 1404 804 1436
rect 836 1404 840 1436
rect 800 1356 840 1404
rect 800 1324 804 1356
rect 836 1324 840 1356
rect 800 1276 840 1324
rect 800 1244 804 1276
rect 836 1244 840 1276
rect 800 1196 840 1244
rect 800 1164 804 1196
rect 836 1164 840 1196
rect 800 1116 840 1164
rect 800 1084 804 1116
rect 836 1084 840 1116
rect 800 1036 840 1084
rect 800 1004 804 1036
rect 836 1004 840 1036
rect 800 956 840 1004
rect 800 924 804 956
rect 836 924 840 956
rect 800 920 840 924
rect 880 1676 920 1680
rect 880 1644 884 1676
rect 916 1644 920 1676
rect 880 1596 920 1644
rect 880 1564 884 1596
rect 916 1564 920 1596
rect 880 1516 920 1564
rect 880 1484 884 1516
rect 916 1484 920 1516
rect 880 1436 920 1484
rect 880 1404 884 1436
rect 916 1404 920 1436
rect 880 1356 920 1404
rect 880 1324 884 1356
rect 916 1324 920 1356
rect 880 1276 920 1324
rect 880 1244 884 1276
rect 916 1244 920 1276
rect 880 1196 920 1244
rect 880 1164 884 1196
rect 916 1164 920 1196
rect 880 1116 920 1164
rect 880 1084 884 1116
rect 916 1084 920 1116
rect 880 1036 920 1084
rect 880 1004 884 1036
rect 916 1004 920 1036
rect 880 956 920 1004
rect 880 924 884 956
rect 916 924 920 956
rect 880 920 920 924
rect 960 1676 1000 1680
rect 960 1644 964 1676
rect 996 1644 1000 1676
rect 960 1596 1000 1644
rect 960 1564 964 1596
rect 996 1564 1000 1596
rect 960 1516 1000 1564
rect 960 1484 964 1516
rect 996 1484 1000 1516
rect 960 1436 1000 1484
rect 960 1404 964 1436
rect 996 1404 1000 1436
rect 960 1356 1000 1404
rect 960 1324 964 1356
rect 996 1324 1000 1356
rect 960 1276 1000 1324
rect 960 1244 964 1276
rect 996 1244 1000 1276
rect 960 1196 1000 1244
rect 960 1164 964 1196
rect 996 1164 1000 1196
rect 960 1116 1000 1164
rect 960 1084 964 1116
rect 996 1084 1000 1116
rect 960 1036 1000 1084
rect 960 1004 964 1036
rect 996 1004 1000 1036
rect 960 956 1000 1004
rect 960 924 964 956
rect 996 924 1000 956
rect 960 920 1000 924
rect 1040 1676 1080 1680
rect 1040 1644 1044 1676
rect 1076 1644 1080 1676
rect 1040 1596 1080 1644
rect 1040 1564 1044 1596
rect 1076 1564 1080 1596
rect 1040 1516 1080 1564
rect 1040 1484 1044 1516
rect 1076 1484 1080 1516
rect 1040 1436 1080 1484
rect 1040 1404 1044 1436
rect 1076 1404 1080 1436
rect 1040 1356 1080 1404
rect 1040 1324 1044 1356
rect 1076 1324 1080 1356
rect 1040 1276 1080 1324
rect 1040 1244 1044 1276
rect 1076 1244 1080 1276
rect 1040 1196 1080 1244
rect 1040 1164 1044 1196
rect 1076 1164 1080 1196
rect 1040 1116 1080 1164
rect 1040 1084 1044 1116
rect 1076 1084 1080 1116
rect 1040 1036 1080 1084
rect 1040 1004 1044 1036
rect 1076 1004 1080 1036
rect 1040 956 1080 1004
rect 1040 924 1044 956
rect 1076 924 1080 956
rect 1040 920 1080 924
rect 1120 1676 1160 1680
rect 1120 1644 1124 1676
rect 1156 1644 1160 1676
rect 1120 1596 1160 1644
rect 1120 1564 1124 1596
rect 1156 1564 1160 1596
rect 1120 1516 1160 1564
rect 1120 1484 1124 1516
rect 1156 1484 1160 1516
rect 1120 1436 1160 1484
rect 1120 1404 1124 1436
rect 1156 1404 1160 1436
rect 1120 1356 1160 1404
rect 1120 1324 1124 1356
rect 1156 1324 1160 1356
rect 1120 1276 1160 1324
rect 1120 1244 1124 1276
rect 1156 1244 1160 1276
rect 1120 1196 1160 1244
rect 1120 1164 1124 1196
rect 1156 1164 1160 1196
rect 1120 1116 1160 1164
rect 1120 1084 1124 1116
rect 1156 1084 1160 1116
rect 1120 1036 1160 1084
rect 1120 1004 1124 1036
rect 1156 1004 1160 1036
rect 1120 956 1160 1004
rect 1120 924 1124 956
rect 1156 924 1160 956
rect 1120 920 1160 924
rect 1200 1676 1240 1680
rect 1200 1644 1204 1676
rect 1236 1644 1240 1676
rect 1200 1596 1240 1644
rect 1200 1564 1204 1596
rect 1236 1564 1240 1596
rect 1200 1516 1240 1564
rect 1200 1484 1204 1516
rect 1236 1484 1240 1516
rect 1200 1436 1240 1484
rect 1200 1404 1204 1436
rect 1236 1404 1240 1436
rect 1200 1356 1240 1404
rect 1200 1324 1204 1356
rect 1236 1324 1240 1356
rect 1200 1276 1240 1324
rect 1200 1244 1204 1276
rect 1236 1244 1240 1276
rect 1200 1196 1240 1244
rect 1200 1164 1204 1196
rect 1236 1164 1240 1196
rect 1200 1116 1240 1164
rect 1200 1084 1204 1116
rect 1236 1084 1240 1116
rect 1200 1036 1240 1084
rect 1200 1004 1204 1036
rect 1236 1004 1240 1036
rect 1200 956 1240 1004
rect 1200 924 1204 956
rect 1236 924 1240 956
rect 1200 920 1240 924
rect 1280 1676 1320 1680
rect 1280 1644 1284 1676
rect 1316 1644 1320 1676
rect 1280 1596 1320 1644
rect 1280 1564 1284 1596
rect 1316 1564 1320 1596
rect 1280 1516 1320 1564
rect 1280 1484 1284 1516
rect 1316 1484 1320 1516
rect 1280 1436 1320 1484
rect 1280 1404 1284 1436
rect 1316 1404 1320 1436
rect 1280 1356 1320 1404
rect 1280 1324 1284 1356
rect 1316 1324 1320 1356
rect 1280 1276 1320 1324
rect 1280 1244 1284 1276
rect 1316 1244 1320 1276
rect 1280 1196 1320 1244
rect 1280 1164 1284 1196
rect 1316 1164 1320 1196
rect 1280 1116 1320 1164
rect 1280 1084 1284 1116
rect 1316 1084 1320 1116
rect 1280 1036 1320 1084
rect 1280 1004 1284 1036
rect 1316 1004 1320 1036
rect 1280 956 1320 1004
rect 1280 924 1284 956
rect 1316 924 1320 956
rect 1280 920 1320 924
rect 1360 1676 1400 1680
rect 1360 1644 1364 1676
rect 1396 1644 1400 1676
rect 1360 1596 1400 1644
rect 1360 1564 1364 1596
rect 1396 1564 1400 1596
rect 1360 1516 1400 1564
rect 1360 1484 1364 1516
rect 1396 1484 1400 1516
rect 1360 1436 1400 1484
rect 1360 1404 1364 1436
rect 1396 1404 1400 1436
rect 1360 1356 1400 1404
rect 1360 1324 1364 1356
rect 1396 1324 1400 1356
rect 1360 1276 1400 1324
rect 1360 1244 1364 1276
rect 1396 1244 1400 1276
rect 1360 1196 1400 1244
rect 1360 1164 1364 1196
rect 1396 1164 1400 1196
rect 1360 1116 1400 1164
rect 1360 1084 1364 1116
rect 1396 1084 1400 1116
rect 1360 1036 1400 1084
rect 1360 1004 1364 1036
rect 1396 1004 1400 1036
rect 1360 956 1400 1004
rect 1360 924 1364 956
rect 1396 924 1400 956
rect 1360 920 1400 924
rect 1440 1676 1480 1680
rect 1440 1644 1444 1676
rect 1476 1644 1480 1676
rect 1440 1596 1480 1644
rect 1440 1564 1444 1596
rect 1476 1564 1480 1596
rect 1440 1516 1480 1564
rect 1440 1484 1444 1516
rect 1476 1484 1480 1516
rect 1440 1436 1480 1484
rect 1440 1404 1444 1436
rect 1476 1404 1480 1436
rect 1440 1356 1480 1404
rect 1440 1324 1444 1356
rect 1476 1324 1480 1356
rect 1440 1276 1480 1324
rect 1440 1244 1444 1276
rect 1476 1244 1480 1276
rect 1440 1196 1480 1244
rect 1440 1164 1444 1196
rect 1476 1164 1480 1196
rect 1440 1116 1480 1164
rect 1440 1084 1444 1116
rect 1476 1084 1480 1116
rect 1440 1036 1480 1084
rect 1440 1004 1444 1036
rect 1476 1004 1480 1036
rect 1440 956 1480 1004
rect 1440 924 1444 956
rect 1476 924 1480 956
rect 1440 920 1480 924
rect 1520 1676 1560 1680
rect 1520 1644 1524 1676
rect 1556 1644 1560 1676
rect 1520 1596 1560 1644
rect 1520 1564 1524 1596
rect 1556 1564 1560 1596
rect 1520 1516 1560 1564
rect 1520 1484 1524 1516
rect 1556 1484 1560 1516
rect 1520 1436 1560 1484
rect 1520 1404 1524 1436
rect 1556 1404 1560 1436
rect 1520 1356 1560 1404
rect 1520 1324 1524 1356
rect 1556 1324 1560 1356
rect 1520 1276 1560 1324
rect 1520 1244 1524 1276
rect 1556 1244 1560 1276
rect 1520 1196 1560 1244
rect 1520 1164 1524 1196
rect 1556 1164 1560 1196
rect 1520 1116 1560 1164
rect 1520 1084 1524 1116
rect 1556 1084 1560 1116
rect 1520 1036 1560 1084
rect 1520 1004 1524 1036
rect 1556 1004 1560 1036
rect 1520 956 1560 1004
rect 1520 924 1524 956
rect 1556 924 1560 956
rect 1520 920 1560 924
rect 1600 1676 1640 1680
rect 1600 1644 1604 1676
rect 1636 1644 1640 1676
rect 1600 1596 1640 1644
rect 1600 1564 1604 1596
rect 1636 1564 1640 1596
rect 1600 1516 1640 1564
rect 1600 1484 1604 1516
rect 1636 1484 1640 1516
rect 1600 1436 1640 1484
rect 1600 1404 1604 1436
rect 1636 1404 1640 1436
rect 1600 1356 1640 1404
rect 1600 1324 1604 1356
rect 1636 1324 1640 1356
rect 1600 1276 1640 1324
rect 1600 1244 1604 1276
rect 1636 1244 1640 1276
rect 1600 1196 1640 1244
rect 1600 1164 1604 1196
rect 1636 1164 1640 1196
rect 1600 1116 1640 1164
rect 1600 1084 1604 1116
rect 1636 1084 1640 1116
rect 1600 1036 1640 1084
rect 1600 1004 1604 1036
rect 1636 1004 1640 1036
rect 1600 956 1640 1004
rect 1600 924 1604 956
rect 1636 924 1640 956
rect 1600 920 1640 924
rect 1680 1676 1720 1680
rect 1680 1644 1684 1676
rect 1716 1644 1720 1676
rect 1680 1596 1720 1644
rect 1680 1564 1684 1596
rect 1716 1564 1720 1596
rect 1680 1516 1720 1564
rect 1680 1484 1684 1516
rect 1716 1484 1720 1516
rect 1680 1436 1720 1484
rect 1680 1404 1684 1436
rect 1716 1404 1720 1436
rect 1680 1356 1720 1404
rect 1680 1324 1684 1356
rect 1716 1324 1720 1356
rect 1680 1276 1720 1324
rect 1680 1244 1684 1276
rect 1716 1244 1720 1276
rect 1680 1196 1720 1244
rect 1680 1164 1684 1196
rect 1716 1164 1720 1196
rect 1680 1116 1720 1164
rect 1680 1084 1684 1116
rect 1716 1084 1720 1116
rect 1680 1036 1720 1084
rect 1680 1004 1684 1036
rect 1716 1004 1720 1036
rect 1680 956 1720 1004
rect 1680 924 1684 956
rect 1716 924 1720 956
rect 1680 920 1720 924
rect 1760 1676 1800 1680
rect 1760 1644 1764 1676
rect 1796 1644 1800 1676
rect 1760 1596 1800 1644
rect 1760 1564 1764 1596
rect 1796 1564 1800 1596
rect 1760 1516 1800 1564
rect 1760 1484 1764 1516
rect 1796 1484 1800 1516
rect 1760 1436 1800 1484
rect 1760 1404 1764 1436
rect 1796 1404 1800 1436
rect 1760 1356 1800 1404
rect 1760 1324 1764 1356
rect 1796 1324 1800 1356
rect 1760 1276 1800 1324
rect 1760 1244 1764 1276
rect 1796 1244 1800 1276
rect 1760 1196 1800 1244
rect 1760 1164 1764 1196
rect 1796 1164 1800 1196
rect 1760 1116 1800 1164
rect 1760 1084 1764 1116
rect 1796 1084 1800 1116
rect 1760 1036 1800 1084
rect 1760 1004 1764 1036
rect 1796 1004 1800 1036
rect 1760 956 1800 1004
rect 1760 924 1764 956
rect 1796 924 1800 956
rect 1760 920 1800 924
rect 1840 1676 1880 1680
rect 1840 1644 1844 1676
rect 1876 1644 1880 1676
rect 1840 1596 1880 1644
rect 1840 1564 1844 1596
rect 1876 1564 1880 1596
rect 1840 1516 1880 1564
rect 1840 1484 1844 1516
rect 1876 1484 1880 1516
rect 1840 1436 1880 1484
rect 1840 1404 1844 1436
rect 1876 1404 1880 1436
rect 1840 1356 1880 1404
rect 1840 1324 1844 1356
rect 1876 1324 1880 1356
rect 1840 1276 1880 1324
rect 1840 1244 1844 1276
rect 1876 1244 1880 1276
rect 1840 1196 1880 1244
rect 1840 1164 1844 1196
rect 1876 1164 1880 1196
rect 1840 1116 1880 1164
rect 1840 1084 1844 1116
rect 1876 1084 1880 1116
rect 1840 1036 1880 1084
rect 1840 1004 1844 1036
rect 1876 1004 1880 1036
rect 1840 956 1880 1004
rect 1840 924 1844 956
rect 1876 924 1880 956
rect 1840 920 1880 924
rect 1920 1676 1960 1680
rect 1920 1644 1924 1676
rect 1956 1644 1960 1676
rect 1920 1596 1960 1644
rect 1920 1564 1924 1596
rect 1956 1564 1960 1596
rect 1920 1516 1960 1564
rect 1920 1484 1924 1516
rect 1956 1484 1960 1516
rect 1920 1436 1960 1484
rect 1920 1404 1924 1436
rect 1956 1404 1960 1436
rect 1920 1356 1960 1404
rect 1920 1324 1924 1356
rect 1956 1324 1960 1356
rect 1920 1276 1960 1324
rect 1920 1244 1924 1276
rect 1956 1244 1960 1276
rect 1920 1196 1960 1244
rect 1920 1164 1924 1196
rect 1956 1164 1960 1196
rect 1920 1116 1960 1164
rect 1920 1084 1924 1116
rect 1956 1084 1960 1116
rect 1920 1036 1960 1084
rect 1920 1004 1924 1036
rect 1956 1004 1960 1036
rect 1920 956 1960 1004
rect 1920 924 1924 956
rect 1956 924 1960 956
rect 1920 920 1960 924
rect 2000 1676 2040 1680
rect 2000 1644 2004 1676
rect 2036 1644 2040 1676
rect 2000 1596 2040 1644
rect 2000 1564 2004 1596
rect 2036 1564 2040 1596
rect 2000 1516 2040 1564
rect 2000 1484 2004 1516
rect 2036 1484 2040 1516
rect 2000 1436 2040 1484
rect 2000 1404 2004 1436
rect 2036 1404 2040 1436
rect 2000 1356 2040 1404
rect 2000 1324 2004 1356
rect 2036 1324 2040 1356
rect 2000 1276 2040 1324
rect 2000 1244 2004 1276
rect 2036 1244 2040 1276
rect 2000 1196 2040 1244
rect 2000 1164 2004 1196
rect 2036 1164 2040 1196
rect 2000 1116 2040 1164
rect 2000 1084 2004 1116
rect 2036 1084 2040 1116
rect 2000 1036 2040 1084
rect 2000 1004 2004 1036
rect 2036 1004 2040 1036
rect 2000 956 2040 1004
rect 2000 924 2004 956
rect 2036 924 2040 956
rect 2000 920 2040 924
rect 2080 1676 2120 1680
rect 2080 1644 2084 1676
rect 2116 1644 2120 1676
rect 2080 1596 2120 1644
rect 2080 1564 2084 1596
rect 2116 1564 2120 1596
rect 2080 1516 2120 1564
rect 2080 1484 2084 1516
rect 2116 1484 2120 1516
rect 2080 1436 2120 1484
rect 2080 1404 2084 1436
rect 2116 1404 2120 1436
rect 2080 1356 2120 1404
rect 2080 1324 2084 1356
rect 2116 1324 2120 1356
rect 2080 1276 2120 1324
rect 2080 1244 2084 1276
rect 2116 1244 2120 1276
rect 2080 1196 2120 1244
rect 2080 1164 2084 1196
rect 2116 1164 2120 1196
rect 2080 1116 2120 1164
rect 2080 1084 2084 1116
rect 2116 1084 2120 1116
rect 2080 1036 2120 1084
rect 2080 1004 2084 1036
rect 2116 1004 2120 1036
rect 2080 956 2120 1004
rect 2080 924 2084 956
rect 2116 924 2120 956
rect 2080 920 2120 924
rect 2160 1676 2200 1680
rect 2160 1644 2164 1676
rect 2196 1644 2200 1676
rect 2160 1596 2200 1644
rect 2160 1564 2164 1596
rect 2196 1564 2200 1596
rect 2160 1516 2200 1564
rect 2160 1484 2164 1516
rect 2196 1484 2200 1516
rect 2160 1436 2200 1484
rect 2160 1404 2164 1436
rect 2196 1404 2200 1436
rect 2160 1356 2200 1404
rect 2160 1324 2164 1356
rect 2196 1324 2200 1356
rect 2160 1276 2200 1324
rect 2160 1244 2164 1276
rect 2196 1244 2200 1276
rect 2160 1196 2200 1244
rect 2160 1164 2164 1196
rect 2196 1164 2200 1196
rect 2160 1116 2200 1164
rect 2160 1084 2164 1116
rect 2196 1084 2200 1116
rect 2160 1036 2200 1084
rect 2160 1004 2164 1036
rect 2196 1004 2200 1036
rect 2160 956 2200 1004
rect 2160 924 2164 956
rect 2196 924 2200 956
rect 2160 920 2200 924
rect 2240 1676 2280 1680
rect 2240 1644 2244 1676
rect 2276 1644 2280 1676
rect 2240 1596 2280 1644
rect 2240 1564 2244 1596
rect 2276 1564 2280 1596
rect 2240 1516 2280 1564
rect 2240 1484 2244 1516
rect 2276 1484 2280 1516
rect 2240 1436 2280 1484
rect 2240 1404 2244 1436
rect 2276 1404 2280 1436
rect 2240 1356 2280 1404
rect 2240 1324 2244 1356
rect 2276 1324 2280 1356
rect 2240 1276 2280 1324
rect 2240 1244 2244 1276
rect 2276 1244 2280 1276
rect 2240 1196 2280 1244
rect 2240 1164 2244 1196
rect 2276 1164 2280 1196
rect 2240 1116 2280 1164
rect 2240 1084 2244 1116
rect 2276 1084 2280 1116
rect 2240 1036 2280 1084
rect 2240 1004 2244 1036
rect 2276 1004 2280 1036
rect 2240 956 2280 1004
rect 2240 924 2244 956
rect 2276 924 2280 956
rect 2240 920 2280 924
rect 2320 1676 2360 1680
rect 2320 1644 2324 1676
rect 2356 1644 2360 1676
rect 2320 1596 2360 1644
rect 2320 1564 2324 1596
rect 2356 1564 2360 1596
rect 2320 1516 2360 1564
rect 2320 1484 2324 1516
rect 2356 1484 2360 1516
rect 2320 1436 2360 1484
rect 2320 1404 2324 1436
rect 2356 1404 2360 1436
rect 2320 1356 2360 1404
rect 2320 1324 2324 1356
rect 2356 1324 2360 1356
rect 2320 1276 2360 1324
rect 2320 1244 2324 1276
rect 2356 1244 2360 1276
rect 2320 1196 2360 1244
rect 2320 1164 2324 1196
rect 2356 1164 2360 1196
rect 2320 1116 2360 1164
rect 2320 1084 2324 1116
rect 2356 1084 2360 1116
rect 2320 1036 2360 1084
rect 2320 1004 2324 1036
rect 2356 1004 2360 1036
rect 2320 956 2360 1004
rect 2320 924 2324 956
rect 2356 924 2360 956
rect 2320 920 2360 924
rect 2400 1676 2440 1680
rect 2400 1644 2404 1676
rect 2436 1644 2440 1676
rect 2400 1596 2440 1644
rect 2400 1564 2404 1596
rect 2436 1564 2440 1596
rect 2400 1516 2440 1564
rect 2400 1484 2404 1516
rect 2436 1484 2440 1516
rect 2400 1436 2440 1484
rect 2400 1404 2404 1436
rect 2436 1404 2440 1436
rect 2400 1356 2440 1404
rect 2400 1324 2404 1356
rect 2436 1324 2440 1356
rect 2400 1276 2440 1324
rect 2400 1244 2404 1276
rect 2436 1244 2440 1276
rect 2400 1196 2440 1244
rect 2400 1164 2404 1196
rect 2436 1164 2440 1196
rect 2400 1116 2440 1164
rect 2400 1084 2404 1116
rect 2436 1084 2440 1116
rect 2400 1036 2440 1084
rect 2400 1004 2404 1036
rect 2436 1004 2440 1036
rect 2400 956 2440 1004
rect 2400 924 2404 956
rect 2436 924 2440 956
rect 2400 920 2440 924
rect 2480 1676 2520 1680
rect 2480 1644 2484 1676
rect 2516 1644 2520 1676
rect 2480 1596 2520 1644
rect 2480 1564 2484 1596
rect 2516 1564 2520 1596
rect 2480 1516 2520 1564
rect 2480 1484 2484 1516
rect 2516 1484 2520 1516
rect 2480 1436 2520 1484
rect 2480 1404 2484 1436
rect 2516 1404 2520 1436
rect 2480 1356 2520 1404
rect 2480 1324 2484 1356
rect 2516 1324 2520 1356
rect 2480 1276 2520 1324
rect 2480 1244 2484 1276
rect 2516 1244 2520 1276
rect 2480 1196 2520 1244
rect 2480 1164 2484 1196
rect 2516 1164 2520 1196
rect 2480 1116 2520 1164
rect 2480 1084 2484 1116
rect 2516 1084 2520 1116
rect 2480 1036 2520 1084
rect 2480 1004 2484 1036
rect 2516 1004 2520 1036
rect 2480 956 2520 1004
rect 2480 924 2484 956
rect 2516 924 2520 956
rect 2480 920 2520 924
rect 2560 1676 2600 1680
rect 2560 1644 2564 1676
rect 2596 1644 2600 1676
rect 2560 1596 2600 1644
rect 2560 1564 2564 1596
rect 2596 1564 2600 1596
rect 2560 1516 2600 1564
rect 2560 1484 2564 1516
rect 2596 1484 2600 1516
rect 2560 1436 2600 1484
rect 2560 1404 2564 1436
rect 2596 1404 2600 1436
rect 2560 1356 2600 1404
rect 2560 1324 2564 1356
rect 2596 1324 2600 1356
rect 2560 1276 2600 1324
rect 2560 1244 2564 1276
rect 2596 1244 2600 1276
rect 2560 1196 2600 1244
rect 2560 1164 2564 1196
rect 2596 1164 2600 1196
rect 2560 1116 2600 1164
rect 2560 1084 2564 1116
rect 2596 1084 2600 1116
rect 2560 1036 2600 1084
rect 2560 1004 2564 1036
rect 2596 1004 2600 1036
rect 2560 956 2600 1004
rect 2560 924 2564 956
rect 2596 924 2600 956
rect 2560 920 2600 924
rect 2640 1676 2680 1680
rect 2640 1644 2644 1676
rect 2676 1644 2680 1676
rect 2640 1596 2680 1644
rect 2640 1564 2644 1596
rect 2676 1564 2680 1596
rect 2640 1516 2680 1564
rect 2640 1484 2644 1516
rect 2676 1484 2680 1516
rect 2640 1436 2680 1484
rect 2640 1404 2644 1436
rect 2676 1404 2680 1436
rect 2640 1356 2680 1404
rect 2640 1324 2644 1356
rect 2676 1324 2680 1356
rect 2640 1276 2680 1324
rect 2640 1244 2644 1276
rect 2676 1244 2680 1276
rect 2640 1196 2680 1244
rect 2640 1164 2644 1196
rect 2676 1164 2680 1196
rect 2640 1116 2680 1164
rect 2640 1084 2644 1116
rect 2676 1084 2680 1116
rect 2640 1036 2680 1084
rect 2640 1004 2644 1036
rect 2676 1004 2680 1036
rect 2640 956 2680 1004
rect 2640 924 2644 956
rect 2676 924 2680 956
rect 2640 920 2680 924
rect 2720 1676 2760 1680
rect 2720 1644 2724 1676
rect 2756 1644 2760 1676
rect 2720 1596 2760 1644
rect 2720 1564 2724 1596
rect 2756 1564 2760 1596
rect 2720 1516 2760 1564
rect 2720 1484 2724 1516
rect 2756 1484 2760 1516
rect 2720 1436 2760 1484
rect 2720 1404 2724 1436
rect 2756 1404 2760 1436
rect 2720 1356 2760 1404
rect 2720 1324 2724 1356
rect 2756 1324 2760 1356
rect 2720 1276 2760 1324
rect 2720 1244 2724 1276
rect 2756 1244 2760 1276
rect 2720 1196 2760 1244
rect 2720 1164 2724 1196
rect 2756 1164 2760 1196
rect 2720 1116 2760 1164
rect 2720 1084 2724 1116
rect 2756 1084 2760 1116
rect 2720 1036 2760 1084
rect 2720 1004 2724 1036
rect 2756 1004 2760 1036
rect 2720 956 2760 1004
rect 2720 924 2724 956
rect 2756 924 2760 956
rect 2720 920 2760 924
rect 2800 1676 2840 1680
rect 2800 1644 2804 1676
rect 2836 1644 2840 1676
rect 2800 1596 2840 1644
rect 2800 1564 2804 1596
rect 2836 1564 2840 1596
rect 2800 1516 2840 1564
rect 2800 1484 2804 1516
rect 2836 1484 2840 1516
rect 2800 1436 2840 1484
rect 2800 1404 2804 1436
rect 2836 1404 2840 1436
rect 2800 1356 2840 1404
rect 2800 1324 2804 1356
rect 2836 1324 2840 1356
rect 2800 1276 2840 1324
rect 2800 1244 2804 1276
rect 2836 1244 2840 1276
rect 2800 1196 2840 1244
rect 2800 1164 2804 1196
rect 2836 1164 2840 1196
rect 2800 1116 2840 1164
rect 2800 1084 2804 1116
rect 2836 1084 2840 1116
rect 2800 1036 2840 1084
rect 2800 1004 2804 1036
rect 2836 1004 2840 1036
rect 2800 956 2840 1004
rect 2800 924 2804 956
rect 2836 924 2840 956
rect 2800 920 2840 924
rect 2880 1676 2920 1680
rect 2880 1644 2884 1676
rect 2916 1644 2920 1676
rect 2880 1596 2920 1644
rect 2880 1564 2884 1596
rect 2916 1564 2920 1596
rect 2880 1516 2920 1564
rect 2880 1484 2884 1516
rect 2916 1484 2920 1516
rect 2880 1436 2920 1484
rect 2880 1404 2884 1436
rect 2916 1404 2920 1436
rect 2880 1356 2920 1404
rect 2880 1324 2884 1356
rect 2916 1324 2920 1356
rect 2880 1276 2920 1324
rect 2880 1244 2884 1276
rect 2916 1244 2920 1276
rect 2880 1196 2920 1244
rect 2880 1164 2884 1196
rect 2916 1164 2920 1196
rect 2880 1116 2920 1164
rect 2880 1084 2884 1116
rect 2916 1084 2920 1116
rect 2880 1036 2920 1084
rect 2880 1004 2884 1036
rect 2916 1004 2920 1036
rect 2880 956 2920 1004
rect 2880 924 2884 956
rect 2916 924 2920 956
rect 2880 920 2920 924
rect 2960 1676 3000 1680
rect 2960 1644 2964 1676
rect 2996 1644 3000 1676
rect 2960 1596 3000 1644
rect 2960 1564 2964 1596
rect 2996 1564 3000 1596
rect 2960 1516 3000 1564
rect 2960 1484 2964 1516
rect 2996 1484 3000 1516
rect 2960 1436 3000 1484
rect 2960 1404 2964 1436
rect 2996 1404 3000 1436
rect 2960 1356 3000 1404
rect 2960 1324 2964 1356
rect 2996 1324 3000 1356
rect 2960 1276 3000 1324
rect 2960 1244 2964 1276
rect 2996 1244 3000 1276
rect 2960 1196 3000 1244
rect 2960 1164 2964 1196
rect 2996 1164 3000 1196
rect 2960 1116 3000 1164
rect 2960 1084 2964 1116
rect 2996 1084 3000 1116
rect 2960 1036 3000 1084
rect 2960 1004 2964 1036
rect 2996 1004 3000 1036
rect 2960 956 3000 1004
rect 2960 924 2964 956
rect 2996 924 3000 956
rect 2960 920 3000 924
rect 3040 1676 3080 1680
rect 3040 1644 3044 1676
rect 3076 1644 3080 1676
rect 3040 1596 3080 1644
rect 3040 1564 3044 1596
rect 3076 1564 3080 1596
rect 3040 1516 3080 1564
rect 3040 1484 3044 1516
rect 3076 1484 3080 1516
rect 3040 1436 3080 1484
rect 3040 1404 3044 1436
rect 3076 1404 3080 1436
rect 3040 1356 3080 1404
rect 3040 1324 3044 1356
rect 3076 1324 3080 1356
rect 3040 1276 3080 1324
rect 3040 1244 3044 1276
rect 3076 1244 3080 1276
rect 3040 1196 3080 1244
rect 3040 1164 3044 1196
rect 3076 1164 3080 1196
rect 3040 1116 3080 1164
rect 3040 1084 3044 1116
rect 3076 1084 3080 1116
rect 3040 1036 3080 1084
rect 3040 1004 3044 1036
rect 3076 1004 3080 1036
rect 3040 956 3080 1004
rect 3040 924 3044 956
rect 3076 924 3080 956
rect 3040 920 3080 924
rect 3120 1676 3160 1680
rect 3120 1644 3124 1676
rect 3156 1644 3160 1676
rect 3120 1596 3160 1644
rect 3120 1564 3124 1596
rect 3156 1564 3160 1596
rect 3120 1516 3160 1564
rect 3120 1484 3124 1516
rect 3156 1484 3160 1516
rect 3120 1436 3160 1484
rect 3120 1404 3124 1436
rect 3156 1404 3160 1436
rect 3120 1356 3160 1404
rect 3120 1324 3124 1356
rect 3156 1324 3160 1356
rect 3120 1276 3160 1324
rect 3120 1244 3124 1276
rect 3156 1244 3160 1276
rect 3120 1196 3160 1244
rect 3120 1164 3124 1196
rect 3156 1164 3160 1196
rect 3120 1116 3160 1164
rect 3120 1084 3124 1116
rect 3156 1084 3160 1116
rect 3120 1036 3160 1084
rect 3120 1004 3124 1036
rect 3156 1004 3160 1036
rect 3120 956 3160 1004
rect 3120 924 3124 956
rect 3156 924 3160 956
rect 3120 920 3160 924
rect 3200 1676 3240 1680
rect 3200 1644 3204 1676
rect 3236 1644 3240 1676
rect 3200 1596 3240 1644
rect 3200 1564 3204 1596
rect 3236 1564 3240 1596
rect 3200 1516 3240 1564
rect 3200 1484 3204 1516
rect 3236 1484 3240 1516
rect 3200 1436 3240 1484
rect 3200 1404 3204 1436
rect 3236 1404 3240 1436
rect 3200 1356 3240 1404
rect 3200 1324 3204 1356
rect 3236 1324 3240 1356
rect 3200 1276 3240 1324
rect 3200 1244 3204 1276
rect 3236 1244 3240 1276
rect 3200 1196 3240 1244
rect 3200 1164 3204 1196
rect 3236 1164 3240 1196
rect 3200 1116 3240 1164
rect 3200 1084 3204 1116
rect 3236 1084 3240 1116
rect 3200 1036 3240 1084
rect 3200 1004 3204 1036
rect 3236 1004 3240 1036
rect 3200 956 3240 1004
rect 3200 924 3204 956
rect 3236 924 3240 956
rect 3200 920 3240 924
rect 3280 1676 3320 1680
rect 3280 1644 3284 1676
rect 3316 1644 3320 1676
rect 3280 1596 3320 1644
rect 3280 1564 3284 1596
rect 3316 1564 3320 1596
rect 3280 1516 3320 1564
rect 3280 1484 3284 1516
rect 3316 1484 3320 1516
rect 3280 1436 3320 1484
rect 3280 1404 3284 1436
rect 3316 1404 3320 1436
rect 3280 1356 3320 1404
rect 3280 1324 3284 1356
rect 3316 1324 3320 1356
rect 3280 1276 3320 1324
rect 3280 1244 3284 1276
rect 3316 1244 3320 1276
rect 3280 1196 3320 1244
rect 3280 1164 3284 1196
rect 3316 1164 3320 1196
rect 3280 1116 3320 1164
rect 3280 1084 3284 1116
rect 3316 1084 3320 1116
rect 3280 1036 3320 1084
rect 3280 1004 3284 1036
rect 3316 1004 3320 1036
rect 3280 956 3320 1004
rect 3280 924 3284 956
rect 3316 924 3320 956
rect 3280 920 3320 924
rect 3360 1676 3400 1680
rect 3360 1644 3364 1676
rect 3396 1644 3400 1676
rect 3360 1596 3400 1644
rect 3360 1564 3364 1596
rect 3396 1564 3400 1596
rect 3360 1516 3400 1564
rect 3360 1484 3364 1516
rect 3396 1484 3400 1516
rect 3360 1436 3400 1484
rect 3360 1404 3364 1436
rect 3396 1404 3400 1436
rect 3360 1356 3400 1404
rect 3360 1324 3364 1356
rect 3396 1324 3400 1356
rect 3360 1276 3400 1324
rect 3360 1244 3364 1276
rect 3396 1244 3400 1276
rect 3360 1196 3400 1244
rect 3360 1164 3364 1196
rect 3396 1164 3400 1196
rect 3360 1116 3400 1164
rect 3360 1084 3364 1116
rect 3396 1084 3400 1116
rect 3360 1036 3400 1084
rect 3360 1004 3364 1036
rect 3396 1004 3400 1036
rect 3360 956 3400 1004
rect 3360 924 3364 956
rect 3396 924 3400 956
rect 3360 920 3400 924
rect 3440 1676 3480 1680
rect 3440 1644 3444 1676
rect 3476 1644 3480 1676
rect 3440 1596 3480 1644
rect 3440 1564 3444 1596
rect 3476 1564 3480 1596
rect 3440 1516 3480 1564
rect 3440 1484 3444 1516
rect 3476 1484 3480 1516
rect 3440 1436 3480 1484
rect 3440 1404 3444 1436
rect 3476 1404 3480 1436
rect 3440 1356 3480 1404
rect 3440 1324 3444 1356
rect 3476 1324 3480 1356
rect 3440 1276 3480 1324
rect 3440 1244 3444 1276
rect 3476 1244 3480 1276
rect 3440 1196 3480 1244
rect 3440 1164 3444 1196
rect 3476 1164 3480 1196
rect 3440 1116 3480 1164
rect 3440 1084 3444 1116
rect 3476 1084 3480 1116
rect 3440 1036 3480 1084
rect 3440 1004 3444 1036
rect 3476 1004 3480 1036
rect 3440 956 3480 1004
rect 3440 924 3444 956
rect 3476 924 3480 956
rect 3440 920 3480 924
rect 3520 1676 3560 1680
rect 3520 1644 3524 1676
rect 3556 1644 3560 1676
rect 3520 1596 3560 1644
rect 3520 1564 3524 1596
rect 3556 1564 3560 1596
rect 3520 1516 3560 1564
rect 3520 1484 3524 1516
rect 3556 1484 3560 1516
rect 3520 1436 3560 1484
rect 3520 1404 3524 1436
rect 3556 1404 3560 1436
rect 3520 1356 3560 1404
rect 3520 1324 3524 1356
rect 3556 1324 3560 1356
rect 3520 1276 3560 1324
rect 3520 1244 3524 1276
rect 3556 1244 3560 1276
rect 3520 1196 3560 1244
rect 3520 1164 3524 1196
rect 3556 1164 3560 1196
rect 3520 1116 3560 1164
rect 3520 1084 3524 1116
rect 3556 1084 3560 1116
rect 3520 1036 3560 1084
rect 3520 1004 3524 1036
rect 3556 1004 3560 1036
rect 3520 956 3560 1004
rect 3520 924 3524 956
rect 3556 924 3560 956
rect 3520 920 3560 924
rect 3600 1676 3640 1680
rect 3600 1644 3604 1676
rect 3636 1644 3640 1676
rect 3600 1596 3640 1644
rect 3600 1564 3604 1596
rect 3636 1564 3640 1596
rect 3600 1516 3640 1564
rect 3600 1484 3604 1516
rect 3636 1484 3640 1516
rect 3600 1436 3640 1484
rect 3600 1404 3604 1436
rect 3636 1404 3640 1436
rect 3600 1356 3640 1404
rect 3600 1324 3604 1356
rect 3636 1324 3640 1356
rect 3600 1276 3640 1324
rect 3600 1244 3604 1276
rect 3636 1244 3640 1276
rect 3600 1196 3640 1244
rect 3600 1164 3604 1196
rect 3636 1164 3640 1196
rect 3600 1116 3640 1164
rect 3600 1084 3604 1116
rect 3636 1084 3640 1116
rect 3600 1036 3640 1084
rect 3600 1004 3604 1036
rect 3636 1004 3640 1036
rect 3600 956 3640 1004
rect 3600 924 3604 956
rect 3636 924 3640 956
rect 3600 920 3640 924
rect 3680 1676 3720 1680
rect 3680 1644 3684 1676
rect 3716 1644 3720 1676
rect 3680 1596 3720 1644
rect 3680 1564 3684 1596
rect 3716 1564 3720 1596
rect 3680 1516 3720 1564
rect 3680 1484 3684 1516
rect 3716 1484 3720 1516
rect 3680 1436 3720 1484
rect 3680 1404 3684 1436
rect 3716 1404 3720 1436
rect 3680 1356 3720 1404
rect 3680 1324 3684 1356
rect 3716 1324 3720 1356
rect 3680 1276 3720 1324
rect 3680 1244 3684 1276
rect 3716 1244 3720 1276
rect 3680 1196 3720 1244
rect 3680 1164 3684 1196
rect 3716 1164 3720 1196
rect 3680 1116 3720 1164
rect 3680 1084 3684 1116
rect 3716 1084 3720 1116
rect 3680 1036 3720 1084
rect 3680 1004 3684 1036
rect 3716 1004 3720 1036
rect 3680 956 3720 1004
rect 3680 924 3684 956
rect 3716 924 3720 956
rect 3680 920 3720 924
rect 3760 1676 3800 1680
rect 3760 1644 3764 1676
rect 3796 1644 3800 1676
rect 3760 1596 3800 1644
rect 3760 1564 3764 1596
rect 3796 1564 3800 1596
rect 3760 1516 3800 1564
rect 3760 1484 3764 1516
rect 3796 1484 3800 1516
rect 3760 1436 3800 1484
rect 3760 1404 3764 1436
rect 3796 1404 3800 1436
rect 3760 1356 3800 1404
rect 3760 1324 3764 1356
rect 3796 1324 3800 1356
rect 3760 1276 3800 1324
rect 3760 1244 3764 1276
rect 3796 1244 3800 1276
rect 3760 1196 3800 1244
rect 3760 1164 3764 1196
rect 3796 1164 3800 1196
rect 3760 1116 3800 1164
rect 3760 1084 3764 1116
rect 3796 1084 3800 1116
rect 3760 1036 3800 1084
rect 3760 1004 3764 1036
rect 3796 1004 3800 1036
rect 3760 956 3800 1004
rect 3760 924 3764 956
rect 3796 924 3800 956
rect 3760 920 3800 924
rect 3840 1676 3880 1680
rect 3840 1644 3844 1676
rect 3876 1644 3880 1676
rect 3840 1596 3880 1644
rect 3840 1564 3844 1596
rect 3876 1564 3880 1596
rect 3840 1516 3880 1564
rect 3840 1484 3844 1516
rect 3876 1484 3880 1516
rect 3840 1436 3880 1484
rect 3840 1404 3844 1436
rect 3876 1404 3880 1436
rect 3840 1356 3880 1404
rect 3840 1324 3844 1356
rect 3876 1324 3880 1356
rect 3840 1276 3880 1324
rect 3840 1244 3844 1276
rect 3876 1244 3880 1276
rect 3840 1196 3880 1244
rect 3840 1164 3844 1196
rect 3876 1164 3880 1196
rect 3840 1116 3880 1164
rect 3840 1084 3844 1116
rect 3876 1084 3880 1116
rect 3840 1036 3880 1084
rect 3840 1004 3844 1036
rect 3876 1004 3880 1036
rect 3840 956 3880 1004
rect 3840 924 3844 956
rect 3876 924 3880 956
rect 3840 920 3880 924
rect 3920 1676 3960 1680
rect 3920 1644 3924 1676
rect 3956 1644 3960 1676
rect 3920 1596 3960 1644
rect 3920 1564 3924 1596
rect 3956 1564 3960 1596
rect 3920 1516 3960 1564
rect 3920 1484 3924 1516
rect 3956 1484 3960 1516
rect 3920 1436 3960 1484
rect 3920 1404 3924 1436
rect 3956 1404 3960 1436
rect 3920 1356 3960 1404
rect 3920 1324 3924 1356
rect 3956 1324 3960 1356
rect 3920 1276 3960 1324
rect 3920 1244 3924 1276
rect 3956 1244 3960 1276
rect 3920 1196 3960 1244
rect 3920 1164 3924 1196
rect 3956 1164 3960 1196
rect 3920 1116 3960 1164
rect 3920 1084 3924 1116
rect 3956 1084 3960 1116
rect 3920 1036 3960 1084
rect 3920 1004 3924 1036
rect 3956 1004 3960 1036
rect 3920 956 3960 1004
rect 3920 924 3924 956
rect 3956 924 3960 956
rect 3920 920 3960 924
rect 4000 1676 4040 1680
rect 4000 1644 4004 1676
rect 4036 1644 4040 1676
rect 4000 1596 4040 1644
rect 4000 1564 4004 1596
rect 4036 1564 4040 1596
rect 4000 1516 4040 1564
rect 4000 1484 4004 1516
rect 4036 1484 4040 1516
rect 4000 1436 4040 1484
rect 4000 1404 4004 1436
rect 4036 1404 4040 1436
rect 4000 1356 4040 1404
rect 4000 1324 4004 1356
rect 4036 1324 4040 1356
rect 4000 1276 4040 1324
rect 4000 1244 4004 1276
rect 4036 1244 4040 1276
rect 4000 1196 4040 1244
rect 4000 1164 4004 1196
rect 4036 1164 4040 1196
rect 4000 1116 4040 1164
rect 4000 1084 4004 1116
rect 4036 1084 4040 1116
rect 4000 1036 4040 1084
rect 4000 1004 4004 1036
rect 4036 1004 4040 1036
rect 4000 956 4040 1004
rect 4000 924 4004 956
rect 4036 924 4040 956
rect 4000 920 4040 924
rect 4080 1676 4120 1680
rect 4080 1644 4084 1676
rect 4116 1644 4120 1676
rect 4080 1596 4120 1644
rect 4080 1564 4084 1596
rect 4116 1564 4120 1596
rect 4080 1516 4120 1564
rect 4080 1484 4084 1516
rect 4116 1484 4120 1516
rect 4080 1436 4120 1484
rect 4080 1404 4084 1436
rect 4116 1404 4120 1436
rect 4080 1356 4120 1404
rect 4080 1324 4084 1356
rect 4116 1324 4120 1356
rect 4080 1276 4120 1324
rect 4080 1244 4084 1276
rect 4116 1244 4120 1276
rect 4080 1196 4120 1244
rect 4080 1164 4084 1196
rect 4116 1164 4120 1196
rect 4080 1116 4120 1164
rect 4080 1084 4084 1116
rect 4116 1084 4120 1116
rect 4080 1036 4120 1084
rect 4080 1004 4084 1036
rect 4116 1004 4120 1036
rect 4080 956 4120 1004
rect 4080 924 4084 956
rect 4116 924 4120 956
rect 4080 920 4120 924
rect 4160 1676 4200 1680
rect 4160 1644 4164 1676
rect 4196 1644 4200 1676
rect 4160 1596 4200 1644
rect 4160 1564 4164 1596
rect 4196 1564 4200 1596
rect 4160 1516 4200 1564
rect 4160 1484 4164 1516
rect 4196 1484 4200 1516
rect 4160 1436 4200 1484
rect 4160 1404 4164 1436
rect 4196 1404 4200 1436
rect 4160 1356 4200 1404
rect 4160 1324 4164 1356
rect 4196 1324 4200 1356
rect 4160 1276 4200 1324
rect 4160 1244 4164 1276
rect 4196 1244 4200 1276
rect 4160 1196 4200 1244
rect 4160 1164 4164 1196
rect 4196 1164 4200 1196
rect 4160 1116 4200 1164
rect 4160 1084 4164 1116
rect 4196 1084 4200 1116
rect 4160 1036 4200 1084
rect 4160 1004 4164 1036
rect 4196 1004 4200 1036
rect 4160 956 4200 1004
rect 4160 924 4164 956
rect 4196 924 4200 956
rect 4160 920 4200 924
rect 4240 1676 4280 1680
rect 4240 1644 4244 1676
rect 4276 1644 4280 1676
rect 4240 1596 4280 1644
rect 4240 1564 4244 1596
rect 4276 1564 4280 1596
rect 4240 1516 4280 1564
rect 4240 1484 4244 1516
rect 4276 1484 4280 1516
rect 4240 1436 4280 1484
rect 4240 1404 4244 1436
rect 4276 1404 4280 1436
rect 4240 1356 4280 1404
rect 4240 1324 4244 1356
rect 4276 1324 4280 1356
rect 4240 1276 4280 1324
rect 4240 1244 4244 1276
rect 4276 1244 4280 1276
rect 4240 1196 4280 1244
rect 4240 1164 4244 1196
rect 4276 1164 4280 1196
rect 4240 1116 4280 1164
rect 4240 1084 4244 1116
rect 4276 1084 4280 1116
rect 4240 1036 4280 1084
rect 4240 1004 4244 1036
rect 4276 1004 4280 1036
rect 4240 956 4280 1004
rect 4240 924 4244 956
rect 4276 924 4280 956
rect 4240 920 4280 924
rect 4320 1676 4360 1680
rect 4320 1644 4324 1676
rect 4356 1644 4360 1676
rect 4320 1596 4360 1644
rect 4320 1564 4324 1596
rect 4356 1564 4360 1596
rect 4320 1516 4360 1564
rect 4320 1484 4324 1516
rect 4356 1484 4360 1516
rect 4320 1436 4360 1484
rect 4320 1404 4324 1436
rect 4356 1404 4360 1436
rect 4320 1356 4360 1404
rect 4320 1324 4324 1356
rect 4356 1324 4360 1356
rect 4320 1276 4360 1324
rect 4320 1244 4324 1276
rect 4356 1244 4360 1276
rect 4320 1196 4360 1244
rect 4320 1164 4324 1196
rect 4356 1164 4360 1196
rect 4320 1116 4360 1164
rect 4320 1084 4324 1116
rect 4356 1084 4360 1116
rect 4320 1036 4360 1084
rect 4320 1004 4324 1036
rect 4356 1004 4360 1036
rect 4320 956 4360 1004
rect 4320 924 4324 956
rect 4356 924 4360 956
rect 4320 920 4360 924
rect 4400 1676 4440 1680
rect 4400 1644 4404 1676
rect 4436 1644 4440 1676
rect 4400 1596 4440 1644
rect 4400 1564 4404 1596
rect 4436 1564 4440 1596
rect 4400 1516 4440 1564
rect 4400 1484 4404 1516
rect 4436 1484 4440 1516
rect 4400 1436 4440 1484
rect 4400 1404 4404 1436
rect 4436 1404 4440 1436
rect 4400 1356 4440 1404
rect 4400 1324 4404 1356
rect 4436 1324 4440 1356
rect 4400 1276 4440 1324
rect 4400 1244 4404 1276
rect 4436 1244 4440 1276
rect 4400 1196 4440 1244
rect 4400 1164 4404 1196
rect 4436 1164 4440 1196
rect 4400 1116 4440 1164
rect 4400 1084 4404 1116
rect 4436 1084 4440 1116
rect 4400 1036 4440 1084
rect 4400 1004 4404 1036
rect 4436 1004 4440 1036
rect 4400 956 4440 1004
rect 4400 924 4404 956
rect 4436 924 4440 956
rect 4400 920 4440 924
rect 4480 1676 4520 1680
rect 4480 1644 4484 1676
rect 4516 1644 4520 1676
rect 4480 1596 4520 1644
rect 4480 1564 4484 1596
rect 4516 1564 4520 1596
rect 4480 1516 4520 1564
rect 4480 1484 4484 1516
rect 4516 1484 4520 1516
rect 4480 1436 4520 1484
rect 4480 1404 4484 1436
rect 4516 1404 4520 1436
rect 4480 1356 4520 1404
rect 4480 1324 4484 1356
rect 4516 1324 4520 1356
rect 4480 1276 4520 1324
rect 4480 1244 4484 1276
rect 4516 1244 4520 1276
rect 4480 1196 4520 1244
rect 4480 1164 4484 1196
rect 4516 1164 4520 1196
rect 4480 1116 4520 1164
rect 4480 1084 4484 1116
rect 4516 1084 4520 1116
rect 4480 1036 4520 1084
rect 4480 1004 4484 1036
rect 4516 1004 4520 1036
rect 4480 956 4520 1004
rect 4480 924 4484 956
rect 4516 924 4520 956
rect 4480 920 4520 924
rect 4560 1676 4600 1680
rect 4560 1644 4564 1676
rect 4596 1644 4600 1676
rect 4560 1596 4600 1644
rect 4560 1564 4564 1596
rect 4596 1564 4600 1596
rect 4560 1516 4600 1564
rect 4560 1484 4564 1516
rect 4596 1484 4600 1516
rect 4560 1436 4600 1484
rect 4560 1404 4564 1436
rect 4596 1404 4600 1436
rect 4560 1356 4600 1404
rect 4560 1324 4564 1356
rect 4596 1324 4600 1356
rect 4560 1276 4600 1324
rect 4560 1244 4564 1276
rect 4596 1244 4600 1276
rect 4560 1196 4600 1244
rect 4560 1164 4564 1196
rect 4596 1164 4600 1196
rect 4560 1116 4600 1164
rect 4560 1084 4564 1116
rect 4596 1084 4600 1116
rect 4560 1036 4600 1084
rect 4560 1004 4564 1036
rect 4596 1004 4600 1036
rect 4560 956 4600 1004
rect 4560 924 4564 956
rect 4596 924 4600 956
rect 4560 920 4600 924
rect 4640 1676 4680 1680
rect 4640 1644 4644 1676
rect 4676 1644 4680 1676
rect 4640 1596 4680 1644
rect 4640 1564 4644 1596
rect 4676 1564 4680 1596
rect 4640 1516 4680 1564
rect 4640 1484 4644 1516
rect 4676 1484 4680 1516
rect 4640 1436 4680 1484
rect 4640 1404 4644 1436
rect 4676 1404 4680 1436
rect 4640 1356 4680 1404
rect 4640 1324 4644 1356
rect 4676 1324 4680 1356
rect 4640 1276 4680 1324
rect 4640 1244 4644 1276
rect 4676 1244 4680 1276
rect 4640 1196 4680 1244
rect 4640 1164 4644 1196
rect 4676 1164 4680 1196
rect 4640 1116 4680 1164
rect 4640 1084 4644 1116
rect 4676 1084 4680 1116
rect 4640 1036 4680 1084
rect 4640 1004 4644 1036
rect 4676 1004 4680 1036
rect 4640 956 4680 1004
rect 4640 924 4644 956
rect 4676 924 4680 956
rect 4640 920 4680 924
rect 4720 1676 4760 1680
rect 4720 1644 4724 1676
rect 4756 1644 4760 1676
rect 4720 1596 4760 1644
rect 4720 1564 4724 1596
rect 4756 1564 4760 1596
rect 4720 1516 4760 1564
rect 4720 1484 4724 1516
rect 4756 1484 4760 1516
rect 4720 1436 4760 1484
rect 4720 1404 4724 1436
rect 4756 1404 4760 1436
rect 4720 1356 4760 1404
rect 4720 1324 4724 1356
rect 4756 1324 4760 1356
rect 4720 1276 4760 1324
rect 4720 1244 4724 1276
rect 4756 1244 4760 1276
rect 4720 1196 4760 1244
rect 4720 1164 4724 1196
rect 4756 1164 4760 1196
rect 4720 1116 4760 1164
rect 4720 1084 4724 1116
rect 4756 1084 4760 1116
rect 4720 1036 4760 1084
rect 4720 1004 4724 1036
rect 4756 1004 4760 1036
rect 4720 956 4760 1004
rect 4720 924 4724 956
rect 4756 924 4760 956
rect 4720 920 4760 924
rect 4800 1676 4840 1680
rect 4800 1644 4804 1676
rect 4836 1644 4840 1676
rect 4800 1596 4840 1644
rect 4800 1564 4804 1596
rect 4836 1564 4840 1596
rect 4800 1516 4840 1564
rect 4800 1484 4804 1516
rect 4836 1484 4840 1516
rect 4800 1436 4840 1484
rect 4800 1404 4804 1436
rect 4836 1404 4840 1436
rect 4800 1356 4840 1404
rect 4800 1324 4804 1356
rect 4836 1324 4840 1356
rect 4800 1276 4840 1324
rect 4800 1244 4804 1276
rect 4836 1244 4840 1276
rect 4800 1196 4840 1244
rect 4800 1164 4804 1196
rect 4836 1164 4840 1196
rect 4800 1116 4840 1164
rect 4800 1084 4804 1116
rect 4836 1084 4840 1116
rect 4800 1036 4840 1084
rect 4800 1004 4804 1036
rect 4836 1004 4840 1036
rect 4800 956 4840 1004
rect 4800 924 4804 956
rect 4836 924 4840 956
rect 4800 920 4840 924
rect 4880 1676 4920 1724
rect 4880 1644 4884 1676
rect 4916 1644 4920 1676
rect 4880 1596 4920 1644
rect 4880 1564 4884 1596
rect 4916 1564 4920 1596
rect 4880 1516 4920 1564
rect 4880 1484 4884 1516
rect 4916 1484 4920 1516
rect 4880 1436 4920 1484
rect 4880 1404 4884 1436
rect 4916 1404 4920 1436
rect 4880 1356 4920 1404
rect 4880 1324 4884 1356
rect 4916 1324 4920 1356
rect 4880 1276 4920 1324
rect 4880 1244 4884 1276
rect 4916 1244 4920 1276
rect 4880 1196 4920 1244
rect 4880 1164 4884 1196
rect 4916 1164 4920 1196
rect 4880 1116 4920 1164
rect 4880 1084 4884 1116
rect 4916 1084 4920 1116
rect 4880 1036 4920 1084
rect 4880 1004 4884 1036
rect 4916 1004 4920 1036
rect 4880 956 4920 1004
rect 4880 924 4884 956
rect 4916 924 4920 956
rect -880 844 -876 876
rect -844 844 -840 876
rect -880 796 -840 844
rect -880 764 -876 796
rect -844 764 -840 796
rect -880 716 -840 764
rect -880 684 -876 716
rect -844 684 -840 716
rect -880 636 -840 684
rect -880 604 -876 636
rect -844 604 -840 636
rect -880 556 -840 604
rect -880 524 -876 556
rect -844 524 -840 556
rect -880 476 -840 524
rect -880 444 -876 476
rect -844 444 -840 476
rect -880 396 -840 444
rect -880 364 -876 396
rect -844 364 -840 396
rect -880 316 -840 364
rect -880 284 -876 316
rect -844 284 -840 316
rect -880 236 -840 284
rect -880 204 -876 236
rect -844 204 -840 236
rect -880 156 -840 204
rect -880 124 -876 156
rect -844 124 -840 156
rect -880 76 -840 124
rect -880 44 -876 76
rect -844 44 -840 76
rect -880 -4 -840 44
rect -880 -36 -876 -4
rect -844 -36 -840 -4
rect -880 -84 -840 -36
rect -880 -116 -876 -84
rect -844 -116 -840 -84
rect -880 -120 -840 -116
rect -800 876 -760 880
rect -800 844 -796 876
rect -764 844 -760 876
rect -800 796 -760 844
rect -800 764 -796 796
rect -764 764 -760 796
rect -800 716 -760 764
rect -800 684 -796 716
rect -764 684 -760 716
rect -800 636 -760 684
rect -800 604 -796 636
rect -764 604 -760 636
rect -800 556 -760 604
rect -800 524 -796 556
rect -764 524 -760 556
rect -800 476 -760 524
rect -800 444 -796 476
rect -764 444 -760 476
rect -800 396 -760 444
rect -800 364 -796 396
rect -764 364 -760 396
rect -800 316 -760 364
rect -800 284 -796 316
rect -764 284 -760 316
rect -800 236 -760 284
rect -800 204 -796 236
rect -764 204 -760 236
rect -800 156 -760 204
rect -800 124 -796 156
rect -764 124 -760 156
rect -800 76 -760 124
rect -800 44 -796 76
rect -764 44 -760 76
rect -800 -4 -760 44
rect -800 -36 -796 -4
rect -764 -36 -760 -4
rect -800 -84 -760 -36
rect -800 -116 -796 -84
rect -764 -116 -760 -84
rect -800 -120 -760 -116
rect -720 876 -680 880
rect -720 844 -716 876
rect -684 844 -680 876
rect -720 796 -680 844
rect -720 764 -716 796
rect -684 764 -680 796
rect -720 716 -680 764
rect -720 684 -716 716
rect -684 684 -680 716
rect -720 636 -680 684
rect -720 604 -716 636
rect -684 604 -680 636
rect -720 556 -680 604
rect -720 524 -716 556
rect -684 524 -680 556
rect -720 476 -680 524
rect -720 444 -716 476
rect -684 444 -680 476
rect -720 396 -680 444
rect -720 364 -716 396
rect -684 364 -680 396
rect -720 316 -680 364
rect -720 284 -716 316
rect -684 284 -680 316
rect -720 236 -680 284
rect -720 204 -716 236
rect -684 204 -680 236
rect -720 156 -680 204
rect -720 124 -716 156
rect -684 124 -680 156
rect -720 76 -680 124
rect -720 44 -716 76
rect -684 44 -680 76
rect -720 -4 -680 44
rect -720 -36 -716 -4
rect -684 -36 -680 -4
rect -720 -84 -680 -36
rect -720 -116 -716 -84
rect -684 -116 -680 -84
rect -720 -120 -680 -116
rect -640 876 -600 880
rect -640 844 -636 876
rect -604 844 -600 876
rect -640 796 -600 844
rect -640 764 -636 796
rect -604 764 -600 796
rect -640 716 -600 764
rect -640 684 -636 716
rect -604 684 -600 716
rect -640 636 -600 684
rect -640 604 -636 636
rect -604 604 -600 636
rect -640 556 -600 604
rect -640 524 -636 556
rect -604 524 -600 556
rect -640 476 -600 524
rect -640 444 -636 476
rect -604 444 -600 476
rect -640 396 -600 444
rect -640 364 -636 396
rect -604 364 -600 396
rect -640 316 -600 364
rect -640 284 -636 316
rect -604 284 -600 316
rect -640 236 -600 284
rect -640 204 -636 236
rect -604 204 -600 236
rect -640 156 -600 204
rect -640 124 -636 156
rect -604 124 -600 156
rect -640 76 -600 124
rect -640 44 -636 76
rect -604 44 -600 76
rect -640 -4 -600 44
rect -640 -36 -636 -4
rect -604 -36 -600 -4
rect -640 -84 -600 -36
rect -640 -116 -636 -84
rect -604 -116 -600 -84
rect -640 -120 -600 -116
rect -560 876 -520 880
rect -560 844 -556 876
rect -524 844 -520 876
rect -560 796 -520 844
rect -560 764 -556 796
rect -524 764 -520 796
rect -560 716 -520 764
rect -560 684 -556 716
rect -524 684 -520 716
rect -560 636 -520 684
rect -560 604 -556 636
rect -524 604 -520 636
rect -560 556 -520 604
rect -560 524 -556 556
rect -524 524 -520 556
rect -560 476 -520 524
rect -560 444 -556 476
rect -524 444 -520 476
rect -560 396 -520 444
rect -560 364 -556 396
rect -524 364 -520 396
rect -560 316 -520 364
rect -560 284 -556 316
rect -524 284 -520 316
rect -560 236 -520 284
rect -560 204 -556 236
rect -524 204 -520 236
rect -560 156 -520 204
rect -560 124 -556 156
rect -524 124 -520 156
rect -560 76 -520 124
rect -560 44 -556 76
rect -524 44 -520 76
rect -560 -4 -520 44
rect -560 -36 -556 -4
rect -524 -36 -520 -4
rect -560 -84 -520 -36
rect -560 -116 -556 -84
rect -524 -116 -520 -84
rect -560 -120 -520 -116
rect -480 876 -440 880
rect -480 844 -476 876
rect -444 844 -440 876
rect -480 796 -440 844
rect -480 764 -476 796
rect -444 764 -440 796
rect -480 716 -440 764
rect -480 684 -476 716
rect -444 684 -440 716
rect -480 636 -440 684
rect -480 604 -476 636
rect -444 604 -440 636
rect -480 556 -440 604
rect -480 524 -476 556
rect -444 524 -440 556
rect -480 476 -440 524
rect -480 444 -476 476
rect -444 444 -440 476
rect -480 396 -440 444
rect -480 364 -476 396
rect -444 364 -440 396
rect -480 316 -440 364
rect -480 284 -476 316
rect -444 284 -440 316
rect -480 236 -440 284
rect -480 204 -476 236
rect -444 204 -440 236
rect -480 156 -440 204
rect -480 124 -476 156
rect -444 124 -440 156
rect -480 76 -440 124
rect -480 44 -476 76
rect -444 44 -440 76
rect -480 -4 -440 44
rect -480 -36 -476 -4
rect -444 -36 -440 -4
rect -480 -84 -440 -36
rect -480 -116 -476 -84
rect -444 -116 -440 -84
rect -480 -120 -440 -116
rect -400 876 -360 880
rect -400 844 -396 876
rect -364 844 -360 876
rect -400 796 -360 844
rect -400 764 -396 796
rect -364 764 -360 796
rect -400 716 -360 764
rect -400 684 -396 716
rect -364 684 -360 716
rect -400 636 -360 684
rect -400 604 -396 636
rect -364 604 -360 636
rect -400 556 -360 604
rect -400 524 -396 556
rect -364 524 -360 556
rect -400 476 -360 524
rect -400 444 -396 476
rect -364 444 -360 476
rect -400 396 -360 444
rect -400 364 -396 396
rect -364 364 -360 396
rect -400 316 -360 364
rect -400 284 -396 316
rect -364 284 -360 316
rect -400 236 -360 284
rect -400 204 -396 236
rect -364 204 -360 236
rect -400 156 -360 204
rect -400 124 -396 156
rect -364 124 -360 156
rect -400 76 -360 124
rect -400 44 -396 76
rect -364 44 -360 76
rect -400 -4 -360 44
rect -400 -36 -396 -4
rect -364 -36 -360 -4
rect -400 -84 -360 -36
rect -400 -116 -396 -84
rect -364 -116 -360 -84
rect -400 -120 -360 -116
rect -320 876 -280 880
rect -320 844 -316 876
rect -284 844 -280 876
rect -320 796 -280 844
rect -320 764 -316 796
rect -284 764 -280 796
rect -320 716 -280 764
rect -320 684 -316 716
rect -284 684 -280 716
rect -320 636 -280 684
rect -320 604 -316 636
rect -284 604 -280 636
rect -320 556 -280 604
rect -320 524 -316 556
rect -284 524 -280 556
rect -320 476 -280 524
rect -320 444 -316 476
rect -284 444 -280 476
rect -320 396 -280 444
rect -320 364 -316 396
rect -284 364 -280 396
rect -320 316 -280 364
rect -320 284 -316 316
rect -284 284 -280 316
rect -320 236 -280 284
rect -320 204 -316 236
rect -284 204 -280 236
rect -320 156 -280 204
rect -320 124 -316 156
rect -284 124 -280 156
rect -320 76 -280 124
rect -320 44 -316 76
rect -284 44 -280 76
rect -320 -4 -280 44
rect -320 -36 -316 -4
rect -284 -36 -280 -4
rect -320 -84 -280 -36
rect -320 -116 -316 -84
rect -284 -116 -280 -84
rect -320 -120 -280 -116
rect -240 876 -200 880
rect -240 844 -236 876
rect -204 844 -200 876
rect -240 796 -200 844
rect -240 764 -236 796
rect -204 764 -200 796
rect -240 716 -200 764
rect -240 684 -236 716
rect -204 684 -200 716
rect -240 636 -200 684
rect -240 604 -236 636
rect -204 604 -200 636
rect -240 556 -200 604
rect -240 524 -236 556
rect -204 524 -200 556
rect -240 476 -200 524
rect -240 444 -236 476
rect -204 444 -200 476
rect -240 396 -200 444
rect -240 364 -236 396
rect -204 364 -200 396
rect -240 316 -200 364
rect -240 284 -236 316
rect -204 284 -200 316
rect -240 236 -200 284
rect -240 204 -236 236
rect -204 204 -200 236
rect -240 156 -200 204
rect -240 124 -236 156
rect -204 124 -200 156
rect -240 76 -200 124
rect -240 44 -236 76
rect -204 44 -200 76
rect -240 -4 -200 44
rect -240 -36 -236 -4
rect -204 -36 -200 -4
rect -240 -84 -200 -36
rect -240 -116 -236 -84
rect -204 -116 -200 -84
rect -240 -120 -200 -116
rect -160 876 -120 880
rect -160 844 -156 876
rect -124 844 -120 876
rect -160 796 -120 844
rect -160 764 -156 796
rect -124 764 -120 796
rect -160 716 -120 764
rect -160 684 -156 716
rect -124 684 -120 716
rect -160 636 -120 684
rect -160 604 -156 636
rect -124 604 -120 636
rect -160 556 -120 604
rect -160 524 -156 556
rect -124 524 -120 556
rect -160 476 -120 524
rect -160 444 -156 476
rect -124 444 -120 476
rect -160 396 -120 444
rect -160 364 -156 396
rect -124 364 -120 396
rect -160 316 -120 364
rect -160 284 -156 316
rect -124 284 -120 316
rect -160 236 -120 284
rect -160 204 -156 236
rect -124 204 -120 236
rect -160 156 -120 204
rect -160 124 -156 156
rect -124 124 -120 156
rect -160 76 -120 124
rect -160 44 -156 76
rect -124 44 -120 76
rect -160 -4 -120 44
rect -160 -36 -156 -4
rect -124 -36 -120 -4
rect -160 -84 -120 -36
rect -160 -116 -156 -84
rect -124 -116 -120 -84
rect -160 -120 -120 -116
rect -80 876 -40 880
rect -80 844 -76 876
rect -44 844 -40 876
rect -80 796 -40 844
rect -80 764 -76 796
rect -44 764 -40 796
rect -80 716 -40 764
rect -80 684 -76 716
rect -44 684 -40 716
rect -80 636 -40 684
rect -80 604 -76 636
rect -44 604 -40 636
rect -80 556 -40 604
rect -80 524 -76 556
rect -44 524 -40 556
rect -80 476 -40 524
rect -80 444 -76 476
rect -44 444 -40 476
rect -80 396 -40 444
rect -80 364 -76 396
rect -44 364 -40 396
rect -80 316 -40 364
rect -80 284 -76 316
rect -44 284 -40 316
rect -80 236 -40 284
rect -80 204 -76 236
rect -44 204 -40 236
rect -80 156 -40 204
rect -80 124 -76 156
rect -44 124 -40 156
rect -80 76 -40 124
rect -80 44 -76 76
rect -44 44 -40 76
rect -80 -4 -40 44
rect -80 -36 -76 -4
rect -44 -36 -40 -4
rect -80 -84 -40 -36
rect -80 -116 -76 -84
rect -44 -116 -40 -84
rect -80 -120 -40 -116
rect 0 876 40 880
rect 0 844 4 876
rect 36 844 40 876
rect 0 796 40 844
rect 0 764 4 796
rect 36 764 40 796
rect 0 716 40 764
rect 0 684 4 716
rect 36 684 40 716
rect 0 636 40 684
rect 0 604 4 636
rect 36 604 40 636
rect 0 556 40 604
rect 0 524 4 556
rect 36 524 40 556
rect 0 476 40 524
rect 0 444 4 476
rect 36 444 40 476
rect 0 396 40 444
rect 0 364 4 396
rect 36 364 40 396
rect 0 316 40 364
rect 0 284 4 316
rect 36 284 40 316
rect 0 236 40 284
rect 0 204 4 236
rect 36 204 40 236
rect 0 156 40 204
rect 0 124 4 156
rect 36 124 40 156
rect 0 76 40 124
rect 0 44 4 76
rect 36 44 40 76
rect 0 -4 40 44
rect 0 -36 4 -4
rect 36 -36 40 -4
rect 0 -84 40 -36
rect 0 -116 4 -84
rect 36 -116 40 -84
rect 0 -120 40 -116
rect 80 876 120 880
rect 80 844 84 876
rect 116 844 120 876
rect 80 796 120 844
rect 80 764 84 796
rect 116 764 120 796
rect 80 716 120 764
rect 80 684 84 716
rect 116 684 120 716
rect 80 636 120 684
rect 80 604 84 636
rect 116 604 120 636
rect 80 556 120 604
rect 80 524 84 556
rect 116 524 120 556
rect 80 476 120 524
rect 80 444 84 476
rect 116 444 120 476
rect 80 396 120 444
rect 80 364 84 396
rect 116 364 120 396
rect 80 316 120 364
rect 80 284 84 316
rect 116 284 120 316
rect 80 236 120 284
rect 80 204 84 236
rect 116 204 120 236
rect 80 156 120 204
rect 80 124 84 156
rect 116 124 120 156
rect 80 76 120 124
rect 80 44 84 76
rect 116 44 120 76
rect 80 -4 120 44
rect 80 -36 84 -4
rect 116 -36 120 -4
rect 80 -84 120 -36
rect 80 -116 84 -84
rect 116 -116 120 -84
rect 80 -120 120 -116
rect 160 876 200 880
rect 160 844 164 876
rect 196 844 200 876
rect 160 796 200 844
rect 160 764 164 796
rect 196 764 200 796
rect 160 716 200 764
rect 160 684 164 716
rect 196 684 200 716
rect 160 636 200 684
rect 160 604 164 636
rect 196 604 200 636
rect 160 556 200 604
rect 160 524 164 556
rect 196 524 200 556
rect 160 476 200 524
rect 160 444 164 476
rect 196 444 200 476
rect 160 396 200 444
rect 160 364 164 396
rect 196 364 200 396
rect 160 316 200 364
rect 160 284 164 316
rect 196 284 200 316
rect 160 236 200 284
rect 160 204 164 236
rect 196 204 200 236
rect 160 156 200 204
rect 160 124 164 156
rect 196 124 200 156
rect 160 76 200 124
rect 160 44 164 76
rect 196 44 200 76
rect 160 -4 200 44
rect 160 -36 164 -4
rect 196 -36 200 -4
rect 160 -84 200 -36
rect 160 -116 164 -84
rect 196 -116 200 -84
rect 160 -120 200 -116
rect 240 876 280 880
rect 240 844 244 876
rect 276 844 280 876
rect 240 796 280 844
rect 240 764 244 796
rect 276 764 280 796
rect 240 716 280 764
rect 240 684 244 716
rect 276 684 280 716
rect 240 636 280 684
rect 240 604 244 636
rect 276 604 280 636
rect 240 556 280 604
rect 240 524 244 556
rect 276 524 280 556
rect 240 476 280 524
rect 240 444 244 476
rect 276 444 280 476
rect 240 396 280 444
rect 240 364 244 396
rect 276 364 280 396
rect 240 316 280 364
rect 240 284 244 316
rect 276 284 280 316
rect 240 236 280 284
rect 240 204 244 236
rect 276 204 280 236
rect 240 156 280 204
rect 240 124 244 156
rect 276 124 280 156
rect 240 76 280 124
rect 240 44 244 76
rect 276 44 280 76
rect 240 -4 280 44
rect 240 -36 244 -4
rect 276 -36 280 -4
rect 240 -84 280 -36
rect 240 -116 244 -84
rect 276 -116 280 -84
rect 240 -120 280 -116
rect 320 876 360 880
rect 320 844 324 876
rect 356 844 360 876
rect 320 796 360 844
rect 320 764 324 796
rect 356 764 360 796
rect 320 716 360 764
rect 320 684 324 716
rect 356 684 360 716
rect 320 636 360 684
rect 320 604 324 636
rect 356 604 360 636
rect 320 556 360 604
rect 320 524 324 556
rect 356 524 360 556
rect 320 476 360 524
rect 320 444 324 476
rect 356 444 360 476
rect 320 396 360 444
rect 320 364 324 396
rect 356 364 360 396
rect 320 316 360 364
rect 320 284 324 316
rect 356 284 360 316
rect 320 236 360 284
rect 320 204 324 236
rect 356 204 360 236
rect 320 156 360 204
rect 320 124 324 156
rect 356 124 360 156
rect 320 76 360 124
rect 320 44 324 76
rect 356 44 360 76
rect 320 -4 360 44
rect 320 -36 324 -4
rect 356 -36 360 -4
rect 320 -84 360 -36
rect 320 -116 324 -84
rect 356 -116 360 -84
rect 320 -120 360 -116
rect 400 876 440 880
rect 400 844 404 876
rect 436 844 440 876
rect 400 796 440 844
rect 400 764 404 796
rect 436 764 440 796
rect 400 716 440 764
rect 400 684 404 716
rect 436 684 440 716
rect 400 636 440 684
rect 400 604 404 636
rect 436 604 440 636
rect 400 556 440 604
rect 400 524 404 556
rect 436 524 440 556
rect 400 476 440 524
rect 400 444 404 476
rect 436 444 440 476
rect 400 396 440 444
rect 400 364 404 396
rect 436 364 440 396
rect 400 316 440 364
rect 400 284 404 316
rect 436 284 440 316
rect 400 236 440 284
rect 400 204 404 236
rect 436 204 440 236
rect 400 156 440 204
rect 400 124 404 156
rect 436 124 440 156
rect 400 76 440 124
rect 400 44 404 76
rect 436 44 440 76
rect 400 -4 440 44
rect 400 -36 404 -4
rect 436 -36 440 -4
rect 400 -84 440 -36
rect 400 -116 404 -84
rect 436 -116 440 -84
rect 400 -120 440 -116
rect 480 876 520 880
rect 480 844 484 876
rect 516 844 520 876
rect 480 796 520 844
rect 480 764 484 796
rect 516 764 520 796
rect 480 716 520 764
rect 480 684 484 716
rect 516 684 520 716
rect 480 636 520 684
rect 480 604 484 636
rect 516 604 520 636
rect 480 556 520 604
rect 480 524 484 556
rect 516 524 520 556
rect 480 476 520 524
rect 480 444 484 476
rect 516 444 520 476
rect 480 396 520 444
rect 480 364 484 396
rect 516 364 520 396
rect 480 316 520 364
rect 480 284 484 316
rect 516 284 520 316
rect 480 236 520 284
rect 480 204 484 236
rect 516 204 520 236
rect 480 156 520 204
rect 480 124 484 156
rect 516 124 520 156
rect 480 76 520 124
rect 480 44 484 76
rect 516 44 520 76
rect 480 -4 520 44
rect 480 -36 484 -4
rect 516 -36 520 -4
rect 480 -84 520 -36
rect 480 -116 484 -84
rect 516 -116 520 -84
rect 480 -120 520 -116
rect 560 876 600 880
rect 560 844 564 876
rect 596 844 600 876
rect 560 796 600 844
rect 560 764 564 796
rect 596 764 600 796
rect 560 716 600 764
rect 560 684 564 716
rect 596 684 600 716
rect 560 636 600 684
rect 560 604 564 636
rect 596 604 600 636
rect 560 556 600 604
rect 560 524 564 556
rect 596 524 600 556
rect 560 476 600 524
rect 560 444 564 476
rect 596 444 600 476
rect 560 396 600 444
rect 560 364 564 396
rect 596 364 600 396
rect 560 316 600 364
rect 560 284 564 316
rect 596 284 600 316
rect 560 236 600 284
rect 560 204 564 236
rect 596 204 600 236
rect 560 156 600 204
rect 560 124 564 156
rect 596 124 600 156
rect 560 76 600 124
rect 560 44 564 76
rect 596 44 600 76
rect 560 -4 600 44
rect 560 -36 564 -4
rect 596 -36 600 -4
rect 560 -84 600 -36
rect 560 -116 564 -84
rect 596 -116 600 -84
rect 560 -120 600 -116
rect 640 876 680 880
rect 640 844 644 876
rect 676 844 680 876
rect 640 796 680 844
rect 640 764 644 796
rect 676 764 680 796
rect 640 716 680 764
rect 640 684 644 716
rect 676 684 680 716
rect 640 636 680 684
rect 640 604 644 636
rect 676 604 680 636
rect 640 556 680 604
rect 640 524 644 556
rect 676 524 680 556
rect 640 476 680 524
rect 640 444 644 476
rect 676 444 680 476
rect 640 396 680 444
rect 640 364 644 396
rect 676 364 680 396
rect 640 316 680 364
rect 640 284 644 316
rect 676 284 680 316
rect 640 236 680 284
rect 640 204 644 236
rect 676 204 680 236
rect 640 156 680 204
rect 640 124 644 156
rect 676 124 680 156
rect 640 76 680 124
rect 640 44 644 76
rect 676 44 680 76
rect 640 -4 680 44
rect 640 -36 644 -4
rect 676 -36 680 -4
rect 640 -84 680 -36
rect 640 -116 644 -84
rect 676 -116 680 -84
rect 640 -120 680 -116
rect 720 876 760 880
rect 720 844 724 876
rect 756 844 760 876
rect 720 796 760 844
rect 720 764 724 796
rect 756 764 760 796
rect 720 716 760 764
rect 720 684 724 716
rect 756 684 760 716
rect 720 636 760 684
rect 720 604 724 636
rect 756 604 760 636
rect 720 556 760 604
rect 720 524 724 556
rect 756 524 760 556
rect 720 476 760 524
rect 720 444 724 476
rect 756 444 760 476
rect 720 396 760 444
rect 720 364 724 396
rect 756 364 760 396
rect 720 316 760 364
rect 720 284 724 316
rect 756 284 760 316
rect 720 236 760 284
rect 720 204 724 236
rect 756 204 760 236
rect 720 156 760 204
rect 720 124 724 156
rect 756 124 760 156
rect 720 76 760 124
rect 720 44 724 76
rect 756 44 760 76
rect 720 -4 760 44
rect 720 -36 724 -4
rect 756 -36 760 -4
rect 720 -84 760 -36
rect 720 -116 724 -84
rect 756 -116 760 -84
rect 720 -120 760 -116
rect 800 876 840 880
rect 800 844 804 876
rect 836 844 840 876
rect 800 796 840 844
rect 800 764 804 796
rect 836 764 840 796
rect 800 716 840 764
rect 800 684 804 716
rect 836 684 840 716
rect 800 636 840 684
rect 800 604 804 636
rect 836 604 840 636
rect 800 556 840 604
rect 800 524 804 556
rect 836 524 840 556
rect 800 476 840 524
rect 800 444 804 476
rect 836 444 840 476
rect 800 396 840 444
rect 800 364 804 396
rect 836 364 840 396
rect 800 316 840 364
rect 800 284 804 316
rect 836 284 840 316
rect 800 236 840 284
rect 800 204 804 236
rect 836 204 840 236
rect 800 156 840 204
rect 800 124 804 156
rect 836 124 840 156
rect 800 76 840 124
rect 800 44 804 76
rect 836 44 840 76
rect 800 -4 840 44
rect 800 -36 804 -4
rect 836 -36 840 -4
rect 800 -84 840 -36
rect 800 -116 804 -84
rect 836 -116 840 -84
rect 800 -120 840 -116
rect 880 876 920 880
rect 880 844 884 876
rect 916 844 920 876
rect 880 796 920 844
rect 880 764 884 796
rect 916 764 920 796
rect 880 716 920 764
rect 880 684 884 716
rect 916 684 920 716
rect 880 636 920 684
rect 880 604 884 636
rect 916 604 920 636
rect 880 556 920 604
rect 880 524 884 556
rect 916 524 920 556
rect 880 476 920 524
rect 880 444 884 476
rect 916 444 920 476
rect 880 396 920 444
rect 880 364 884 396
rect 916 364 920 396
rect 880 316 920 364
rect 880 284 884 316
rect 916 284 920 316
rect 880 236 920 284
rect 880 204 884 236
rect 916 204 920 236
rect 880 156 920 204
rect 880 124 884 156
rect 916 124 920 156
rect 880 76 920 124
rect 880 44 884 76
rect 916 44 920 76
rect 880 -4 920 44
rect 880 -36 884 -4
rect 916 -36 920 -4
rect 880 -84 920 -36
rect 880 -116 884 -84
rect 916 -116 920 -84
rect 880 -120 920 -116
rect 960 876 1000 880
rect 960 844 964 876
rect 996 844 1000 876
rect 960 796 1000 844
rect 960 764 964 796
rect 996 764 1000 796
rect 960 716 1000 764
rect 960 684 964 716
rect 996 684 1000 716
rect 960 636 1000 684
rect 960 604 964 636
rect 996 604 1000 636
rect 960 556 1000 604
rect 960 524 964 556
rect 996 524 1000 556
rect 960 476 1000 524
rect 960 444 964 476
rect 996 444 1000 476
rect 960 396 1000 444
rect 960 364 964 396
rect 996 364 1000 396
rect 960 316 1000 364
rect 960 284 964 316
rect 996 284 1000 316
rect 960 236 1000 284
rect 960 204 964 236
rect 996 204 1000 236
rect 960 156 1000 204
rect 960 124 964 156
rect 996 124 1000 156
rect 960 76 1000 124
rect 960 44 964 76
rect 996 44 1000 76
rect 960 -4 1000 44
rect 960 -36 964 -4
rect 996 -36 1000 -4
rect 960 -84 1000 -36
rect 960 -116 964 -84
rect 996 -116 1000 -84
rect 960 -120 1000 -116
rect 1040 876 1080 880
rect 1040 844 1044 876
rect 1076 844 1080 876
rect 1040 796 1080 844
rect 1040 764 1044 796
rect 1076 764 1080 796
rect 1040 716 1080 764
rect 1040 684 1044 716
rect 1076 684 1080 716
rect 1040 636 1080 684
rect 1040 604 1044 636
rect 1076 604 1080 636
rect 1040 556 1080 604
rect 1040 524 1044 556
rect 1076 524 1080 556
rect 1040 476 1080 524
rect 1040 444 1044 476
rect 1076 444 1080 476
rect 1040 396 1080 444
rect 1040 364 1044 396
rect 1076 364 1080 396
rect 1040 316 1080 364
rect 1040 284 1044 316
rect 1076 284 1080 316
rect 1040 236 1080 284
rect 1040 204 1044 236
rect 1076 204 1080 236
rect 1040 156 1080 204
rect 1040 124 1044 156
rect 1076 124 1080 156
rect 1040 76 1080 124
rect 1040 44 1044 76
rect 1076 44 1080 76
rect 1040 -4 1080 44
rect 1040 -36 1044 -4
rect 1076 -36 1080 -4
rect 1040 -84 1080 -36
rect 1040 -116 1044 -84
rect 1076 -116 1080 -84
rect 1040 -120 1080 -116
rect 1120 876 1160 880
rect 1120 844 1124 876
rect 1156 844 1160 876
rect 1120 796 1160 844
rect 1120 764 1124 796
rect 1156 764 1160 796
rect 1120 716 1160 764
rect 1120 684 1124 716
rect 1156 684 1160 716
rect 1120 636 1160 684
rect 1120 604 1124 636
rect 1156 604 1160 636
rect 1120 556 1160 604
rect 1120 524 1124 556
rect 1156 524 1160 556
rect 1120 476 1160 524
rect 1120 444 1124 476
rect 1156 444 1160 476
rect 1120 396 1160 444
rect 1120 364 1124 396
rect 1156 364 1160 396
rect 1120 316 1160 364
rect 1120 284 1124 316
rect 1156 284 1160 316
rect 1120 236 1160 284
rect 1120 204 1124 236
rect 1156 204 1160 236
rect 1120 156 1160 204
rect 1120 124 1124 156
rect 1156 124 1160 156
rect 1120 76 1160 124
rect 1120 44 1124 76
rect 1156 44 1160 76
rect 1120 -4 1160 44
rect 1120 -36 1124 -4
rect 1156 -36 1160 -4
rect 1120 -84 1160 -36
rect 1120 -116 1124 -84
rect 1156 -116 1160 -84
rect 1120 -120 1160 -116
rect 1200 876 1240 880
rect 1200 844 1204 876
rect 1236 844 1240 876
rect 1200 796 1240 844
rect 1200 764 1204 796
rect 1236 764 1240 796
rect 1200 716 1240 764
rect 1200 684 1204 716
rect 1236 684 1240 716
rect 1200 636 1240 684
rect 1200 604 1204 636
rect 1236 604 1240 636
rect 1200 556 1240 604
rect 1200 524 1204 556
rect 1236 524 1240 556
rect 1200 476 1240 524
rect 1200 444 1204 476
rect 1236 444 1240 476
rect 1200 396 1240 444
rect 1200 364 1204 396
rect 1236 364 1240 396
rect 1200 316 1240 364
rect 1200 284 1204 316
rect 1236 284 1240 316
rect 1200 236 1240 284
rect 1200 204 1204 236
rect 1236 204 1240 236
rect 1200 156 1240 204
rect 1200 124 1204 156
rect 1236 124 1240 156
rect 1200 76 1240 124
rect 1200 44 1204 76
rect 1236 44 1240 76
rect 1200 -4 1240 44
rect 1200 -36 1204 -4
rect 1236 -36 1240 -4
rect 1200 -84 1240 -36
rect 1200 -116 1204 -84
rect 1236 -116 1240 -84
rect 1200 -120 1240 -116
rect 1280 876 1320 880
rect 1280 844 1284 876
rect 1316 844 1320 876
rect 1280 796 1320 844
rect 1280 764 1284 796
rect 1316 764 1320 796
rect 1280 716 1320 764
rect 1280 684 1284 716
rect 1316 684 1320 716
rect 1280 636 1320 684
rect 1280 604 1284 636
rect 1316 604 1320 636
rect 1280 556 1320 604
rect 1280 524 1284 556
rect 1316 524 1320 556
rect 1280 476 1320 524
rect 1280 444 1284 476
rect 1316 444 1320 476
rect 1280 396 1320 444
rect 1280 364 1284 396
rect 1316 364 1320 396
rect 1280 316 1320 364
rect 1280 284 1284 316
rect 1316 284 1320 316
rect 1280 236 1320 284
rect 1280 204 1284 236
rect 1316 204 1320 236
rect 1280 156 1320 204
rect 1280 124 1284 156
rect 1316 124 1320 156
rect 1280 76 1320 124
rect 1280 44 1284 76
rect 1316 44 1320 76
rect 1280 -4 1320 44
rect 1280 -36 1284 -4
rect 1316 -36 1320 -4
rect 1280 -84 1320 -36
rect 1280 -116 1284 -84
rect 1316 -116 1320 -84
rect 1280 -120 1320 -116
rect 1360 876 1400 880
rect 1360 844 1364 876
rect 1396 844 1400 876
rect 1360 796 1400 844
rect 1360 764 1364 796
rect 1396 764 1400 796
rect 1360 716 1400 764
rect 1360 684 1364 716
rect 1396 684 1400 716
rect 1360 636 1400 684
rect 1360 604 1364 636
rect 1396 604 1400 636
rect 1360 556 1400 604
rect 1360 524 1364 556
rect 1396 524 1400 556
rect 1360 476 1400 524
rect 1360 444 1364 476
rect 1396 444 1400 476
rect 1360 396 1400 444
rect 1360 364 1364 396
rect 1396 364 1400 396
rect 1360 316 1400 364
rect 1360 284 1364 316
rect 1396 284 1400 316
rect 1360 236 1400 284
rect 1360 204 1364 236
rect 1396 204 1400 236
rect 1360 156 1400 204
rect 1360 124 1364 156
rect 1396 124 1400 156
rect 1360 76 1400 124
rect 1360 44 1364 76
rect 1396 44 1400 76
rect 1360 -4 1400 44
rect 1360 -36 1364 -4
rect 1396 -36 1400 -4
rect 1360 -84 1400 -36
rect 1360 -116 1364 -84
rect 1396 -116 1400 -84
rect 1360 -120 1400 -116
rect 1440 876 1480 880
rect 1440 844 1444 876
rect 1476 844 1480 876
rect 1440 796 1480 844
rect 1440 764 1444 796
rect 1476 764 1480 796
rect 1440 716 1480 764
rect 1440 684 1444 716
rect 1476 684 1480 716
rect 1440 636 1480 684
rect 1440 604 1444 636
rect 1476 604 1480 636
rect 1440 556 1480 604
rect 1440 524 1444 556
rect 1476 524 1480 556
rect 1440 476 1480 524
rect 1440 444 1444 476
rect 1476 444 1480 476
rect 1440 396 1480 444
rect 1440 364 1444 396
rect 1476 364 1480 396
rect 1440 316 1480 364
rect 1440 284 1444 316
rect 1476 284 1480 316
rect 1440 236 1480 284
rect 1440 204 1444 236
rect 1476 204 1480 236
rect 1440 156 1480 204
rect 1440 124 1444 156
rect 1476 124 1480 156
rect 1440 76 1480 124
rect 1440 44 1444 76
rect 1476 44 1480 76
rect 1440 -4 1480 44
rect 1440 -36 1444 -4
rect 1476 -36 1480 -4
rect 1440 -84 1480 -36
rect 1440 -116 1444 -84
rect 1476 -116 1480 -84
rect 1440 -120 1480 -116
rect 1520 876 1560 880
rect 1520 844 1524 876
rect 1556 844 1560 876
rect 1520 796 1560 844
rect 1520 764 1524 796
rect 1556 764 1560 796
rect 1520 716 1560 764
rect 1520 684 1524 716
rect 1556 684 1560 716
rect 1520 636 1560 684
rect 1520 604 1524 636
rect 1556 604 1560 636
rect 1520 556 1560 604
rect 1520 524 1524 556
rect 1556 524 1560 556
rect 1520 476 1560 524
rect 1520 444 1524 476
rect 1556 444 1560 476
rect 1520 396 1560 444
rect 1520 364 1524 396
rect 1556 364 1560 396
rect 1520 316 1560 364
rect 1520 284 1524 316
rect 1556 284 1560 316
rect 1520 236 1560 284
rect 1520 204 1524 236
rect 1556 204 1560 236
rect 1520 156 1560 204
rect 1520 124 1524 156
rect 1556 124 1560 156
rect 1520 76 1560 124
rect 1520 44 1524 76
rect 1556 44 1560 76
rect 1520 -4 1560 44
rect 1520 -36 1524 -4
rect 1556 -36 1560 -4
rect 1520 -84 1560 -36
rect 1520 -116 1524 -84
rect 1556 -116 1560 -84
rect 1520 -120 1560 -116
rect 1600 876 1640 880
rect 1600 844 1604 876
rect 1636 844 1640 876
rect 1600 796 1640 844
rect 1600 764 1604 796
rect 1636 764 1640 796
rect 1600 716 1640 764
rect 1600 684 1604 716
rect 1636 684 1640 716
rect 1600 636 1640 684
rect 1600 604 1604 636
rect 1636 604 1640 636
rect 1600 556 1640 604
rect 1600 524 1604 556
rect 1636 524 1640 556
rect 1600 476 1640 524
rect 1600 444 1604 476
rect 1636 444 1640 476
rect 1600 396 1640 444
rect 1600 364 1604 396
rect 1636 364 1640 396
rect 1600 316 1640 364
rect 1600 284 1604 316
rect 1636 284 1640 316
rect 1600 236 1640 284
rect 1600 204 1604 236
rect 1636 204 1640 236
rect 1600 156 1640 204
rect 1600 124 1604 156
rect 1636 124 1640 156
rect 1600 76 1640 124
rect 1600 44 1604 76
rect 1636 44 1640 76
rect 1600 -4 1640 44
rect 1600 -36 1604 -4
rect 1636 -36 1640 -4
rect 1600 -84 1640 -36
rect 1600 -116 1604 -84
rect 1636 -116 1640 -84
rect 1600 -120 1640 -116
rect 1680 876 1720 880
rect 1680 844 1684 876
rect 1716 844 1720 876
rect 1680 796 1720 844
rect 1680 764 1684 796
rect 1716 764 1720 796
rect 1680 716 1720 764
rect 1680 684 1684 716
rect 1716 684 1720 716
rect 1680 636 1720 684
rect 1680 604 1684 636
rect 1716 604 1720 636
rect 1680 556 1720 604
rect 1680 524 1684 556
rect 1716 524 1720 556
rect 1680 476 1720 524
rect 1680 444 1684 476
rect 1716 444 1720 476
rect 1680 396 1720 444
rect 1680 364 1684 396
rect 1716 364 1720 396
rect 1680 316 1720 364
rect 1680 284 1684 316
rect 1716 284 1720 316
rect 1680 236 1720 284
rect 1680 204 1684 236
rect 1716 204 1720 236
rect 1680 156 1720 204
rect 1680 124 1684 156
rect 1716 124 1720 156
rect 1680 76 1720 124
rect 1680 44 1684 76
rect 1716 44 1720 76
rect 1680 -4 1720 44
rect 1680 -36 1684 -4
rect 1716 -36 1720 -4
rect 1680 -84 1720 -36
rect 1680 -116 1684 -84
rect 1716 -116 1720 -84
rect 1680 -120 1720 -116
rect 1760 876 1800 880
rect 1760 844 1764 876
rect 1796 844 1800 876
rect 1760 796 1800 844
rect 1760 764 1764 796
rect 1796 764 1800 796
rect 1760 716 1800 764
rect 1760 684 1764 716
rect 1796 684 1800 716
rect 1760 636 1800 684
rect 1760 604 1764 636
rect 1796 604 1800 636
rect 1760 556 1800 604
rect 1760 524 1764 556
rect 1796 524 1800 556
rect 1760 476 1800 524
rect 1760 444 1764 476
rect 1796 444 1800 476
rect 1760 396 1800 444
rect 1760 364 1764 396
rect 1796 364 1800 396
rect 1760 316 1800 364
rect 1760 284 1764 316
rect 1796 284 1800 316
rect 1760 236 1800 284
rect 1760 204 1764 236
rect 1796 204 1800 236
rect 1760 156 1800 204
rect 1760 124 1764 156
rect 1796 124 1800 156
rect 1760 76 1800 124
rect 1760 44 1764 76
rect 1796 44 1800 76
rect 1760 -4 1800 44
rect 1760 -36 1764 -4
rect 1796 -36 1800 -4
rect 1760 -84 1800 -36
rect 1760 -116 1764 -84
rect 1796 -116 1800 -84
rect 1760 -120 1800 -116
rect 1840 876 1880 880
rect 1840 844 1844 876
rect 1876 844 1880 876
rect 1840 796 1880 844
rect 1840 764 1844 796
rect 1876 764 1880 796
rect 1840 716 1880 764
rect 1840 684 1844 716
rect 1876 684 1880 716
rect 1840 636 1880 684
rect 1840 604 1844 636
rect 1876 604 1880 636
rect 1840 556 1880 604
rect 1840 524 1844 556
rect 1876 524 1880 556
rect 1840 476 1880 524
rect 1840 444 1844 476
rect 1876 444 1880 476
rect 1840 396 1880 444
rect 1840 364 1844 396
rect 1876 364 1880 396
rect 1840 316 1880 364
rect 1840 284 1844 316
rect 1876 284 1880 316
rect 1840 236 1880 284
rect 1840 204 1844 236
rect 1876 204 1880 236
rect 1840 156 1880 204
rect 1840 124 1844 156
rect 1876 124 1880 156
rect 1840 76 1880 124
rect 1840 44 1844 76
rect 1876 44 1880 76
rect 1840 -4 1880 44
rect 1840 -36 1844 -4
rect 1876 -36 1880 -4
rect 1840 -84 1880 -36
rect 1840 -116 1844 -84
rect 1876 -116 1880 -84
rect 1840 -120 1880 -116
rect 1920 876 1960 880
rect 1920 844 1924 876
rect 1956 844 1960 876
rect 1920 796 1960 844
rect 1920 764 1924 796
rect 1956 764 1960 796
rect 1920 716 1960 764
rect 1920 684 1924 716
rect 1956 684 1960 716
rect 1920 636 1960 684
rect 1920 604 1924 636
rect 1956 604 1960 636
rect 1920 556 1960 604
rect 1920 524 1924 556
rect 1956 524 1960 556
rect 1920 476 1960 524
rect 1920 444 1924 476
rect 1956 444 1960 476
rect 1920 396 1960 444
rect 1920 364 1924 396
rect 1956 364 1960 396
rect 1920 316 1960 364
rect 1920 284 1924 316
rect 1956 284 1960 316
rect 1920 236 1960 284
rect 1920 204 1924 236
rect 1956 204 1960 236
rect 1920 156 1960 204
rect 1920 124 1924 156
rect 1956 124 1960 156
rect 1920 76 1960 124
rect 1920 44 1924 76
rect 1956 44 1960 76
rect 1920 -4 1960 44
rect 1920 -36 1924 -4
rect 1956 -36 1960 -4
rect 1920 -84 1960 -36
rect 1920 -116 1924 -84
rect 1956 -116 1960 -84
rect 1920 -120 1960 -116
rect 2000 876 2040 880
rect 2000 844 2004 876
rect 2036 844 2040 876
rect 2000 796 2040 844
rect 2000 764 2004 796
rect 2036 764 2040 796
rect 2000 716 2040 764
rect 2000 684 2004 716
rect 2036 684 2040 716
rect 2000 636 2040 684
rect 2000 604 2004 636
rect 2036 604 2040 636
rect 2000 556 2040 604
rect 2000 524 2004 556
rect 2036 524 2040 556
rect 2000 476 2040 524
rect 2000 444 2004 476
rect 2036 444 2040 476
rect 2000 396 2040 444
rect 2000 364 2004 396
rect 2036 364 2040 396
rect 2000 316 2040 364
rect 2000 284 2004 316
rect 2036 284 2040 316
rect 2000 236 2040 284
rect 2000 204 2004 236
rect 2036 204 2040 236
rect 2000 156 2040 204
rect 2000 124 2004 156
rect 2036 124 2040 156
rect 2000 76 2040 124
rect 2000 44 2004 76
rect 2036 44 2040 76
rect 2000 -4 2040 44
rect 2000 -36 2004 -4
rect 2036 -36 2040 -4
rect 2000 -84 2040 -36
rect 2000 -116 2004 -84
rect 2036 -116 2040 -84
rect 2000 -120 2040 -116
rect 2080 876 2120 880
rect 2080 844 2084 876
rect 2116 844 2120 876
rect 2080 796 2120 844
rect 2080 764 2084 796
rect 2116 764 2120 796
rect 2080 716 2120 764
rect 2080 684 2084 716
rect 2116 684 2120 716
rect 2080 636 2120 684
rect 2080 604 2084 636
rect 2116 604 2120 636
rect 2080 556 2120 604
rect 2080 524 2084 556
rect 2116 524 2120 556
rect 2080 476 2120 524
rect 2080 444 2084 476
rect 2116 444 2120 476
rect 2080 396 2120 444
rect 2080 364 2084 396
rect 2116 364 2120 396
rect 2080 316 2120 364
rect 2080 284 2084 316
rect 2116 284 2120 316
rect 2080 236 2120 284
rect 2080 204 2084 236
rect 2116 204 2120 236
rect 2080 156 2120 204
rect 2080 124 2084 156
rect 2116 124 2120 156
rect 2080 76 2120 124
rect 2080 44 2084 76
rect 2116 44 2120 76
rect 2080 -4 2120 44
rect 2080 -36 2084 -4
rect 2116 -36 2120 -4
rect 2080 -84 2120 -36
rect 2080 -116 2084 -84
rect 2116 -116 2120 -84
rect 2080 -120 2120 -116
rect 2160 876 2200 880
rect 2160 844 2164 876
rect 2196 844 2200 876
rect 2160 796 2200 844
rect 2160 764 2164 796
rect 2196 764 2200 796
rect 2160 716 2200 764
rect 2160 684 2164 716
rect 2196 684 2200 716
rect 2160 636 2200 684
rect 2160 604 2164 636
rect 2196 604 2200 636
rect 2160 556 2200 604
rect 2160 524 2164 556
rect 2196 524 2200 556
rect 2160 476 2200 524
rect 2160 444 2164 476
rect 2196 444 2200 476
rect 2160 396 2200 444
rect 2160 364 2164 396
rect 2196 364 2200 396
rect 2160 316 2200 364
rect 2160 284 2164 316
rect 2196 284 2200 316
rect 2160 236 2200 284
rect 2160 204 2164 236
rect 2196 204 2200 236
rect 2160 156 2200 204
rect 2160 124 2164 156
rect 2196 124 2200 156
rect 2160 76 2200 124
rect 2160 44 2164 76
rect 2196 44 2200 76
rect 2160 -4 2200 44
rect 2160 -36 2164 -4
rect 2196 -36 2200 -4
rect 2160 -84 2200 -36
rect 2160 -116 2164 -84
rect 2196 -116 2200 -84
rect 2160 -120 2200 -116
rect 2240 876 2280 880
rect 2240 844 2244 876
rect 2276 844 2280 876
rect 2240 796 2280 844
rect 2240 764 2244 796
rect 2276 764 2280 796
rect 2240 716 2280 764
rect 2240 684 2244 716
rect 2276 684 2280 716
rect 2240 636 2280 684
rect 2240 604 2244 636
rect 2276 604 2280 636
rect 2240 556 2280 604
rect 2240 524 2244 556
rect 2276 524 2280 556
rect 2240 476 2280 524
rect 2240 444 2244 476
rect 2276 444 2280 476
rect 2240 396 2280 444
rect 2240 364 2244 396
rect 2276 364 2280 396
rect 2240 316 2280 364
rect 2240 284 2244 316
rect 2276 284 2280 316
rect 2240 236 2280 284
rect 2240 204 2244 236
rect 2276 204 2280 236
rect 2240 156 2280 204
rect 2240 124 2244 156
rect 2276 124 2280 156
rect 2240 76 2280 124
rect 2240 44 2244 76
rect 2276 44 2280 76
rect 2240 -4 2280 44
rect 2240 -36 2244 -4
rect 2276 -36 2280 -4
rect 2240 -84 2280 -36
rect 2240 -116 2244 -84
rect 2276 -116 2280 -84
rect 2240 -120 2280 -116
rect 2320 876 2360 880
rect 2320 844 2324 876
rect 2356 844 2360 876
rect 2320 796 2360 844
rect 2320 764 2324 796
rect 2356 764 2360 796
rect 2320 716 2360 764
rect 2320 684 2324 716
rect 2356 684 2360 716
rect 2320 636 2360 684
rect 2320 604 2324 636
rect 2356 604 2360 636
rect 2320 556 2360 604
rect 2320 524 2324 556
rect 2356 524 2360 556
rect 2320 476 2360 524
rect 2320 444 2324 476
rect 2356 444 2360 476
rect 2320 396 2360 444
rect 2320 364 2324 396
rect 2356 364 2360 396
rect 2320 316 2360 364
rect 2320 284 2324 316
rect 2356 284 2360 316
rect 2320 236 2360 284
rect 2320 204 2324 236
rect 2356 204 2360 236
rect 2320 156 2360 204
rect 2320 124 2324 156
rect 2356 124 2360 156
rect 2320 76 2360 124
rect 2320 44 2324 76
rect 2356 44 2360 76
rect 2320 -4 2360 44
rect 2320 -36 2324 -4
rect 2356 -36 2360 -4
rect 2320 -84 2360 -36
rect 2320 -116 2324 -84
rect 2356 -116 2360 -84
rect 2320 -120 2360 -116
rect 2400 876 2440 880
rect 2400 844 2404 876
rect 2436 844 2440 876
rect 2400 796 2440 844
rect 2400 764 2404 796
rect 2436 764 2440 796
rect 2400 716 2440 764
rect 2400 684 2404 716
rect 2436 684 2440 716
rect 2400 636 2440 684
rect 2400 604 2404 636
rect 2436 604 2440 636
rect 2400 556 2440 604
rect 2400 524 2404 556
rect 2436 524 2440 556
rect 2400 476 2440 524
rect 2400 444 2404 476
rect 2436 444 2440 476
rect 2400 396 2440 444
rect 2400 364 2404 396
rect 2436 364 2440 396
rect 2400 316 2440 364
rect 2400 284 2404 316
rect 2436 284 2440 316
rect 2400 236 2440 284
rect 2400 204 2404 236
rect 2436 204 2440 236
rect 2400 156 2440 204
rect 2400 124 2404 156
rect 2436 124 2440 156
rect 2400 76 2440 124
rect 2400 44 2404 76
rect 2436 44 2440 76
rect 2400 -4 2440 44
rect 2400 -36 2404 -4
rect 2436 -36 2440 -4
rect 2400 -84 2440 -36
rect 2400 -116 2404 -84
rect 2436 -116 2440 -84
rect 2400 -120 2440 -116
rect 2480 876 2520 880
rect 2480 844 2484 876
rect 2516 844 2520 876
rect 2480 796 2520 844
rect 2480 764 2484 796
rect 2516 764 2520 796
rect 2480 716 2520 764
rect 2480 684 2484 716
rect 2516 684 2520 716
rect 2480 636 2520 684
rect 2480 604 2484 636
rect 2516 604 2520 636
rect 2480 556 2520 604
rect 2480 524 2484 556
rect 2516 524 2520 556
rect 2480 476 2520 524
rect 2480 444 2484 476
rect 2516 444 2520 476
rect 2480 396 2520 444
rect 2480 364 2484 396
rect 2516 364 2520 396
rect 2480 316 2520 364
rect 2480 284 2484 316
rect 2516 284 2520 316
rect 2480 236 2520 284
rect 2480 204 2484 236
rect 2516 204 2520 236
rect 2480 156 2520 204
rect 2480 124 2484 156
rect 2516 124 2520 156
rect 2480 76 2520 124
rect 2480 44 2484 76
rect 2516 44 2520 76
rect 2480 -4 2520 44
rect 2480 -36 2484 -4
rect 2516 -36 2520 -4
rect 2480 -84 2520 -36
rect 2480 -116 2484 -84
rect 2516 -116 2520 -84
rect 2480 -120 2520 -116
rect 2560 876 2600 880
rect 2560 844 2564 876
rect 2596 844 2600 876
rect 2560 796 2600 844
rect 2560 764 2564 796
rect 2596 764 2600 796
rect 2560 716 2600 764
rect 2560 684 2564 716
rect 2596 684 2600 716
rect 2560 636 2600 684
rect 2560 604 2564 636
rect 2596 604 2600 636
rect 2560 556 2600 604
rect 2560 524 2564 556
rect 2596 524 2600 556
rect 2560 476 2600 524
rect 2560 444 2564 476
rect 2596 444 2600 476
rect 2560 396 2600 444
rect 2560 364 2564 396
rect 2596 364 2600 396
rect 2560 316 2600 364
rect 2560 284 2564 316
rect 2596 284 2600 316
rect 2560 236 2600 284
rect 2560 204 2564 236
rect 2596 204 2600 236
rect 2560 156 2600 204
rect 2560 124 2564 156
rect 2596 124 2600 156
rect 2560 76 2600 124
rect 2560 44 2564 76
rect 2596 44 2600 76
rect 2560 -4 2600 44
rect 2560 -36 2564 -4
rect 2596 -36 2600 -4
rect 2560 -84 2600 -36
rect 2560 -116 2564 -84
rect 2596 -116 2600 -84
rect 2560 -120 2600 -116
rect 2640 876 2680 880
rect 2640 844 2644 876
rect 2676 844 2680 876
rect 2640 796 2680 844
rect 2640 764 2644 796
rect 2676 764 2680 796
rect 2640 716 2680 764
rect 2640 684 2644 716
rect 2676 684 2680 716
rect 2640 636 2680 684
rect 2640 604 2644 636
rect 2676 604 2680 636
rect 2640 556 2680 604
rect 2640 524 2644 556
rect 2676 524 2680 556
rect 2640 476 2680 524
rect 2640 444 2644 476
rect 2676 444 2680 476
rect 2640 396 2680 444
rect 2640 364 2644 396
rect 2676 364 2680 396
rect 2640 316 2680 364
rect 2640 284 2644 316
rect 2676 284 2680 316
rect 2640 236 2680 284
rect 2640 204 2644 236
rect 2676 204 2680 236
rect 2640 156 2680 204
rect 2640 124 2644 156
rect 2676 124 2680 156
rect 2640 76 2680 124
rect 2640 44 2644 76
rect 2676 44 2680 76
rect 2640 -4 2680 44
rect 2640 -36 2644 -4
rect 2676 -36 2680 -4
rect 2640 -84 2680 -36
rect 2640 -116 2644 -84
rect 2676 -116 2680 -84
rect 2640 -120 2680 -116
rect 2720 876 2760 880
rect 2720 844 2724 876
rect 2756 844 2760 876
rect 2720 796 2760 844
rect 2720 764 2724 796
rect 2756 764 2760 796
rect 2720 716 2760 764
rect 2720 684 2724 716
rect 2756 684 2760 716
rect 2720 636 2760 684
rect 2720 604 2724 636
rect 2756 604 2760 636
rect 2720 556 2760 604
rect 2720 524 2724 556
rect 2756 524 2760 556
rect 2720 476 2760 524
rect 2720 444 2724 476
rect 2756 444 2760 476
rect 2720 396 2760 444
rect 2720 364 2724 396
rect 2756 364 2760 396
rect 2720 316 2760 364
rect 2720 284 2724 316
rect 2756 284 2760 316
rect 2720 236 2760 284
rect 2720 204 2724 236
rect 2756 204 2760 236
rect 2720 156 2760 204
rect 2720 124 2724 156
rect 2756 124 2760 156
rect 2720 76 2760 124
rect 2720 44 2724 76
rect 2756 44 2760 76
rect 2720 -4 2760 44
rect 2720 -36 2724 -4
rect 2756 -36 2760 -4
rect 2720 -84 2760 -36
rect 2720 -116 2724 -84
rect 2756 -116 2760 -84
rect 2720 -120 2760 -116
rect 2800 876 2840 880
rect 2800 844 2804 876
rect 2836 844 2840 876
rect 2800 796 2840 844
rect 2800 764 2804 796
rect 2836 764 2840 796
rect 2800 716 2840 764
rect 2800 684 2804 716
rect 2836 684 2840 716
rect 2800 636 2840 684
rect 2800 604 2804 636
rect 2836 604 2840 636
rect 2800 556 2840 604
rect 2800 524 2804 556
rect 2836 524 2840 556
rect 2800 476 2840 524
rect 2800 444 2804 476
rect 2836 444 2840 476
rect 2800 396 2840 444
rect 2800 364 2804 396
rect 2836 364 2840 396
rect 2800 316 2840 364
rect 2800 284 2804 316
rect 2836 284 2840 316
rect 2800 236 2840 284
rect 2800 204 2804 236
rect 2836 204 2840 236
rect 2800 156 2840 204
rect 2800 124 2804 156
rect 2836 124 2840 156
rect 2800 76 2840 124
rect 2800 44 2804 76
rect 2836 44 2840 76
rect 2800 -4 2840 44
rect 2800 -36 2804 -4
rect 2836 -36 2840 -4
rect 2800 -84 2840 -36
rect 2800 -116 2804 -84
rect 2836 -116 2840 -84
rect 2800 -120 2840 -116
rect 2880 876 2920 880
rect 2880 844 2884 876
rect 2916 844 2920 876
rect 2880 796 2920 844
rect 2880 764 2884 796
rect 2916 764 2920 796
rect 2880 716 2920 764
rect 2880 684 2884 716
rect 2916 684 2920 716
rect 2880 636 2920 684
rect 2880 604 2884 636
rect 2916 604 2920 636
rect 2880 556 2920 604
rect 2880 524 2884 556
rect 2916 524 2920 556
rect 2880 476 2920 524
rect 2880 444 2884 476
rect 2916 444 2920 476
rect 2880 396 2920 444
rect 2880 364 2884 396
rect 2916 364 2920 396
rect 2880 316 2920 364
rect 2880 284 2884 316
rect 2916 284 2920 316
rect 2880 236 2920 284
rect 2880 204 2884 236
rect 2916 204 2920 236
rect 2880 156 2920 204
rect 2880 124 2884 156
rect 2916 124 2920 156
rect 2880 76 2920 124
rect 2880 44 2884 76
rect 2916 44 2920 76
rect 2880 -4 2920 44
rect 2880 -36 2884 -4
rect 2916 -36 2920 -4
rect 2880 -84 2920 -36
rect 2880 -116 2884 -84
rect 2916 -116 2920 -84
rect 2880 -120 2920 -116
rect 2960 876 3000 880
rect 2960 844 2964 876
rect 2996 844 3000 876
rect 2960 796 3000 844
rect 2960 764 2964 796
rect 2996 764 3000 796
rect 2960 716 3000 764
rect 2960 684 2964 716
rect 2996 684 3000 716
rect 2960 636 3000 684
rect 2960 604 2964 636
rect 2996 604 3000 636
rect 2960 556 3000 604
rect 2960 524 2964 556
rect 2996 524 3000 556
rect 2960 476 3000 524
rect 2960 444 2964 476
rect 2996 444 3000 476
rect 2960 396 3000 444
rect 2960 364 2964 396
rect 2996 364 3000 396
rect 2960 316 3000 364
rect 2960 284 2964 316
rect 2996 284 3000 316
rect 2960 236 3000 284
rect 2960 204 2964 236
rect 2996 204 3000 236
rect 2960 156 3000 204
rect 2960 124 2964 156
rect 2996 124 3000 156
rect 2960 76 3000 124
rect 2960 44 2964 76
rect 2996 44 3000 76
rect 2960 -4 3000 44
rect 2960 -36 2964 -4
rect 2996 -36 3000 -4
rect 2960 -84 3000 -36
rect 2960 -116 2964 -84
rect 2996 -116 3000 -84
rect 2960 -120 3000 -116
rect 3040 876 3080 880
rect 3040 844 3044 876
rect 3076 844 3080 876
rect 3040 796 3080 844
rect 3040 764 3044 796
rect 3076 764 3080 796
rect 3040 716 3080 764
rect 3040 684 3044 716
rect 3076 684 3080 716
rect 3040 636 3080 684
rect 3040 604 3044 636
rect 3076 604 3080 636
rect 3040 556 3080 604
rect 3040 524 3044 556
rect 3076 524 3080 556
rect 3040 476 3080 524
rect 3040 444 3044 476
rect 3076 444 3080 476
rect 3040 396 3080 444
rect 3040 364 3044 396
rect 3076 364 3080 396
rect 3040 316 3080 364
rect 3040 284 3044 316
rect 3076 284 3080 316
rect 3040 236 3080 284
rect 3040 204 3044 236
rect 3076 204 3080 236
rect 3040 156 3080 204
rect 3040 124 3044 156
rect 3076 124 3080 156
rect 3040 76 3080 124
rect 3040 44 3044 76
rect 3076 44 3080 76
rect 3040 -4 3080 44
rect 3040 -36 3044 -4
rect 3076 -36 3080 -4
rect 3040 -84 3080 -36
rect 3040 -116 3044 -84
rect 3076 -116 3080 -84
rect 3040 -120 3080 -116
rect 3120 876 3160 880
rect 3120 844 3124 876
rect 3156 844 3160 876
rect 3120 796 3160 844
rect 3120 764 3124 796
rect 3156 764 3160 796
rect 3120 716 3160 764
rect 3120 684 3124 716
rect 3156 684 3160 716
rect 3120 636 3160 684
rect 3120 604 3124 636
rect 3156 604 3160 636
rect 3120 556 3160 604
rect 3120 524 3124 556
rect 3156 524 3160 556
rect 3120 476 3160 524
rect 3120 444 3124 476
rect 3156 444 3160 476
rect 3120 396 3160 444
rect 3120 364 3124 396
rect 3156 364 3160 396
rect 3120 316 3160 364
rect 3120 284 3124 316
rect 3156 284 3160 316
rect 3120 236 3160 284
rect 3120 204 3124 236
rect 3156 204 3160 236
rect 3120 156 3160 204
rect 3120 124 3124 156
rect 3156 124 3160 156
rect 3120 76 3160 124
rect 3120 44 3124 76
rect 3156 44 3160 76
rect 3120 -4 3160 44
rect 3120 -36 3124 -4
rect 3156 -36 3160 -4
rect 3120 -84 3160 -36
rect 3120 -116 3124 -84
rect 3156 -116 3160 -84
rect 3120 -120 3160 -116
rect 3200 876 3240 880
rect 3200 844 3204 876
rect 3236 844 3240 876
rect 3200 796 3240 844
rect 3200 764 3204 796
rect 3236 764 3240 796
rect 3200 716 3240 764
rect 3200 684 3204 716
rect 3236 684 3240 716
rect 3200 636 3240 684
rect 3200 604 3204 636
rect 3236 604 3240 636
rect 3200 556 3240 604
rect 3200 524 3204 556
rect 3236 524 3240 556
rect 3200 476 3240 524
rect 3200 444 3204 476
rect 3236 444 3240 476
rect 3200 396 3240 444
rect 3200 364 3204 396
rect 3236 364 3240 396
rect 3200 316 3240 364
rect 3200 284 3204 316
rect 3236 284 3240 316
rect 3200 236 3240 284
rect 3200 204 3204 236
rect 3236 204 3240 236
rect 3200 156 3240 204
rect 3200 124 3204 156
rect 3236 124 3240 156
rect 3200 76 3240 124
rect 3200 44 3204 76
rect 3236 44 3240 76
rect 3200 -4 3240 44
rect 3200 -36 3204 -4
rect 3236 -36 3240 -4
rect 3200 -84 3240 -36
rect 3200 -116 3204 -84
rect 3236 -116 3240 -84
rect 3200 -120 3240 -116
rect 3280 876 3320 880
rect 3280 844 3284 876
rect 3316 844 3320 876
rect 3280 796 3320 844
rect 3280 764 3284 796
rect 3316 764 3320 796
rect 3280 716 3320 764
rect 3280 684 3284 716
rect 3316 684 3320 716
rect 3280 636 3320 684
rect 3280 604 3284 636
rect 3316 604 3320 636
rect 3280 556 3320 604
rect 3280 524 3284 556
rect 3316 524 3320 556
rect 3280 476 3320 524
rect 3280 444 3284 476
rect 3316 444 3320 476
rect 3280 396 3320 444
rect 3280 364 3284 396
rect 3316 364 3320 396
rect 3280 316 3320 364
rect 3280 284 3284 316
rect 3316 284 3320 316
rect 3280 236 3320 284
rect 3280 204 3284 236
rect 3316 204 3320 236
rect 3280 156 3320 204
rect 3280 124 3284 156
rect 3316 124 3320 156
rect 3280 76 3320 124
rect 3280 44 3284 76
rect 3316 44 3320 76
rect 3280 -4 3320 44
rect 3280 -36 3284 -4
rect 3316 -36 3320 -4
rect 3280 -84 3320 -36
rect 3280 -116 3284 -84
rect 3316 -116 3320 -84
rect 3280 -120 3320 -116
rect 3360 876 3400 880
rect 3360 844 3364 876
rect 3396 844 3400 876
rect 3360 796 3400 844
rect 3360 764 3364 796
rect 3396 764 3400 796
rect 3360 716 3400 764
rect 3360 684 3364 716
rect 3396 684 3400 716
rect 3360 636 3400 684
rect 3360 604 3364 636
rect 3396 604 3400 636
rect 3360 556 3400 604
rect 3360 524 3364 556
rect 3396 524 3400 556
rect 3360 476 3400 524
rect 3360 444 3364 476
rect 3396 444 3400 476
rect 3360 396 3400 444
rect 3360 364 3364 396
rect 3396 364 3400 396
rect 3360 316 3400 364
rect 3360 284 3364 316
rect 3396 284 3400 316
rect 3360 236 3400 284
rect 3360 204 3364 236
rect 3396 204 3400 236
rect 3360 156 3400 204
rect 3360 124 3364 156
rect 3396 124 3400 156
rect 3360 76 3400 124
rect 3360 44 3364 76
rect 3396 44 3400 76
rect 3360 -4 3400 44
rect 3360 -36 3364 -4
rect 3396 -36 3400 -4
rect 3360 -84 3400 -36
rect 3360 -116 3364 -84
rect 3396 -116 3400 -84
rect 3360 -120 3400 -116
rect 3440 876 3480 880
rect 3440 844 3444 876
rect 3476 844 3480 876
rect 3440 796 3480 844
rect 3440 764 3444 796
rect 3476 764 3480 796
rect 3440 716 3480 764
rect 3440 684 3444 716
rect 3476 684 3480 716
rect 3440 636 3480 684
rect 3440 604 3444 636
rect 3476 604 3480 636
rect 3440 556 3480 604
rect 3440 524 3444 556
rect 3476 524 3480 556
rect 3440 476 3480 524
rect 3440 444 3444 476
rect 3476 444 3480 476
rect 3440 396 3480 444
rect 3440 364 3444 396
rect 3476 364 3480 396
rect 3440 316 3480 364
rect 3440 284 3444 316
rect 3476 284 3480 316
rect 3440 236 3480 284
rect 3440 204 3444 236
rect 3476 204 3480 236
rect 3440 156 3480 204
rect 3440 124 3444 156
rect 3476 124 3480 156
rect 3440 76 3480 124
rect 3440 44 3444 76
rect 3476 44 3480 76
rect 3440 -4 3480 44
rect 3440 -36 3444 -4
rect 3476 -36 3480 -4
rect 3440 -84 3480 -36
rect 3440 -116 3444 -84
rect 3476 -116 3480 -84
rect 3440 -120 3480 -116
rect 3520 876 3560 880
rect 3520 844 3524 876
rect 3556 844 3560 876
rect 3520 796 3560 844
rect 3520 764 3524 796
rect 3556 764 3560 796
rect 3520 716 3560 764
rect 3520 684 3524 716
rect 3556 684 3560 716
rect 3520 636 3560 684
rect 3520 604 3524 636
rect 3556 604 3560 636
rect 3520 556 3560 604
rect 3520 524 3524 556
rect 3556 524 3560 556
rect 3520 476 3560 524
rect 3520 444 3524 476
rect 3556 444 3560 476
rect 3520 396 3560 444
rect 3520 364 3524 396
rect 3556 364 3560 396
rect 3520 316 3560 364
rect 3520 284 3524 316
rect 3556 284 3560 316
rect 3520 236 3560 284
rect 3520 204 3524 236
rect 3556 204 3560 236
rect 3520 156 3560 204
rect 3520 124 3524 156
rect 3556 124 3560 156
rect 3520 76 3560 124
rect 3520 44 3524 76
rect 3556 44 3560 76
rect 3520 -4 3560 44
rect 3520 -36 3524 -4
rect 3556 -36 3560 -4
rect 3520 -84 3560 -36
rect 3520 -116 3524 -84
rect 3556 -116 3560 -84
rect 3520 -120 3560 -116
rect 3600 876 3640 880
rect 3600 844 3604 876
rect 3636 844 3640 876
rect 3600 796 3640 844
rect 3600 764 3604 796
rect 3636 764 3640 796
rect 3600 716 3640 764
rect 3600 684 3604 716
rect 3636 684 3640 716
rect 3600 636 3640 684
rect 3600 604 3604 636
rect 3636 604 3640 636
rect 3600 556 3640 604
rect 3600 524 3604 556
rect 3636 524 3640 556
rect 3600 476 3640 524
rect 3600 444 3604 476
rect 3636 444 3640 476
rect 3600 396 3640 444
rect 3600 364 3604 396
rect 3636 364 3640 396
rect 3600 316 3640 364
rect 3600 284 3604 316
rect 3636 284 3640 316
rect 3600 236 3640 284
rect 3600 204 3604 236
rect 3636 204 3640 236
rect 3600 156 3640 204
rect 3600 124 3604 156
rect 3636 124 3640 156
rect 3600 76 3640 124
rect 3600 44 3604 76
rect 3636 44 3640 76
rect 3600 -4 3640 44
rect 3600 -36 3604 -4
rect 3636 -36 3640 -4
rect 3600 -84 3640 -36
rect 3600 -116 3604 -84
rect 3636 -116 3640 -84
rect 3600 -120 3640 -116
rect 3680 876 3720 880
rect 3680 844 3684 876
rect 3716 844 3720 876
rect 3680 796 3720 844
rect 3680 764 3684 796
rect 3716 764 3720 796
rect 3680 716 3720 764
rect 3680 684 3684 716
rect 3716 684 3720 716
rect 3680 636 3720 684
rect 3680 604 3684 636
rect 3716 604 3720 636
rect 3680 556 3720 604
rect 3680 524 3684 556
rect 3716 524 3720 556
rect 3680 476 3720 524
rect 3680 444 3684 476
rect 3716 444 3720 476
rect 3680 396 3720 444
rect 3680 364 3684 396
rect 3716 364 3720 396
rect 3680 316 3720 364
rect 3680 284 3684 316
rect 3716 284 3720 316
rect 3680 236 3720 284
rect 3680 204 3684 236
rect 3716 204 3720 236
rect 3680 156 3720 204
rect 3680 124 3684 156
rect 3716 124 3720 156
rect 3680 76 3720 124
rect 3680 44 3684 76
rect 3716 44 3720 76
rect 3680 -4 3720 44
rect 3680 -36 3684 -4
rect 3716 -36 3720 -4
rect 3680 -84 3720 -36
rect 3680 -116 3684 -84
rect 3716 -116 3720 -84
rect 3680 -120 3720 -116
rect 3760 876 3800 880
rect 3760 844 3764 876
rect 3796 844 3800 876
rect 3760 796 3800 844
rect 3760 764 3764 796
rect 3796 764 3800 796
rect 3760 716 3800 764
rect 3760 684 3764 716
rect 3796 684 3800 716
rect 3760 636 3800 684
rect 3760 604 3764 636
rect 3796 604 3800 636
rect 3760 556 3800 604
rect 3760 524 3764 556
rect 3796 524 3800 556
rect 3760 476 3800 524
rect 3760 444 3764 476
rect 3796 444 3800 476
rect 3760 396 3800 444
rect 3760 364 3764 396
rect 3796 364 3800 396
rect 3760 316 3800 364
rect 3760 284 3764 316
rect 3796 284 3800 316
rect 3760 236 3800 284
rect 3760 204 3764 236
rect 3796 204 3800 236
rect 3760 156 3800 204
rect 3760 124 3764 156
rect 3796 124 3800 156
rect 3760 76 3800 124
rect 3760 44 3764 76
rect 3796 44 3800 76
rect 3760 -4 3800 44
rect 3760 -36 3764 -4
rect 3796 -36 3800 -4
rect 3760 -84 3800 -36
rect 3760 -116 3764 -84
rect 3796 -116 3800 -84
rect 3760 -120 3800 -116
rect 3840 876 3880 880
rect 3840 844 3844 876
rect 3876 844 3880 876
rect 3840 796 3880 844
rect 3840 764 3844 796
rect 3876 764 3880 796
rect 3840 716 3880 764
rect 3840 684 3844 716
rect 3876 684 3880 716
rect 3840 636 3880 684
rect 3840 604 3844 636
rect 3876 604 3880 636
rect 3840 556 3880 604
rect 3840 524 3844 556
rect 3876 524 3880 556
rect 3840 476 3880 524
rect 3840 444 3844 476
rect 3876 444 3880 476
rect 3840 396 3880 444
rect 3840 364 3844 396
rect 3876 364 3880 396
rect 3840 316 3880 364
rect 3840 284 3844 316
rect 3876 284 3880 316
rect 3840 236 3880 284
rect 3840 204 3844 236
rect 3876 204 3880 236
rect 3840 156 3880 204
rect 3840 124 3844 156
rect 3876 124 3880 156
rect 3840 76 3880 124
rect 3840 44 3844 76
rect 3876 44 3880 76
rect 3840 -4 3880 44
rect 3840 -36 3844 -4
rect 3876 -36 3880 -4
rect 3840 -84 3880 -36
rect 3840 -116 3844 -84
rect 3876 -116 3880 -84
rect 3840 -120 3880 -116
rect 3920 876 3960 880
rect 3920 844 3924 876
rect 3956 844 3960 876
rect 3920 796 3960 844
rect 3920 764 3924 796
rect 3956 764 3960 796
rect 3920 716 3960 764
rect 3920 684 3924 716
rect 3956 684 3960 716
rect 3920 636 3960 684
rect 3920 604 3924 636
rect 3956 604 3960 636
rect 3920 556 3960 604
rect 3920 524 3924 556
rect 3956 524 3960 556
rect 3920 476 3960 524
rect 3920 444 3924 476
rect 3956 444 3960 476
rect 3920 396 3960 444
rect 3920 364 3924 396
rect 3956 364 3960 396
rect 3920 316 3960 364
rect 3920 284 3924 316
rect 3956 284 3960 316
rect 3920 236 3960 284
rect 3920 204 3924 236
rect 3956 204 3960 236
rect 3920 156 3960 204
rect 3920 124 3924 156
rect 3956 124 3960 156
rect 3920 76 3960 124
rect 3920 44 3924 76
rect 3956 44 3960 76
rect 3920 -4 3960 44
rect 3920 -36 3924 -4
rect 3956 -36 3960 -4
rect 3920 -84 3960 -36
rect 3920 -116 3924 -84
rect 3956 -116 3960 -84
rect 3920 -120 3960 -116
rect 4000 876 4040 880
rect 4000 844 4004 876
rect 4036 844 4040 876
rect 4000 796 4040 844
rect 4000 764 4004 796
rect 4036 764 4040 796
rect 4000 716 4040 764
rect 4000 684 4004 716
rect 4036 684 4040 716
rect 4000 636 4040 684
rect 4000 604 4004 636
rect 4036 604 4040 636
rect 4000 556 4040 604
rect 4000 524 4004 556
rect 4036 524 4040 556
rect 4000 476 4040 524
rect 4000 444 4004 476
rect 4036 444 4040 476
rect 4000 396 4040 444
rect 4000 364 4004 396
rect 4036 364 4040 396
rect 4000 316 4040 364
rect 4000 284 4004 316
rect 4036 284 4040 316
rect 4000 236 4040 284
rect 4000 204 4004 236
rect 4036 204 4040 236
rect 4000 156 4040 204
rect 4000 124 4004 156
rect 4036 124 4040 156
rect 4000 76 4040 124
rect 4000 44 4004 76
rect 4036 44 4040 76
rect 4000 -4 4040 44
rect 4000 -36 4004 -4
rect 4036 -36 4040 -4
rect 4000 -84 4040 -36
rect 4000 -116 4004 -84
rect 4036 -116 4040 -84
rect 4000 -120 4040 -116
rect 4080 876 4120 880
rect 4080 844 4084 876
rect 4116 844 4120 876
rect 4080 796 4120 844
rect 4080 764 4084 796
rect 4116 764 4120 796
rect 4080 716 4120 764
rect 4080 684 4084 716
rect 4116 684 4120 716
rect 4080 636 4120 684
rect 4080 604 4084 636
rect 4116 604 4120 636
rect 4080 556 4120 604
rect 4080 524 4084 556
rect 4116 524 4120 556
rect 4080 476 4120 524
rect 4080 444 4084 476
rect 4116 444 4120 476
rect 4080 396 4120 444
rect 4080 364 4084 396
rect 4116 364 4120 396
rect 4080 316 4120 364
rect 4080 284 4084 316
rect 4116 284 4120 316
rect 4080 236 4120 284
rect 4080 204 4084 236
rect 4116 204 4120 236
rect 4080 156 4120 204
rect 4080 124 4084 156
rect 4116 124 4120 156
rect 4080 76 4120 124
rect 4080 44 4084 76
rect 4116 44 4120 76
rect 4080 -4 4120 44
rect 4080 -36 4084 -4
rect 4116 -36 4120 -4
rect 4080 -84 4120 -36
rect 4080 -116 4084 -84
rect 4116 -116 4120 -84
rect 4080 -120 4120 -116
rect 4160 876 4200 880
rect 4160 844 4164 876
rect 4196 844 4200 876
rect 4160 796 4200 844
rect 4160 764 4164 796
rect 4196 764 4200 796
rect 4160 716 4200 764
rect 4160 684 4164 716
rect 4196 684 4200 716
rect 4160 636 4200 684
rect 4160 604 4164 636
rect 4196 604 4200 636
rect 4160 556 4200 604
rect 4160 524 4164 556
rect 4196 524 4200 556
rect 4160 476 4200 524
rect 4160 444 4164 476
rect 4196 444 4200 476
rect 4160 396 4200 444
rect 4160 364 4164 396
rect 4196 364 4200 396
rect 4160 316 4200 364
rect 4160 284 4164 316
rect 4196 284 4200 316
rect 4160 236 4200 284
rect 4160 204 4164 236
rect 4196 204 4200 236
rect 4160 156 4200 204
rect 4160 124 4164 156
rect 4196 124 4200 156
rect 4160 76 4200 124
rect 4160 44 4164 76
rect 4196 44 4200 76
rect 4160 -4 4200 44
rect 4160 -36 4164 -4
rect 4196 -36 4200 -4
rect 4160 -84 4200 -36
rect 4160 -116 4164 -84
rect 4196 -116 4200 -84
rect 4160 -120 4200 -116
rect 4240 876 4280 880
rect 4240 844 4244 876
rect 4276 844 4280 876
rect 4240 796 4280 844
rect 4240 764 4244 796
rect 4276 764 4280 796
rect 4240 716 4280 764
rect 4240 684 4244 716
rect 4276 684 4280 716
rect 4240 636 4280 684
rect 4240 604 4244 636
rect 4276 604 4280 636
rect 4240 556 4280 604
rect 4240 524 4244 556
rect 4276 524 4280 556
rect 4240 476 4280 524
rect 4240 444 4244 476
rect 4276 444 4280 476
rect 4240 396 4280 444
rect 4240 364 4244 396
rect 4276 364 4280 396
rect 4240 316 4280 364
rect 4240 284 4244 316
rect 4276 284 4280 316
rect 4240 236 4280 284
rect 4240 204 4244 236
rect 4276 204 4280 236
rect 4240 156 4280 204
rect 4240 124 4244 156
rect 4276 124 4280 156
rect 4240 76 4280 124
rect 4240 44 4244 76
rect 4276 44 4280 76
rect 4240 -4 4280 44
rect 4240 -36 4244 -4
rect 4276 -36 4280 -4
rect 4240 -84 4280 -36
rect 4240 -116 4244 -84
rect 4276 -116 4280 -84
rect 4240 -120 4280 -116
rect 4320 876 4360 880
rect 4320 844 4324 876
rect 4356 844 4360 876
rect 4320 796 4360 844
rect 4320 764 4324 796
rect 4356 764 4360 796
rect 4320 716 4360 764
rect 4320 684 4324 716
rect 4356 684 4360 716
rect 4320 636 4360 684
rect 4320 604 4324 636
rect 4356 604 4360 636
rect 4320 556 4360 604
rect 4320 524 4324 556
rect 4356 524 4360 556
rect 4320 476 4360 524
rect 4320 444 4324 476
rect 4356 444 4360 476
rect 4320 396 4360 444
rect 4320 364 4324 396
rect 4356 364 4360 396
rect 4320 316 4360 364
rect 4320 284 4324 316
rect 4356 284 4360 316
rect 4320 236 4360 284
rect 4320 204 4324 236
rect 4356 204 4360 236
rect 4320 156 4360 204
rect 4320 124 4324 156
rect 4356 124 4360 156
rect 4320 76 4360 124
rect 4320 44 4324 76
rect 4356 44 4360 76
rect 4320 -4 4360 44
rect 4320 -36 4324 -4
rect 4356 -36 4360 -4
rect 4320 -84 4360 -36
rect 4320 -116 4324 -84
rect 4356 -116 4360 -84
rect 4320 -120 4360 -116
rect 4400 876 4440 880
rect 4400 844 4404 876
rect 4436 844 4440 876
rect 4400 796 4440 844
rect 4400 764 4404 796
rect 4436 764 4440 796
rect 4400 716 4440 764
rect 4400 684 4404 716
rect 4436 684 4440 716
rect 4400 636 4440 684
rect 4400 604 4404 636
rect 4436 604 4440 636
rect 4400 556 4440 604
rect 4400 524 4404 556
rect 4436 524 4440 556
rect 4400 476 4440 524
rect 4400 444 4404 476
rect 4436 444 4440 476
rect 4400 396 4440 444
rect 4400 364 4404 396
rect 4436 364 4440 396
rect 4400 316 4440 364
rect 4400 284 4404 316
rect 4436 284 4440 316
rect 4400 236 4440 284
rect 4400 204 4404 236
rect 4436 204 4440 236
rect 4400 156 4440 204
rect 4400 124 4404 156
rect 4436 124 4440 156
rect 4400 76 4440 124
rect 4400 44 4404 76
rect 4436 44 4440 76
rect 4400 -4 4440 44
rect 4400 -36 4404 -4
rect 4436 -36 4440 -4
rect 4400 -84 4440 -36
rect 4400 -116 4404 -84
rect 4436 -116 4440 -84
rect 4400 -120 4440 -116
rect 4480 876 4520 880
rect 4480 844 4484 876
rect 4516 844 4520 876
rect 4480 796 4520 844
rect 4480 764 4484 796
rect 4516 764 4520 796
rect 4480 716 4520 764
rect 4480 684 4484 716
rect 4516 684 4520 716
rect 4480 636 4520 684
rect 4480 604 4484 636
rect 4516 604 4520 636
rect 4480 556 4520 604
rect 4480 524 4484 556
rect 4516 524 4520 556
rect 4480 476 4520 524
rect 4480 444 4484 476
rect 4516 444 4520 476
rect 4480 396 4520 444
rect 4480 364 4484 396
rect 4516 364 4520 396
rect 4480 316 4520 364
rect 4480 284 4484 316
rect 4516 284 4520 316
rect 4480 236 4520 284
rect 4480 204 4484 236
rect 4516 204 4520 236
rect 4480 156 4520 204
rect 4480 124 4484 156
rect 4516 124 4520 156
rect 4480 76 4520 124
rect 4480 44 4484 76
rect 4516 44 4520 76
rect 4480 -4 4520 44
rect 4480 -36 4484 -4
rect 4516 -36 4520 -4
rect 4480 -84 4520 -36
rect 4480 -116 4484 -84
rect 4516 -116 4520 -84
rect 4480 -120 4520 -116
rect 4560 876 4600 880
rect 4560 844 4564 876
rect 4596 844 4600 876
rect 4560 796 4600 844
rect 4560 764 4564 796
rect 4596 764 4600 796
rect 4560 716 4600 764
rect 4560 684 4564 716
rect 4596 684 4600 716
rect 4560 636 4600 684
rect 4560 604 4564 636
rect 4596 604 4600 636
rect 4560 556 4600 604
rect 4560 524 4564 556
rect 4596 524 4600 556
rect 4560 476 4600 524
rect 4560 444 4564 476
rect 4596 444 4600 476
rect 4560 396 4600 444
rect 4560 364 4564 396
rect 4596 364 4600 396
rect 4560 316 4600 364
rect 4560 284 4564 316
rect 4596 284 4600 316
rect 4560 236 4600 284
rect 4560 204 4564 236
rect 4596 204 4600 236
rect 4560 156 4600 204
rect 4560 124 4564 156
rect 4596 124 4600 156
rect 4560 76 4600 124
rect 4560 44 4564 76
rect 4596 44 4600 76
rect 4560 -4 4600 44
rect 4560 -36 4564 -4
rect 4596 -36 4600 -4
rect 4560 -84 4600 -36
rect 4560 -116 4564 -84
rect 4596 -116 4600 -84
rect 4560 -120 4600 -116
rect 4640 876 4680 880
rect 4640 844 4644 876
rect 4676 844 4680 876
rect 4640 796 4680 844
rect 4640 764 4644 796
rect 4676 764 4680 796
rect 4640 716 4680 764
rect 4640 684 4644 716
rect 4676 684 4680 716
rect 4640 636 4680 684
rect 4640 604 4644 636
rect 4676 604 4680 636
rect 4640 556 4680 604
rect 4640 524 4644 556
rect 4676 524 4680 556
rect 4640 476 4680 524
rect 4640 444 4644 476
rect 4676 444 4680 476
rect 4640 396 4680 444
rect 4640 364 4644 396
rect 4676 364 4680 396
rect 4640 316 4680 364
rect 4640 284 4644 316
rect 4676 284 4680 316
rect 4640 236 4680 284
rect 4640 204 4644 236
rect 4676 204 4680 236
rect 4640 156 4680 204
rect 4640 124 4644 156
rect 4676 124 4680 156
rect 4640 76 4680 124
rect 4640 44 4644 76
rect 4676 44 4680 76
rect 4640 -4 4680 44
rect 4640 -36 4644 -4
rect 4676 -36 4680 -4
rect 4640 -84 4680 -36
rect 4640 -116 4644 -84
rect 4676 -116 4680 -84
rect 4640 -120 4680 -116
rect 4720 876 4760 880
rect 4720 844 4724 876
rect 4756 844 4760 876
rect 4720 796 4760 844
rect 4720 764 4724 796
rect 4756 764 4760 796
rect 4720 716 4760 764
rect 4720 684 4724 716
rect 4756 684 4760 716
rect 4720 636 4760 684
rect 4720 604 4724 636
rect 4756 604 4760 636
rect 4720 556 4760 604
rect 4720 524 4724 556
rect 4756 524 4760 556
rect 4720 476 4760 524
rect 4720 444 4724 476
rect 4756 444 4760 476
rect 4720 396 4760 444
rect 4720 364 4724 396
rect 4756 364 4760 396
rect 4720 316 4760 364
rect 4720 284 4724 316
rect 4756 284 4760 316
rect 4720 236 4760 284
rect 4720 204 4724 236
rect 4756 204 4760 236
rect 4720 156 4760 204
rect 4720 124 4724 156
rect 4756 124 4760 156
rect 4720 76 4760 124
rect 4720 44 4724 76
rect 4756 44 4760 76
rect 4720 -4 4760 44
rect 4720 -36 4724 -4
rect 4756 -36 4760 -4
rect 4720 -84 4760 -36
rect 4720 -116 4724 -84
rect 4756 -116 4760 -84
rect 4720 -120 4760 -116
rect 4800 876 4840 880
rect 4800 844 4804 876
rect 4836 844 4840 876
rect 4800 796 4840 844
rect 4800 764 4804 796
rect 4836 764 4840 796
rect 4800 716 4840 764
rect 4800 684 4804 716
rect 4836 684 4840 716
rect 4800 636 4840 684
rect 4800 604 4804 636
rect 4836 604 4840 636
rect 4800 556 4840 604
rect 4800 524 4804 556
rect 4836 524 4840 556
rect 4800 476 4840 524
rect 4800 444 4804 476
rect 4836 444 4840 476
rect 4800 396 4840 444
rect 4800 364 4804 396
rect 4836 364 4840 396
rect 4800 316 4840 364
rect 4800 284 4804 316
rect 4836 284 4840 316
rect 4800 236 4840 284
rect 4800 204 4804 236
rect 4836 204 4840 236
rect 4800 156 4840 204
rect 4800 124 4804 156
rect 4836 124 4840 156
rect 4800 76 4840 124
rect 4800 44 4804 76
rect 4836 44 4840 76
rect 4800 -4 4840 44
rect 4800 -36 4804 -4
rect 4836 -36 4840 -4
rect 4800 -84 4840 -36
rect 4800 -116 4804 -84
rect 4836 -116 4840 -84
rect 4800 -120 4840 -116
rect 4880 876 4920 924
rect 4880 844 4884 876
rect 4916 844 4920 876
rect 4880 796 4920 844
rect 4880 764 4884 796
rect 4916 764 4920 796
rect 4880 716 4920 764
rect 4880 684 4884 716
rect 4916 684 4920 716
rect 4880 636 4920 684
rect 4880 604 4884 636
rect 4916 604 4920 636
rect 4880 556 4920 604
rect 4880 524 4884 556
rect 4916 524 4920 556
rect 4880 476 4920 524
rect 4880 444 4884 476
rect 4916 444 4920 476
rect 4880 396 4920 444
rect 4880 364 4884 396
rect 4916 364 4920 396
rect 4880 316 4920 364
rect 4880 284 4884 316
rect 4916 284 4920 316
rect 4880 236 4920 284
rect 4880 204 4884 236
rect 4916 204 4920 236
rect 4880 156 4920 204
rect 4880 124 4884 156
rect 4916 124 4920 156
rect 4880 76 4920 124
rect 4880 44 4884 76
rect 4916 44 4920 76
rect 4880 -4 4920 44
rect 4880 -36 4884 -4
rect 4916 -36 4920 -4
rect 4880 -84 4920 -36
rect 4880 -116 4884 -84
rect 4916 -116 4920 -84
rect 4880 -120 4920 -116
rect 4960 4155 5000 5640
rect 4960 4125 4965 4155
rect 4995 4125 5000 4155
rect 4960 2235 5000 4125
rect 4960 2205 4965 2235
rect 4995 2205 5000 2235
rect 4960 315 5000 2205
rect 4960 285 4965 315
rect 4995 285 5000 315
rect 4960 -120 5000 285
rect 5040 5596 5080 5640
rect 5040 5564 5044 5596
rect 5076 5564 5080 5596
rect 5040 5516 5080 5564
rect 5040 5484 5044 5516
rect 5076 5484 5080 5516
rect 5040 5436 5080 5484
rect 5040 5404 5044 5436
rect 5076 5404 5080 5436
rect 5040 5356 5080 5404
rect 5040 5324 5044 5356
rect 5076 5324 5080 5356
rect 5040 5276 5080 5324
rect 5040 5244 5044 5276
rect 5076 5244 5080 5276
rect 5040 5196 5080 5244
rect 5040 5164 5044 5196
rect 5076 5164 5080 5196
rect 5040 5116 5080 5164
rect 5040 5084 5044 5116
rect 5076 5084 5080 5116
rect 5040 5036 5080 5084
rect 5040 5004 5044 5036
rect 5076 5004 5080 5036
rect 5040 4956 5080 5004
rect 5040 4924 5044 4956
rect 5076 4924 5080 4956
rect 5040 4876 5080 4924
rect 5040 4844 5044 4876
rect 5076 4844 5080 4876
rect 5040 4796 5080 4844
rect 5040 4764 5044 4796
rect 5076 4764 5080 4796
rect 5040 4716 5080 4764
rect 5040 4684 5044 4716
rect 5076 4684 5080 4716
rect 5040 4636 5080 4684
rect 5040 4604 5044 4636
rect 5076 4604 5080 4636
rect 5040 4556 5080 4604
rect 5040 4524 5044 4556
rect 5076 4524 5080 4556
rect 5040 4476 5080 4524
rect 5040 4444 5044 4476
rect 5076 4444 5080 4476
rect 5040 4396 5080 4444
rect 5040 4364 5044 4396
rect 5076 4364 5080 4396
rect 5040 4316 5080 4364
rect 5040 4284 5044 4316
rect 5076 4284 5080 4316
rect 5040 4236 5080 4284
rect 5040 4204 5044 4236
rect 5076 4204 5080 4236
rect 5040 4156 5080 4204
rect 5040 4124 5044 4156
rect 5076 4124 5080 4156
rect 5040 4076 5080 4124
rect 5040 4044 5044 4076
rect 5076 4044 5080 4076
rect 5040 3996 5080 4044
rect 5040 3964 5044 3996
rect 5076 3964 5080 3996
rect 5040 3916 5080 3964
rect 5040 3884 5044 3916
rect 5076 3884 5080 3916
rect 5040 3836 5080 3884
rect 5040 3804 5044 3836
rect 5076 3804 5080 3836
rect 5040 3756 5080 3804
rect 5040 3724 5044 3756
rect 5076 3724 5080 3756
rect 5040 3676 5080 3724
rect 5040 3644 5044 3676
rect 5076 3644 5080 3676
rect 5040 3596 5080 3644
rect 5040 3564 5044 3596
rect 5076 3564 5080 3596
rect 5040 3516 5080 3564
rect 5040 3484 5044 3516
rect 5076 3484 5080 3516
rect 5040 3436 5080 3484
rect 5040 3404 5044 3436
rect 5076 3404 5080 3436
rect 5040 3356 5080 3404
rect 5040 3324 5044 3356
rect 5076 3324 5080 3356
rect 5040 3276 5080 3324
rect 5040 3244 5044 3276
rect 5076 3244 5080 3276
rect 5040 3196 5080 3244
rect 5040 3164 5044 3196
rect 5076 3164 5080 3196
rect 5040 3116 5080 3164
rect 5040 3084 5044 3116
rect 5076 3084 5080 3116
rect 5040 3036 5080 3084
rect 5040 3004 5044 3036
rect 5076 3004 5080 3036
rect 5040 2956 5080 3004
rect 5040 2924 5044 2956
rect 5076 2924 5080 2956
rect 5040 2876 5080 2924
rect 5040 2844 5044 2876
rect 5076 2844 5080 2876
rect 5040 2796 5080 2844
rect 5040 2764 5044 2796
rect 5076 2764 5080 2796
rect 5040 2716 5080 2764
rect 5040 2684 5044 2716
rect 5076 2684 5080 2716
rect 5040 2636 5080 2684
rect 5040 2604 5044 2636
rect 5076 2604 5080 2636
rect 5040 2556 5080 2604
rect 5040 2524 5044 2556
rect 5076 2524 5080 2556
rect 5040 2476 5080 2524
rect 5040 2444 5044 2476
rect 5076 2444 5080 2476
rect 5040 2396 5080 2444
rect 5040 2364 5044 2396
rect 5076 2364 5080 2396
rect 5040 2316 5080 2364
rect 5040 2284 5044 2316
rect 5076 2284 5080 2316
rect 5040 2236 5080 2284
rect 5040 2204 5044 2236
rect 5076 2204 5080 2236
rect 5040 2156 5080 2204
rect 5040 2124 5044 2156
rect 5076 2124 5080 2156
rect 5040 2076 5080 2124
rect 5040 2044 5044 2076
rect 5076 2044 5080 2076
rect 5040 1996 5080 2044
rect 5040 1964 5044 1996
rect 5076 1964 5080 1996
rect 5040 1916 5080 1964
rect 5040 1884 5044 1916
rect 5076 1884 5080 1916
rect 5040 1836 5080 1884
rect 5040 1804 5044 1836
rect 5076 1804 5080 1836
rect 5040 1756 5080 1804
rect 5040 1724 5044 1756
rect 5076 1724 5080 1756
rect 5040 1676 5080 1724
rect 5040 1644 5044 1676
rect 5076 1644 5080 1676
rect 5040 1596 5080 1644
rect 5040 1564 5044 1596
rect 5076 1564 5080 1596
rect 5040 1516 5080 1564
rect 5040 1484 5044 1516
rect 5076 1484 5080 1516
rect 5040 1436 5080 1484
rect 5040 1404 5044 1436
rect 5076 1404 5080 1436
rect 5040 1356 5080 1404
rect 5040 1324 5044 1356
rect 5076 1324 5080 1356
rect 5040 1276 5080 1324
rect 5040 1244 5044 1276
rect 5076 1244 5080 1276
rect 5040 1196 5080 1244
rect 5040 1164 5044 1196
rect 5076 1164 5080 1196
rect 5040 1116 5080 1164
rect 5040 1084 5044 1116
rect 5076 1084 5080 1116
rect 5040 1036 5080 1084
rect 5040 1004 5044 1036
rect 5076 1004 5080 1036
rect 5040 956 5080 1004
rect 5040 924 5044 956
rect 5076 924 5080 956
rect 5040 876 5080 924
rect 5040 844 5044 876
rect 5076 844 5080 876
rect 5040 796 5080 844
rect 5040 764 5044 796
rect 5076 764 5080 796
rect 5040 716 5080 764
rect 5040 684 5044 716
rect 5076 684 5080 716
rect 5040 636 5080 684
rect 5040 604 5044 636
rect 5076 604 5080 636
rect 5040 556 5080 604
rect 5040 524 5044 556
rect 5076 524 5080 556
rect 5040 476 5080 524
rect 5040 444 5044 476
rect 5076 444 5080 476
rect 5040 396 5080 444
rect 5040 364 5044 396
rect 5076 364 5080 396
rect 5040 316 5080 364
rect 5040 284 5044 316
rect 5076 284 5080 316
rect 5040 236 5080 284
rect 5040 204 5044 236
rect 5076 204 5080 236
rect 5040 156 5080 204
rect 5040 124 5044 156
rect 5076 124 5080 156
rect 5040 76 5080 124
rect 5040 44 5044 76
rect 5076 44 5080 76
rect 5040 -4 5080 44
rect 5040 -36 5044 -4
rect 5076 -36 5080 -4
rect 5040 -84 5080 -36
rect 5040 -116 5044 -84
rect 5076 -116 5080 -84
rect 5040 -120 5080 -116
rect 5120 475 5160 5640
rect 5120 445 5125 475
rect 5155 445 5160 475
rect 5120 -120 5160 445
rect 5200 5596 5240 5640
rect 5200 5564 5204 5596
rect 5236 5564 5240 5596
rect 5200 5516 5240 5564
rect 5200 5484 5204 5516
rect 5236 5484 5240 5516
rect 5200 5436 5240 5484
rect 5200 5404 5204 5436
rect 5236 5404 5240 5436
rect 5200 5356 5240 5404
rect 5200 5324 5204 5356
rect 5236 5324 5240 5356
rect 5200 5276 5240 5324
rect 5200 5244 5204 5276
rect 5236 5244 5240 5276
rect 5200 5196 5240 5244
rect 5200 5164 5204 5196
rect 5236 5164 5240 5196
rect 5200 5116 5240 5164
rect 5200 5084 5204 5116
rect 5236 5084 5240 5116
rect 5200 5036 5240 5084
rect 5200 5004 5204 5036
rect 5236 5004 5240 5036
rect 5200 4956 5240 5004
rect 5200 4924 5204 4956
rect 5236 4924 5240 4956
rect 5200 4876 5240 4924
rect 5200 4844 5204 4876
rect 5236 4844 5240 4876
rect 5200 4796 5240 4844
rect 5200 4764 5204 4796
rect 5236 4764 5240 4796
rect 5200 4716 5240 4764
rect 5200 4684 5204 4716
rect 5236 4684 5240 4716
rect 5200 4636 5240 4684
rect 5200 4604 5204 4636
rect 5236 4604 5240 4636
rect 5200 4556 5240 4604
rect 5200 4524 5204 4556
rect 5236 4524 5240 4556
rect 5200 4476 5240 4524
rect 5200 4444 5204 4476
rect 5236 4444 5240 4476
rect 5200 4396 5240 4444
rect 5200 4364 5204 4396
rect 5236 4364 5240 4396
rect 5200 4316 5240 4364
rect 5200 4284 5204 4316
rect 5236 4284 5240 4316
rect 5200 4236 5240 4284
rect 5200 4204 5204 4236
rect 5236 4204 5240 4236
rect 5200 4156 5240 4204
rect 5200 4124 5204 4156
rect 5236 4124 5240 4156
rect 5200 4076 5240 4124
rect 5200 4044 5204 4076
rect 5236 4044 5240 4076
rect 5200 3996 5240 4044
rect 5200 3964 5204 3996
rect 5236 3964 5240 3996
rect 5200 3916 5240 3964
rect 5200 3884 5204 3916
rect 5236 3884 5240 3916
rect 5200 3836 5240 3884
rect 5200 3804 5204 3836
rect 5236 3804 5240 3836
rect 5200 3756 5240 3804
rect 5200 3724 5204 3756
rect 5236 3724 5240 3756
rect 5200 3676 5240 3724
rect 5200 3644 5204 3676
rect 5236 3644 5240 3676
rect 5200 3596 5240 3644
rect 5200 3564 5204 3596
rect 5236 3564 5240 3596
rect 5200 3516 5240 3564
rect 5200 3484 5204 3516
rect 5236 3484 5240 3516
rect 5200 3436 5240 3484
rect 5200 3404 5204 3436
rect 5236 3404 5240 3436
rect 5200 3356 5240 3404
rect 5200 3324 5204 3356
rect 5236 3324 5240 3356
rect 5200 3276 5240 3324
rect 5200 3244 5204 3276
rect 5236 3244 5240 3276
rect 5200 3196 5240 3244
rect 5200 3164 5204 3196
rect 5236 3164 5240 3196
rect 5200 3116 5240 3164
rect 5200 3084 5204 3116
rect 5236 3084 5240 3116
rect 5200 3036 5240 3084
rect 5200 3004 5204 3036
rect 5236 3004 5240 3036
rect 5200 2956 5240 3004
rect 5200 2924 5204 2956
rect 5236 2924 5240 2956
rect 5200 2876 5240 2924
rect 5200 2844 5204 2876
rect 5236 2844 5240 2876
rect 5200 2796 5240 2844
rect 5200 2764 5204 2796
rect 5236 2764 5240 2796
rect 5200 2716 5240 2764
rect 5200 2684 5204 2716
rect 5236 2684 5240 2716
rect 5200 2636 5240 2684
rect 5200 2604 5204 2636
rect 5236 2604 5240 2636
rect 5200 2556 5240 2604
rect 5200 2524 5204 2556
rect 5236 2524 5240 2556
rect 5200 2476 5240 2524
rect 5200 2444 5204 2476
rect 5236 2444 5240 2476
rect 5200 2396 5240 2444
rect 5200 2364 5204 2396
rect 5236 2364 5240 2396
rect 5200 2316 5240 2364
rect 5200 2284 5204 2316
rect 5236 2284 5240 2316
rect 5200 2236 5240 2284
rect 5200 2204 5204 2236
rect 5236 2204 5240 2236
rect 5200 2156 5240 2204
rect 5200 2124 5204 2156
rect 5236 2124 5240 2156
rect 5200 2076 5240 2124
rect 5200 2044 5204 2076
rect 5236 2044 5240 2076
rect 5200 1996 5240 2044
rect 5200 1964 5204 1996
rect 5236 1964 5240 1996
rect 5200 1916 5240 1964
rect 5200 1884 5204 1916
rect 5236 1884 5240 1916
rect 5200 1836 5240 1884
rect 5200 1804 5204 1836
rect 5236 1804 5240 1836
rect 5200 1756 5240 1804
rect 5200 1724 5204 1756
rect 5236 1724 5240 1756
rect 5200 1676 5240 1724
rect 5200 1644 5204 1676
rect 5236 1644 5240 1676
rect 5200 1596 5240 1644
rect 5200 1564 5204 1596
rect 5236 1564 5240 1596
rect 5200 1516 5240 1564
rect 5200 1484 5204 1516
rect 5236 1484 5240 1516
rect 5200 1436 5240 1484
rect 5200 1404 5204 1436
rect 5236 1404 5240 1436
rect 5200 1356 5240 1404
rect 5200 1324 5204 1356
rect 5236 1324 5240 1356
rect 5200 1276 5240 1324
rect 5200 1244 5204 1276
rect 5236 1244 5240 1276
rect 5200 1196 5240 1244
rect 5200 1164 5204 1196
rect 5236 1164 5240 1196
rect 5200 1116 5240 1164
rect 5200 1084 5204 1116
rect 5236 1084 5240 1116
rect 5200 1036 5240 1084
rect 5200 1004 5204 1036
rect 5236 1004 5240 1036
rect 5200 956 5240 1004
rect 5200 924 5204 956
rect 5236 924 5240 956
rect 5200 876 5240 924
rect 5200 844 5204 876
rect 5236 844 5240 876
rect 5200 796 5240 844
rect 5200 764 5204 796
rect 5236 764 5240 796
rect 5200 716 5240 764
rect 5200 684 5204 716
rect 5236 684 5240 716
rect 5200 636 5240 684
rect 5200 604 5204 636
rect 5236 604 5240 636
rect 5200 556 5240 604
rect 5200 524 5204 556
rect 5236 524 5240 556
rect 5200 476 5240 524
rect 5200 444 5204 476
rect 5236 444 5240 476
rect 5200 396 5240 444
rect 5200 364 5204 396
rect 5236 364 5240 396
rect 5200 316 5240 364
rect 5200 284 5204 316
rect 5236 284 5240 316
rect 5200 236 5240 284
rect 5200 204 5204 236
rect 5236 204 5240 236
rect 5200 156 5240 204
rect 5200 124 5204 156
rect 5236 124 5240 156
rect 5200 76 5240 124
rect 5200 44 5204 76
rect 5236 44 5240 76
rect 5200 -4 5240 44
rect 5200 -36 5204 -4
rect 5236 -36 5240 -4
rect 5200 -84 5240 -36
rect 5200 -116 5204 -84
rect 5236 -116 5240 -84
rect 5200 -120 5240 -116
rect 5280 2395 5320 5640
rect 5280 2365 5285 2395
rect 5315 2365 5320 2395
rect 5280 635 5320 2365
rect 5280 605 5285 635
rect 5315 605 5320 635
rect 5280 -120 5320 605
rect 5360 5596 5400 5640
rect 5360 5564 5364 5596
rect 5396 5564 5400 5596
rect 5360 5516 5400 5564
rect 5360 5484 5364 5516
rect 5396 5484 5400 5516
rect 5360 5436 5400 5484
rect 5360 5404 5364 5436
rect 5396 5404 5400 5436
rect 5360 5356 5400 5404
rect 5360 5324 5364 5356
rect 5396 5324 5400 5356
rect 5360 5276 5400 5324
rect 5360 5244 5364 5276
rect 5396 5244 5400 5276
rect 5360 5196 5400 5244
rect 5360 5164 5364 5196
rect 5396 5164 5400 5196
rect 5360 5116 5400 5164
rect 5360 5084 5364 5116
rect 5396 5084 5400 5116
rect 5360 5036 5400 5084
rect 5360 5004 5364 5036
rect 5396 5004 5400 5036
rect 5360 4956 5400 5004
rect 5360 4924 5364 4956
rect 5396 4924 5400 4956
rect 5360 4876 5400 4924
rect 5360 4844 5364 4876
rect 5396 4844 5400 4876
rect 5360 4796 5400 4844
rect 5360 4764 5364 4796
rect 5396 4764 5400 4796
rect 5360 4716 5400 4764
rect 5360 4684 5364 4716
rect 5396 4684 5400 4716
rect 5360 4636 5400 4684
rect 5360 4604 5364 4636
rect 5396 4604 5400 4636
rect 5360 4556 5400 4604
rect 5360 4524 5364 4556
rect 5396 4524 5400 4556
rect 5360 4476 5400 4524
rect 5360 4444 5364 4476
rect 5396 4444 5400 4476
rect 5360 4396 5400 4444
rect 5360 4364 5364 4396
rect 5396 4364 5400 4396
rect 5360 4316 5400 4364
rect 5360 4284 5364 4316
rect 5396 4284 5400 4316
rect 5360 4236 5400 4284
rect 5360 4204 5364 4236
rect 5396 4204 5400 4236
rect 5360 4156 5400 4204
rect 5360 4124 5364 4156
rect 5396 4124 5400 4156
rect 5360 4076 5400 4124
rect 5360 4044 5364 4076
rect 5396 4044 5400 4076
rect 5360 3996 5400 4044
rect 5360 3964 5364 3996
rect 5396 3964 5400 3996
rect 5360 3916 5400 3964
rect 5360 3884 5364 3916
rect 5396 3884 5400 3916
rect 5360 3836 5400 3884
rect 5360 3804 5364 3836
rect 5396 3804 5400 3836
rect 5360 3756 5400 3804
rect 5360 3724 5364 3756
rect 5396 3724 5400 3756
rect 5360 3676 5400 3724
rect 5360 3644 5364 3676
rect 5396 3644 5400 3676
rect 5360 3596 5400 3644
rect 5360 3564 5364 3596
rect 5396 3564 5400 3596
rect 5360 3516 5400 3564
rect 5360 3484 5364 3516
rect 5396 3484 5400 3516
rect 5360 3436 5400 3484
rect 5360 3404 5364 3436
rect 5396 3404 5400 3436
rect 5360 3356 5400 3404
rect 5360 3324 5364 3356
rect 5396 3324 5400 3356
rect 5360 3276 5400 3324
rect 5360 3244 5364 3276
rect 5396 3244 5400 3276
rect 5360 3196 5400 3244
rect 5360 3164 5364 3196
rect 5396 3164 5400 3196
rect 5360 3116 5400 3164
rect 5360 3084 5364 3116
rect 5396 3084 5400 3116
rect 5360 3036 5400 3084
rect 5360 3004 5364 3036
rect 5396 3004 5400 3036
rect 5360 2956 5400 3004
rect 5360 2924 5364 2956
rect 5396 2924 5400 2956
rect 5360 2876 5400 2924
rect 5360 2844 5364 2876
rect 5396 2844 5400 2876
rect 5360 2796 5400 2844
rect 5360 2764 5364 2796
rect 5396 2764 5400 2796
rect 5360 2716 5400 2764
rect 5360 2684 5364 2716
rect 5396 2684 5400 2716
rect 5360 2636 5400 2684
rect 5360 2604 5364 2636
rect 5396 2604 5400 2636
rect 5360 2556 5400 2604
rect 5360 2524 5364 2556
rect 5396 2524 5400 2556
rect 5360 2476 5400 2524
rect 5360 2444 5364 2476
rect 5396 2444 5400 2476
rect 5360 2396 5400 2444
rect 5360 2364 5364 2396
rect 5396 2364 5400 2396
rect 5360 2316 5400 2364
rect 5360 2284 5364 2316
rect 5396 2284 5400 2316
rect 5360 2236 5400 2284
rect 5360 2204 5364 2236
rect 5396 2204 5400 2236
rect 5360 2156 5400 2204
rect 5360 2124 5364 2156
rect 5396 2124 5400 2156
rect 5360 2076 5400 2124
rect 5360 2044 5364 2076
rect 5396 2044 5400 2076
rect 5360 1996 5400 2044
rect 5360 1964 5364 1996
rect 5396 1964 5400 1996
rect 5360 1916 5400 1964
rect 5360 1884 5364 1916
rect 5396 1884 5400 1916
rect 5360 1836 5400 1884
rect 5360 1804 5364 1836
rect 5396 1804 5400 1836
rect 5360 1756 5400 1804
rect 5360 1724 5364 1756
rect 5396 1724 5400 1756
rect 5360 1676 5400 1724
rect 5360 1644 5364 1676
rect 5396 1644 5400 1676
rect 5360 1596 5400 1644
rect 5360 1564 5364 1596
rect 5396 1564 5400 1596
rect 5360 1516 5400 1564
rect 5360 1484 5364 1516
rect 5396 1484 5400 1516
rect 5360 1436 5400 1484
rect 5360 1404 5364 1436
rect 5396 1404 5400 1436
rect 5360 1356 5400 1404
rect 5360 1324 5364 1356
rect 5396 1324 5400 1356
rect 5360 1276 5400 1324
rect 5360 1244 5364 1276
rect 5396 1244 5400 1276
rect 5360 1196 5400 1244
rect 5360 1164 5364 1196
rect 5396 1164 5400 1196
rect 5360 1116 5400 1164
rect 5360 1084 5364 1116
rect 5396 1084 5400 1116
rect 5360 1036 5400 1084
rect 5360 1004 5364 1036
rect 5396 1004 5400 1036
rect 5360 956 5400 1004
rect 5360 924 5364 956
rect 5396 924 5400 956
rect 5360 876 5400 924
rect 5360 844 5364 876
rect 5396 844 5400 876
rect 5360 796 5400 844
rect 5360 764 5364 796
rect 5396 764 5400 796
rect 5360 716 5400 764
rect 5360 684 5364 716
rect 5396 684 5400 716
rect 5360 636 5400 684
rect 5360 604 5364 636
rect 5396 604 5400 636
rect 5360 556 5400 604
rect 5360 524 5364 556
rect 5396 524 5400 556
rect 5360 476 5400 524
rect 5360 444 5364 476
rect 5396 444 5400 476
rect 5360 396 5400 444
rect 5360 364 5364 396
rect 5396 364 5400 396
rect 5360 316 5400 364
rect 5360 284 5364 316
rect 5396 284 5400 316
rect 5360 236 5400 284
rect 5360 204 5364 236
rect 5396 204 5400 236
rect 5360 156 5400 204
rect 5360 124 5364 156
rect 5396 124 5400 156
rect 5360 76 5400 124
rect 5360 44 5364 76
rect 5396 44 5400 76
rect 5360 -4 5400 44
rect 5360 -36 5364 -4
rect 5396 -36 5400 -4
rect 5360 -84 5400 -36
rect 5360 -116 5364 -84
rect 5396 -116 5400 -84
rect 5360 -120 5400 -116
rect 5440 795 5480 5640
rect 5440 765 5445 795
rect 5475 765 5480 795
rect 5440 -120 5480 765
rect 5520 5596 5560 5640
rect 5520 5564 5524 5596
rect 5556 5564 5560 5596
rect 5520 5516 5560 5564
rect 5520 5484 5524 5516
rect 5556 5484 5560 5516
rect 5520 5436 5560 5484
rect 5520 5404 5524 5436
rect 5556 5404 5560 5436
rect 5520 5356 5560 5404
rect 5520 5324 5524 5356
rect 5556 5324 5560 5356
rect 5520 5276 5560 5324
rect 5520 5244 5524 5276
rect 5556 5244 5560 5276
rect 5520 5196 5560 5244
rect 5520 5164 5524 5196
rect 5556 5164 5560 5196
rect 5520 5116 5560 5164
rect 5520 5084 5524 5116
rect 5556 5084 5560 5116
rect 5520 5036 5560 5084
rect 5520 5004 5524 5036
rect 5556 5004 5560 5036
rect 5520 4956 5560 5004
rect 5520 4924 5524 4956
rect 5556 4924 5560 4956
rect 5520 4876 5560 4924
rect 5520 4844 5524 4876
rect 5556 4844 5560 4876
rect 5520 4796 5560 4844
rect 5520 4764 5524 4796
rect 5556 4764 5560 4796
rect 5520 4716 5560 4764
rect 5520 4684 5524 4716
rect 5556 4684 5560 4716
rect 5520 4636 5560 4684
rect 5520 4604 5524 4636
rect 5556 4604 5560 4636
rect 5520 4556 5560 4604
rect 5520 4524 5524 4556
rect 5556 4524 5560 4556
rect 5520 4476 5560 4524
rect 5520 4444 5524 4476
rect 5556 4444 5560 4476
rect 5520 4396 5560 4444
rect 5520 4364 5524 4396
rect 5556 4364 5560 4396
rect 5520 4316 5560 4364
rect 5520 4284 5524 4316
rect 5556 4284 5560 4316
rect 5520 4236 5560 4284
rect 5520 4204 5524 4236
rect 5556 4204 5560 4236
rect 5520 4156 5560 4204
rect 5520 4124 5524 4156
rect 5556 4124 5560 4156
rect 5520 4076 5560 4124
rect 5520 4044 5524 4076
rect 5556 4044 5560 4076
rect 5520 3996 5560 4044
rect 5520 3964 5524 3996
rect 5556 3964 5560 3996
rect 5520 3916 5560 3964
rect 5520 3884 5524 3916
rect 5556 3884 5560 3916
rect 5520 3836 5560 3884
rect 5520 3804 5524 3836
rect 5556 3804 5560 3836
rect 5520 3756 5560 3804
rect 5520 3724 5524 3756
rect 5556 3724 5560 3756
rect 5520 3676 5560 3724
rect 5520 3644 5524 3676
rect 5556 3644 5560 3676
rect 5520 3596 5560 3644
rect 5520 3564 5524 3596
rect 5556 3564 5560 3596
rect 5520 3516 5560 3564
rect 5520 3484 5524 3516
rect 5556 3484 5560 3516
rect 5520 3436 5560 3484
rect 5520 3404 5524 3436
rect 5556 3404 5560 3436
rect 5520 3356 5560 3404
rect 5520 3324 5524 3356
rect 5556 3324 5560 3356
rect 5520 3276 5560 3324
rect 5520 3244 5524 3276
rect 5556 3244 5560 3276
rect 5520 3196 5560 3244
rect 5520 3164 5524 3196
rect 5556 3164 5560 3196
rect 5520 3116 5560 3164
rect 5520 3084 5524 3116
rect 5556 3084 5560 3116
rect 5520 3036 5560 3084
rect 5520 3004 5524 3036
rect 5556 3004 5560 3036
rect 5520 2956 5560 3004
rect 5520 2924 5524 2956
rect 5556 2924 5560 2956
rect 5520 2876 5560 2924
rect 5520 2844 5524 2876
rect 5556 2844 5560 2876
rect 5520 2796 5560 2844
rect 5520 2764 5524 2796
rect 5556 2764 5560 2796
rect 5520 2716 5560 2764
rect 5520 2684 5524 2716
rect 5556 2684 5560 2716
rect 5520 2636 5560 2684
rect 5520 2604 5524 2636
rect 5556 2604 5560 2636
rect 5520 2556 5560 2604
rect 5520 2524 5524 2556
rect 5556 2524 5560 2556
rect 5520 2476 5560 2524
rect 5520 2444 5524 2476
rect 5556 2444 5560 2476
rect 5520 2396 5560 2444
rect 5520 2364 5524 2396
rect 5556 2364 5560 2396
rect 5520 2316 5560 2364
rect 5520 2284 5524 2316
rect 5556 2284 5560 2316
rect 5520 2236 5560 2284
rect 5520 2204 5524 2236
rect 5556 2204 5560 2236
rect 5520 2156 5560 2204
rect 5520 2124 5524 2156
rect 5556 2124 5560 2156
rect 5520 2076 5560 2124
rect 5520 2044 5524 2076
rect 5556 2044 5560 2076
rect 5520 1996 5560 2044
rect 5520 1964 5524 1996
rect 5556 1964 5560 1996
rect 5520 1916 5560 1964
rect 5520 1884 5524 1916
rect 5556 1884 5560 1916
rect 5520 1836 5560 1884
rect 5520 1804 5524 1836
rect 5556 1804 5560 1836
rect 5520 1756 5560 1804
rect 5520 1724 5524 1756
rect 5556 1724 5560 1756
rect 5520 1676 5560 1724
rect 5520 1644 5524 1676
rect 5556 1644 5560 1676
rect 5520 1596 5560 1644
rect 5520 1564 5524 1596
rect 5556 1564 5560 1596
rect 5520 1516 5560 1564
rect 5520 1484 5524 1516
rect 5556 1484 5560 1516
rect 5520 1436 5560 1484
rect 5520 1404 5524 1436
rect 5556 1404 5560 1436
rect 5520 1356 5560 1404
rect 5520 1324 5524 1356
rect 5556 1324 5560 1356
rect 5520 1276 5560 1324
rect 5520 1244 5524 1276
rect 5556 1244 5560 1276
rect 5520 1196 5560 1244
rect 5520 1164 5524 1196
rect 5556 1164 5560 1196
rect 5520 1116 5560 1164
rect 5520 1084 5524 1116
rect 5556 1084 5560 1116
rect 5520 1036 5560 1084
rect 5520 1004 5524 1036
rect 5556 1004 5560 1036
rect 5520 956 5560 1004
rect 5520 924 5524 956
rect 5556 924 5560 956
rect 5520 876 5560 924
rect 5520 844 5524 876
rect 5556 844 5560 876
rect 5520 796 5560 844
rect 5520 764 5524 796
rect 5556 764 5560 796
rect 5520 716 5560 764
rect 5520 684 5524 716
rect 5556 684 5560 716
rect 5520 636 5560 684
rect 5520 604 5524 636
rect 5556 604 5560 636
rect 5520 556 5560 604
rect 5520 524 5524 556
rect 5556 524 5560 556
rect 5520 476 5560 524
rect 5520 444 5524 476
rect 5556 444 5560 476
rect 5520 396 5560 444
rect 5520 364 5524 396
rect 5556 364 5560 396
rect 5520 316 5560 364
rect 5520 284 5524 316
rect 5556 284 5560 316
rect 5520 236 5560 284
rect 5520 204 5524 236
rect 5556 204 5560 236
rect 5520 156 5560 204
rect 5520 124 5524 156
rect 5556 124 5560 156
rect 5520 76 5560 124
rect 5520 44 5524 76
rect 5556 44 5560 76
rect 5520 -4 5560 44
rect 5520 -36 5524 -4
rect 5556 -36 5560 -4
rect 5520 -84 5560 -36
rect 5520 -116 5524 -84
rect 5556 -116 5560 -84
rect 5520 -120 5560 -116
rect 5600 4315 5640 5640
rect 5600 4285 5605 4315
rect 5635 4285 5640 4315
rect 5600 -120 5640 4285
rect 5680 5596 5720 5640
rect 5680 5564 5684 5596
rect 5716 5564 5720 5596
rect 5680 5516 5720 5564
rect 5680 5484 5684 5516
rect 5716 5484 5720 5516
rect 5680 5436 5720 5484
rect 5680 5404 5684 5436
rect 5716 5404 5720 5436
rect 5680 5356 5720 5404
rect 5680 5324 5684 5356
rect 5716 5324 5720 5356
rect 5680 5276 5720 5324
rect 5680 5244 5684 5276
rect 5716 5244 5720 5276
rect 5680 5196 5720 5244
rect 5680 5164 5684 5196
rect 5716 5164 5720 5196
rect 5680 5116 5720 5164
rect 5680 5084 5684 5116
rect 5716 5084 5720 5116
rect 5680 5036 5720 5084
rect 5680 5004 5684 5036
rect 5716 5004 5720 5036
rect 5680 4956 5720 5004
rect 5680 4924 5684 4956
rect 5716 4924 5720 4956
rect 5680 4876 5720 4924
rect 5680 4844 5684 4876
rect 5716 4844 5720 4876
rect 5680 4796 5720 4844
rect 5680 4764 5684 4796
rect 5716 4764 5720 4796
rect 5680 4716 5720 4764
rect 5680 4684 5684 4716
rect 5716 4684 5720 4716
rect 5680 4636 5720 4684
rect 5680 4604 5684 4636
rect 5716 4604 5720 4636
rect 5680 4556 5720 4604
rect 5680 4524 5684 4556
rect 5716 4524 5720 4556
rect 5680 4476 5720 4524
rect 5680 4444 5684 4476
rect 5716 4444 5720 4476
rect 5680 4396 5720 4444
rect 5680 4364 5684 4396
rect 5716 4364 5720 4396
rect 5680 4316 5720 4364
rect 5680 4284 5684 4316
rect 5716 4284 5720 4316
rect 5680 4236 5720 4284
rect 5680 4204 5684 4236
rect 5716 4204 5720 4236
rect 5680 4156 5720 4204
rect 5680 4124 5684 4156
rect 5716 4124 5720 4156
rect 5680 4076 5720 4124
rect 5680 4044 5684 4076
rect 5716 4044 5720 4076
rect 5680 3996 5720 4044
rect 5680 3964 5684 3996
rect 5716 3964 5720 3996
rect 5680 3916 5720 3964
rect 5680 3884 5684 3916
rect 5716 3884 5720 3916
rect 5680 3836 5720 3884
rect 5680 3804 5684 3836
rect 5716 3804 5720 3836
rect 5680 3756 5720 3804
rect 5680 3724 5684 3756
rect 5716 3724 5720 3756
rect 5680 3676 5720 3724
rect 5680 3644 5684 3676
rect 5716 3644 5720 3676
rect 5680 3596 5720 3644
rect 5680 3564 5684 3596
rect 5716 3564 5720 3596
rect 5680 3516 5720 3564
rect 5680 3484 5684 3516
rect 5716 3484 5720 3516
rect 5680 3436 5720 3484
rect 5680 3404 5684 3436
rect 5716 3404 5720 3436
rect 5680 3356 5720 3404
rect 5680 3324 5684 3356
rect 5716 3324 5720 3356
rect 5680 3276 5720 3324
rect 5680 3244 5684 3276
rect 5716 3244 5720 3276
rect 5680 3196 5720 3244
rect 5680 3164 5684 3196
rect 5716 3164 5720 3196
rect 5680 3116 5720 3164
rect 5680 3084 5684 3116
rect 5716 3084 5720 3116
rect 5680 3036 5720 3084
rect 5680 3004 5684 3036
rect 5716 3004 5720 3036
rect 5680 2956 5720 3004
rect 5680 2924 5684 2956
rect 5716 2924 5720 2956
rect 5680 2876 5720 2924
rect 5680 2844 5684 2876
rect 5716 2844 5720 2876
rect 5680 2796 5720 2844
rect 5680 2764 5684 2796
rect 5716 2764 5720 2796
rect 5680 2716 5720 2764
rect 5680 2684 5684 2716
rect 5716 2684 5720 2716
rect 5680 2636 5720 2684
rect 5680 2604 5684 2636
rect 5716 2604 5720 2636
rect 5680 2556 5720 2604
rect 5680 2524 5684 2556
rect 5716 2524 5720 2556
rect 5680 2476 5720 2524
rect 5680 2444 5684 2476
rect 5716 2444 5720 2476
rect 5680 2396 5720 2444
rect 5680 2364 5684 2396
rect 5716 2364 5720 2396
rect 5680 2316 5720 2364
rect 5680 2284 5684 2316
rect 5716 2284 5720 2316
rect 5680 2236 5720 2284
rect 5680 2204 5684 2236
rect 5716 2204 5720 2236
rect 5680 2156 5720 2204
rect 5680 2124 5684 2156
rect 5716 2124 5720 2156
rect 5680 2076 5720 2124
rect 5680 2044 5684 2076
rect 5716 2044 5720 2076
rect 5680 1996 5720 2044
rect 5680 1964 5684 1996
rect 5716 1964 5720 1996
rect 5680 1916 5720 1964
rect 5680 1884 5684 1916
rect 5716 1884 5720 1916
rect 5680 1836 5720 1884
rect 5680 1804 5684 1836
rect 5716 1804 5720 1836
rect 5680 1756 5720 1804
rect 5680 1724 5684 1756
rect 5716 1724 5720 1756
rect 5680 1676 5720 1724
rect 5680 1644 5684 1676
rect 5716 1644 5720 1676
rect 5680 1596 5720 1644
rect 5680 1564 5684 1596
rect 5716 1564 5720 1596
rect 5680 1516 5720 1564
rect 5680 1484 5684 1516
rect 5716 1484 5720 1516
rect 5680 1436 5720 1484
rect 5680 1404 5684 1436
rect 5716 1404 5720 1436
rect 5680 1356 5720 1404
rect 5680 1324 5684 1356
rect 5716 1324 5720 1356
rect 5680 1276 5720 1324
rect 5680 1244 5684 1276
rect 5716 1244 5720 1276
rect 5680 1196 5720 1244
rect 5680 1164 5684 1196
rect 5716 1164 5720 1196
rect 5680 1116 5720 1164
rect 5680 1084 5684 1116
rect 5716 1084 5720 1116
rect 5680 1036 5720 1084
rect 5680 1004 5684 1036
rect 5716 1004 5720 1036
rect 5680 956 5720 1004
rect 5680 924 5684 956
rect 5716 924 5720 956
rect 5680 876 5720 924
rect 5680 844 5684 876
rect 5716 844 5720 876
rect 5680 796 5720 844
rect 5680 764 5684 796
rect 5716 764 5720 796
rect 5680 716 5720 764
rect 5680 684 5684 716
rect 5716 684 5720 716
rect 5680 636 5720 684
rect 5680 604 5684 636
rect 5716 604 5720 636
rect 5680 556 5720 604
rect 5680 524 5684 556
rect 5716 524 5720 556
rect 5680 476 5720 524
rect 5680 444 5684 476
rect 5716 444 5720 476
rect 5680 396 5720 444
rect 5680 364 5684 396
rect 5716 364 5720 396
rect 5680 316 5720 364
rect 5680 284 5684 316
rect 5716 284 5720 316
rect 5680 236 5720 284
rect 5680 204 5684 236
rect 5716 204 5720 236
rect 5680 156 5720 204
rect 5680 124 5684 156
rect 5716 124 5720 156
rect 5680 76 5720 124
rect 5680 44 5684 76
rect 5716 44 5720 76
rect 5680 -4 5720 44
rect 5680 -36 5684 -4
rect 5716 -36 5720 -4
rect 5680 -84 5720 -36
rect 5680 -116 5684 -84
rect 5716 -116 5720 -84
rect 5680 -120 5720 -116
<< via3 >>
rect -1516 5595 -1484 5596
rect -1516 5565 -1515 5595
rect -1515 5565 -1485 5595
rect -1485 5565 -1484 5595
rect -1516 5564 -1484 5565
rect -1516 5515 -1484 5516
rect -1516 5485 -1515 5515
rect -1515 5485 -1485 5515
rect -1485 5485 -1484 5515
rect -1516 5484 -1484 5485
rect -1516 5435 -1484 5436
rect -1516 5405 -1515 5435
rect -1515 5405 -1485 5435
rect -1485 5405 -1484 5435
rect -1516 5404 -1484 5405
rect -1516 5355 -1484 5356
rect -1516 5325 -1515 5355
rect -1515 5325 -1485 5355
rect -1485 5325 -1484 5355
rect -1516 5324 -1484 5325
rect -1516 5275 -1484 5276
rect -1516 5245 -1515 5275
rect -1515 5245 -1485 5275
rect -1485 5245 -1484 5275
rect -1516 5244 -1484 5245
rect -1516 5195 -1484 5196
rect -1516 5165 -1515 5195
rect -1515 5165 -1485 5195
rect -1485 5165 -1484 5195
rect -1516 5164 -1484 5165
rect -1516 5115 -1484 5116
rect -1516 5085 -1515 5115
rect -1515 5085 -1485 5115
rect -1485 5085 -1484 5115
rect -1516 5084 -1484 5085
rect -1516 5035 -1484 5036
rect -1516 5005 -1515 5035
rect -1515 5005 -1485 5035
rect -1485 5005 -1484 5035
rect -1516 5004 -1484 5005
rect -1516 4955 -1484 4956
rect -1516 4925 -1515 4955
rect -1515 4925 -1485 4955
rect -1485 4925 -1484 4955
rect -1516 4924 -1484 4925
rect -1516 4875 -1484 4876
rect -1516 4845 -1515 4875
rect -1515 4845 -1485 4875
rect -1485 4845 -1484 4875
rect -1516 4844 -1484 4845
rect -1516 4764 -1484 4796
rect -1516 4715 -1484 4716
rect -1516 4685 -1515 4715
rect -1515 4685 -1485 4715
rect -1485 4685 -1484 4715
rect -1516 4684 -1484 4685
rect -1516 4635 -1484 4636
rect -1516 4605 -1515 4635
rect -1515 4605 -1485 4635
rect -1485 4605 -1484 4635
rect -1516 4604 -1484 4605
rect -1516 4555 -1484 4556
rect -1516 4525 -1515 4555
rect -1515 4525 -1485 4555
rect -1485 4525 -1484 4555
rect -1516 4524 -1484 4525
rect -1516 4475 -1484 4476
rect -1516 4445 -1515 4475
rect -1515 4445 -1485 4475
rect -1485 4445 -1484 4475
rect -1516 4444 -1484 4445
rect -1516 4395 -1484 4396
rect -1516 4365 -1515 4395
rect -1515 4365 -1485 4395
rect -1485 4365 -1484 4395
rect -1516 4364 -1484 4365
rect -1516 4315 -1484 4316
rect -1516 4285 -1515 4315
rect -1515 4285 -1485 4315
rect -1485 4285 -1484 4315
rect -1516 4284 -1484 4285
rect -1516 4235 -1484 4236
rect -1516 4205 -1515 4235
rect -1515 4205 -1485 4235
rect -1485 4205 -1484 4235
rect -1516 4204 -1484 4205
rect -1516 4155 -1484 4156
rect -1516 4125 -1515 4155
rect -1515 4125 -1485 4155
rect -1485 4125 -1484 4155
rect -1516 4124 -1484 4125
rect -1516 4075 -1484 4076
rect -1516 4045 -1515 4075
rect -1515 4045 -1485 4075
rect -1485 4045 -1484 4075
rect -1516 4044 -1484 4045
rect -1516 3995 -1484 3996
rect -1516 3965 -1515 3995
rect -1515 3965 -1485 3995
rect -1485 3965 -1484 3995
rect -1516 3964 -1484 3965
rect -1516 3915 -1484 3916
rect -1516 3885 -1515 3915
rect -1515 3885 -1485 3915
rect -1485 3885 -1484 3915
rect -1516 3884 -1484 3885
rect -1516 3835 -1484 3836
rect -1516 3805 -1515 3835
rect -1515 3805 -1485 3835
rect -1485 3805 -1484 3835
rect -1516 3804 -1484 3805
rect -1516 3755 -1484 3756
rect -1516 3725 -1515 3755
rect -1515 3725 -1485 3755
rect -1485 3725 -1484 3755
rect -1516 3724 -1484 3725
rect -1516 3675 -1484 3676
rect -1516 3645 -1515 3675
rect -1515 3645 -1485 3675
rect -1485 3645 -1484 3675
rect -1516 3644 -1484 3645
rect -1516 3595 -1484 3596
rect -1516 3565 -1515 3595
rect -1515 3565 -1485 3595
rect -1485 3565 -1484 3595
rect -1516 3564 -1484 3565
rect -1516 3515 -1484 3516
rect -1516 3485 -1515 3515
rect -1515 3485 -1485 3515
rect -1485 3485 -1484 3515
rect -1516 3484 -1484 3485
rect -1516 3435 -1484 3436
rect -1516 3405 -1515 3435
rect -1515 3405 -1485 3435
rect -1485 3405 -1484 3435
rect -1516 3404 -1484 3405
rect -1516 3355 -1484 3356
rect -1516 3325 -1515 3355
rect -1515 3325 -1485 3355
rect -1485 3325 -1484 3355
rect -1516 3324 -1484 3325
rect -1516 3275 -1484 3276
rect -1516 3245 -1515 3275
rect -1515 3245 -1485 3275
rect -1485 3245 -1484 3275
rect -1516 3244 -1484 3245
rect -1516 3195 -1484 3196
rect -1516 3165 -1515 3195
rect -1515 3165 -1485 3195
rect -1485 3165 -1484 3195
rect -1516 3164 -1484 3165
rect -1516 3115 -1484 3116
rect -1516 3085 -1515 3115
rect -1515 3085 -1485 3115
rect -1485 3085 -1484 3115
rect -1516 3084 -1484 3085
rect -1516 3035 -1484 3036
rect -1516 3005 -1515 3035
rect -1515 3005 -1485 3035
rect -1485 3005 -1484 3035
rect -1516 3004 -1484 3005
rect -1516 2955 -1484 2956
rect -1516 2925 -1515 2955
rect -1515 2925 -1485 2955
rect -1485 2925 -1484 2955
rect -1516 2924 -1484 2925
rect -1516 2875 -1484 2876
rect -1516 2845 -1515 2875
rect -1515 2845 -1485 2875
rect -1485 2845 -1484 2875
rect -1516 2844 -1484 2845
rect -1516 2795 -1484 2796
rect -1516 2765 -1515 2795
rect -1515 2765 -1485 2795
rect -1485 2765 -1484 2795
rect -1516 2764 -1484 2765
rect -1516 2715 -1484 2716
rect -1516 2685 -1515 2715
rect -1515 2685 -1485 2715
rect -1485 2685 -1484 2715
rect -1516 2684 -1484 2685
rect -1516 2635 -1484 2636
rect -1516 2605 -1515 2635
rect -1515 2605 -1485 2635
rect -1485 2605 -1484 2635
rect -1516 2604 -1484 2605
rect -1516 2555 -1484 2556
rect -1516 2525 -1515 2555
rect -1515 2525 -1485 2555
rect -1485 2525 -1484 2555
rect -1516 2524 -1484 2525
rect -1516 2475 -1484 2476
rect -1516 2445 -1515 2475
rect -1515 2445 -1485 2475
rect -1485 2445 -1484 2475
rect -1516 2444 -1484 2445
rect -1516 2395 -1484 2396
rect -1516 2365 -1515 2395
rect -1515 2365 -1485 2395
rect -1485 2365 -1484 2395
rect -1516 2364 -1484 2365
rect -1516 2315 -1484 2316
rect -1516 2285 -1515 2315
rect -1515 2285 -1485 2315
rect -1485 2285 -1484 2315
rect -1516 2284 -1484 2285
rect -1516 2235 -1484 2236
rect -1516 2205 -1515 2235
rect -1515 2205 -1485 2235
rect -1485 2205 -1484 2235
rect -1516 2204 -1484 2205
rect -1516 2155 -1484 2156
rect -1516 2125 -1515 2155
rect -1515 2125 -1485 2155
rect -1485 2125 -1484 2155
rect -1516 2124 -1484 2125
rect -1516 2075 -1484 2076
rect -1516 2045 -1515 2075
rect -1515 2045 -1485 2075
rect -1485 2045 -1484 2075
rect -1516 2044 -1484 2045
rect -1516 1995 -1484 1996
rect -1516 1965 -1515 1995
rect -1515 1965 -1485 1995
rect -1485 1965 -1484 1995
rect -1516 1964 -1484 1965
rect -1516 1915 -1484 1916
rect -1516 1885 -1515 1915
rect -1515 1885 -1485 1915
rect -1485 1885 -1484 1915
rect -1516 1884 -1484 1885
rect -1516 1835 -1484 1836
rect -1516 1805 -1515 1835
rect -1515 1805 -1485 1835
rect -1485 1805 -1484 1835
rect -1516 1804 -1484 1805
rect -1516 1755 -1484 1756
rect -1516 1725 -1515 1755
rect -1515 1725 -1485 1755
rect -1485 1725 -1484 1755
rect -1516 1724 -1484 1725
rect -1516 1675 -1484 1676
rect -1516 1645 -1515 1675
rect -1515 1645 -1485 1675
rect -1485 1645 -1484 1675
rect -1516 1644 -1484 1645
rect -1516 1595 -1484 1596
rect -1516 1565 -1515 1595
rect -1515 1565 -1485 1595
rect -1485 1565 -1484 1595
rect -1516 1564 -1484 1565
rect -1516 1515 -1484 1516
rect -1516 1485 -1515 1515
rect -1515 1485 -1485 1515
rect -1485 1485 -1484 1515
rect -1516 1484 -1484 1485
rect -1516 1435 -1484 1436
rect -1516 1405 -1515 1435
rect -1515 1405 -1485 1435
rect -1485 1405 -1484 1435
rect -1516 1404 -1484 1405
rect -1516 1355 -1484 1356
rect -1516 1325 -1515 1355
rect -1515 1325 -1485 1355
rect -1485 1325 -1484 1355
rect -1516 1324 -1484 1325
rect -1516 1275 -1484 1276
rect -1516 1245 -1515 1275
rect -1515 1245 -1485 1275
rect -1485 1245 -1484 1275
rect -1516 1244 -1484 1245
rect -1516 1195 -1484 1196
rect -1516 1165 -1515 1195
rect -1515 1165 -1485 1195
rect -1485 1165 -1484 1195
rect -1516 1164 -1484 1165
rect -1516 1115 -1484 1116
rect -1516 1085 -1515 1115
rect -1515 1085 -1485 1115
rect -1485 1085 -1484 1115
rect -1516 1084 -1484 1085
rect -1516 1035 -1484 1036
rect -1516 1005 -1515 1035
rect -1515 1005 -1485 1035
rect -1485 1005 -1484 1035
rect -1516 1004 -1484 1005
rect -1516 955 -1484 956
rect -1516 925 -1515 955
rect -1515 925 -1485 955
rect -1485 925 -1484 955
rect -1516 924 -1484 925
rect -1516 875 -1484 876
rect -1516 845 -1515 875
rect -1515 845 -1485 875
rect -1485 845 -1484 875
rect -1516 844 -1484 845
rect -1516 795 -1484 796
rect -1516 765 -1515 795
rect -1515 765 -1485 795
rect -1485 765 -1484 795
rect -1516 764 -1484 765
rect -1516 715 -1484 716
rect -1516 685 -1515 715
rect -1515 685 -1485 715
rect -1485 685 -1484 715
rect -1516 684 -1484 685
rect -1516 635 -1484 636
rect -1516 605 -1515 635
rect -1515 605 -1485 635
rect -1485 605 -1484 635
rect -1516 604 -1484 605
rect -1516 555 -1484 556
rect -1516 525 -1515 555
rect -1515 525 -1485 555
rect -1485 525 -1484 555
rect -1516 524 -1484 525
rect -1516 475 -1484 476
rect -1516 445 -1515 475
rect -1515 445 -1485 475
rect -1485 445 -1484 475
rect -1516 444 -1484 445
rect -1516 395 -1484 396
rect -1516 365 -1515 395
rect -1515 365 -1485 395
rect -1485 365 -1484 395
rect -1516 364 -1484 365
rect -1516 315 -1484 316
rect -1516 285 -1515 315
rect -1515 285 -1485 315
rect -1485 285 -1484 315
rect -1516 284 -1484 285
rect -1516 235 -1484 236
rect -1516 205 -1515 235
rect -1515 205 -1485 235
rect -1485 205 -1484 235
rect -1516 204 -1484 205
rect -1516 155 -1484 156
rect -1516 125 -1515 155
rect -1515 125 -1485 155
rect -1485 125 -1484 155
rect -1516 124 -1484 125
rect -1516 75 -1484 76
rect -1516 45 -1515 75
rect -1515 45 -1485 75
rect -1485 45 -1484 75
rect -1516 44 -1484 45
rect -1516 -5 -1484 -4
rect -1516 -35 -1515 -5
rect -1515 -35 -1485 -5
rect -1485 -35 -1484 -5
rect -1516 -36 -1484 -35
rect -1516 -85 -1484 -84
rect -1516 -115 -1515 -85
rect -1515 -115 -1485 -85
rect -1485 -115 -1484 -85
rect -1516 -116 -1484 -115
rect -1356 5595 -1324 5596
rect -1356 5565 -1355 5595
rect -1355 5565 -1325 5595
rect -1325 5565 -1324 5595
rect -1356 5564 -1324 5565
rect -1356 5515 -1324 5516
rect -1356 5485 -1355 5515
rect -1355 5485 -1325 5515
rect -1325 5485 -1324 5515
rect -1356 5484 -1324 5485
rect -1356 5435 -1324 5436
rect -1356 5405 -1355 5435
rect -1355 5405 -1325 5435
rect -1325 5405 -1324 5435
rect -1356 5404 -1324 5405
rect -1356 5355 -1324 5356
rect -1356 5325 -1355 5355
rect -1355 5325 -1325 5355
rect -1325 5325 -1324 5355
rect -1356 5324 -1324 5325
rect -1356 5275 -1324 5276
rect -1356 5245 -1355 5275
rect -1355 5245 -1325 5275
rect -1325 5245 -1324 5275
rect -1356 5244 -1324 5245
rect -1356 5195 -1324 5196
rect -1356 5165 -1355 5195
rect -1355 5165 -1325 5195
rect -1325 5165 -1324 5195
rect -1356 5164 -1324 5165
rect -1356 5115 -1324 5116
rect -1356 5085 -1355 5115
rect -1355 5085 -1325 5115
rect -1325 5085 -1324 5115
rect -1356 5084 -1324 5085
rect -1356 5035 -1324 5036
rect -1356 5005 -1355 5035
rect -1355 5005 -1325 5035
rect -1325 5005 -1324 5035
rect -1356 5004 -1324 5005
rect -1356 4955 -1324 4956
rect -1356 4925 -1355 4955
rect -1355 4925 -1325 4955
rect -1325 4925 -1324 4955
rect -1356 4924 -1324 4925
rect -1356 4875 -1324 4876
rect -1356 4845 -1355 4875
rect -1355 4845 -1325 4875
rect -1325 4845 -1324 4875
rect -1356 4844 -1324 4845
rect -1356 4764 -1324 4796
rect -1356 4715 -1324 4716
rect -1356 4685 -1355 4715
rect -1355 4685 -1325 4715
rect -1325 4685 -1324 4715
rect -1356 4684 -1324 4685
rect -1356 4635 -1324 4636
rect -1356 4605 -1355 4635
rect -1355 4605 -1325 4635
rect -1325 4605 -1324 4635
rect -1356 4604 -1324 4605
rect -1356 4555 -1324 4556
rect -1356 4525 -1355 4555
rect -1355 4525 -1325 4555
rect -1325 4525 -1324 4555
rect -1356 4524 -1324 4525
rect -1356 4475 -1324 4476
rect -1356 4445 -1355 4475
rect -1355 4445 -1325 4475
rect -1325 4445 -1324 4475
rect -1356 4444 -1324 4445
rect -1356 4395 -1324 4396
rect -1356 4365 -1355 4395
rect -1355 4365 -1325 4395
rect -1325 4365 -1324 4395
rect -1356 4364 -1324 4365
rect -1356 4315 -1324 4316
rect -1356 4285 -1355 4315
rect -1355 4285 -1325 4315
rect -1325 4285 -1324 4315
rect -1356 4284 -1324 4285
rect -1356 4235 -1324 4236
rect -1356 4205 -1355 4235
rect -1355 4205 -1325 4235
rect -1325 4205 -1324 4235
rect -1356 4204 -1324 4205
rect -1356 4155 -1324 4156
rect -1356 4125 -1355 4155
rect -1355 4125 -1325 4155
rect -1325 4125 -1324 4155
rect -1356 4124 -1324 4125
rect -1356 4075 -1324 4076
rect -1356 4045 -1355 4075
rect -1355 4045 -1325 4075
rect -1325 4045 -1324 4075
rect -1356 4044 -1324 4045
rect -1356 3995 -1324 3996
rect -1356 3965 -1355 3995
rect -1355 3965 -1325 3995
rect -1325 3965 -1324 3995
rect -1356 3964 -1324 3965
rect -1356 3915 -1324 3916
rect -1356 3885 -1355 3915
rect -1355 3885 -1325 3915
rect -1325 3885 -1324 3915
rect -1356 3884 -1324 3885
rect -1356 3835 -1324 3836
rect -1356 3805 -1355 3835
rect -1355 3805 -1325 3835
rect -1325 3805 -1324 3835
rect -1356 3804 -1324 3805
rect -1356 3755 -1324 3756
rect -1356 3725 -1355 3755
rect -1355 3725 -1325 3755
rect -1325 3725 -1324 3755
rect -1356 3724 -1324 3725
rect -1356 3675 -1324 3676
rect -1356 3645 -1355 3675
rect -1355 3645 -1325 3675
rect -1325 3645 -1324 3675
rect -1356 3644 -1324 3645
rect -1356 3595 -1324 3596
rect -1356 3565 -1355 3595
rect -1355 3565 -1325 3595
rect -1325 3565 -1324 3595
rect -1356 3564 -1324 3565
rect -1356 3515 -1324 3516
rect -1356 3485 -1355 3515
rect -1355 3485 -1325 3515
rect -1325 3485 -1324 3515
rect -1356 3484 -1324 3485
rect -1356 3435 -1324 3436
rect -1356 3405 -1355 3435
rect -1355 3405 -1325 3435
rect -1325 3405 -1324 3435
rect -1356 3404 -1324 3405
rect -1356 3355 -1324 3356
rect -1356 3325 -1355 3355
rect -1355 3325 -1325 3355
rect -1325 3325 -1324 3355
rect -1356 3324 -1324 3325
rect -1356 3275 -1324 3276
rect -1356 3245 -1355 3275
rect -1355 3245 -1325 3275
rect -1325 3245 -1324 3275
rect -1356 3244 -1324 3245
rect -1356 3195 -1324 3196
rect -1356 3165 -1355 3195
rect -1355 3165 -1325 3195
rect -1325 3165 -1324 3195
rect -1356 3164 -1324 3165
rect -1356 3115 -1324 3116
rect -1356 3085 -1355 3115
rect -1355 3085 -1325 3115
rect -1325 3085 -1324 3115
rect -1356 3084 -1324 3085
rect -1356 3035 -1324 3036
rect -1356 3005 -1355 3035
rect -1355 3005 -1325 3035
rect -1325 3005 -1324 3035
rect -1356 3004 -1324 3005
rect -1356 2955 -1324 2956
rect -1356 2925 -1355 2955
rect -1355 2925 -1325 2955
rect -1325 2925 -1324 2955
rect -1356 2924 -1324 2925
rect -1356 2875 -1324 2876
rect -1356 2845 -1355 2875
rect -1355 2845 -1325 2875
rect -1325 2845 -1324 2875
rect -1356 2844 -1324 2845
rect -1356 2795 -1324 2796
rect -1356 2765 -1355 2795
rect -1355 2765 -1325 2795
rect -1325 2765 -1324 2795
rect -1356 2764 -1324 2765
rect -1356 2715 -1324 2716
rect -1356 2685 -1355 2715
rect -1355 2685 -1325 2715
rect -1325 2685 -1324 2715
rect -1356 2684 -1324 2685
rect -1356 2635 -1324 2636
rect -1356 2605 -1355 2635
rect -1355 2605 -1325 2635
rect -1325 2605 -1324 2635
rect -1356 2604 -1324 2605
rect -1356 2555 -1324 2556
rect -1356 2525 -1355 2555
rect -1355 2525 -1325 2555
rect -1325 2525 -1324 2555
rect -1356 2524 -1324 2525
rect -1356 2475 -1324 2476
rect -1356 2445 -1355 2475
rect -1355 2445 -1325 2475
rect -1325 2445 -1324 2475
rect -1356 2444 -1324 2445
rect -1356 2395 -1324 2396
rect -1356 2365 -1355 2395
rect -1355 2365 -1325 2395
rect -1325 2365 -1324 2395
rect -1356 2364 -1324 2365
rect -1356 2315 -1324 2316
rect -1356 2285 -1355 2315
rect -1355 2285 -1325 2315
rect -1325 2285 -1324 2315
rect -1356 2284 -1324 2285
rect -1356 2235 -1324 2236
rect -1356 2205 -1355 2235
rect -1355 2205 -1325 2235
rect -1325 2205 -1324 2235
rect -1356 2204 -1324 2205
rect -1356 2155 -1324 2156
rect -1356 2125 -1355 2155
rect -1355 2125 -1325 2155
rect -1325 2125 -1324 2155
rect -1356 2124 -1324 2125
rect -1356 2075 -1324 2076
rect -1356 2045 -1355 2075
rect -1355 2045 -1325 2075
rect -1325 2045 -1324 2075
rect -1356 2044 -1324 2045
rect -1356 1995 -1324 1996
rect -1356 1965 -1355 1995
rect -1355 1965 -1325 1995
rect -1325 1965 -1324 1995
rect -1356 1964 -1324 1965
rect -1356 1915 -1324 1916
rect -1356 1885 -1355 1915
rect -1355 1885 -1325 1915
rect -1325 1885 -1324 1915
rect -1356 1884 -1324 1885
rect -1356 1835 -1324 1836
rect -1356 1805 -1355 1835
rect -1355 1805 -1325 1835
rect -1325 1805 -1324 1835
rect -1356 1804 -1324 1805
rect -1356 1755 -1324 1756
rect -1356 1725 -1355 1755
rect -1355 1725 -1325 1755
rect -1325 1725 -1324 1755
rect -1356 1724 -1324 1725
rect -1356 1675 -1324 1676
rect -1356 1645 -1355 1675
rect -1355 1645 -1325 1675
rect -1325 1645 -1324 1675
rect -1356 1644 -1324 1645
rect -1356 1595 -1324 1596
rect -1356 1565 -1355 1595
rect -1355 1565 -1325 1595
rect -1325 1565 -1324 1595
rect -1356 1564 -1324 1565
rect -1356 1515 -1324 1516
rect -1356 1485 -1355 1515
rect -1355 1485 -1325 1515
rect -1325 1485 -1324 1515
rect -1356 1484 -1324 1485
rect -1356 1435 -1324 1436
rect -1356 1405 -1355 1435
rect -1355 1405 -1325 1435
rect -1325 1405 -1324 1435
rect -1356 1404 -1324 1405
rect -1356 1355 -1324 1356
rect -1356 1325 -1355 1355
rect -1355 1325 -1325 1355
rect -1325 1325 -1324 1355
rect -1356 1324 -1324 1325
rect -1356 1275 -1324 1276
rect -1356 1245 -1355 1275
rect -1355 1245 -1325 1275
rect -1325 1245 -1324 1275
rect -1356 1244 -1324 1245
rect -1356 1195 -1324 1196
rect -1356 1165 -1355 1195
rect -1355 1165 -1325 1195
rect -1325 1165 -1324 1195
rect -1356 1164 -1324 1165
rect -1356 1115 -1324 1116
rect -1356 1085 -1355 1115
rect -1355 1085 -1325 1115
rect -1325 1085 -1324 1115
rect -1356 1084 -1324 1085
rect -1356 1035 -1324 1036
rect -1356 1005 -1355 1035
rect -1355 1005 -1325 1035
rect -1325 1005 -1324 1035
rect -1356 1004 -1324 1005
rect -1356 955 -1324 956
rect -1356 925 -1355 955
rect -1355 925 -1325 955
rect -1325 925 -1324 955
rect -1356 924 -1324 925
rect -1356 875 -1324 876
rect -1356 845 -1355 875
rect -1355 845 -1325 875
rect -1325 845 -1324 875
rect -1356 844 -1324 845
rect -1356 795 -1324 796
rect -1356 765 -1355 795
rect -1355 765 -1325 795
rect -1325 765 -1324 795
rect -1356 764 -1324 765
rect -1356 715 -1324 716
rect -1356 685 -1355 715
rect -1355 685 -1325 715
rect -1325 685 -1324 715
rect -1356 684 -1324 685
rect -1356 635 -1324 636
rect -1356 605 -1355 635
rect -1355 605 -1325 635
rect -1325 605 -1324 635
rect -1356 604 -1324 605
rect -1356 555 -1324 556
rect -1356 525 -1355 555
rect -1355 525 -1325 555
rect -1325 525 -1324 555
rect -1356 524 -1324 525
rect -1356 475 -1324 476
rect -1356 445 -1355 475
rect -1355 445 -1325 475
rect -1325 445 -1324 475
rect -1356 444 -1324 445
rect -1356 395 -1324 396
rect -1356 365 -1355 395
rect -1355 365 -1325 395
rect -1325 365 -1324 395
rect -1356 364 -1324 365
rect -1356 315 -1324 316
rect -1356 285 -1355 315
rect -1355 285 -1325 315
rect -1325 285 -1324 315
rect -1356 284 -1324 285
rect -1356 235 -1324 236
rect -1356 205 -1355 235
rect -1355 205 -1325 235
rect -1325 205 -1324 235
rect -1356 204 -1324 205
rect -1356 155 -1324 156
rect -1356 125 -1355 155
rect -1355 125 -1325 155
rect -1325 125 -1324 155
rect -1356 124 -1324 125
rect -1356 75 -1324 76
rect -1356 45 -1355 75
rect -1355 45 -1325 75
rect -1325 45 -1324 75
rect -1356 44 -1324 45
rect -1356 -5 -1324 -4
rect -1356 -35 -1355 -5
rect -1355 -35 -1325 -5
rect -1325 -35 -1324 -5
rect -1356 -36 -1324 -35
rect -1356 -85 -1324 -84
rect -1356 -115 -1355 -85
rect -1355 -115 -1325 -85
rect -1325 -115 -1324 -85
rect -1356 -116 -1324 -115
rect -1196 5595 -1164 5596
rect -1196 5565 -1195 5595
rect -1195 5565 -1165 5595
rect -1165 5565 -1164 5595
rect -1196 5564 -1164 5565
rect -1196 5515 -1164 5516
rect -1196 5485 -1195 5515
rect -1195 5485 -1165 5515
rect -1165 5485 -1164 5515
rect -1196 5484 -1164 5485
rect -1196 5435 -1164 5436
rect -1196 5405 -1195 5435
rect -1195 5405 -1165 5435
rect -1165 5405 -1164 5435
rect -1196 5404 -1164 5405
rect -1196 5355 -1164 5356
rect -1196 5325 -1195 5355
rect -1195 5325 -1165 5355
rect -1165 5325 -1164 5355
rect -1196 5324 -1164 5325
rect -1196 5275 -1164 5276
rect -1196 5245 -1195 5275
rect -1195 5245 -1165 5275
rect -1165 5245 -1164 5275
rect -1196 5244 -1164 5245
rect -1196 5195 -1164 5196
rect -1196 5165 -1195 5195
rect -1195 5165 -1165 5195
rect -1165 5165 -1164 5195
rect -1196 5164 -1164 5165
rect -1196 5115 -1164 5116
rect -1196 5085 -1195 5115
rect -1195 5085 -1165 5115
rect -1165 5085 -1164 5115
rect -1196 5084 -1164 5085
rect -1196 5035 -1164 5036
rect -1196 5005 -1195 5035
rect -1195 5005 -1165 5035
rect -1165 5005 -1164 5035
rect -1196 5004 -1164 5005
rect -1196 4955 -1164 4956
rect -1196 4925 -1195 4955
rect -1195 4925 -1165 4955
rect -1165 4925 -1164 4955
rect -1196 4924 -1164 4925
rect -1196 4875 -1164 4876
rect -1196 4845 -1195 4875
rect -1195 4845 -1165 4875
rect -1165 4845 -1164 4875
rect -1196 4844 -1164 4845
rect -1196 4764 -1164 4796
rect -1196 4715 -1164 4716
rect -1196 4685 -1195 4715
rect -1195 4685 -1165 4715
rect -1165 4685 -1164 4715
rect -1196 4684 -1164 4685
rect -1196 4635 -1164 4636
rect -1196 4605 -1195 4635
rect -1195 4605 -1165 4635
rect -1165 4605 -1164 4635
rect -1196 4604 -1164 4605
rect -1196 4555 -1164 4556
rect -1196 4525 -1195 4555
rect -1195 4525 -1165 4555
rect -1165 4525 -1164 4555
rect -1196 4524 -1164 4525
rect -1196 4475 -1164 4476
rect -1196 4445 -1195 4475
rect -1195 4445 -1165 4475
rect -1165 4445 -1164 4475
rect -1196 4444 -1164 4445
rect -1196 4395 -1164 4396
rect -1196 4365 -1195 4395
rect -1195 4365 -1165 4395
rect -1165 4365 -1164 4395
rect -1196 4364 -1164 4365
rect -1196 4315 -1164 4316
rect -1196 4285 -1195 4315
rect -1195 4285 -1165 4315
rect -1165 4285 -1164 4315
rect -1196 4284 -1164 4285
rect -1196 4235 -1164 4236
rect -1196 4205 -1195 4235
rect -1195 4205 -1165 4235
rect -1165 4205 -1164 4235
rect -1196 4204 -1164 4205
rect -1196 4155 -1164 4156
rect -1196 4125 -1195 4155
rect -1195 4125 -1165 4155
rect -1165 4125 -1164 4155
rect -1196 4124 -1164 4125
rect -1196 4075 -1164 4076
rect -1196 4045 -1195 4075
rect -1195 4045 -1165 4075
rect -1165 4045 -1164 4075
rect -1196 4044 -1164 4045
rect -1196 3995 -1164 3996
rect -1196 3965 -1195 3995
rect -1195 3965 -1165 3995
rect -1165 3965 -1164 3995
rect -1196 3964 -1164 3965
rect -1196 3915 -1164 3916
rect -1196 3885 -1195 3915
rect -1195 3885 -1165 3915
rect -1165 3885 -1164 3915
rect -1196 3884 -1164 3885
rect -1196 3835 -1164 3836
rect -1196 3805 -1195 3835
rect -1195 3805 -1165 3835
rect -1165 3805 -1164 3835
rect -1196 3804 -1164 3805
rect -1196 3755 -1164 3756
rect -1196 3725 -1195 3755
rect -1195 3725 -1165 3755
rect -1165 3725 -1164 3755
rect -1196 3724 -1164 3725
rect -1196 3675 -1164 3676
rect -1196 3645 -1195 3675
rect -1195 3645 -1165 3675
rect -1165 3645 -1164 3675
rect -1196 3644 -1164 3645
rect -1196 3595 -1164 3596
rect -1196 3565 -1195 3595
rect -1195 3565 -1165 3595
rect -1165 3565 -1164 3595
rect -1196 3564 -1164 3565
rect -1196 3515 -1164 3516
rect -1196 3485 -1195 3515
rect -1195 3485 -1165 3515
rect -1165 3485 -1164 3515
rect -1196 3484 -1164 3485
rect -1196 3404 -1164 3436
rect -1196 3355 -1164 3356
rect -1196 3325 -1195 3355
rect -1195 3325 -1165 3355
rect -1165 3325 -1164 3355
rect -1196 3324 -1164 3325
rect -1196 3275 -1164 3276
rect -1196 3245 -1195 3275
rect -1195 3245 -1165 3275
rect -1165 3245 -1164 3275
rect -1196 3244 -1164 3245
rect -1196 3195 -1164 3196
rect -1196 3165 -1195 3195
rect -1195 3165 -1165 3195
rect -1165 3165 -1164 3195
rect -1196 3164 -1164 3165
rect -1196 3115 -1164 3116
rect -1196 3085 -1195 3115
rect -1195 3085 -1165 3115
rect -1165 3085 -1164 3115
rect -1196 3084 -1164 3085
rect -1196 3035 -1164 3036
rect -1196 3005 -1195 3035
rect -1195 3005 -1165 3035
rect -1165 3005 -1164 3035
rect -1196 3004 -1164 3005
rect -1196 2955 -1164 2956
rect -1196 2925 -1195 2955
rect -1195 2925 -1165 2955
rect -1165 2925 -1164 2955
rect -1196 2924 -1164 2925
rect -1196 2875 -1164 2876
rect -1196 2845 -1195 2875
rect -1195 2845 -1165 2875
rect -1165 2845 -1164 2875
rect -1196 2844 -1164 2845
rect -1196 2795 -1164 2796
rect -1196 2765 -1195 2795
rect -1195 2765 -1165 2795
rect -1165 2765 -1164 2795
rect -1196 2764 -1164 2765
rect -1196 2715 -1164 2716
rect -1196 2685 -1195 2715
rect -1195 2685 -1165 2715
rect -1165 2685 -1164 2715
rect -1196 2684 -1164 2685
rect -1196 2604 -1164 2636
rect -1196 2555 -1164 2556
rect -1196 2525 -1195 2555
rect -1195 2525 -1165 2555
rect -1165 2525 -1164 2555
rect -1196 2524 -1164 2525
rect -1196 2475 -1164 2476
rect -1196 2445 -1195 2475
rect -1195 2445 -1165 2475
rect -1165 2445 -1164 2475
rect -1196 2444 -1164 2445
rect -1196 2395 -1164 2396
rect -1196 2365 -1195 2395
rect -1195 2365 -1165 2395
rect -1165 2365 -1164 2395
rect -1196 2364 -1164 2365
rect -1196 2315 -1164 2316
rect -1196 2285 -1195 2315
rect -1195 2285 -1165 2315
rect -1165 2285 -1164 2315
rect -1196 2284 -1164 2285
rect -1196 2235 -1164 2236
rect -1196 2205 -1195 2235
rect -1195 2205 -1165 2235
rect -1165 2205 -1164 2235
rect -1196 2204 -1164 2205
rect -1196 2155 -1164 2156
rect -1196 2125 -1195 2155
rect -1195 2125 -1165 2155
rect -1165 2125 -1164 2155
rect -1196 2124 -1164 2125
rect -1196 2075 -1164 2076
rect -1196 2045 -1195 2075
rect -1195 2045 -1165 2075
rect -1165 2045 -1164 2075
rect -1196 2044 -1164 2045
rect -1196 1995 -1164 1996
rect -1196 1965 -1195 1995
rect -1195 1965 -1165 1995
rect -1165 1965 -1164 1995
rect -1196 1964 -1164 1965
rect -1196 1915 -1164 1916
rect -1196 1885 -1195 1915
rect -1195 1885 -1165 1915
rect -1165 1885 -1164 1915
rect -1196 1884 -1164 1885
rect -1196 1835 -1164 1836
rect -1196 1805 -1195 1835
rect -1195 1805 -1165 1835
rect -1165 1805 -1164 1835
rect -1196 1804 -1164 1805
rect -1196 1755 -1164 1756
rect -1196 1725 -1195 1755
rect -1195 1725 -1165 1755
rect -1165 1725 -1164 1755
rect -1196 1724 -1164 1725
rect -1196 1675 -1164 1676
rect -1196 1645 -1195 1675
rect -1195 1645 -1165 1675
rect -1165 1645 -1164 1675
rect -1196 1644 -1164 1645
rect -1196 1595 -1164 1596
rect -1196 1565 -1195 1595
rect -1195 1565 -1165 1595
rect -1165 1565 -1164 1595
rect -1196 1564 -1164 1565
rect -1196 1515 -1164 1516
rect -1196 1485 -1195 1515
rect -1195 1485 -1165 1515
rect -1165 1485 -1164 1515
rect -1196 1484 -1164 1485
rect -1196 1435 -1164 1436
rect -1196 1405 -1195 1435
rect -1195 1405 -1165 1435
rect -1165 1405 -1164 1435
rect -1196 1404 -1164 1405
rect -1196 1355 -1164 1356
rect -1196 1325 -1195 1355
rect -1195 1325 -1165 1355
rect -1165 1325 -1164 1355
rect -1196 1324 -1164 1325
rect -1196 1275 -1164 1276
rect -1196 1245 -1195 1275
rect -1195 1245 -1165 1275
rect -1165 1245 -1164 1275
rect -1196 1244 -1164 1245
rect -1196 1195 -1164 1196
rect -1196 1165 -1195 1195
rect -1195 1165 -1165 1195
rect -1165 1165 -1164 1195
rect -1196 1164 -1164 1165
rect -1196 1115 -1164 1116
rect -1196 1085 -1195 1115
rect -1195 1085 -1165 1115
rect -1165 1085 -1164 1115
rect -1196 1084 -1164 1085
rect -1196 1035 -1164 1036
rect -1196 1005 -1195 1035
rect -1195 1005 -1165 1035
rect -1165 1005 -1164 1035
rect -1196 1004 -1164 1005
rect -1196 955 -1164 956
rect -1196 925 -1195 955
rect -1195 925 -1165 955
rect -1165 925 -1164 955
rect -1196 924 -1164 925
rect -1196 875 -1164 876
rect -1196 845 -1195 875
rect -1195 845 -1165 875
rect -1165 845 -1164 875
rect -1196 844 -1164 845
rect -1196 795 -1164 796
rect -1196 765 -1195 795
rect -1195 765 -1165 795
rect -1165 765 -1164 795
rect -1196 764 -1164 765
rect -1196 715 -1164 716
rect -1196 685 -1195 715
rect -1195 685 -1165 715
rect -1165 685 -1164 715
rect -1196 684 -1164 685
rect -1196 635 -1164 636
rect -1196 605 -1195 635
rect -1195 605 -1165 635
rect -1165 605 -1164 635
rect -1196 604 -1164 605
rect -1196 555 -1164 556
rect -1196 525 -1195 555
rect -1195 525 -1165 555
rect -1165 525 -1164 555
rect -1196 524 -1164 525
rect -1196 475 -1164 476
rect -1196 445 -1195 475
rect -1195 445 -1165 475
rect -1165 445 -1164 475
rect -1196 444 -1164 445
rect -1196 395 -1164 396
rect -1196 365 -1195 395
rect -1195 365 -1165 395
rect -1165 365 -1164 395
rect -1196 364 -1164 365
rect -1196 315 -1164 316
rect -1196 285 -1195 315
rect -1195 285 -1165 315
rect -1165 285 -1164 315
rect -1196 284 -1164 285
rect -1196 235 -1164 236
rect -1196 205 -1195 235
rect -1195 205 -1165 235
rect -1165 205 -1164 235
rect -1196 204 -1164 205
rect -1196 155 -1164 156
rect -1196 125 -1195 155
rect -1195 125 -1165 155
rect -1165 125 -1164 155
rect -1196 124 -1164 125
rect -1196 75 -1164 76
rect -1196 45 -1195 75
rect -1195 45 -1165 75
rect -1165 45 -1164 75
rect -1196 44 -1164 45
rect -1196 -5 -1164 -4
rect -1196 -35 -1195 -5
rect -1195 -35 -1165 -5
rect -1165 -35 -1164 -5
rect -1196 -36 -1164 -35
rect -1196 -85 -1164 -84
rect -1196 -115 -1195 -85
rect -1195 -115 -1165 -85
rect -1165 -115 -1164 -85
rect -1196 -116 -1164 -115
rect -1036 5595 -1004 5596
rect -1036 5565 -1035 5595
rect -1035 5565 -1005 5595
rect -1005 5565 -1004 5595
rect -1036 5564 -1004 5565
rect -1036 5515 -1004 5516
rect -1036 5485 -1035 5515
rect -1035 5485 -1005 5515
rect -1005 5485 -1004 5515
rect -1036 5484 -1004 5485
rect -1036 5435 -1004 5436
rect -1036 5405 -1035 5435
rect -1035 5405 -1005 5435
rect -1005 5405 -1004 5435
rect -1036 5404 -1004 5405
rect -1036 5355 -1004 5356
rect -1036 5325 -1035 5355
rect -1035 5325 -1005 5355
rect -1005 5325 -1004 5355
rect -1036 5324 -1004 5325
rect -1036 5275 -1004 5276
rect -1036 5245 -1035 5275
rect -1035 5245 -1005 5275
rect -1005 5245 -1004 5275
rect -1036 5244 -1004 5245
rect -1036 5195 -1004 5196
rect -1036 5165 -1035 5195
rect -1035 5165 -1005 5195
rect -1005 5165 -1004 5195
rect -1036 5164 -1004 5165
rect -1036 5115 -1004 5116
rect -1036 5085 -1035 5115
rect -1035 5085 -1005 5115
rect -1005 5085 -1004 5115
rect -1036 5084 -1004 5085
rect -1036 5035 -1004 5036
rect -1036 5005 -1035 5035
rect -1035 5005 -1005 5035
rect -1005 5005 -1004 5035
rect -1036 5004 -1004 5005
rect -1036 4924 -1004 4956
rect -1036 4875 -1004 4876
rect -1036 4845 -1035 4875
rect -1035 4845 -1005 4875
rect -1005 4845 -1004 4875
rect -1036 4844 -1004 4845
rect -1036 4764 -1004 4796
rect -1036 4715 -1004 4716
rect -1036 4685 -1035 4715
rect -1035 4685 -1005 4715
rect -1005 4685 -1004 4715
rect -1036 4684 -1004 4685
rect -1036 4635 -1004 4636
rect -1036 4605 -1035 4635
rect -1035 4605 -1005 4635
rect -1005 4605 -1004 4635
rect -1036 4604 -1004 4605
rect -1036 4555 -1004 4556
rect -1036 4525 -1035 4555
rect -1035 4525 -1005 4555
rect -1005 4525 -1004 4555
rect -1036 4524 -1004 4525
rect -1036 4475 -1004 4476
rect -1036 4445 -1035 4475
rect -1035 4445 -1005 4475
rect -1005 4445 -1004 4475
rect -1036 4444 -1004 4445
rect -1036 4395 -1004 4396
rect -1036 4365 -1035 4395
rect -1035 4365 -1005 4395
rect -1005 4365 -1004 4395
rect -1036 4364 -1004 4365
rect -1036 4315 -1004 4316
rect -1036 4285 -1035 4315
rect -1035 4285 -1005 4315
rect -1005 4285 -1004 4315
rect -1036 4284 -1004 4285
rect -1036 4235 -1004 4236
rect -1036 4205 -1035 4235
rect -1035 4205 -1005 4235
rect -1005 4205 -1004 4235
rect -1036 4204 -1004 4205
rect -1036 4155 -1004 4156
rect -1036 4125 -1035 4155
rect -1035 4125 -1005 4155
rect -1005 4125 -1004 4155
rect -1036 4124 -1004 4125
rect -1036 4075 -1004 4076
rect -1036 4045 -1035 4075
rect -1035 4045 -1005 4075
rect -1005 4045 -1004 4075
rect -1036 4044 -1004 4045
rect -1036 3995 -1004 3996
rect -1036 3965 -1035 3995
rect -1035 3965 -1005 3995
rect -1005 3965 -1004 3995
rect -1036 3964 -1004 3965
rect -1036 3915 -1004 3916
rect -1036 3885 -1035 3915
rect -1035 3885 -1005 3915
rect -1005 3885 -1004 3915
rect -1036 3884 -1004 3885
rect -1036 3835 -1004 3836
rect -1036 3805 -1035 3835
rect -1035 3805 -1005 3835
rect -1005 3805 -1004 3835
rect -1036 3804 -1004 3805
rect -1036 3755 -1004 3756
rect -1036 3725 -1035 3755
rect -1035 3725 -1005 3755
rect -1005 3725 -1004 3755
rect -1036 3724 -1004 3725
rect -1036 3675 -1004 3676
rect -1036 3645 -1035 3675
rect -1035 3645 -1005 3675
rect -1005 3645 -1004 3675
rect -1036 3644 -1004 3645
rect -1036 3595 -1004 3596
rect -1036 3565 -1035 3595
rect -1035 3565 -1005 3595
rect -1005 3565 -1004 3595
rect -1036 3564 -1004 3565
rect -1036 3515 -1004 3516
rect -1036 3485 -1035 3515
rect -1035 3485 -1005 3515
rect -1005 3485 -1004 3515
rect -1036 3484 -1004 3485
rect -1036 3404 -1004 3436
rect -1036 3355 -1004 3356
rect -1036 3325 -1035 3355
rect -1035 3325 -1005 3355
rect -1005 3325 -1004 3355
rect -1036 3324 -1004 3325
rect -1036 3275 -1004 3276
rect -1036 3245 -1035 3275
rect -1035 3245 -1005 3275
rect -1005 3245 -1004 3275
rect -1036 3244 -1004 3245
rect -1036 3195 -1004 3196
rect -1036 3165 -1035 3195
rect -1035 3165 -1005 3195
rect -1005 3165 -1004 3195
rect -1036 3164 -1004 3165
rect -1036 3115 -1004 3116
rect -1036 3085 -1035 3115
rect -1035 3085 -1005 3115
rect -1005 3085 -1004 3115
rect -1036 3084 -1004 3085
rect -1036 3004 -1004 3036
rect -1036 2955 -1004 2956
rect -1036 2925 -1035 2955
rect -1035 2925 -1005 2955
rect -1005 2925 -1004 2955
rect -1036 2924 -1004 2925
rect -1036 2875 -1004 2876
rect -1036 2845 -1035 2875
rect -1035 2845 -1005 2875
rect -1005 2845 -1004 2875
rect -1036 2844 -1004 2845
rect -1036 2795 -1004 2796
rect -1036 2765 -1035 2795
rect -1035 2765 -1005 2795
rect -1005 2765 -1004 2795
rect -1036 2764 -1004 2765
rect -1036 2715 -1004 2716
rect -1036 2685 -1035 2715
rect -1035 2685 -1005 2715
rect -1005 2685 -1004 2715
rect -1036 2684 -1004 2685
rect -1036 2604 -1004 2636
rect -1036 2555 -1004 2556
rect -1036 2525 -1035 2555
rect -1035 2525 -1005 2555
rect -1005 2525 -1004 2555
rect -1036 2524 -1004 2525
rect -1036 2475 -1004 2476
rect -1036 2445 -1035 2475
rect -1035 2445 -1005 2475
rect -1005 2445 -1004 2475
rect -1036 2444 -1004 2445
rect -1036 2395 -1004 2396
rect -1036 2365 -1035 2395
rect -1035 2365 -1005 2395
rect -1005 2365 -1004 2395
rect -1036 2364 -1004 2365
rect -1036 2315 -1004 2316
rect -1036 2285 -1035 2315
rect -1035 2285 -1005 2315
rect -1005 2285 -1004 2315
rect -1036 2284 -1004 2285
rect -1036 2235 -1004 2236
rect -1036 2205 -1035 2235
rect -1035 2205 -1005 2235
rect -1005 2205 -1004 2235
rect -1036 2204 -1004 2205
rect -1036 2155 -1004 2156
rect -1036 2125 -1035 2155
rect -1035 2125 -1005 2155
rect -1005 2125 -1004 2155
rect -1036 2124 -1004 2125
rect -1036 2075 -1004 2076
rect -1036 2045 -1035 2075
rect -1035 2045 -1005 2075
rect -1005 2045 -1004 2075
rect -1036 2044 -1004 2045
rect -1036 1995 -1004 1996
rect -1036 1965 -1035 1995
rect -1035 1965 -1005 1995
rect -1005 1965 -1004 1995
rect -1036 1964 -1004 1965
rect -1036 1915 -1004 1916
rect -1036 1885 -1035 1915
rect -1035 1885 -1005 1915
rect -1005 1885 -1004 1915
rect -1036 1884 -1004 1885
rect -1036 1835 -1004 1836
rect -1036 1805 -1035 1835
rect -1035 1805 -1005 1835
rect -1005 1805 -1004 1835
rect -1036 1804 -1004 1805
rect -1036 1755 -1004 1756
rect -1036 1725 -1035 1755
rect -1035 1725 -1005 1755
rect -1005 1725 -1004 1755
rect -1036 1724 -1004 1725
rect -1036 1675 -1004 1676
rect -1036 1645 -1035 1675
rect -1035 1645 -1005 1675
rect -1005 1645 -1004 1675
rect -1036 1644 -1004 1645
rect -1036 1595 -1004 1596
rect -1036 1565 -1035 1595
rect -1035 1565 -1005 1595
rect -1005 1565 -1004 1595
rect -1036 1564 -1004 1565
rect -1036 1515 -1004 1516
rect -1036 1485 -1035 1515
rect -1035 1485 -1005 1515
rect -1005 1485 -1004 1515
rect -1036 1484 -1004 1485
rect -1036 1435 -1004 1436
rect -1036 1405 -1035 1435
rect -1035 1405 -1005 1435
rect -1005 1405 -1004 1435
rect -1036 1404 -1004 1405
rect -1036 1355 -1004 1356
rect -1036 1325 -1035 1355
rect -1035 1325 -1005 1355
rect -1005 1325 -1004 1355
rect -1036 1324 -1004 1325
rect -1036 1275 -1004 1276
rect -1036 1245 -1035 1275
rect -1035 1245 -1005 1275
rect -1005 1245 -1004 1275
rect -1036 1244 -1004 1245
rect -1036 1195 -1004 1196
rect -1036 1165 -1035 1195
rect -1035 1165 -1005 1195
rect -1005 1165 -1004 1195
rect -1036 1164 -1004 1165
rect -1036 1084 -1004 1116
rect -1036 1035 -1004 1036
rect -1036 1005 -1035 1035
rect -1035 1005 -1005 1035
rect -1005 1005 -1004 1035
rect -1036 1004 -1004 1005
rect -1036 955 -1004 956
rect -1036 925 -1035 955
rect -1035 925 -1005 955
rect -1005 925 -1004 955
rect -1036 924 -1004 925
rect -1036 875 -1004 876
rect -1036 845 -1035 875
rect -1035 845 -1005 875
rect -1005 845 -1004 875
rect -1036 844 -1004 845
rect -1036 795 -1004 796
rect -1036 765 -1035 795
rect -1035 765 -1005 795
rect -1005 765 -1004 795
rect -1036 764 -1004 765
rect -1036 715 -1004 716
rect -1036 685 -1035 715
rect -1035 685 -1005 715
rect -1005 685 -1004 715
rect -1036 684 -1004 685
rect -1036 635 -1004 636
rect -1036 605 -1035 635
rect -1035 605 -1005 635
rect -1005 605 -1004 635
rect -1036 604 -1004 605
rect -1036 555 -1004 556
rect -1036 525 -1035 555
rect -1035 525 -1005 555
rect -1005 525 -1004 555
rect -1036 524 -1004 525
rect -1036 475 -1004 476
rect -1036 445 -1035 475
rect -1035 445 -1005 475
rect -1005 445 -1004 475
rect -1036 444 -1004 445
rect -1036 395 -1004 396
rect -1036 365 -1035 395
rect -1035 365 -1005 395
rect -1005 365 -1004 395
rect -1036 364 -1004 365
rect -1036 315 -1004 316
rect -1036 285 -1035 315
rect -1035 285 -1005 315
rect -1005 285 -1004 315
rect -1036 284 -1004 285
rect -1036 235 -1004 236
rect -1036 205 -1035 235
rect -1035 205 -1005 235
rect -1005 205 -1004 235
rect -1036 204 -1004 205
rect -1036 155 -1004 156
rect -1036 125 -1035 155
rect -1035 125 -1005 155
rect -1005 125 -1004 155
rect -1036 124 -1004 125
rect -1036 75 -1004 76
rect -1036 45 -1035 75
rect -1035 45 -1005 75
rect -1005 45 -1004 75
rect -1036 44 -1004 45
rect -1036 -5 -1004 -4
rect -1036 -35 -1035 -5
rect -1035 -35 -1005 -5
rect -1005 -35 -1004 -5
rect -1036 -36 -1004 -35
rect -1036 -85 -1004 -84
rect -1036 -115 -1035 -85
rect -1035 -115 -1005 -85
rect -1005 -115 -1004 -85
rect -1036 -116 -1004 -115
rect -876 5595 -844 5596
rect -876 5565 -875 5595
rect -875 5565 -845 5595
rect -845 5565 -844 5595
rect -876 5564 -844 5565
rect 4884 5595 4916 5596
rect 4884 5565 4885 5595
rect 4885 5565 4915 5595
rect 4915 5565 4916 5595
rect 4884 5564 4916 5565
rect -876 5515 -844 5516
rect -876 5485 -875 5515
rect -875 5485 -845 5515
rect -845 5485 -844 5515
rect -876 5484 -844 5485
rect -876 5435 -844 5436
rect -876 5405 -875 5435
rect -875 5405 -845 5435
rect -845 5405 -844 5435
rect -876 5404 -844 5405
rect -876 5324 -844 5356
rect -876 5275 -844 5276
rect -876 5245 -875 5275
rect -875 5245 -845 5275
rect -845 5245 -844 5275
rect -876 5244 -844 5245
rect -876 5195 -844 5196
rect -876 5165 -875 5195
rect -875 5165 -845 5195
rect -845 5165 -844 5195
rect -876 5164 -844 5165
rect -876 5115 -844 5116
rect -876 5085 -875 5115
rect -875 5085 -845 5115
rect -845 5085 -844 5115
rect -876 5084 -844 5085
rect -876 5035 -844 5036
rect -876 5005 -875 5035
rect -875 5005 -845 5035
rect -845 5005 -844 5035
rect -876 5004 -844 5005
rect -876 4924 -844 4956
rect -876 4875 -844 4876
rect -876 4845 -875 4875
rect -875 4845 -845 4875
rect -845 4845 -844 4875
rect -876 4844 -844 4845
rect -876 4764 -844 4796
rect -876 4715 -844 4716
rect -876 4685 -875 4715
rect -875 4685 -845 4715
rect -845 4685 -844 4715
rect -876 4684 -844 4685
rect -876 4635 -844 4636
rect -876 4605 -875 4635
rect -875 4605 -845 4635
rect -845 4605 -844 4635
rect -876 4604 -844 4605
rect -876 4524 -844 4556
rect -876 4475 -844 4476
rect -876 4445 -875 4475
rect -875 4445 -845 4475
rect -845 4445 -844 4475
rect -876 4444 -844 4445
rect -796 5515 -764 5516
rect -796 5485 -795 5515
rect -795 5485 -765 5515
rect -765 5485 -764 5515
rect -796 5484 -764 5485
rect -796 5435 -764 5436
rect -796 5405 -795 5435
rect -795 5405 -765 5435
rect -765 5405 -764 5435
rect -796 5404 -764 5405
rect -796 5324 -764 5356
rect -796 5275 -764 5276
rect -796 5245 -795 5275
rect -795 5245 -765 5275
rect -765 5245 -764 5275
rect -796 5244 -764 5245
rect -796 5195 -764 5196
rect -796 5165 -795 5195
rect -795 5165 -765 5195
rect -765 5165 -764 5195
rect -796 5164 -764 5165
rect -796 5115 -764 5116
rect -796 5085 -795 5115
rect -795 5085 -765 5115
rect -765 5085 -764 5115
rect -796 5084 -764 5085
rect -796 5035 -764 5036
rect -796 5005 -795 5035
rect -795 5005 -765 5035
rect -765 5005 -764 5035
rect -796 5004 -764 5005
rect -796 4924 -764 4956
rect -796 4875 -764 4876
rect -796 4845 -795 4875
rect -795 4845 -765 4875
rect -765 4845 -764 4875
rect -796 4844 -764 4845
rect -796 4764 -764 4796
rect -796 4715 -764 4716
rect -796 4685 -795 4715
rect -795 4685 -765 4715
rect -765 4685 -764 4715
rect -796 4684 -764 4685
rect -796 4635 -764 4636
rect -796 4605 -795 4635
rect -795 4605 -765 4635
rect -765 4605 -764 4635
rect -796 4604 -764 4605
rect -796 4524 -764 4556
rect -796 4475 -764 4476
rect -796 4445 -795 4475
rect -795 4445 -765 4475
rect -765 4445 -764 4475
rect -796 4444 -764 4445
rect -716 5515 -684 5516
rect -716 5485 -715 5515
rect -715 5485 -685 5515
rect -685 5485 -684 5515
rect -716 5484 -684 5485
rect -716 5435 -684 5436
rect -716 5405 -715 5435
rect -715 5405 -685 5435
rect -685 5405 -684 5435
rect -716 5404 -684 5405
rect -716 5324 -684 5356
rect -716 5275 -684 5276
rect -716 5245 -715 5275
rect -715 5245 -685 5275
rect -685 5245 -684 5275
rect -716 5244 -684 5245
rect -716 5195 -684 5196
rect -716 5165 -715 5195
rect -715 5165 -685 5195
rect -685 5165 -684 5195
rect -716 5164 -684 5165
rect -716 5115 -684 5116
rect -716 5085 -715 5115
rect -715 5085 -685 5115
rect -685 5085 -684 5115
rect -716 5084 -684 5085
rect -716 5035 -684 5036
rect -716 5005 -715 5035
rect -715 5005 -685 5035
rect -685 5005 -684 5035
rect -716 5004 -684 5005
rect -716 4924 -684 4956
rect -716 4875 -684 4876
rect -716 4845 -715 4875
rect -715 4845 -685 4875
rect -685 4845 -684 4875
rect -716 4844 -684 4845
rect -716 4764 -684 4796
rect -716 4715 -684 4716
rect -716 4685 -715 4715
rect -715 4685 -685 4715
rect -685 4685 -684 4715
rect -716 4684 -684 4685
rect -716 4635 -684 4636
rect -716 4605 -715 4635
rect -715 4605 -685 4635
rect -685 4605 -684 4635
rect -716 4604 -684 4605
rect -716 4524 -684 4556
rect -716 4475 -684 4476
rect -716 4445 -715 4475
rect -715 4445 -685 4475
rect -685 4445 -684 4475
rect -716 4444 -684 4445
rect -636 5515 -604 5516
rect -636 5485 -635 5515
rect -635 5485 -605 5515
rect -605 5485 -604 5515
rect -636 5484 -604 5485
rect -636 5435 -604 5436
rect -636 5405 -635 5435
rect -635 5405 -605 5435
rect -605 5405 -604 5435
rect -636 5404 -604 5405
rect -636 5324 -604 5356
rect -636 5275 -604 5276
rect -636 5245 -635 5275
rect -635 5245 -605 5275
rect -605 5245 -604 5275
rect -636 5244 -604 5245
rect -636 5195 -604 5196
rect -636 5165 -635 5195
rect -635 5165 -605 5195
rect -605 5165 -604 5195
rect -636 5164 -604 5165
rect -636 5115 -604 5116
rect -636 5085 -635 5115
rect -635 5085 -605 5115
rect -605 5085 -604 5115
rect -636 5084 -604 5085
rect -636 5035 -604 5036
rect -636 5005 -635 5035
rect -635 5005 -605 5035
rect -605 5005 -604 5035
rect -636 5004 -604 5005
rect -636 4924 -604 4956
rect -636 4875 -604 4876
rect -636 4845 -635 4875
rect -635 4845 -605 4875
rect -605 4845 -604 4875
rect -636 4844 -604 4845
rect -636 4764 -604 4796
rect -636 4715 -604 4716
rect -636 4685 -635 4715
rect -635 4685 -605 4715
rect -605 4685 -604 4715
rect -636 4684 -604 4685
rect -636 4635 -604 4636
rect -636 4605 -635 4635
rect -635 4605 -605 4635
rect -605 4605 -604 4635
rect -636 4604 -604 4605
rect -636 4524 -604 4556
rect -636 4475 -604 4476
rect -636 4445 -635 4475
rect -635 4445 -605 4475
rect -605 4445 -604 4475
rect -636 4444 -604 4445
rect -556 5515 -524 5516
rect -556 5485 -555 5515
rect -555 5485 -525 5515
rect -525 5485 -524 5515
rect -556 5484 -524 5485
rect -556 5435 -524 5436
rect -556 5405 -555 5435
rect -555 5405 -525 5435
rect -525 5405 -524 5435
rect -556 5404 -524 5405
rect -556 5324 -524 5356
rect -556 5275 -524 5276
rect -556 5245 -555 5275
rect -555 5245 -525 5275
rect -525 5245 -524 5275
rect -556 5244 -524 5245
rect -556 5195 -524 5196
rect -556 5165 -555 5195
rect -555 5165 -525 5195
rect -525 5165 -524 5195
rect -556 5164 -524 5165
rect -556 5115 -524 5116
rect -556 5085 -555 5115
rect -555 5085 -525 5115
rect -525 5085 -524 5115
rect -556 5084 -524 5085
rect -556 5035 -524 5036
rect -556 5005 -555 5035
rect -555 5005 -525 5035
rect -525 5005 -524 5035
rect -556 5004 -524 5005
rect -556 4924 -524 4956
rect -556 4875 -524 4876
rect -556 4845 -555 4875
rect -555 4845 -525 4875
rect -525 4845 -524 4875
rect -556 4844 -524 4845
rect -556 4764 -524 4796
rect -556 4715 -524 4716
rect -556 4685 -555 4715
rect -555 4685 -525 4715
rect -525 4685 -524 4715
rect -556 4684 -524 4685
rect -556 4635 -524 4636
rect -556 4605 -555 4635
rect -555 4605 -525 4635
rect -525 4605 -524 4635
rect -556 4604 -524 4605
rect -556 4524 -524 4556
rect -556 4475 -524 4476
rect -556 4445 -555 4475
rect -555 4445 -525 4475
rect -525 4445 -524 4475
rect -556 4444 -524 4445
rect -476 5515 -444 5516
rect -476 5485 -475 5515
rect -475 5485 -445 5515
rect -445 5485 -444 5515
rect -476 5484 -444 5485
rect -476 5435 -444 5436
rect -476 5405 -475 5435
rect -475 5405 -445 5435
rect -445 5405 -444 5435
rect -476 5404 -444 5405
rect -476 5324 -444 5356
rect -476 5275 -444 5276
rect -476 5245 -475 5275
rect -475 5245 -445 5275
rect -445 5245 -444 5275
rect -476 5244 -444 5245
rect -476 5195 -444 5196
rect -476 5165 -475 5195
rect -475 5165 -445 5195
rect -445 5165 -444 5195
rect -476 5164 -444 5165
rect -476 5115 -444 5116
rect -476 5085 -475 5115
rect -475 5085 -445 5115
rect -445 5085 -444 5115
rect -476 5084 -444 5085
rect -476 5035 -444 5036
rect -476 5005 -475 5035
rect -475 5005 -445 5035
rect -445 5005 -444 5035
rect -476 5004 -444 5005
rect -476 4924 -444 4956
rect -476 4875 -444 4876
rect -476 4845 -475 4875
rect -475 4845 -445 4875
rect -445 4845 -444 4875
rect -476 4844 -444 4845
rect -476 4764 -444 4796
rect -476 4715 -444 4716
rect -476 4685 -475 4715
rect -475 4685 -445 4715
rect -445 4685 -444 4715
rect -476 4684 -444 4685
rect -476 4635 -444 4636
rect -476 4605 -475 4635
rect -475 4605 -445 4635
rect -445 4605 -444 4635
rect -476 4604 -444 4605
rect -476 4524 -444 4556
rect -476 4475 -444 4476
rect -476 4445 -475 4475
rect -475 4445 -445 4475
rect -445 4445 -444 4475
rect -476 4444 -444 4445
rect -396 5515 -364 5516
rect -396 5485 -395 5515
rect -395 5485 -365 5515
rect -365 5485 -364 5515
rect -396 5484 -364 5485
rect -396 5435 -364 5436
rect -396 5405 -395 5435
rect -395 5405 -365 5435
rect -365 5405 -364 5435
rect -396 5404 -364 5405
rect -396 5324 -364 5356
rect -396 5275 -364 5276
rect -396 5245 -395 5275
rect -395 5245 -365 5275
rect -365 5245 -364 5275
rect -396 5244 -364 5245
rect -396 5195 -364 5196
rect -396 5165 -395 5195
rect -395 5165 -365 5195
rect -365 5165 -364 5195
rect -396 5164 -364 5165
rect -396 5115 -364 5116
rect -396 5085 -395 5115
rect -395 5085 -365 5115
rect -365 5085 -364 5115
rect -396 5084 -364 5085
rect -396 5035 -364 5036
rect -396 5005 -395 5035
rect -395 5005 -365 5035
rect -365 5005 -364 5035
rect -396 5004 -364 5005
rect -396 4924 -364 4956
rect -396 4875 -364 4876
rect -396 4845 -395 4875
rect -395 4845 -365 4875
rect -365 4845 -364 4875
rect -396 4844 -364 4845
rect -396 4764 -364 4796
rect -396 4715 -364 4716
rect -396 4685 -395 4715
rect -395 4685 -365 4715
rect -365 4685 -364 4715
rect -396 4684 -364 4685
rect -396 4635 -364 4636
rect -396 4605 -395 4635
rect -395 4605 -365 4635
rect -365 4605 -364 4635
rect -396 4604 -364 4605
rect -396 4524 -364 4556
rect -396 4475 -364 4476
rect -396 4445 -395 4475
rect -395 4445 -365 4475
rect -365 4445 -364 4475
rect -396 4444 -364 4445
rect -316 5515 -284 5516
rect -316 5485 -315 5515
rect -315 5485 -285 5515
rect -285 5485 -284 5515
rect -316 5484 -284 5485
rect -316 5435 -284 5436
rect -316 5405 -315 5435
rect -315 5405 -285 5435
rect -285 5405 -284 5435
rect -316 5404 -284 5405
rect -316 5324 -284 5356
rect -316 5275 -284 5276
rect -316 5245 -315 5275
rect -315 5245 -285 5275
rect -285 5245 -284 5275
rect -316 5244 -284 5245
rect -316 5195 -284 5196
rect -316 5165 -315 5195
rect -315 5165 -285 5195
rect -285 5165 -284 5195
rect -316 5164 -284 5165
rect -316 5115 -284 5116
rect -316 5085 -315 5115
rect -315 5085 -285 5115
rect -285 5085 -284 5115
rect -316 5084 -284 5085
rect -316 5035 -284 5036
rect -316 5005 -315 5035
rect -315 5005 -285 5035
rect -285 5005 -284 5035
rect -316 5004 -284 5005
rect -316 4924 -284 4956
rect -316 4875 -284 4876
rect -316 4845 -315 4875
rect -315 4845 -285 4875
rect -285 4845 -284 4875
rect -316 4844 -284 4845
rect -316 4764 -284 4796
rect -316 4715 -284 4716
rect -316 4685 -315 4715
rect -315 4685 -285 4715
rect -285 4685 -284 4715
rect -316 4684 -284 4685
rect -316 4635 -284 4636
rect -316 4605 -315 4635
rect -315 4605 -285 4635
rect -285 4605 -284 4635
rect -316 4604 -284 4605
rect -316 4524 -284 4556
rect -316 4475 -284 4476
rect -316 4445 -315 4475
rect -315 4445 -285 4475
rect -285 4445 -284 4475
rect -316 4444 -284 4445
rect -236 5515 -204 5516
rect -236 5485 -235 5515
rect -235 5485 -205 5515
rect -205 5485 -204 5515
rect -236 5484 -204 5485
rect -236 5435 -204 5436
rect -236 5405 -235 5435
rect -235 5405 -205 5435
rect -205 5405 -204 5435
rect -236 5404 -204 5405
rect -236 5324 -204 5356
rect -236 5275 -204 5276
rect -236 5245 -235 5275
rect -235 5245 -205 5275
rect -205 5245 -204 5275
rect -236 5244 -204 5245
rect -236 5195 -204 5196
rect -236 5165 -235 5195
rect -235 5165 -205 5195
rect -205 5165 -204 5195
rect -236 5164 -204 5165
rect -236 5115 -204 5116
rect -236 5085 -235 5115
rect -235 5085 -205 5115
rect -205 5085 -204 5115
rect -236 5084 -204 5085
rect -236 5035 -204 5036
rect -236 5005 -235 5035
rect -235 5005 -205 5035
rect -205 5005 -204 5035
rect -236 5004 -204 5005
rect -236 4924 -204 4956
rect -236 4875 -204 4876
rect -236 4845 -235 4875
rect -235 4845 -205 4875
rect -205 4845 -204 4875
rect -236 4844 -204 4845
rect -236 4764 -204 4796
rect -236 4715 -204 4716
rect -236 4685 -235 4715
rect -235 4685 -205 4715
rect -205 4685 -204 4715
rect -236 4684 -204 4685
rect -236 4635 -204 4636
rect -236 4605 -235 4635
rect -235 4605 -205 4635
rect -205 4605 -204 4635
rect -236 4604 -204 4605
rect -236 4524 -204 4556
rect -236 4475 -204 4476
rect -236 4445 -235 4475
rect -235 4445 -205 4475
rect -205 4445 -204 4475
rect -236 4444 -204 4445
rect -156 5515 -124 5516
rect -156 5485 -155 5515
rect -155 5485 -125 5515
rect -125 5485 -124 5515
rect -156 5484 -124 5485
rect -156 5435 -124 5436
rect -156 5405 -155 5435
rect -155 5405 -125 5435
rect -125 5405 -124 5435
rect -156 5404 -124 5405
rect -156 5324 -124 5356
rect -156 5275 -124 5276
rect -156 5245 -155 5275
rect -155 5245 -125 5275
rect -125 5245 -124 5275
rect -156 5244 -124 5245
rect -156 5195 -124 5196
rect -156 5165 -155 5195
rect -155 5165 -125 5195
rect -125 5165 -124 5195
rect -156 5164 -124 5165
rect -156 5115 -124 5116
rect -156 5085 -155 5115
rect -155 5085 -125 5115
rect -125 5085 -124 5115
rect -156 5084 -124 5085
rect -156 5035 -124 5036
rect -156 5005 -155 5035
rect -155 5005 -125 5035
rect -125 5005 -124 5035
rect -156 5004 -124 5005
rect -156 4924 -124 4956
rect -156 4875 -124 4876
rect -156 4845 -155 4875
rect -155 4845 -125 4875
rect -125 4845 -124 4875
rect -156 4844 -124 4845
rect -156 4764 -124 4796
rect -156 4715 -124 4716
rect -156 4685 -155 4715
rect -155 4685 -125 4715
rect -125 4685 -124 4715
rect -156 4684 -124 4685
rect -156 4635 -124 4636
rect -156 4605 -155 4635
rect -155 4605 -125 4635
rect -125 4605 -124 4635
rect -156 4604 -124 4605
rect -156 4524 -124 4556
rect -156 4475 -124 4476
rect -156 4445 -155 4475
rect -155 4445 -125 4475
rect -125 4445 -124 4475
rect -156 4444 -124 4445
rect -76 5515 -44 5516
rect -76 5485 -75 5515
rect -75 5485 -45 5515
rect -45 5485 -44 5515
rect -76 5484 -44 5485
rect -76 5435 -44 5436
rect -76 5405 -75 5435
rect -75 5405 -45 5435
rect -45 5405 -44 5435
rect -76 5404 -44 5405
rect -76 5324 -44 5356
rect -76 5275 -44 5276
rect -76 5245 -75 5275
rect -75 5245 -45 5275
rect -45 5245 -44 5275
rect -76 5244 -44 5245
rect -76 5195 -44 5196
rect -76 5165 -75 5195
rect -75 5165 -45 5195
rect -45 5165 -44 5195
rect -76 5164 -44 5165
rect -76 5115 -44 5116
rect -76 5085 -75 5115
rect -75 5085 -45 5115
rect -45 5085 -44 5115
rect -76 5084 -44 5085
rect -76 5035 -44 5036
rect -76 5005 -75 5035
rect -75 5005 -45 5035
rect -45 5005 -44 5035
rect -76 5004 -44 5005
rect -76 4924 -44 4956
rect -76 4875 -44 4876
rect -76 4845 -75 4875
rect -75 4845 -45 4875
rect -45 4845 -44 4875
rect -76 4844 -44 4845
rect -76 4764 -44 4796
rect -76 4715 -44 4716
rect -76 4685 -75 4715
rect -75 4685 -45 4715
rect -45 4685 -44 4715
rect -76 4684 -44 4685
rect -76 4635 -44 4636
rect -76 4605 -75 4635
rect -75 4605 -45 4635
rect -45 4605 -44 4635
rect -76 4604 -44 4605
rect -76 4524 -44 4556
rect -76 4475 -44 4476
rect -76 4445 -75 4475
rect -75 4445 -45 4475
rect -45 4445 -44 4475
rect -76 4444 -44 4445
rect 4 5515 36 5516
rect 4 5485 5 5515
rect 5 5485 35 5515
rect 35 5485 36 5515
rect 4 5484 36 5485
rect 4 5435 36 5436
rect 4 5405 5 5435
rect 5 5405 35 5435
rect 35 5405 36 5435
rect 4 5404 36 5405
rect 4 5324 36 5356
rect 4 5275 36 5276
rect 4 5245 5 5275
rect 5 5245 35 5275
rect 35 5245 36 5275
rect 4 5244 36 5245
rect 4 5195 36 5196
rect 4 5165 5 5195
rect 5 5165 35 5195
rect 35 5165 36 5195
rect 4 5164 36 5165
rect 4 5115 36 5116
rect 4 5085 5 5115
rect 5 5085 35 5115
rect 35 5085 36 5115
rect 4 5084 36 5085
rect 4 5035 36 5036
rect 4 5005 5 5035
rect 5 5005 35 5035
rect 35 5005 36 5035
rect 4 5004 36 5005
rect 4 4924 36 4956
rect 4 4875 36 4876
rect 4 4845 5 4875
rect 5 4845 35 4875
rect 35 4845 36 4875
rect 4 4844 36 4845
rect 4 4764 36 4796
rect 4 4715 36 4716
rect 4 4685 5 4715
rect 5 4685 35 4715
rect 35 4685 36 4715
rect 4 4684 36 4685
rect 4 4635 36 4636
rect 4 4605 5 4635
rect 5 4605 35 4635
rect 35 4605 36 4635
rect 4 4604 36 4605
rect 4 4524 36 4556
rect 4 4475 36 4476
rect 4 4445 5 4475
rect 5 4445 35 4475
rect 35 4445 36 4475
rect 4 4444 36 4445
rect 84 5515 116 5516
rect 84 5485 85 5515
rect 85 5485 115 5515
rect 115 5485 116 5515
rect 84 5484 116 5485
rect 84 5435 116 5436
rect 84 5405 85 5435
rect 85 5405 115 5435
rect 115 5405 116 5435
rect 84 5404 116 5405
rect 84 5324 116 5356
rect 84 5275 116 5276
rect 84 5245 85 5275
rect 85 5245 115 5275
rect 115 5245 116 5275
rect 84 5244 116 5245
rect 84 5195 116 5196
rect 84 5165 85 5195
rect 85 5165 115 5195
rect 115 5165 116 5195
rect 84 5164 116 5165
rect 84 5115 116 5116
rect 84 5085 85 5115
rect 85 5085 115 5115
rect 115 5085 116 5115
rect 84 5084 116 5085
rect 84 5035 116 5036
rect 84 5005 85 5035
rect 85 5005 115 5035
rect 115 5005 116 5035
rect 84 5004 116 5005
rect 84 4924 116 4956
rect 84 4875 116 4876
rect 84 4845 85 4875
rect 85 4845 115 4875
rect 115 4845 116 4875
rect 84 4844 116 4845
rect 84 4764 116 4796
rect 84 4715 116 4716
rect 84 4685 85 4715
rect 85 4685 115 4715
rect 115 4685 116 4715
rect 84 4684 116 4685
rect 84 4635 116 4636
rect 84 4605 85 4635
rect 85 4605 115 4635
rect 115 4605 116 4635
rect 84 4604 116 4605
rect 84 4524 116 4556
rect 84 4475 116 4476
rect 84 4445 85 4475
rect 85 4445 115 4475
rect 115 4445 116 4475
rect 84 4444 116 4445
rect 164 5515 196 5516
rect 164 5485 165 5515
rect 165 5485 195 5515
rect 195 5485 196 5515
rect 164 5484 196 5485
rect 164 5435 196 5436
rect 164 5405 165 5435
rect 165 5405 195 5435
rect 195 5405 196 5435
rect 164 5404 196 5405
rect 164 5324 196 5356
rect 164 5275 196 5276
rect 164 5245 165 5275
rect 165 5245 195 5275
rect 195 5245 196 5275
rect 164 5244 196 5245
rect 164 5195 196 5196
rect 164 5165 165 5195
rect 165 5165 195 5195
rect 195 5165 196 5195
rect 164 5164 196 5165
rect 164 5115 196 5116
rect 164 5085 165 5115
rect 165 5085 195 5115
rect 195 5085 196 5115
rect 164 5084 196 5085
rect 164 5035 196 5036
rect 164 5005 165 5035
rect 165 5005 195 5035
rect 195 5005 196 5035
rect 164 5004 196 5005
rect 164 4924 196 4956
rect 164 4875 196 4876
rect 164 4845 165 4875
rect 165 4845 195 4875
rect 195 4845 196 4875
rect 164 4844 196 4845
rect 164 4764 196 4796
rect 164 4715 196 4716
rect 164 4685 165 4715
rect 165 4685 195 4715
rect 195 4685 196 4715
rect 164 4684 196 4685
rect 164 4635 196 4636
rect 164 4605 165 4635
rect 165 4605 195 4635
rect 195 4605 196 4635
rect 164 4604 196 4605
rect 164 4524 196 4556
rect 164 4475 196 4476
rect 164 4445 165 4475
rect 165 4445 195 4475
rect 195 4445 196 4475
rect 164 4444 196 4445
rect 244 5515 276 5516
rect 244 5485 245 5515
rect 245 5485 275 5515
rect 275 5485 276 5515
rect 244 5484 276 5485
rect 244 5435 276 5436
rect 244 5405 245 5435
rect 245 5405 275 5435
rect 275 5405 276 5435
rect 244 5404 276 5405
rect 244 5324 276 5356
rect 244 5275 276 5276
rect 244 5245 245 5275
rect 245 5245 275 5275
rect 275 5245 276 5275
rect 244 5244 276 5245
rect 244 5195 276 5196
rect 244 5165 245 5195
rect 245 5165 275 5195
rect 275 5165 276 5195
rect 244 5164 276 5165
rect 244 5115 276 5116
rect 244 5085 245 5115
rect 245 5085 275 5115
rect 275 5085 276 5115
rect 244 5084 276 5085
rect 244 5035 276 5036
rect 244 5005 245 5035
rect 245 5005 275 5035
rect 275 5005 276 5035
rect 244 5004 276 5005
rect 244 4924 276 4956
rect 244 4875 276 4876
rect 244 4845 245 4875
rect 245 4845 275 4875
rect 275 4845 276 4875
rect 244 4844 276 4845
rect 244 4764 276 4796
rect 244 4715 276 4716
rect 244 4685 245 4715
rect 245 4685 275 4715
rect 275 4685 276 4715
rect 244 4684 276 4685
rect 244 4635 276 4636
rect 244 4605 245 4635
rect 245 4605 275 4635
rect 275 4605 276 4635
rect 244 4604 276 4605
rect 244 4524 276 4556
rect 244 4475 276 4476
rect 244 4445 245 4475
rect 245 4445 275 4475
rect 275 4445 276 4475
rect 244 4444 276 4445
rect 324 5515 356 5516
rect 324 5485 325 5515
rect 325 5485 355 5515
rect 355 5485 356 5515
rect 324 5484 356 5485
rect 324 5435 356 5436
rect 324 5405 325 5435
rect 325 5405 355 5435
rect 355 5405 356 5435
rect 324 5404 356 5405
rect 324 5324 356 5356
rect 324 5275 356 5276
rect 324 5245 325 5275
rect 325 5245 355 5275
rect 355 5245 356 5275
rect 324 5244 356 5245
rect 324 5195 356 5196
rect 324 5165 325 5195
rect 325 5165 355 5195
rect 355 5165 356 5195
rect 324 5164 356 5165
rect 324 5115 356 5116
rect 324 5085 325 5115
rect 325 5085 355 5115
rect 355 5085 356 5115
rect 324 5084 356 5085
rect 324 5035 356 5036
rect 324 5005 325 5035
rect 325 5005 355 5035
rect 355 5005 356 5035
rect 324 5004 356 5005
rect 324 4924 356 4956
rect 324 4875 356 4876
rect 324 4845 325 4875
rect 325 4845 355 4875
rect 355 4845 356 4875
rect 324 4844 356 4845
rect 324 4764 356 4796
rect 324 4715 356 4716
rect 324 4685 325 4715
rect 325 4685 355 4715
rect 355 4685 356 4715
rect 324 4684 356 4685
rect 324 4635 356 4636
rect 324 4605 325 4635
rect 325 4605 355 4635
rect 355 4605 356 4635
rect 324 4604 356 4605
rect 324 4524 356 4556
rect 324 4475 356 4476
rect 324 4445 325 4475
rect 325 4445 355 4475
rect 355 4445 356 4475
rect 324 4444 356 4445
rect 404 5515 436 5516
rect 404 5485 405 5515
rect 405 5485 435 5515
rect 435 5485 436 5515
rect 404 5484 436 5485
rect 404 5435 436 5436
rect 404 5405 405 5435
rect 405 5405 435 5435
rect 435 5405 436 5435
rect 404 5404 436 5405
rect 404 5324 436 5356
rect 404 5275 436 5276
rect 404 5245 405 5275
rect 405 5245 435 5275
rect 435 5245 436 5275
rect 404 5244 436 5245
rect 404 5195 436 5196
rect 404 5165 405 5195
rect 405 5165 435 5195
rect 435 5165 436 5195
rect 404 5164 436 5165
rect 404 5115 436 5116
rect 404 5085 405 5115
rect 405 5085 435 5115
rect 435 5085 436 5115
rect 404 5084 436 5085
rect 404 5035 436 5036
rect 404 5005 405 5035
rect 405 5005 435 5035
rect 435 5005 436 5035
rect 404 5004 436 5005
rect 404 4924 436 4956
rect 404 4875 436 4876
rect 404 4845 405 4875
rect 405 4845 435 4875
rect 435 4845 436 4875
rect 404 4844 436 4845
rect 404 4764 436 4796
rect 404 4715 436 4716
rect 404 4685 405 4715
rect 405 4685 435 4715
rect 435 4685 436 4715
rect 404 4684 436 4685
rect 404 4635 436 4636
rect 404 4605 405 4635
rect 405 4605 435 4635
rect 435 4605 436 4635
rect 404 4604 436 4605
rect 404 4524 436 4556
rect 404 4475 436 4476
rect 404 4445 405 4475
rect 405 4445 435 4475
rect 435 4445 436 4475
rect 404 4444 436 4445
rect 484 5515 516 5516
rect 484 5485 485 5515
rect 485 5485 515 5515
rect 515 5485 516 5515
rect 484 5484 516 5485
rect 484 5435 516 5436
rect 484 5405 485 5435
rect 485 5405 515 5435
rect 515 5405 516 5435
rect 484 5404 516 5405
rect 484 5324 516 5356
rect 484 5275 516 5276
rect 484 5245 485 5275
rect 485 5245 515 5275
rect 515 5245 516 5275
rect 484 5244 516 5245
rect 484 5195 516 5196
rect 484 5165 485 5195
rect 485 5165 515 5195
rect 515 5165 516 5195
rect 484 5164 516 5165
rect 484 5115 516 5116
rect 484 5085 485 5115
rect 485 5085 515 5115
rect 515 5085 516 5115
rect 484 5084 516 5085
rect 484 5035 516 5036
rect 484 5005 485 5035
rect 485 5005 515 5035
rect 515 5005 516 5035
rect 484 5004 516 5005
rect 484 4924 516 4956
rect 484 4875 516 4876
rect 484 4845 485 4875
rect 485 4845 515 4875
rect 515 4845 516 4875
rect 484 4844 516 4845
rect 484 4764 516 4796
rect 484 4715 516 4716
rect 484 4685 485 4715
rect 485 4685 515 4715
rect 515 4685 516 4715
rect 484 4684 516 4685
rect 484 4635 516 4636
rect 484 4605 485 4635
rect 485 4605 515 4635
rect 515 4605 516 4635
rect 484 4604 516 4605
rect 484 4524 516 4556
rect 484 4475 516 4476
rect 484 4445 485 4475
rect 485 4445 515 4475
rect 515 4445 516 4475
rect 484 4444 516 4445
rect 564 5515 596 5516
rect 564 5485 565 5515
rect 565 5485 595 5515
rect 595 5485 596 5515
rect 564 5484 596 5485
rect 564 5435 596 5436
rect 564 5405 565 5435
rect 565 5405 595 5435
rect 595 5405 596 5435
rect 564 5404 596 5405
rect 564 5324 596 5356
rect 564 5275 596 5276
rect 564 5245 565 5275
rect 565 5245 595 5275
rect 595 5245 596 5275
rect 564 5244 596 5245
rect 564 5195 596 5196
rect 564 5165 565 5195
rect 565 5165 595 5195
rect 595 5165 596 5195
rect 564 5164 596 5165
rect 564 5115 596 5116
rect 564 5085 565 5115
rect 565 5085 595 5115
rect 595 5085 596 5115
rect 564 5084 596 5085
rect 564 5035 596 5036
rect 564 5005 565 5035
rect 565 5005 595 5035
rect 595 5005 596 5035
rect 564 5004 596 5005
rect 564 4924 596 4956
rect 564 4875 596 4876
rect 564 4845 565 4875
rect 565 4845 595 4875
rect 595 4845 596 4875
rect 564 4844 596 4845
rect 564 4764 596 4796
rect 564 4715 596 4716
rect 564 4685 565 4715
rect 565 4685 595 4715
rect 595 4685 596 4715
rect 564 4684 596 4685
rect 564 4635 596 4636
rect 564 4605 565 4635
rect 565 4605 595 4635
rect 595 4605 596 4635
rect 564 4604 596 4605
rect 564 4524 596 4556
rect 564 4475 596 4476
rect 564 4445 565 4475
rect 565 4445 595 4475
rect 595 4445 596 4475
rect 564 4444 596 4445
rect 644 5515 676 5516
rect 644 5485 645 5515
rect 645 5485 675 5515
rect 675 5485 676 5515
rect 644 5484 676 5485
rect 644 5435 676 5436
rect 644 5405 645 5435
rect 645 5405 675 5435
rect 675 5405 676 5435
rect 644 5404 676 5405
rect 644 5324 676 5356
rect 644 5275 676 5276
rect 644 5245 645 5275
rect 645 5245 675 5275
rect 675 5245 676 5275
rect 644 5244 676 5245
rect 644 5195 676 5196
rect 644 5165 645 5195
rect 645 5165 675 5195
rect 675 5165 676 5195
rect 644 5164 676 5165
rect 644 5115 676 5116
rect 644 5085 645 5115
rect 645 5085 675 5115
rect 675 5085 676 5115
rect 644 5084 676 5085
rect 644 5035 676 5036
rect 644 5005 645 5035
rect 645 5005 675 5035
rect 675 5005 676 5035
rect 644 5004 676 5005
rect 644 4924 676 4956
rect 644 4875 676 4876
rect 644 4845 645 4875
rect 645 4845 675 4875
rect 675 4845 676 4875
rect 644 4844 676 4845
rect 644 4764 676 4796
rect 644 4715 676 4716
rect 644 4685 645 4715
rect 645 4685 675 4715
rect 675 4685 676 4715
rect 644 4684 676 4685
rect 644 4635 676 4636
rect 644 4605 645 4635
rect 645 4605 675 4635
rect 675 4605 676 4635
rect 644 4604 676 4605
rect 644 4524 676 4556
rect 644 4475 676 4476
rect 644 4445 645 4475
rect 645 4445 675 4475
rect 675 4445 676 4475
rect 644 4444 676 4445
rect 724 5515 756 5516
rect 724 5485 725 5515
rect 725 5485 755 5515
rect 755 5485 756 5515
rect 724 5484 756 5485
rect 724 5435 756 5436
rect 724 5405 725 5435
rect 725 5405 755 5435
rect 755 5405 756 5435
rect 724 5404 756 5405
rect 724 5324 756 5356
rect 724 5275 756 5276
rect 724 5245 725 5275
rect 725 5245 755 5275
rect 755 5245 756 5275
rect 724 5244 756 5245
rect 724 5195 756 5196
rect 724 5165 725 5195
rect 725 5165 755 5195
rect 755 5165 756 5195
rect 724 5164 756 5165
rect 724 5115 756 5116
rect 724 5085 725 5115
rect 725 5085 755 5115
rect 755 5085 756 5115
rect 724 5084 756 5085
rect 724 5035 756 5036
rect 724 5005 725 5035
rect 725 5005 755 5035
rect 755 5005 756 5035
rect 724 5004 756 5005
rect 724 4924 756 4956
rect 724 4875 756 4876
rect 724 4845 725 4875
rect 725 4845 755 4875
rect 755 4845 756 4875
rect 724 4844 756 4845
rect 724 4764 756 4796
rect 724 4715 756 4716
rect 724 4685 725 4715
rect 725 4685 755 4715
rect 755 4685 756 4715
rect 724 4684 756 4685
rect 724 4635 756 4636
rect 724 4605 725 4635
rect 725 4605 755 4635
rect 755 4605 756 4635
rect 724 4604 756 4605
rect 724 4524 756 4556
rect 724 4475 756 4476
rect 724 4445 725 4475
rect 725 4445 755 4475
rect 755 4445 756 4475
rect 724 4444 756 4445
rect 804 5515 836 5516
rect 804 5485 805 5515
rect 805 5485 835 5515
rect 835 5485 836 5515
rect 804 5484 836 5485
rect 804 5435 836 5436
rect 804 5405 805 5435
rect 805 5405 835 5435
rect 835 5405 836 5435
rect 804 5404 836 5405
rect 804 5324 836 5356
rect 804 5275 836 5276
rect 804 5245 805 5275
rect 805 5245 835 5275
rect 835 5245 836 5275
rect 804 5244 836 5245
rect 804 5195 836 5196
rect 804 5165 805 5195
rect 805 5165 835 5195
rect 835 5165 836 5195
rect 804 5164 836 5165
rect 804 5115 836 5116
rect 804 5085 805 5115
rect 805 5085 835 5115
rect 835 5085 836 5115
rect 804 5084 836 5085
rect 804 5035 836 5036
rect 804 5005 805 5035
rect 805 5005 835 5035
rect 835 5005 836 5035
rect 804 5004 836 5005
rect 804 4924 836 4956
rect 804 4875 836 4876
rect 804 4845 805 4875
rect 805 4845 835 4875
rect 835 4845 836 4875
rect 804 4844 836 4845
rect 804 4764 836 4796
rect 804 4715 836 4716
rect 804 4685 805 4715
rect 805 4685 835 4715
rect 835 4685 836 4715
rect 804 4684 836 4685
rect 804 4635 836 4636
rect 804 4605 805 4635
rect 805 4605 835 4635
rect 835 4605 836 4635
rect 804 4604 836 4605
rect 804 4524 836 4556
rect 804 4475 836 4476
rect 804 4445 805 4475
rect 805 4445 835 4475
rect 835 4445 836 4475
rect 804 4444 836 4445
rect 884 5515 916 5516
rect 884 5485 885 5515
rect 885 5485 915 5515
rect 915 5485 916 5515
rect 884 5484 916 5485
rect 884 5435 916 5436
rect 884 5405 885 5435
rect 885 5405 915 5435
rect 915 5405 916 5435
rect 884 5404 916 5405
rect 884 5324 916 5356
rect 884 5275 916 5276
rect 884 5245 885 5275
rect 885 5245 915 5275
rect 915 5245 916 5275
rect 884 5244 916 5245
rect 884 5195 916 5196
rect 884 5165 885 5195
rect 885 5165 915 5195
rect 915 5165 916 5195
rect 884 5164 916 5165
rect 884 5115 916 5116
rect 884 5085 885 5115
rect 885 5085 915 5115
rect 915 5085 916 5115
rect 884 5084 916 5085
rect 884 5035 916 5036
rect 884 5005 885 5035
rect 885 5005 915 5035
rect 915 5005 916 5035
rect 884 5004 916 5005
rect 884 4924 916 4956
rect 884 4875 916 4876
rect 884 4845 885 4875
rect 885 4845 915 4875
rect 915 4845 916 4875
rect 884 4844 916 4845
rect 884 4764 916 4796
rect 884 4715 916 4716
rect 884 4685 885 4715
rect 885 4685 915 4715
rect 915 4685 916 4715
rect 884 4684 916 4685
rect 884 4635 916 4636
rect 884 4605 885 4635
rect 885 4605 915 4635
rect 915 4605 916 4635
rect 884 4604 916 4605
rect 884 4524 916 4556
rect 884 4475 916 4476
rect 884 4445 885 4475
rect 885 4445 915 4475
rect 915 4445 916 4475
rect 884 4444 916 4445
rect 964 5515 996 5516
rect 964 5485 965 5515
rect 965 5485 995 5515
rect 995 5485 996 5515
rect 964 5484 996 5485
rect 964 5435 996 5436
rect 964 5405 965 5435
rect 965 5405 995 5435
rect 995 5405 996 5435
rect 964 5404 996 5405
rect 964 5324 996 5356
rect 964 5275 996 5276
rect 964 5245 965 5275
rect 965 5245 995 5275
rect 995 5245 996 5275
rect 964 5244 996 5245
rect 964 5195 996 5196
rect 964 5165 965 5195
rect 965 5165 995 5195
rect 995 5165 996 5195
rect 964 5164 996 5165
rect 964 5115 996 5116
rect 964 5085 965 5115
rect 965 5085 995 5115
rect 995 5085 996 5115
rect 964 5084 996 5085
rect 964 5035 996 5036
rect 964 5005 965 5035
rect 965 5005 995 5035
rect 995 5005 996 5035
rect 964 5004 996 5005
rect 964 4924 996 4956
rect 964 4875 996 4876
rect 964 4845 965 4875
rect 965 4845 995 4875
rect 995 4845 996 4875
rect 964 4844 996 4845
rect 964 4764 996 4796
rect 964 4715 996 4716
rect 964 4685 965 4715
rect 965 4685 995 4715
rect 995 4685 996 4715
rect 964 4684 996 4685
rect 964 4635 996 4636
rect 964 4605 965 4635
rect 965 4605 995 4635
rect 995 4605 996 4635
rect 964 4604 996 4605
rect 964 4524 996 4556
rect 964 4475 996 4476
rect 964 4445 965 4475
rect 965 4445 995 4475
rect 995 4445 996 4475
rect 964 4444 996 4445
rect 1044 5515 1076 5516
rect 1044 5485 1045 5515
rect 1045 5485 1075 5515
rect 1075 5485 1076 5515
rect 1044 5484 1076 5485
rect 1044 5435 1076 5436
rect 1044 5405 1045 5435
rect 1045 5405 1075 5435
rect 1075 5405 1076 5435
rect 1044 5404 1076 5405
rect 1044 5324 1076 5356
rect 1044 5275 1076 5276
rect 1044 5245 1045 5275
rect 1045 5245 1075 5275
rect 1075 5245 1076 5275
rect 1044 5244 1076 5245
rect 1044 5195 1076 5196
rect 1044 5165 1045 5195
rect 1045 5165 1075 5195
rect 1075 5165 1076 5195
rect 1044 5164 1076 5165
rect 1044 5115 1076 5116
rect 1044 5085 1045 5115
rect 1045 5085 1075 5115
rect 1075 5085 1076 5115
rect 1044 5084 1076 5085
rect 1044 5035 1076 5036
rect 1044 5005 1045 5035
rect 1045 5005 1075 5035
rect 1075 5005 1076 5035
rect 1044 5004 1076 5005
rect 1044 4924 1076 4956
rect 1044 4875 1076 4876
rect 1044 4845 1045 4875
rect 1045 4845 1075 4875
rect 1075 4845 1076 4875
rect 1044 4844 1076 4845
rect 1044 4764 1076 4796
rect 1044 4715 1076 4716
rect 1044 4685 1045 4715
rect 1045 4685 1075 4715
rect 1075 4685 1076 4715
rect 1044 4684 1076 4685
rect 1044 4635 1076 4636
rect 1044 4605 1045 4635
rect 1045 4605 1075 4635
rect 1075 4605 1076 4635
rect 1044 4604 1076 4605
rect 1044 4524 1076 4556
rect 1044 4475 1076 4476
rect 1044 4445 1045 4475
rect 1045 4445 1075 4475
rect 1075 4445 1076 4475
rect 1044 4444 1076 4445
rect 1124 5515 1156 5516
rect 1124 5485 1125 5515
rect 1125 5485 1155 5515
rect 1155 5485 1156 5515
rect 1124 5484 1156 5485
rect 1124 5435 1156 5436
rect 1124 5405 1125 5435
rect 1125 5405 1155 5435
rect 1155 5405 1156 5435
rect 1124 5404 1156 5405
rect 1124 5324 1156 5356
rect 1124 5275 1156 5276
rect 1124 5245 1125 5275
rect 1125 5245 1155 5275
rect 1155 5245 1156 5275
rect 1124 5244 1156 5245
rect 1124 5195 1156 5196
rect 1124 5165 1125 5195
rect 1125 5165 1155 5195
rect 1155 5165 1156 5195
rect 1124 5164 1156 5165
rect 1124 5115 1156 5116
rect 1124 5085 1125 5115
rect 1125 5085 1155 5115
rect 1155 5085 1156 5115
rect 1124 5084 1156 5085
rect 1124 5035 1156 5036
rect 1124 5005 1125 5035
rect 1125 5005 1155 5035
rect 1155 5005 1156 5035
rect 1124 5004 1156 5005
rect 1124 4924 1156 4956
rect 1124 4875 1156 4876
rect 1124 4845 1125 4875
rect 1125 4845 1155 4875
rect 1155 4845 1156 4875
rect 1124 4844 1156 4845
rect 1124 4764 1156 4796
rect 1124 4715 1156 4716
rect 1124 4685 1125 4715
rect 1125 4685 1155 4715
rect 1155 4685 1156 4715
rect 1124 4684 1156 4685
rect 1124 4635 1156 4636
rect 1124 4605 1125 4635
rect 1125 4605 1155 4635
rect 1155 4605 1156 4635
rect 1124 4604 1156 4605
rect 1124 4524 1156 4556
rect 1124 4475 1156 4476
rect 1124 4445 1125 4475
rect 1125 4445 1155 4475
rect 1155 4445 1156 4475
rect 1124 4444 1156 4445
rect 1204 5515 1236 5516
rect 1204 5485 1205 5515
rect 1205 5485 1235 5515
rect 1235 5485 1236 5515
rect 1204 5484 1236 5485
rect 1204 5435 1236 5436
rect 1204 5405 1205 5435
rect 1205 5405 1235 5435
rect 1235 5405 1236 5435
rect 1204 5404 1236 5405
rect 1204 5324 1236 5356
rect 1204 5275 1236 5276
rect 1204 5245 1205 5275
rect 1205 5245 1235 5275
rect 1235 5245 1236 5275
rect 1204 5244 1236 5245
rect 1204 5195 1236 5196
rect 1204 5165 1205 5195
rect 1205 5165 1235 5195
rect 1235 5165 1236 5195
rect 1204 5164 1236 5165
rect 1204 5115 1236 5116
rect 1204 5085 1205 5115
rect 1205 5085 1235 5115
rect 1235 5085 1236 5115
rect 1204 5084 1236 5085
rect 1204 5035 1236 5036
rect 1204 5005 1205 5035
rect 1205 5005 1235 5035
rect 1235 5005 1236 5035
rect 1204 5004 1236 5005
rect 1204 4924 1236 4956
rect 1204 4875 1236 4876
rect 1204 4845 1205 4875
rect 1205 4845 1235 4875
rect 1235 4845 1236 4875
rect 1204 4844 1236 4845
rect 1204 4764 1236 4796
rect 1204 4715 1236 4716
rect 1204 4685 1205 4715
rect 1205 4685 1235 4715
rect 1235 4685 1236 4715
rect 1204 4684 1236 4685
rect 1204 4635 1236 4636
rect 1204 4605 1205 4635
rect 1205 4605 1235 4635
rect 1235 4605 1236 4635
rect 1204 4604 1236 4605
rect 1204 4524 1236 4556
rect 1204 4475 1236 4476
rect 1204 4445 1205 4475
rect 1205 4445 1235 4475
rect 1235 4445 1236 4475
rect 1204 4444 1236 4445
rect 1284 5515 1316 5516
rect 1284 5485 1285 5515
rect 1285 5485 1315 5515
rect 1315 5485 1316 5515
rect 1284 5484 1316 5485
rect 1284 5435 1316 5436
rect 1284 5405 1285 5435
rect 1285 5405 1315 5435
rect 1315 5405 1316 5435
rect 1284 5404 1316 5405
rect 1284 5324 1316 5356
rect 1284 5275 1316 5276
rect 1284 5245 1285 5275
rect 1285 5245 1315 5275
rect 1315 5245 1316 5275
rect 1284 5244 1316 5245
rect 1284 5195 1316 5196
rect 1284 5165 1285 5195
rect 1285 5165 1315 5195
rect 1315 5165 1316 5195
rect 1284 5164 1316 5165
rect 1284 5115 1316 5116
rect 1284 5085 1285 5115
rect 1285 5085 1315 5115
rect 1315 5085 1316 5115
rect 1284 5084 1316 5085
rect 1284 5035 1316 5036
rect 1284 5005 1285 5035
rect 1285 5005 1315 5035
rect 1315 5005 1316 5035
rect 1284 5004 1316 5005
rect 1284 4924 1316 4956
rect 1284 4875 1316 4876
rect 1284 4845 1285 4875
rect 1285 4845 1315 4875
rect 1315 4845 1316 4875
rect 1284 4844 1316 4845
rect 1284 4764 1316 4796
rect 1284 4715 1316 4716
rect 1284 4685 1285 4715
rect 1285 4685 1315 4715
rect 1315 4685 1316 4715
rect 1284 4684 1316 4685
rect 1284 4635 1316 4636
rect 1284 4605 1285 4635
rect 1285 4605 1315 4635
rect 1315 4605 1316 4635
rect 1284 4604 1316 4605
rect 1284 4524 1316 4556
rect 1284 4475 1316 4476
rect 1284 4445 1285 4475
rect 1285 4445 1315 4475
rect 1315 4445 1316 4475
rect 1284 4444 1316 4445
rect 1364 5515 1396 5516
rect 1364 5485 1365 5515
rect 1365 5485 1395 5515
rect 1395 5485 1396 5515
rect 1364 5484 1396 5485
rect 1364 5435 1396 5436
rect 1364 5405 1365 5435
rect 1365 5405 1395 5435
rect 1395 5405 1396 5435
rect 1364 5404 1396 5405
rect 1364 5324 1396 5356
rect 1364 5275 1396 5276
rect 1364 5245 1365 5275
rect 1365 5245 1395 5275
rect 1395 5245 1396 5275
rect 1364 5244 1396 5245
rect 1364 5195 1396 5196
rect 1364 5165 1365 5195
rect 1365 5165 1395 5195
rect 1395 5165 1396 5195
rect 1364 5164 1396 5165
rect 1364 5115 1396 5116
rect 1364 5085 1365 5115
rect 1365 5085 1395 5115
rect 1395 5085 1396 5115
rect 1364 5084 1396 5085
rect 1364 5035 1396 5036
rect 1364 5005 1365 5035
rect 1365 5005 1395 5035
rect 1395 5005 1396 5035
rect 1364 5004 1396 5005
rect 1364 4924 1396 4956
rect 1364 4875 1396 4876
rect 1364 4845 1365 4875
rect 1365 4845 1395 4875
rect 1395 4845 1396 4875
rect 1364 4844 1396 4845
rect 1364 4764 1396 4796
rect 1364 4715 1396 4716
rect 1364 4685 1365 4715
rect 1365 4685 1395 4715
rect 1395 4685 1396 4715
rect 1364 4684 1396 4685
rect 1364 4635 1396 4636
rect 1364 4605 1365 4635
rect 1365 4605 1395 4635
rect 1395 4605 1396 4635
rect 1364 4604 1396 4605
rect 1364 4524 1396 4556
rect 1364 4475 1396 4476
rect 1364 4445 1365 4475
rect 1365 4445 1395 4475
rect 1395 4445 1396 4475
rect 1364 4444 1396 4445
rect 1444 5515 1476 5516
rect 1444 5485 1445 5515
rect 1445 5485 1475 5515
rect 1475 5485 1476 5515
rect 1444 5484 1476 5485
rect 1444 5435 1476 5436
rect 1444 5405 1445 5435
rect 1445 5405 1475 5435
rect 1475 5405 1476 5435
rect 1444 5404 1476 5405
rect 1444 5324 1476 5356
rect 1444 5275 1476 5276
rect 1444 5245 1445 5275
rect 1445 5245 1475 5275
rect 1475 5245 1476 5275
rect 1444 5244 1476 5245
rect 1444 5195 1476 5196
rect 1444 5165 1445 5195
rect 1445 5165 1475 5195
rect 1475 5165 1476 5195
rect 1444 5164 1476 5165
rect 1444 5115 1476 5116
rect 1444 5085 1445 5115
rect 1445 5085 1475 5115
rect 1475 5085 1476 5115
rect 1444 5084 1476 5085
rect 1444 5035 1476 5036
rect 1444 5005 1445 5035
rect 1445 5005 1475 5035
rect 1475 5005 1476 5035
rect 1444 5004 1476 5005
rect 1444 4924 1476 4956
rect 1444 4875 1476 4876
rect 1444 4845 1445 4875
rect 1445 4845 1475 4875
rect 1475 4845 1476 4875
rect 1444 4844 1476 4845
rect 1444 4764 1476 4796
rect 1444 4715 1476 4716
rect 1444 4685 1445 4715
rect 1445 4685 1475 4715
rect 1475 4685 1476 4715
rect 1444 4684 1476 4685
rect 1444 4635 1476 4636
rect 1444 4605 1445 4635
rect 1445 4605 1475 4635
rect 1475 4605 1476 4635
rect 1444 4604 1476 4605
rect 1444 4524 1476 4556
rect 1444 4475 1476 4476
rect 1444 4445 1445 4475
rect 1445 4445 1475 4475
rect 1475 4445 1476 4475
rect 1444 4444 1476 4445
rect 1524 5515 1556 5516
rect 1524 5485 1525 5515
rect 1525 5485 1555 5515
rect 1555 5485 1556 5515
rect 1524 5484 1556 5485
rect 1524 5435 1556 5436
rect 1524 5405 1525 5435
rect 1525 5405 1555 5435
rect 1555 5405 1556 5435
rect 1524 5404 1556 5405
rect 1524 5324 1556 5356
rect 1524 5275 1556 5276
rect 1524 5245 1525 5275
rect 1525 5245 1555 5275
rect 1555 5245 1556 5275
rect 1524 5244 1556 5245
rect 1524 5195 1556 5196
rect 1524 5165 1525 5195
rect 1525 5165 1555 5195
rect 1555 5165 1556 5195
rect 1524 5164 1556 5165
rect 1524 5115 1556 5116
rect 1524 5085 1525 5115
rect 1525 5085 1555 5115
rect 1555 5085 1556 5115
rect 1524 5084 1556 5085
rect 1524 5035 1556 5036
rect 1524 5005 1525 5035
rect 1525 5005 1555 5035
rect 1555 5005 1556 5035
rect 1524 5004 1556 5005
rect 1524 4924 1556 4956
rect 1524 4875 1556 4876
rect 1524 4845 1525 4875
rect 1525 4845 1555 4875
rect 1555 4845 1556 4875
rect 1524 4844 1556 4845
rect 1524 4764 1556 4796
rect 1524 4715 1556 4716
rect 1524 4685 1525 4715
rect 1525 4685 1555 4715
rect 1555 4685 1556 4715
rect 1524 4684 1556 4685
rect 1524 4635 1556 4636
rect 1524 4605 1525 4635
rect 1525 4605 1555 4635
rect 1555 4605 1556 4635
rect 1524 4604 1556 4605
rect 1524 4524 1556 4556
rect 1524 4475 1556 4476
rect 1524 4445 1525 4475
rect 1525 4445 1555 4475
rect 1555 4445 1556 4475
rect 1524 4444 1556 4445
rect 1604 5515 1636 5516
rect 1604 5485 1605 5515
rect 1605 5485 1635 5515
rect 1635 5485 1636 5515
rect 1604 5484 1636 5485
rect 1604 5435 1636 5436
rect 1604 5405 1605 5435
rect 1605 5405 1635 5435
rect 1635 5405 1636 5435
rect 1604 5404 1636 5405
rect 1604 5324 1636 5356
rect 1604 5275 1636 5276
rect 1604 5245 1605 5275
rect 1605 5245 1635 5275
rect 1635 5245 1636 5275
rect 1604 5244 1636 5245
rect 1604 5195 1636 5196
rect 1604 5165 1605 5195
rect 1605 5165 1635 5195
rect 1635 5165 1636 5195
rect 1604 5164 1636 5165
rect 1604 5115 1636 5116
rect 1604 5085 1605 5115
rect 1605 5085 1635 5115
rect 1635 5085 1636 5115
rect 1604 5084 1636 5085
rect 1604 5035 1636 5036
rect 1604 5005 1605 5035
rect 1605 5005 1635 5035
rect 1635 5005 1636 5035
rect 1604 5004 1636 5005
rect 1604 4924 1636 4956
rect 1604 4875 1636 4876
rect 1604 4845 1605 4875
rect 1605 4845 1635 4875
rect 1635 4845 1636 4875
rect 1604 4844 1636 4845
rect 1604 4764 1636 4796
rect 1604 4715 1636 4716
rect 1604 4685 1605 4715
rect 1605 4685 1635 4715
rect 1635 4685 1636 4715
rect 1604 4684 1636 4685
rect 1604 4635 1636 4636
rect 1604 4605 1605 4635
rect 1605 4605 1635 4635
rect 1635 4605 1636 4635
rect 1604 4604 1636 4605
rect 1604 4524 1636 4556
rect 1604 4475 1636 4476
rect 1604 4445 1605 4475
rect 1605 4445 1635 4475
rect 1635 4445 1636 4475
rect 1604 4444 1636 4445
rect 1684 5515 1716 5516
rect 1684 5485 1685 5515
rect 1685 5485 1715 5515
rect 1715 5485 1716 5515
rect 1684 5484 1716 5485
rect 1684 5435 1716 5436
rect 1684 5405 1685 5435
rect 1685 5405 1715 5435
rect 1715 5405 1716 5435
rect 1684 5404 1716 5405
rect 1684 5324 1716 5356
rect 1684 5275 1716 5276
rect 1684 5245 1685 5275
rect 1685 5245 1715 5275
rect 1715 5245 1716 5275
rect 1684 5244 1716 5245
rect 1684 5195 1716 5196
rect 1684 5165 1685 5195
rect 1685 5165 1715 5195
rect 1715 5165 1716 5195
rect 1684 5164 1716 5165
rect 1684 5115 1716 5116
rect 1684 5085 1685 5115
rect 1685 5085 1715 5115
rect 1715 5085 1716 5115
rect 1684 5084 1716 5085
rect 1684 5035 1716 5036
rect 1684 5005 1685 5035
rect 1685 5005 1715 5035
rect 1715 5005 1716 5035
rect 1684 5004 1716 5005
rect 1684 4924 1716 4956
rect 1684 4875 1716 4876
rect 1684 4845 1685 4875
rect 1685 4845 1715 4875
rect 1715 4845 1716 4875
rect 1684 4844 1716 4845
rect 1684 4764 1716 4796
rect 1684 4715 1716 4716
rect 1684 4685 1685 4715
rect 1685 4685 1715 4715
rect 1715 4685 1716 4715
rect 1684 4684 1716 4685
rect 1684 4635 1716 4636
rect 1684 4605 1685 4635
rect 1685 4605 1715 4635
rect 1715 4605 1716 4635
rect 1684 4604 1716 4605
rect 1684 4524 1716 4556
rect 1684 4475 1716 4476
rect 1684 4445 1685 4475
rect 1685 4445 1715 4475
rect 1715 4445 1716 4475
rect 1684 4444 1716 4445
rect 1764 5515 1796 5516
rect 1764 5485 1765 5515
rect 1765 5485 1795 5515
rect 1795 5485 1796 5515
rect 1764 5484 1796 5485
rect 1764 5435 1796 5436
rect 1764 5405 1765 5435
rect 1765 5405 1795 5435
rect 1795 5405 1796 5435
rect 1764 5404 1796 5405
rect 1764 5324 1796 5356
rect 1764 5275 1796 5276
rect 1764 5245 1765 5275
rect 1765 5245 1795 5275
rect 1795 5245 1796 5275
rect 1764 5244 1796 5245
rect 1764 5195 1796 5196
rect 1764 5165 1765 5195
rect 1765 5165 1795 5195
rect 1795 5165 1796 5195
rect 1764 5164 1796 5165
rect 1764 5115 1796 5116
rect 1764 5085 1765 5115
rect 1765 5085 1795 5115
rect 1795 5085 1796 5115
rect 1764 5084 1796 5085
rect 1764 5035 1796 5036
rect 1764 5005 1765 5035
rect 1765 5005 1795 5035
rect 1795 5005 1796 5035
rect 1764 5004 1796 5005
rect 1764 4924 1796 4956
rect 1764 4875 1796 4876
rect 1764 4845 1765 4875
rect 1765 4845 1795 4875
rect 1795 4845 1796 4875
rect 1764 4844 1796 4845
rect 1764 4764 1796 4796
rect 1764 4715 1796 4716
rect 1764 4685 1765 4715
rect 1765 4685 1795 4715
rect 1795 4685 1796 4715
rect 1764 4684 1796 4685
rect 1764 4635 1796 4636
rect 1764 4605 1765 4635
rect 1765 4605 1795 4635
rect 1795 4605 1796 4635
rect 1764 4604 1796 4605
rect 1764 4524 1796 4556
rect 1764 4475 1796 4476
rect 1764 4445 1765 4475
rect 1765 4445 1795 4475
rect 1795 4445 1796 4475
rect 1764 4444 1796 4445
rect 1844 5515 1876 5516
rect 1844 5485 1845 5515
rect 1845 5485 1875 5515
rect 1875 5485 1876 5515
rect 1844 5484 1876 5485
rect 1844 5435 1876 5436
rect 1844 5405 1845 5435
rect 1845 5405 1875 5435
rect 1875 5405 1876 5435
rect 1844 5404 1876 5405
rect 1844 5324 1876 5356
rect 1844 5275 1876 5276
rect 1844 5245 1845 5275
rect 1845 5245 1875 5275
rect 1875 5245 1876 5275
rect 1844 5244 1876 5245
rect 1844 5195 1876 5196
rect 1844 5165 1845 5195
rect 1845 5165 1875 5195
rect 1875 5165 1876 5195
rect 1844 5164 1876 5165
rect 1844 5115 1876 5116
rect 1844 5085 1845 5115
rect 1845 5085 1875 5115
rect 1875 5085 1876 5115
rect 1844 5084 1876 5085
rect 1844 5035 1876 5036
rect 1844 5005 1845 5035
rect 1845 5005 1875 5035
rect 1875 5005 1876 5035
rect 1844 5004 1876 5005
rect 1844 4924 1876 4956
rect 1844 4875 1876 4876
rect 1844 4845 1845 4875
rect 1845 4845 1875 4875
rect 1875 4845 1876 4875
rect 1844 4844 1876 4845
rect 1844 4764 1876 4796
rect 1844 4715 1876 4716
rect 1844 4685 1845 4715
rect 1845 4685 1875 4715
rect 1875 4685 1876 4715
rect 1844 4684 1876 4685
rect 1844 4635 1876 4636
rect 1844 4605 1845 4635
rect 1845 4605 1875 4635
rect 1875 4605 1876 4635
rect 1844 4604 1876 4605
rect 1844 4524 1876 4556
rect 1844 4475 1876 4476
rect 1844 4445 1845 4475
rect 1845 4445 1875 4475
rect 1875 4445 1876 4475
rect 1844 4444 1876 4445
rect 1924 5515 1956 5516
rect 1924 5485 1925 5515
rect 1925 5485 1955 5515
rect 1955 5485 1956 5515
rect 1924 5484 1956 5485
rect 1924 5435 1956 5436
rect 1924 5405 1925 5435
rect 1925 5405 1955 5435
rect 1955 5405 1956 5435
rect 1924 5404 1956 5405
rect 1924 5324 1956 5356
rect 1924 5275 1956 5276
rect 1924 5245 1925 5275
rect 1925 5245 1955 5275
rect 1955 5245 1956 5275
rect 1924 5244 1956 5245
rect 1924 5195 1956 5196
rect 1924 5165 1925 5195
rect 1925 5165 1955 5195
rect 1955 5165 1956 5195
rect 1924 5164 1956 5165
rect 1924 5115 1956 5116
rect 1924 5085 1925 5115
rect 1925 5085 1955 5115
rect 1955 5085 1956 5115
rect 1924 5084 1956 5085
rect 1924 5035 1956 5036
rect 1924 5005 1925 5035
rect 1925 5005 1955 5035
rect 1955 5005 1956 5035
rect 1924 5004 1956 5005
rect 1924 4924 1956 4956
rect 1924 4875 1956 4876
rect 1924 4845 1925 4875
rect 1925 4845 1955 4875
rect 1955 4845 1956 4875
rect 1924 4844 1956 4845
rect 1924 4764 1956 4796
rect 1924 4715 1956 4716
rect 1924 4685 1925 4715
rect 1925 4685 1955 4715
rect 1955 4685 1956 4715
rect 1924 4684 1956 4685
rect 1924 4635 1956 4636
rect 1924 4605 1925 4635
rect 1925 4605 1955 4635
rect 1955 4605 1956 4635
rect 1924 4604 1956 4605
rect 1924 4524 1956 4556
rect 1924 4475 1956 4476
rect 1924 4445 1925 4475
rect 1925 4445 1955 4475
rect 1955 4445 1956 4475
rect 1924 4444 1956 4445
rect 2004 5515 2036 5516
rect 2004 5485 2005 5515
rect 2005 5485 2035 5515
rect 2035 5485 2036 5515
rect 2004 5484 2036 5485
rect 2004 5435 2036 5436
rect 2004 5405 2005 5435
rect 2005 5405 2035 5435
rect 2035 5405 2036 5435
rect 2004 5404 2036 5405
rect 2004 5324 2036 5356
rect 2004 5275 2036 5276
rect 2004 5245 2005 5275
rect 2005 5245 2035 5275
rect 2035 5245 2036 5275
rect 2004 5244 2036 5245
rect 2004 5195 2036 5196
rect 2004 5165 2005 5195
rect 2005 5165 2035 5195
rect 2035 5165 2036 5195
rect 2004 5164 2036 5165
rect 2004 5115 2036 5116
rect 2004 5085 2005 5115
rect 2005 5085 2035 5115
rect 2035 5085 2036 5115
rect 2004 5084 2036 5085
rect 2004 5035 2036 5036
rect 2004 5005 2005 5035
rect 2005 5005 2035 5035
rect 2035 5005 2036 5035
rect 2004 5004 2036 5005
rect 2004 4924 2036 4956
rect 2004 4875 2036 4876
rect 2004 4845 2005 4875
rect 2005 4845 2035 4875
rect 2035 4845 2036 4875
rect 2004 4844 2036 4845
rect 2004 4764 2036 4796
rect 2004 4715 2036 4716
rect 2004 4685 2005 4715
rect 2005 4685 2035 4715
rect 2035 4685 2036 4715
rect 2004 4684 2036 4685
rect 2004 4635 2036 4636
rect 2004 4605 2005 4635
rect 2005 4605 2035 4635
rect 2035 4605 2036 4635
rect 2004 4604 2036 4605
rect 2004 4524 2036 4556
rect 2004 4475 2036 4476
rect 2004 4445 2005 4475
rect 2005 4445 2035 4475
rect 2035 4445 2036 4475
rect 2004 4444 2036 4445
rect 2084 5515 2116 5516
rect 2084 5485 2085 5515
rect 2085 5485 2115 5515
rect 2115 5485 2116 5515
rect 2084 5484 2116 5485
rect 2084 5435 2116 5436
rect 2084 5405 2085 5435
rect 2085 5405 2115 5435
rect 2115 5405 2116 5435
rect 2084 5404 2116 5405
rect 2084 5324 2116 5356
rect 2084 5275 2116 5276
rect 2084 5245 2085 5275
rect 2085 5245 2115 5275
rect 2115 5245 2116 5275
rect 2084 5244 2116 5245
rect 2084 5195 2116 5196
rect 2084 5165 2085 5195
rect 2085 5165 2115 5195
rect 2115 5165 2116 5195
rect 2084 5164 2116 5165
rect 2084 5115 2116 5116
rect 2084 5085 2085 5115
rect 2085 5085 2115 5115
rect 2115 5085 2116 5115
rect 2084 5084 2116 5085
rect 2084 5035 2116 5036
rect 2084 5005 2085 5035
rect 2085 5005 2115 5035
rect 2115 5005 2116 5035
rect 2084 5004 2116 5005
rect 2084 4924 2116 4956
rect 2084 4875 2116 4876
rect 2084 4845 2085 4875
rect 2085 4845 2115 4875
rect 2115 4845 2116 4875
rect 2084 4844 2116 4845
rect 2084 4764 2116 4796
rect 2084 4715 2116 4716
rect 2084 4685 2085 4715
rect 2085 4685 2115 4715
rect 2115 4685 2116 4715
rect 2084 4684 2116 4685
rect 2084 4635 2116 4636
rect 2084 4605 2085 4635
rect 2085 4605 2115 4635
rect 2115 4605 2116 4635
rect 2084 4604 2116 4605
rect 2084 4524 2116 4556
rect 2084 4475 2116 4476
rect 2084 4445 2085 4475
rect 2085 4445 2115 4475
rect 2115 4445 2116 4475
rect 2084 4444 2116 4445
rect 2164 5515 2196 5516
rect 2164 5485 2165 5515
rect 2165 5485 2195 5515
rect 2195 5485 2196 5515
rect 2164 5484 2196 5485
rect 2164 5435 2196 5436
rect 2164 5405 2165 5435
rect 2165 5405 2195 5435
rect 2195 5405 2196 5435
rect 2164 5404 2196 5405
rect 2164 5324 2196 5356
rect 2164 5275 2196 5276
rect 2164 5245 2165 5275
rect 2165 5245 2195 5275
rect 2195 5245 2196 5275
rect 2164 5244 2196 5245
rect 2164 5195 2196 5196
rect 2164 5165 2165 5195
rect 2165 5165 2195 5195
rect 2195 5165 2196 5195
rect 2164 5164 2196 5165
rect 2164 5115 2196 5116
rect 2164 5085 2165 5115
rect 2165 5085 2195 5115
rect 2195 5085 2196 5115
rect 2164 5084 2196 5085
rect 2164 5035 2196 5036
rect 2164 5005 2165 5035
rect 2165 5005 2195 5035
rect 2195 5005 2196 5035
rect 2164 5004 2196 5005
rect 2164 4924 2196 4956
rect 2164 4875 2196 4876
rect 2164 4845 2165 4875
rect 2165 4845 2195 4875
rect 2195 4845 2196 4875
rect 2164 4844 2196 4845
rect 2164 4764 2196 4796
rect 2164 4715 2196 4716
rect 2164 4685 2165 4715
rect 2165 4685 2195 4715
rect 2195 4685 2196 4715
rect 2164 4684 2196 4685
rect 2164 4635 2196 4636
rect 2164 4605 2165 4635
rect 2165 4605 2195 4635
rect 2195 4605 2196 4635
rect 2164 4604 2196 4605
rect 2164 4524 2196 4556
rect 2164 4475 2196 4476
rect 2164 4445 2165 4475
rect 2165 4445 2195 4475
rect 2195 4445 2196 4475
rect 2164 4444 2196 4445
rect 2244 5515 2276 5516
rect 2244 5485 2245 5515
rect 2245 5485 2275 5515
rect 2275 5485 2276 5515
rect 2244 5484 2276 5485
rect 2244 5435 2276 5436
rect 2244 5405 2245 5435
rect 2245 5405 2275 5435
rect 2275 5405 2276 5435
rect 2244 5404 2276 5405
rect 2244 5324 2276 5356
rect 2244 5275 2276 5276
rect 2244 5245 2245 5275
rect 2245 5245 2275 5275
rect 2275 5245 2276 5275
rect 2244 5244 2276 5245
rect 2244 5195 2276 5196
rect 2244 5165 2245 5195
rect 2245 5165 2275 5195
rect 2275 5165 2276 5195
rect 2244 5164 2276 5165
rect 2244 5115 2276 5116
rect 2244 5085 2245 5115
rect 2245 5085 2275 5115
rect 2275 5085 2276 5115
rect 2244 5084 2276 5085
rect 2244 5035 2276 5036
rect 2244 5005 2245 5035
rect 2245 5005 2275 5035
rect 2275 5005 2276 5035
rect 2244 5004 2276 5005
rect 2244 4924 2276 4956
rect 2244 4875 2276 4876
rect 2244 4845 2245 4875
rect 2245 4845 2275 4875
rect 2275 4845 2276 4875
rect 2244 4844 2276 4845
rect 2244 4764 2276 4796
rect 2244 4715 2276 4716
rect 2244 4685 2245 4715
rect 2245 4685 2275 4715
rect 2275 4685 2276 4715
rect 2244 4684 2276 4685
rect 2244 4635 2276 4636
rect 2244 4605 2245 4635
rect 2245 4605 2275 4635
rect 2275 4605 2276 4635
rect 2244 4604 2276 4605
rect 2244 4524 2276 4556
rect 2244 4475 2276 4476
rect 2244 4445 2245 4475
rect 2245 4445 2275 4475
rect 2275 4445 2276 4475
rect 2244 4444 2276 4445
rect 2324 5515 2356 5516
rect 2324 5485 2325 5515
rect 2325 5485 2355 5515
rect 2355 5485 2356 5515
rect 2324 5484 2356 5485
rect 2324 5435 2356 5436
rect 2324 5405 2325 5435
rect 2325 5405 2355 5435
rect 2355 5405 2356 5435
rect 2324 5404 2356 5405
rect 2324 5324 2356 5356
rect 2324 5275 2356 5276
rect 2324 5245 2325 5275
rect 2325 5245 2355 5275
rect 2355 5245 2356 5275
rect 2324 5244 2356 5245
rect 2324 5195 2356 5196
rect 2324 5165 2325 5195
rect 2325 5165 2355 5195
rect 2355 5165 2356 5195
rect 2324 5164 2356 5165
rect 2324 5115 2356 5116
rect 2324 5085 2325 5115
rect 2325 5085 2355 5115
rect 2355 5085 2356 5115
rect 2324 5084 2356 5085
rect 2324 5035 2356 5036
rect 2324 5005 2325 5035
rect 2325 5005 2355 5035
rect 2355 5005 2356 5035
rect 2324 5004 2356 5005
rect 2324 4924 2356 4956
rect 2324 4875 2356 4876
rect 2324 4845 2325 4875
rect 2325 4845 2355 4875
rect 2355 4845 2356 4875
rect 2324 4844 2356 4845
rect 2324 4764 2356 4796
rect 2324 4715 2356 4716
rect 2324 4685 2325 4715
rect 2325 4685 2355 4715
rect 2355 4685 2356 4715
rect 2324 4684 2356 4685
rect 2324 4635 2356 4636
rect 2324 4605 2325 4635
rect 2325 4605 2355 4635
rect 2355 4605 2356 4635
rect 2324 4604 2356 4605
rect 2324 4524 2356 4556
rect 2324 4475 2356 4476
rect 2324 4445 2325 4475
rect 2325 4445 2355 4475
rect 2355 4445 2356 4475
rect 2324 4444 2356 4445
rect 2404 5515 2436 5516
rect 2404 5485 2405 5515
rect 2405 5485 2435 5515
rect 2435 5485 2436 5515
rect 2404 5484 2436 5485
rect 2404 5435 2436 5436
rect 2404 5405 2405 5435
rect 2405 5405 2435 5435
rect 2435 5405 2436 5435
rect 2404 5404 2436 5405
rect 2404 5324 2436 5356
rect 2404 5275 2436 5276
rect 2404 5245 2405 5275
rect 2405 5245 2435 5275
rect 2435 5245 2436 5275
rect 2404 5244 2436 5245
rect 2404 5195 2436 5196
rect 2404 5165 2405 5195
rect 2405 5165 2435 5195
rect 2435 5165 2436 5195
rect 2404 5164 2436 5165
rect 2404 5115 2436 5116
rect 2404 5085 2405 5115
rect 2405 5085 2435 5115
rect 2435 5085 2436 5115
rect 2404 5084 2436 5085
rect 2404 5035 2436 5036
rect 2404 5005 2405 5035
rect 2405 5005 2435 5035
rect 2435 5005 2436 5035
rect 2404 5004 2436 5005
rect 2404 4924 2436 4956
rect 2404 4875 2436 4876
rect 2404 4845 2405 4875
rect 2405 4845 2435 4875
rect 2435 4845 2436 4875
rect 2404 4844 2436 4845
rect 2404 4764 2436 4796
rect 2404 4715 2436 4716
rect 2404 4685 2405 4715
rect 2405 4685 2435 4715
rect 2435 4685 2436 4715
rect 2404 4684 2436 4685
rect 2404 4635 2436 4636
rect 2404 4605 2405 4635
rect 2405 4605 2435 4635
rect 2435 4605 2436 4635
rect 2404 4604 2436 4605
rect 2404 4524 2436 4556
rect 2404 4475 2436 4476
rect 2404 4445 2405 4475
rect 2405 4445 2435 4475
rect 2435 4445 2436 4475
rect 2404 4444 2436 4445
rect 2484 5515 2516 5516
rect 2484 5485 2485 5515
rect 2485 5485 2515 5515
rect 2515 5485 2516 5515
rect 2484 5484 2516 5485
rect 2484 5435 2516 5436
rect 2484 5405 2485 5435
rect 2485 5405 2515 5435
rect 2515 5405 2516 5435
rect 2484 5404 2516 5405
rect 2484 5324 2516 5356
rect 2484 5275 2516 5276
rect 2484 5245 2485 5275
rect 2485 5245 2515 5275
rect 2515 5245 2516 5275
rect 2484 5244 2516 5245
rect 2484 5195 2516 5196
rect 2484 5165 2485 5195
rect 2485 5165 2515 5195
rect 2515 5165 2516 5195
rect 2484 5164 2516 5165
rect 2484 5115 2516 5116
rect 2484 5085 2485 5115
rect 2485 5085 2515 5115
rect 2515 5085 2516 5115
rect 2484 5084 2516 5085
rect 2484 5035 2516 5036
rect 2484 5005 2485 5035
rect 2485 5005 2515 5035
rect 2515 5005 2516 5035
rect 2484 5004 2516 5005
rect 2484 4924 2516 4956
rect 2484 4875 2516 4876
rect 2484 4845 2485 4875
rect 2485 4845 2515 4875
rect 2515 4845 2516 4875
rect 2484 4844 2516 4845
rect 2484 4764 2516 4796
rect 2484 4715 2516 4716
rect 2484 4685 2485 4715
rect 2485 4685 2515 4715
rect 2515 4685 2516 4715
rect 2484 4684 2516 4685
rect 2484 4635 2516 4636
rect 2484 4605 2485 4635
rect 2485 4605 2515 4635
rect 2515 4605 2516 4635
rect 2484 4604 2516 4605
rect 2484 4524 2516 4556
rect 2484 4475 2516 4476
rect 2484 4445 2485 4475
rect 2485 4445 2515 4475
rect 2515 4445 2516 4475
rect 2484 4444 2516 4445
rect 2564 5515 2596 5516
rect 2564 5485 2565 5515
rect 2565 5485 2595 5515
rect 2595 5485 2596 5515
rect 2564 5484 2596 5485
rect 2564 5435 2596 5436
rect 2564 5405 2565 5435
rect 2565 5405 2595 5435
rect 2595 5405 2596 5435
rect 2564 5404 2596 5405
rect 2564 5324 2596 5356
rect 2564 5275 2596 5276
rect 2564 5245 2565 5275
rect 2565 5245 2595 5275
rect 2595 5245 2596 5275
rect 2564 5244 2596 5245
rect 2564 5195 2596 5196
rect 2564 5165 2565 5195
rect 2565 5165 2595 5195
rect 2595 5165 2596 5195
rect 2564 5164 2596 5165
rect 2564 5115 2596 5116
rect 2564 5085 2565 5115
rect 2565 5085 2595 5115
rect 2595 5085 2596 5115
rect 2564 5084 2596 5085
rect 2564 5035 2596 5036
rect 2564 5005 2565 5035
rect 2565 5005 2595 5035
rect 2595 5005 2596 5035
rect 2564 5004 2596 5005
rect 2564 4924 2596 4956
rect 2564 4875 2596 4876
rect 2564 4845 2565 4875
rect 2565 4845 2595 4875
rect 2595 4845 2596 4875
rect 2564 4844 2596 4845
rect 2564 4764 2596 4796
rect 2564 4715 2596 4716
rect 2564 4685 2565 4715
rect 2565 4685 2595 4715
rect 2595 4685 2596 4715
rect 2564 4684 2596 4685
rect 2564 4635 2596 4636
rect 2564 4605 2565 4635
rect 2565 4605 2595 4635
rect 2595 4605 2596 4635
rect 2564 4604 2596 4605
rect 2564 4524 2596 4556
rect 2564 4475 2596 4476
rect 2564 4445 2565 4475
rect 2565 4445 2595 4475
rect 2595 4445 2596 4475
rect 2564 4444 2596 4445
rect 2644 5515 2676 5516
rect 2644 5485 2645 5515
rect 2645 5485 2675 5515
rect 2675 5485 2676 5515
rect 2644 5484 2676 5485
rect 2644 5435 2676 5436
rect 2644 5405 2645 5435
rect 2645 5405 2675 5435
rect 2675 5405 2676 5435
rect 2644 5404 2676 5405
rect 2644 5324 2676 5356
rect 2644 5275 2676 5276
rect 2644 5245 2645 5275
rect 2645 5245 2675 5275
rect 2675 5245 2676 5275
rect 2644 5244 2676 5245
rect 2644 5195 2676 5196
rect 2644 5165 2645 5195
rect 2645 5165 2675 5195
rect 2675 5165 2676 5195
rect 2644 5164 2676 5165
rect 2644 5115 2676 5116
rect 2644 5085 2645 5115
rect 2645 5085 2675 5115
rect 2675 5085 2676 5115
rect 2644 5084 2676 5085
rect 2644 5035 2676 5036
rect 2644 5005 2645 5035
rect 2645 5005 2675 5035
rect 2675 5005 2676 5035
rect 2644 5004 2676 5005
rect 2644 4924 2676 4956
rect 2644 4875 2676 4876
rect 2644 4845 2645 4875
rect 2645 4845 2675 4875
rect 2675 4845 2676 4875
rect 2644 4844 2676 4845
rect 2644 4764 2676 4796
rect 2644 4715 2676 4716
rect 2644 4685 2645 4715
rect 2645 4685 2675 4715
rect 2675 4685 2676 4715
rect 2644 4684 2676 4685
rect 2644 4635 2676 4636
rect 2644 4605 2645 4635
rect 2645 4605 2675 4635
rect 2675 4605 2676 4635
rect 2644 4604 2676 4605
rect 2644 4524 2676 4556
rect 2644 4475 2676 4476
rect 2644 4445 2645 4475
rect 2645 4445 2675 4475
rect 2675 4445 2676 4475
rect 2644 4444 2676 4445
rect 2724 5515 2756 5516
rect 2724 5485 2725 5515
rect 2725 5485 2755 5515
rect 2755 5485 2756 5515
rect 2724 5484 2756 5485
rect 2724 5435 2756 5436
rect 2724 5405 2725 5435
rect 2725 5405 2755 5435
rect 2755 5405 2756 5435
rect 2724 5404 2756 5405
rect 2724 5324 2756 5356
rect 2724 5275 2756 5276
rect 2724 5245 2725 5275
rect 2725 5245 2755 5275
rect 2755 5245 2756 5275
rect 2724 5244 2756 5245
rect 2724 5195 2756 5196
rect 2724 5165 2725 5195
rect 2725 5165 2755 5195
rect 2755 5165 2756 5195
rect 2724 5164 2756 5165
rect 2724 5115 2756 5116
rect 2724 5085 2725 5115
rect 2725 5085 2755 5115
rect 2755 5085 2756 5115
rect 2724 5084 2756 5085
rect 2724 5035 2756 5036
rect 2724 5005 2725 5035
rect 2725 5005 2755 5035
rect 2755 5005 2756 5035
rect 2724 5004 2756 5005
rect 2724 4924 2756 4956
rect 2724 4875 2756 4876
rect 2724 4845 2725 4875
rect 2725 4845 2755 4875
rect 2755 4845 2756 4875
rect 2724 4844 2756 4845
rect 2724 4764 2756 4796
rect 2724 4715 2756 4716
rect 2724 4685 2725 4715
rect 2725 4685 2755 4715
rect 2755 4685 2756 4715
rect 2724 4684 2756 4685
rect 2724 4635 2756 4636
rect 2724 4605 2725 4635
rect 2725 4605 2755 4635
rect 2755 4605 2756 4635
rect 2724 4604 2756 4605
rect 2724 4524 2756 4556
rect 2724 4475 2756 4476
rect 2724 4445 2725 4475
rect 2725 4445 2755 4475
rect 2755 4445 2756 4475
rect 2724 4444 2756 4445
rect 2804 5515 2836 5516
rect 2804 5485 2805 5515
rect 2805 5485 2835 5515
rect 2835 5485 2836 5515
rect 2804 5484 2836 5485
rect 2804 5435 2836 5436
rect 2804 5405 2805 5435
rect 2805 5405 2835 5435
rect 2835 5405 2836 5435
rect 2804 5404 2836 5405
rect 2804 5324 2836 5356
rect 2804 5275 2836 5276
rect 2804 5245 2805 5275
rect 2805 5245 2835 5275
rect 2835 5245 2836 5275
rect 2804 5244 2836 5245
rect 2804 5195 2836 5196
rect 2804 5165 2805 5195
rect 2805 5165 2835 5195
rect 2835 5165 2836 5195
rect 2804 5164 2836 5165
rect 2804 5115 2836 5116
rect 2804 5085 2805 5115
rect 2805 5085 2835 5115
rect 2835 5085 2836 5115
rect 2804 5084 2836 5085
rect 2804 5035 2836 5036
rect 2804 5005 2805 5035
rect 2805 5005 2835 5035
rect 2835 5005 2836 5035
rect 2804 5004 2836 5005
rect 2804 4924 2836 4956
rect 2804 4875 2836 4876
rect 2804 4845 2805 4875
rect 2805 4845 2835 4875
rect 2835 4845 2836 4875
rect 2804 4844 2836 4845
rect 2804 4764 2836 4796
rect 2804 4715 2836 4716
rect 2804 4685 2805 4715
rect 2805 4685 2835 4715
rect 2835 4685 2836 4715
rect 2804 4684 2836 4685
rect 2804 4635 2836 4636
rect 2804 4605 2805 4635
rect 2805 4605 2835 4635
rect 2835 4605 2836 4635
rect 2804 4604 2836 4605
rect 2804 4524 2836 4556
rect 2804 4475 2836 4476
rect 2804 4445 2805 4475
rect 2805 4445 2835 4475
rect 2835 4445 2836 4475
rect 2804 4444 2836 4445
rect 2884 5515 2916 5516
rect 2884 5485 2885 5515
rect 2885 5485 2915 5515
rect 2915 5485 2916 5515
rect 2884 5484 2916 5485
rect 2884 5435 2916 5436
rect 2884 5405 2885 5435
rect 2885 5405 2915 5435
rect 2915 5405 2916 5435
rect 2884 5404 2916 5405
rect 2884 5324 2916 5356
rect 2884 5275 2916 5276
rect 2884 5245 2885 5275
rect 2885 5245 2915 5275
rect 2915 5245 2916 5275
rect 2884 5244 2916 5245
rect 2884 5195 2916 5196
rect 2884 5165 2885 5195
rect 2885 5165 2915 5195
rect 2915 5165 2916 5195
rect 2884 5164 2916 5165
rect 2884 5115 2916 5116
rect 2884 5085 2885 5115
rect 2885 5085 2915 5115
rect 2915 5085 2916 5115
rect 2884 5084 2916 5085
rect 2884 5035 2916 5036
rect 2884 5005 2885 5035
rect 2885 5005 2915 5035
rect 2915 5005 2916 5035
rect 2884 5004 2916 5005
rect 2884 4924 2916 4956
rect 2884 4875 2916 4876
rect 2884 4845 2885 4875
rect 2885 4845 2915 4875
rect 2915 4845 2916 4875
rect 2884 4844 2916 4845
rect 2884 4764 2916 4796
rect 2884 4715 2916 4716
rect 2884 4685 2885 4715
rect 2885 4685 2915 4715
rect 2915 4685 2916 4715
rect 2884 4684 2916 4685
rect 2884 4635 2916 4636
rect 2884 4605 2885 4635
rect 2885 4605 2915 4635
rect 2915 4605 2916 4635
rect 2884 4604 2916 4605
rect 2884 4524 2916 4556
rect 2884 4475 2916 4476
rect 2884 4445 2885 4475
rect 2885 4445 2915 4475
rect 2915 4445 2916 4475
rect 2884 4444 2916 4445
rect 2964 5515 2996 5516
rect 2964 5485 2965 5515
rect 2965 5485 2995 5515
rect 2995 5485 2996 5515
rect 2964 5484 2996 5485
rect 2964 5435 2996 5436
rect 2964 5405 2965 5435
rect 2965 5405 2995 5435
rect 2995 5405 2996 5435
rect 2964 5404 2996 5405
rect 2964 5324 2996 5356
rect 2964 5275 2996 5276
rect 2964 5245 2965 5275
rect 2965 5245 2995 5275
rect 2995 5245 2996 5275
rect 2964 5244 2996 5245
rect 2964 5195 2996 5196
rect 2964 5165 2965 5195
rect 2965 5165 2995 5195
rect 2995 5165 2996 5195
rect 2964 5164 2996 5165
rect 2964 5115 2996 5116
rect 2964 5085 2965 5115
rect 2965 5085 2995 5115
rect 2995 5085 2996 5115
rect 2964 5084 2996 5085
rect 2964 5035 2996 5036
rect 2964 5005 2965 5035
rect 2965 5005 2995 5035
rect 2995 5005 2996 5035
rect 2964 5004 2996 5005
rect 2964 4924 2996 4956
rect 2964 4875 2996 4876
rect 2964 4845 2965 4875
rect 2965 4845 2995 4875
rect 2995 4845 2996 4875
rect 2964 4844 2996 4845
rect 2964 4764 2996 4796
rect 2964 4715 2996 4716
rect 2964 4685 2965 4715
rect 2965 4685 2995 4715
rect 2995 4685 2996 4715
rect 2964 4684 2996 4685
rect 2964 4635 2996 4636
rect 2964 4605 2965 4635
rect 2965 4605 2995 4635
rect 2995 4605 2996 4635
rect 2964 4604 2996 4605
rect 2964 4524 2996 4556
rect 2964 4475 2996 4476
rect 2964 4445 2965 4475
rect 2965 4445 2995 4475
rect 2995 4445 2996 4475
rect 2964 4444 2996 4445
rect 3044 5515 3076 5516
rect 3044 5485 3045 5515
rect 3045 5485 3075 5515
rect 3075 5485 3076 5515
rect 3044 5484 3076 5485
rect 3044 5435 3076 5436
rect 3044 5405 3045 5435
rect 3045 5405 3075 5435
rect 3075 5405 3076 5435
rect 3044 5404 3076 5405
rect 3044 5324 3076 5356
rect 3044 5275 3076 5276
rect 3044 5245 3045 5275
rect 3045 5245 3075 5275
rect 3075 5245 3076 5275
rect 3044 5244 3076 5245
rect 3044 5195 3076 5196
rect 3044 5165 3045 5195
rect 3045 5165 3075 5195
rect 3075 5165 3076 5195
rect 3044 5164 3076 5165
rect 3044 5115 3076 5116
rect 3044 5085 3045 5115
rect 3045 5085 3075 5115
rect 3075 5085 3076 5115
rect 3044 5084 3076 5085
rect 3044 5035 3076 5036
rect 3044 5005 3045 5035
rect 3045 5005 3075 5035
rect 3075 5005 3076 5035
rect 3044 5004 3076 5005
rect 3044 4924 3076 4956
rect 3044 4875 3076 4876
rect 3044 4845 3045 4875
rect 3045 4845 3075 4875
rect 3075 4845 3076 4875
rect 3044 4844 3076 4845
rect 3044 4764 3076 4796
rect 3044 4715 3076 4716
rect 3044 4685 3045 4715
rect 3045 4685 3075 4715
rect 3075 4685 3076 4715
rect 3044 4684 3076 4685
rect 3044 4635 3076 4636
rect 3044 4605 3045 4635
rect 3045 4605 3075 4635
rect 3075 4605 3076 4635
rect 3044 4604 3076 4605
rect 3044 4524 3076 4556
rect 3044 4475 3076 4476
rect 3044 4445 3045 4475
rect 3045 4445 3075 4475
rect 3075 4445 3076 4475
rect 3044 4444 3076 4445
rect 3124 5515 3156 5516
rect 3124 5485 3125 5515
rect 3125 5485 3155 5515
rect 3155 5485 3156 5515
rect 3124 5484 3156 5485
rect 3124 5435 3156 5436
rect 3124 5405 3125 5435
rect 3125 5405 3155 5435
rect 3155 5405 3156 5435
rect 3124 5404 3156 5405
rect 3124 5324 3156 5356
rect 3124 5275 3156 5276
rect 3124 5245 3125 5275
rect 3125 5245 3155 5275
rect 3155 5245 3156 5275
rect 3124 5244 3156 5245
rect 3124 5195 3156 5196
rect 3124 5165 3125 5195
rect 3125 5165 3155 5195
rect 3155 5165 3156 5195
rect 3124 5164 3156 5165
rect 3124 5115 3156 5116
rect 3124 5085 3125 5115
rect 3125 5085 3155 5115
rect 3155 5085 3156 5115
rect 3124 5084 3156 5085
rect 3124 5035 3156 5036
rect 3124 5005 3125 5035
rect 3125 5005 3155 5035
rect 3155 5005 3156 5035
rect 3124 5004 3156 5005
rect 3124 4924 3156 4956
rect 3124 4875 3156 4876
rect 3124 4845 3125 4875
rect 3125 4845 3155 4875
rect 3155 4845 3156 4875
rect 3124 4844 3156 4845
rect 3124 4764 3156 4796
rect 3124 4715 3156 4716
rect 3124 4685 3125 4715
rect 3125 4685 3155 4715
rect 3155 4685 3156 4715
rect 3124 4684 3156 4685
rect 3124 4635 3156 4636
rect 3124 4605 3125 4635
rect 3125 4605 3155 4635
rect 3155 4605 3156 4635
rect 3124 4604 3156 4605
rect 3124 4524 3156 4556
rect 3124 4475 3156 4476
rect 3124 4445 3125 4475
rect 3125 4445 3155 4475
rect 3155 4445 3156 4475
rect 3124 4444 3156 4445
rect 3204 5515 3236 5516
rect 3204 5485 3205 5515
rect 3205 5485 3235 5515
rect 3235 5485 3236 5515
rect 3204 5484 3236 5485
rect 3204 5435 3236 5436
rect 3204 5405 3205 5435
rect 3205 5405 3235 5435
rect 3235 5405 3236 5435
rect 3204 5404 3236 5405
rect 3204 5324 3236 5356
rect 3204 5275 3236 5276
rect 3204 5245 3205 5275
rect 3205 5245 3235 5275
rect 3235 5245 3236 5275
rect 3204 5244 3236 5245
rect 3204 5195 3236 5196
rect 3204 5165 3205 5195
rect 3205 5165 3235 5195
rect 3235 5165 3236 5195
rect 3204 5164 3236 5165
rect 3204 5115 3236 5116
rect 3204 5085 3205 5115
rect 3205 5085 3235 5115
rect 3235 5085 3236 5115
rect 3204 5084 3236 5085
rect 3204 5035 3236 5036
rect 3204 5005 3205 5035
rect 3205 5005 3235 5035
rect 3235 5005 3236 5035
rect 3204 5004 3236 5005
rect 3204 4924 3236 4956
rect 3204 4875 3236 4876
rect 3204 4845 3205 4875
rect 3205 4845 3235 4875
rect 3235 4845 3236 4875
rect 3204 4844 3236 4845
rect 3204 4764 3236 4796
rect 3204 4715 3236 4716
rect 3204 4685 3205 4715
rect 3205 4685 3235 4715
rect 3235 4685 3236 4715
rect 3204 4684 3236 4685
rect 3204 4635 3236 4636
rect 3204 4605 3205 4635
rect 3205 4605 3235 4635
rect 3235 4605 3236 4635
rect 3204 4604 3236 4605
rect 3204 4524 3236 4556
rect 3204 4475 3236 4476
rect 3204 4445 3205 4475
rect 3205 4445 3235 4475
rect 3235 4445 3236 4475
rect 3204 4444 3236 4445
rect 3284 5515 3316 5516
rect 3284 5485 3285 5515
rect 3285 5485 3315 5515
rect 3315 5485 3316 5515
rect 3284 5484 3316 5485
rect 3284 5435 3316 5436
rect 3284 5405 3285 5435
rect 3285 5405 3315 5435
rect 3315 5405 3316 5435
rect 3284 5404 3316 5405
rect 3284 5324 3316 5356
rect 3284 5275 3316 5276
rect 3284 5245 3285 5275
rect 3285 5245 3315 5275
rect 3315 5245 3316 5275
rect 3284 5244 3316 5245
rect 3284 5195 3316 5196
rect 3284 5165 3285 5195
rect 3285 5165 3315 5195
rect 3315 5165 3316 5195
rect 3284 5164 3316 5165
rect 3284 5115 3316 5116
rect 3284 5085 3285 5115
rect 3285 5085 3315 5115
rect 3315 5085 3316 5115
rect 3284 5084 3316 5085
rect 3284 5035 3316 5036
rect 3284 5005 3285 5035
rect 3285 5005 3315 5035
rect 3315 5005 3316 5035
rect 3284 5004 3316 5005
rect 3284 4924 3316 4956
rect 3284 4875 3316 4876
rect 3284 4845 3285 4875
rect 3285 4845 3315 4875
rect 3315 4845 3316 4875
rect 3284 4844 3316 4845
rect 3284 4764 3316 4796
rect 3284 4715 3316 4716
rect 3284 4685 3285 4715
rect 3285 4685 3315 4715
rect 3315 4685 3316 4715
rect 3284 4684 3316 4685
rect 3284 4635 3316 4636
rect 3284 4605 3285 4635
rect 3285 4605 3315 4635
rect 3315 4605 3316 4635
rect 3284 4604 3316 4605
rect 3284 4524 3316 4556
rect 3284 4475 3316 4476
rect 3284 4445 3285 4475
rect 3285 4445 3315 4475
rect 3315 4445 3316 4475
rect 3284 4444 3316 4445
rect 3364 5515 3396 5516
rect 3364 5485 3365 5515
rect 3365 5485 3395 5515
rect 3395 5485 3396 5515
rect 3364 5484 3396 5485
rect 3364 5435 3396 5436
rect 3364 5405 3365 5435
rect 3365 5405 3395 5435
rect 3395 5405 3396 5435
rect 3364 5404 3396 5405
rect 3364 5324 3396 5356
rect 3364 5275 3396 5276
rect 3364 5245 3365 5275
rect 3365 5245 3395 5275
rect 3395 5245 3396 5275
rect 3364 5244 3396 5245
rect 3364 5195 3396 5196
rect 3364 5165 3365 5195
rect 3365 5165 3395 5195
rect 3395 5165 3396 5195
rect 3364 5164 3396 5165
rect 3364 5115 3396 5116
rect 3364 5085 3365 5115
rect 3365 5085 3395 5115
rect 3395 5085 3396 5115
rect 3364 5084 3396 5085
rect 3364 5035 3396 5036
rect 3364 5005 3365 5035
rect 3365 5005 3395 5035
rect 3395 5005 3396 5035
rect 3364 5004 3396 5005
rect 3364 4924 3396 4956
rect 3364 4875 3396 4876
rect 3364 4845 3365 4875
rect 3365 4845 3395 4875
rect 3395 4845 3396 4875
rect 3364 4844 3396 4845
rect 3364 4764 3396 4796
rect 3364 4715 3396 4716
rect 3364 4685 3365 4715
rect 3365 4685 3395 4715
rect 3395 4685 3396 4715
rect 3364 4684 3396 4685
rect 3364 4635 3396 4636
rect 3364 4605 3365 4635
rect 3365 4605 3395 4635
rect 3395 4605 3396 4635
rect 3364 4604 3396 4605
rect 3364 4524 3396 4556
rect 3364 4475 3396 4476
rect 3364 4445 3365 4475
rect 3365 4445 3395 4475
rect 3395 4445 3396 4475
rect 3364 4444 3396 4445
rect 3444 5515 3476 5516
rect 3444 5485 3445 5515
rect 3445 5485 3475 5515
rect 3475 5485 3476 5515
rect 3444 5484 3476 5485
rect 3444 5435 3476 5436
rect 3444 5405 3445 5435
rect 3445 5405 3475 5435
rect 3475 5405 3476 5435
rect 3444 5404 3476 5405
rect 3444 5324 3476 5356
rect 3444 5275 3476 5276
rect 3444 5245 3445 5275
rect 3445 5245 3475 5275
rect 3475 5245 3476 5275
rect 3444 5244 3476 5245
rect 3444 5195 3476 5196
rect 3444 5165 3445 5195
rect 3445 5165 3475 5195
rect 3475 5165 3476 5195
rect 3444 5164 3476 5165
rect 3444 5115 3476 5116
rect 3444 5085 3445 5115
rect 3445 5085 3475 5115
rect 3475 5085 3476 5115
rect 3444 5084 3476 5085
rect 3444 5035 3476 5036
rect 3444 5005 3445 5035
rect 3445 5005 3475 5035
rect 3475 5005 3476 5035
rect 3444 5004 3476 5005
rect 3444 4924 3476 4956
rect 3444 4875 3476 4876
rect 3444 4845 3445 4875
rect 3445 4845 3475 4875
rect 3475 4845 3476 4875
rect 3444 4844 3476 4845
rect 3444 4764 3476 4796
rect 3444 4715 3476 4716
rect 3444 4685 3445 4715
rect 3445 4685 3475 4715
rect 3475 4685 3476 4715
rect 3444 4684 3476 4685
rect 3444 4635 3476 4636
rect 3444 4605 3445 4635
rect 3445 4605 3475 4635
rect 3475 4605 3476 4635
rect 3444 4604 3476 4605
rect 3444 4524 3476 4556
rect 3444 4475 3476 4476
rect 3444 4445 3445 4475
rect 3445 4445 3475 4475
rect 3475 4445 3476 4475
rect 3444 4444 3476 4445
rect 3524 5515 3556 5516
rect 3524 5485 3525 5515
rect 3525 5485 3555 5515
rect 3555 5485 3556 5515
rect 3524 5484 3556 5485
rect 3524 5435 3556 5436
rect 3524 5405 3525 5435
rect 3525 5405 3555 5435
rect 3555 5405 3556 5435
rect 3524 5404 3556 5405
rect 3524 5324 3556 5356
rect 3524 5275 3556 5276
rect 3524 5245 3525 5275
rect 3525 5245 3555 5275
rect 3555 5245 3556 5275
rect 3524 5244 3556 5245
rect 3524 5195 3556 5196
rect 3524 5165 3525 5195
rect 3525 5165 3555 5195
rect 3555 5165 3556 5195
rect 3524 5164 3556 5165
rect 3524 5115 3556 5116
rect 3524 5085 3525 5115
rect 3525 5085 3555 5115
rect 3555 5085 3556 5115
rect 3524 5084 3556 5085
rect 3524 5035 3556 5036
rect 3524 5005 3525 5035
rect 3525 5005 3555 5035
rect 3555 5005 3556 5035
rect 3524 5004 3556 5005
rect 3524 4924 3556 4956
rect 3524 4875 3556 4876
rect 3524 4845 3525 4875
rect 3525 4845 3555 4875
rect 3555 4845 3556 4875
rect 3524 4844 3556 4845
rect 3524 4764 3556 4796
rect 3524 4715 3556 4716
rect 3524 4685 3525 4715
rect 3525 4685 3555 4715
rect 3555 4685 3556 4715
rect 3524 4684 3556 4685
rect 3524 4635 3556 4636
rect 3524 4605 3525 4635
rect 3525 4605 3555 4635
rect 3555 4605 3556 4635
rect 3524 4604 3556 4605
rect 3524 4524 3556 4556
rect 3524 4475 3556 4476
rect 3524 4445 3525 4475
rect 3525 4445 3555 4475
rect 3555 4445 3556 4475
rect 3524 4444 3556 4445
rect 3604 5515 3636 5516
rect 3604 5485 3605 5515
rect 3605 5485 3635 5515
rect 3635 5485 3636 5515
rect 3604 5484 3636 5485
rect 3604 5435 3636 5436
rect 3604 5405 3605 5435
rect 3605 5405 3635 5435
rect 3635 5405 3636 5435
rect 3604 5404 3636 5405
rect 3604 5324 3636 5356
rect 3604 5275 3636 5276
rect 3604 5245 3605 5275
rect 3605 5245 3635 5275
rect 3635 5245 3636 5275
rect 3604 5244 3636 5245
rect 3604 5195 3636 5196
rect 3604 5165 3605 5195
rect 3605 5165 3635 5195
rect 3635 5165 3636 5195
rect 3604 5164 3636 5165
rect 3604 5115 3636 5116
rect 3604 5085 3605 5115
rect 3605 5085 3635 5115
rect 3635 5085 3636 5115
rect 3604 5084 3636 5085
rect 3604 5035 3636 5036
rect 3604 5005 3605 5035
rect 3605 5005 3635 5035
rect 3635 5005 3636 5035
rect 3604 5004 3636 5005
rect 3604 4924 3636 4956
rect 3604 4875 3636 4876
rect 3604 4845 3605 4875
rect 3605 4845 3635 4875
rect 3635 4845 3636 4875
rect 3604 4844 3636 4845
rect 3604 4764 3636 4796
rect 3604 4715 3636 4716
rect 3604 4685 3605 4715
rect 3605 4685 3635 4715
rect 3635 4685 3636 4715
rect 3604 4684 3636 4685
rect 3604 4635 3636 4636
rect 3604 4605 3605 4635
rect 3605 4605 3635 4635
rect 3635 4605 3636 4635
rect 3604 4604 3636 4605
rect 3604 4524 3636 4556
rect 3604 4475 3636 4476
rect 3604 4445 3605 4475
rect 3605 4445 3635 4475
rect 3635 4445 3636 4475
rect 3604 4444 3636 4445
rect 3684 5515 3716 5516
rect 3684 5485 3685 5515
rect 3685 5485 3715 5515
rect 3715 5485 3716 5515
rect 3684 5484 3716 5485
rect 3684 5435 3716 5436
rect 3684 5405 3685 5435
rect 3685 5405 3715 5435
rect 3715 5405 3716 5435
rect 3684 5404 3716 5405
rect 3684 5324 3716 5356
rect 3684 5275 3716 5276
rect 3684 5245 3685 5275
rect 3685 5245 3715 5275
rect 3715 5245 3716 5275
rect 3684 5244 3716 5245
rect 3684 5195 3716 5196
rect 3684 5165 3685 5195
rect 3685 5165 3715 5195
rect 3715 5165 3716 5195
rect 3684 5164 3716 5165
rect 3684 5115 3716 5116
rect 3684 5085 3685 5115
rect 3685 5085 3715 5115
rect 3715 5085 3716 5115
rect 3684 5084 3716 5085
rect 3684 5035 3716 5036
rect 3684 5005 3685 5035
rect 3685 5005 3715 5035
rect 3715 5005 3716 5035
rect 3684 5004 3716 5005
rect 3684 4924 3716 4956
rect 3684 4875 3716 4876
rect 3684 4845 3685 4875
rect 3685 4845 3715 4875
rect 3715 4845 3716 4875
rect 3684 4844 3716 4845
rect 3684 4764 3716 4796
rect 3684 4715 3716 4716
rect 3684 4685 3685 4715
rect 3685 4685 3715 4715
rect 3715 4685 3716 4715
rect 3684 4684 3716 4685
rect 3684 4635 3716 4636
rect 3684 4605 3685 4635
rect 3685 4605 3715 4635
rect 3715 4605 3716 4635
rect 3684 4604 3716 4605
rect 3684 4524 3716 4556
rect 3684 4475 3716 4476
rect 3684 4445 3685 4475
rect 3685 4445 3715 4475
rect 3715 4445 3716 4475
rect 3684 4444 3716 4445
rect 3764 5515 3796 5516
rect 3764 5485 3765 5515
rect 3765 5485 3795 5515
rect 3795 5485 3796 5515
rect 3764 5484 3796 5485
rect 3764 5435 3796 5436
rect 3764 5405 3765 5435
rect 3765 5405 3795 5435
rect 3795 5405 3796 5435
rect 3764 5404 3796 5405
rect 3764 5324 3796 5356
rect 3764 5275 3796 5276
rect 3764 5245 3765 5275
rect 3765 5245 3795 5275
rect 3795 5245 3796 5275
rect 3764 5244 3796 5245
rect 3764 5195 3796 5196
rect 3764 5165 3765 5195
rect 3765 5165 3795 5195
rect 3795 5165 3796 5195
rect 3764 5164 3796 5165
rect 3764 5115 3796 5116
rect 3764 5085 3765 5115
rect 3765 5085 3795 5115
rect 3795 5085 3796 5115
rect 3764 5084 3796 5085
rect 3764 5035 3796 5036
rect 3764 5005 3765 5035
rect 3765 5005 3795 5035
rect 3795 5005 3796 5035
rect 3764 5004 3796 5005
rect 3764 4924 3796 4956
rect 3764 4875 3796 4876
rect 3764 4845 3765 4875
rect 3765 4845 3795 4875
rect 3795 4845 3796 4875
rect 3764 4844 3796 4845
rect 3764 4764 3796 4796
rect 3764 4715 3796 4716
rect 3764 4685 3765 4715
rect 3765 4685 3795 4715
rect 3795 4685 3796 4715
rect 3764 4684 3796 4685
rect 3764 4635 3796 4636
rect 3764 4605 3765 4635
rect 3765 4605 3795 4635
rect 3795 4605 3796 4635
rect 3764 4604 3796 4605
rect 3764 4524 3796 4556
rect 3764 4475 3796 4476
rect 3764 4445 3765 4475
rect 3765 4445 3795 4475
rect 3795 4445 3796 4475
rect 3764 4444 3796 4445
rect 3844 5515 3876 5516
rect 3844 5485 3845 5515
rect 3845 5485 3875 5515
rect 3875 5485 3876 5515
rect 3844 5484 3876 5485
rect 3844 5435 3876 5436
rect 3844 5405 3845 5435
rect 3845 5405 3875 5435
rect 3875 5405 3876 5435
rect 3844 5404 3876 5405
rect 3844 5324 3876 5356
rect 3844 5275 3876 5276
rect 3844 5245 3845 5275
rect 3845 5245 3875 5275
rect 3875 5245 3876 5275
rect 3844 5244 3876 5245
rect 3844 5195 3876 5196
rect 3844 5165 3845 5195
rect 3845 5165 3875 5195
rect 3875 5165 3876 5195
rect 3844 5164 3876 5165
rect 3844 5115 3876 5116
rect 3844 5085 3845 5115
rect 3845 5085 3875 5115
rect 3875 5085 3876 5115
rect 3844 5084 3876 5085
rect 3844 5035 3876 5036
rect 3844 5005 3845 5035
rect 3845 5005 3875 5035
rect 3875 5005 3876 5035
rect 3844 5004 3876 5005
rect 3844 4924 3876 4956
rect 3844 4875 3876 4876
rect 3844 4845 3845 4875
rect 3845 4845 3875 4875
rect 3875 4845 3876 4875
rect 3844 4844 3876 4845
rect 3844 4764 3876 4796
rect 3844 4715 3876 4716
rect 3844 4685 3845 4715
rect 3845 4685 3875 4715
rect 3875 4685 3876 4715
rect 3844 4684 3876 4685
rect 3844 4635 3876 4636
rect 3844 4605 3845 4635
rect 3845 4605 3875 4635
rect 3875 4605 3876 4635
rect 3844 4604 3876 4605
rect 3844 4524 3876 4556
rect 3844 4475 3876 4476
rect 3844 4445 3845 4475
rect 3845 4445 3875 4475
rect 3875 4445 3876 4475
rect 3844 4444 3876 4445
rect 3924 5515 3956 5516
rect 3924 5485 3925 5515
rect 3925 5485 3955 5515
rect 3955 5485 3956 5515
rect 3924 5484 3956 5485
rect 3924 5435 3956 5436
rect 3924 5405 3925 5435
rect 3925 5405 3955 5435
rect 3955 5405 3956 5435
rect 3924 5404 3956 5405
rect 3924 5324 3956 5356
rect 3924 5275 3956 5276
rect 3924 5245 3925 5275
rect 3925 5245 3955 5275
rect 3955 5245 3956 5275
rect 3924 5244 3956 5245
rect 3924 5195 3956 5196
rect 3924 5165 3925 5195
rect 3925 5165 3955 5195
rect 3955 5165 3956 5195
rect 3924 5164 3956 5165
rect 3924 5115 3956 5116
rect 3924 5085 3925 5115
rect 3925 5085 3955 5115
rect 3955 5085 3956 5115
rect 3924 5084 3956 5085
rect 3924 5035 3956 5036
rect 3924 5005 3925 5035
rect 3925 5005 3955 5035
rect 3955 5005 3956 5035
rect 3924 5004 3956 5005
rect 3924 4924 3956 4956
rect 3924 4875 3956 4876
rect 3924 4845 3925 4875
rect 3925 4845 3955 4875
rect 3955 4845 3956 4875
rect 3924 4844 3956 4845
rect 3924 4764 3956 4796
rect 3924 4715 3956 4716
rect 3924 4685 3925 4715
rect 3925 4685 3955 4715
rect 3955 4685 3956 4715
rect 3924 4684 3956 4685
rect 3924 4635 3956 4636
rect 3924 4605 3925 4635
rect 3925 4605 3955 4635
rect 3955 4605 3956 4635
rect 3924 4604 3956 4605
rect 3924 4524 3956 4556
rect 3924 4475 3956 4476
rect 3924 4445 3925 4475
rect 3925 4445 3955 4475
rect 3955 4445 3956 4475
rect 3924 4444 3956 4445
rect 4004 5515 4036 5516
rect 4004 5485 4005 5515
rect 4005 5485 4035 5515
rect 4035 5485 4036 5515
rect 4004 5484 4036 5485
rect 4004 5435 4036 5436
rect 4004 5405 4005 5435
rect 4005 5405 4035 5435
rect 4035 5405 4036 5435
rect 4004 5404 4036 5405
rect 4004 5324 4036 5356
rect 4004 5275 4036 5276
rect 4004 5245 4005 5275
rect 4005 5245 4035 5275
rect 4035 5245 4036 5275
rect 4004 5244 4036 5245
rect 4004 5195 4036 5196
rect 4004 5165 4005 5195
rect 4005 5165 4035 5195
rect 4035 5165 4036 5195
rect 4004 5164 4036 5165
rect 4004 5115 4036 5116
rect 4004 5085 4005 5115
rect 4005 5085 4035 5115
rect 4035 5085 4036 5115
rect 4004 5084 4036 5085
rect 4004 5035 4036 5036
rect 4004 5005 4005 5035
rect 4005 5005 4035 5035
rect 4035 5005 4036 5035
rect 4004 5004 4036 5005
rect 4004 4924 4036 4956
rect 4004 4875 4036 4876
rect 4004 4845 4005 4875
rect 4005 4845 4035 4875
rect 4035 4845 4036 4875
rect 4004 4844 4036 4845
rect 4004 4764 4036 4796
rect 4004 4715 4036 4716
rect 4004 4685 4005 4715
rect 4005 4685 4035 4715
rect 4035 4685 4036 4715
rect 4004 4684 4036 4685
rect 4004 4635 4036 4636
rect 4004 4605 4005 4635
rect 4005 4605 4035 4635
rect 4035 4605 4036 4635
rect 4004 4604 4036 4605
rect 4004 4524 4036 4556
rect 4004 4475 4036 4476
rect 4004 4445 4005 4475
rect 4005 4445 4035 4475
rect 4035 4445 4036 4475
rect 4004 4444 4036 4445
rect 4084 5515 4116 5516
rect 4084 5485 4085 5515
rect 4085 5485 4115 5515
rect 4115 5485 4116 5515
rect 4084 5484 4116 5485
rect 4084 5435 4116 5436
rect 4084 5405 4085 5435
rect 4085 5405 4115 5435
rect 4115 5405 4116 5435
rect 4084 5404 4116 5405
rect 4084 5324 4116 5356
rect 4084 5275 4116 5276
rect 4084 5245 4085 5275
rect 4085 5245 4115 5275
rect 4115 5245 4116 5275
rect 4084 5244 4116 5245
rect 4084 5195 4116 5196
rect 4084 5165 4085 5195
rect 4085 5165 4115 5195
rect 4115 5165 4116 5195
rect 4084 5164 4116 5165
rect 4084 5115 4116 5116
rect 4084 5085 4085 5115
rect 4085 5085 4115 5115
rect 4115 5085 4116 5115
rect 4084 5084 4116 5085
rect 4084 5035 4116 5036
rect 4084 5005 4085 5035
rect 4085 5005 4115 5035
rect 4115 5005 4116 5035
rect 4084 5004 4116 5005
rect 4084 4924 4116 4956
rect 4084 4875 4116 4876
rect 4084 4845 4085 4875
rect 4085 4845 4115 4875
rect 4115 4845 4116 4875
rect 4084 4844 4116 4845
rect 4084 4764 4116 4796
rect 4084 4715 4116 4716
rect 4084 4685 4085 4715
rect 4085 4685 4115 4715
rect 4115 4685 4116 4715
rect 4084 4684 4116 4685
rect 4084 4635 4116 4636
rect 4084 4605 4085 4635
rect 4085 4605 4115 4635
rect 4115 4605 4116 4635
rect 4084 4604 4116 4605
rect 4084 4524 4116 4556
rect 4084 4475 4116 4476
rect 4084 4445 4085 4475
rect 4085 4445 4115 4475
rect 4115 4445 4116 4475
rect 4084 4444 4116 4445
rect 4164 5515 4196 5516
rect 4164 5485 4165 5515
rect 4165 5485 4195 5515
rect 4195 5485 4196 5515
rect 4164 5484 4196 5485
rect 4164 5435 4196 5436
rect 4164 5405 4165 5435
rect 4165 5405 4195 5435
rect 4195 5405 4196 5435
rect 4164 5404 4196 5405
rect 4164 5324 4196 5356
rect 4164 5275 4196 5276
rect 4164 5245 4165 5275
rect 4165 5245 4195 5275
rect 4195 5245 4196 5275
rect 4164 5244 4196 5245
rect 4164 5195 4196 5196
rect 4164 5165 4165 5195
rect 4165 5165 4195 5195
rect 4195 5165 4196 5195
rect 4164 5164 4196 5165
rect 4164 5115 4196 5116
rect 4164 5085 4165 5115
rect 4165 5085 4195 5115
rect 4195 5085 4196 5115
rect 4164 5084 4196 5085
rect 4164 5035 4196 5036
rect 4164 5005 4165 5035
rect 4165 5005 4195 5035
rect 4195 5005 4196 5035
rect 4164 5004 4196 5005
rect 4164 4924 4196 4956
rect 4164 4875 4196 4876
rect 4164 4845 4165 4875
rect 4165 4845 4195 4875
rect 4195 4845 4196 4875
rect 4164 4844 4196 4845
rect 4164 4764 4196 4796
rect 4164 4715 4196 4716
rect 4164 4685 4165 4715
rect 4165 4685 4195 4715
rect 4195 4685 4196 4715
rect 4164 4684 4196 4685
rect 4164 4635 4196 4636
rect 4164 4605 4165 4635
rect 4165 4605 4195 4635
rect 4195 4605 4196 4635
rect 4164 4604 4196 4605
rect 4164 4524 4196 4556
rect 4164 4475 4196 4476
rect 4164 4445 4165 4475
rect 4165 4445 4195 4475
rect 4195 4445 4196 4475
rect 4164 4444 4196 4445
rect 4244 5515 4276 5516
rect 4244 5485 4245 5515
rect 4245 5485 4275 5515
rect 4275 5485 4276 5515
rect 4244 5484 4276 5485
rect 4244 5435 4276 5436
rect 4244 5405 4245 5435
rect 4245 5405 4275 5435
rect 4275 5405 4276 5435
rect 4244 5404 4276 5405
rect 4244 5324 4276 5356
rect 4244 5275 4276 5276
rect 4244 5245 4245 5275
rect 4245 5245 4275 5275
rect 4275 5245 4276 5275
rect 4244 5244 4276 5245
rect 4244 5195 4276 5196
rect 4244 5165 4245 5195
rect 4245 5165 4275 5195
rect 4275 5165 4276 5195
rect 4244 5164 4276 5165
rect 4244 5115 4276 5116
rect 4244 5085 4245 5115
rect 4245 5085 4275 5115
rect 4275 5085 4276 5115
rect 4244 5084 4276 5085
rect 4244 5035 4276 5036
rect 4244 5005 4245 5035
rect 4245 5005 4275 5035
rect 4275 5005 4276 5035
rect 4244 5004 4276 5005
rect 4244 4924 4276 4956
rect 4244 4875 4276 4876
rect 4244 4845 4245 4875
rect 4245 4845 4275 4875
rect 4275 4845 4276 4875
rect 4244 4844 4276 4845
rect 4244 4764 4276 4796
rect 4244 4715 4276 4716
rect 4244 4685 4245 4715
rect 4245 4685 4275 4715
rect 4275 4685 4276 4715
rect 4244 4684 4276 4685
rect 4244 4635 4276 4636
rect 4244 4605 4245 4635
rect 4245 4605 4275 4635
rect 4275 4605 4276 4635
rect 4244 4604 4276 4605
rect 4244 4524 4276 4556
rect 4244 4475 4276 4476
rect 4244 4445 4245 4475
rect 4245 4445 4275 4475
rect 4275 4445 4276 4475
rect 4244 4444 4276 4445
rect 4324 5515 4356 5516
rect 4324 5485 4325 5515
rect 4325 5485 4355 5515
rect 4355 5485 4356 5515
rect 4324 5484 4356 5485
rect 4324 5435 4356 5436
rect 4324 5405 4325 5435
rect 4325 5405 4355 5435
rect 4355 5405 4356 5435
rect 4324 5404 4356 5405
rect 4324 5324 4356 5356
rect 4324 5275 4356 5276
rect 4324 5245 4325 5275
rect 4325 5245 4355 5275
rect 4355 5245 4356 5275
rect 4324 5244 4356 5245
rect 4324 5195 4356 5196
rect 4324 5165 4325 5195
rect 4325 5165 4355 5195
rect 4355 5165 4356 5195
rect 4324 5164 4356 5165
rect 4324 5115 4356 5116
rect 4324 5085 4325 5115
rect 4325 5085 4355 5115
rect 4355 5085 4356 5115
rect 4324 5084 4356 5085
rect 4324 5035 4356 5036
rect 4324 5005 4325 5035
rect 4325 5005 4355 5035
rect 4355 5005 4356 5035
rect 4324 5004 4356 5005
rect 4324 4924 4356 4956
rect 4324 4875 4356 4876
rect 4324 4845 4325 4875
rect 4325 4845 4355 4875
rect 4355 4845 4356 4875
rect 4324 4844 4356 4845
rect 4324 4764 4356 4796
rect 4324 4715 4356 4716
rect 4324 4685 4325 4715
rect 4325 4685 4355 4715
rect 4355 4685 4356 4715
rect 4324 4684 4356 4685
rect 4324 4635 4356 4636
rect 4324 4605 4325 4635
rect 4325 4605 4355 4635
rect 4355 4605 4356 4635
rect 4324 4604 4356 4605
rect 4324 4524 4356 4556
rect 4324 4475 4356 4476
rect 4324 4445 4325 4475
rect 4325 4445 4355 4475
rect 4355 4445 4356 4475
rect 4324 4444 4356 4445
rect 4404 5515 4436 5516
rect 4404 5485 4405 5515
rect 4405 5485 4435 5515
rect 4435 5485 4436 5515
rect 4404 5484 4436 5485
rect 4404 5435 4436 5436
rect 4404 5405 4405 5435
rect 4405 5405 4435 5435
rect 4435 5405 4436 5435
rect 4404 5404 4436 5405
rect 4404 5324 4436 5356
rect 4404 5275 4436 5276
rect 4404 5245 4405 5275
rect 4405 5245 4435 5275
rect 4435 5245 4436 5275
rect 4404 5244 4436 5245
rect 4404 5195 4436 5196
rect 4404 5165 4405 5195
rect 4405 5165 4435 5195
rect 4435 5165 4436 5195
rect 4404 5164 4436 5165
rect 4404 5115 4436 5116
rect 4404 5085 4405 5115
rect 4405 5085 4435 5115
rect 4435 5085 4436 5115
rect 4404 5084 4436 5085
rect 4404 5035 4436 5036
rect 4404 5005 4405 5035
rect 4405 5005 4435 5035
rect 4435 5005 4436 5035
rect 4404 5004 4436 5005
rect 4404 4924 4436 4956
rect 4404 4875 4436 4876
rect 4404 4845 4405 4875
rect 4405 4845 4435 4875
rect 4435 4845 4436 4875
rect 4404 4844 4436 4845
rect 4404 4764 4436 4796
rect 4404 4715 4436 4716
rect 4404 4685 4405 4715
rect 4405 4685 4435 4715
rect 4435 4685 4436 4715
rect 4404 4684 4436 4685
rect 4404 4635 4436 4636
rect 4404 4605 4405 4635
rect 4405 4605 4435 4635
rect 4435 4605 4436 4635
rect 4404 4604 4436 4605
rect 4404 4524 4436 4556
rect 4404 4475 4436 4476
rect 4404 4445 4405 4475
rect 4405 4445 4435 4475
rect 4435 4445 4436 4475
rect 4404 4444 4436 4445
rect 4484 5515 4516 5516
rect 4484 5485 4485 5515
rect 4485 5485 4515 5515
rect 4515 5485 4516 5515
rect 4484 5484 4516 5485
rect 4484 5435 4516 5436
rect 4484 5405 4485 5435
rect 4485 5405 4515 5435
rect 4515 5405 4516 5435
rect 4484 5404 4516 5405
rect 4484 5324 4516 5356
rect 4484 5275 4516 5276
rect 4484 5245 4485 5275
rect 4485 5245 4515 5275
rect 4515 5245 4516 5275
rect 4484 5244 4516 5245
rect 4484 5195 4516 5196
rect 4484 5165 4485 5195
rect 4485 5165 4515 5195
rect 4515 5165 4516 5195
rect 4484 5164 4516 5165
rect 4484 5115 4516 5116
rect 4484 5085 4485 5115
rect 4485 5085 4515 5115
rect 4515 5085 4516 5115
rect 4484 5084 4516 5085
rect 4484 5035 4516 5036
rect 4484 5005 4485 5035
rect 4485 5005 4515 5035
rect 4515 5005 4516 5035
rect 4484 5004 4516 5005
rect 4484 4924 4516 4956
rect 4484 4875 4516 4876
rect 4484 4845 4485 4875
rect 4485 4845 4515 4875
rect 4515 4845 4516 4875
rect 4484 4844 4516 4845
rect 4484 4764 4516 4796
rect 4484 4715 4516 4716
rect 4484 4685 4485 4715
rect 4485 4685 4515 4715
rect 4515 4685 4516 4715
rect 4484 4684 4516 4685
rect 4484 4635 4516 4636
rect 4484 4605 4485 4635
rect 4485 4605 4515 4635
rect 4515 4605 4516 4635
rect 4484 4604 4516 4605
rect 4484 4524 4516 4556
rect 4484 4475 4516 4476
rect 4484 4445 4485 4475
rect 4485 4445 4515 4475
rect 4515 4445 4516 4475
rect 4484 4444 4516 4445
rect 4564 5515 4596 5516
rect 4564 5485 4565 5515
rect 4565 5485 4595 5515
rect 4595 5485 4596 5515
rect 4564 5484 4596 5485
rect 4564 5435 4596 5436
rect 4564 5405 4565 5435
rect 4565 5405 4595 5435
rect 4595 5405 4596 5435
rect 4564 5404 4596 5405
rect 4564 5324 4596 5356
rect 4564 5275 4596 5276
rect 4564 5245 4565 5275
rect 4565 5245 4595 5275
rect 4595 5245 4596 5275
rect 4564 5244 4596 5245
rect 4564 5195 4596 5196
rect 4564 5165 4565 5195
rect 4565 5165 4595 5195
rect 4595 5165 4596 5195
rect 4564 5164 4596 5165
rect 4564 5115 4596 5116
rect 4564 5085 4565 5115
rect 4565 5085 4595 5115
rect 4595 5085 4596 5115
rect 4564 5084 4596 5085
rect 4564 5035 4596 5036
rect 4564 5005 4565 5035
rect 4565 5005 4595 5035
rect 4595 5005 4596 5035
rect 4564 5004 4596 5005
rect 4564 4924 4596 4956
rect 4564 4875 4596 4876
rect 4564 4845 4565 4875
rect 4565 4845 4595 4875
rect 4595 4845 4596 4875
rect 4564 4844 4596 4845
rect 4564 4764 4596 4796
rect 4564 4715 4596 4716
rect 4564 4685 4565 4715
rect 4565 4685 4595 4715
rect 4595 4685 4596 4715
rect 4564 4684 4596 4685
rect 4564 4635 4596 4636
rect 4564 4605 4565 4635
rect 4565 4605 4595 4635
rect 4595 4605 4596 4635
rect 4564 4604 4596 4605
rect 4564 4524 4596 4556
rect 4564 4475 4596 4476
rect 4564 4445 4565 4475
rect 4565 4445 4595 4475
rect 4595 4445 4596 4475
rect 4564 4444 4596 4445
rect 4644 5515 4676 5516
rect 4644 5485 4645 5515
rect 4645 5485 4675 5515
rect 4675 5485 4676 5515
rect 4644 5484 4676 5485
rect 4644 5435 4676 5436
rect 4644 5405 4645 5435
rect 4645 5405 4675 5435
rect 4675 5405 4676 5435
rect 4644 5404 4676 5405
rect 4644 5324 4676 5356
rect 4644 5275 4676 5276
rect 4644 5245 4645 5275
rect 4645 5245 4675 5275
rect 4675 5245 4676 5275
rect 4644 5244 4676 5245
rect 4644 5195 4676 5196
rect 4644 5165 4645 5195
rect 4645 5165 4675 5195
rect 4675 5165 4676 5195
rect 4644 5164 4676 5165
rect 4644 5115 4676 5116
rect 4644 5085 4645 5115
rect 4645 5085 4675 5115
rect 4675 5085 4676 5115
rect 4644 5084 4676 5085
rect 4644 5035 4676 5036
rect 4644 5005 4645 5035
rect 4645 5005 4675 5035
rect 4675 5005 4676 5035
rect 4644 5004 4676 5005
rect 4644 4924 4676 4956
rect 4644 4875 4676 4876
rect 4644 4845 4645 4875
rect 4645 4845 4675 4875
rect 4675 4845 4676 4875
rect 4644 4844 4676 4845
rect 4644 4764 4676 4796
rect 4644 4715 4676 4716
rect 4644 4685 4645 4715
rect 4645 4685 4675 4715
rect 4675 4685 4676 4715
rect 4644 4684 4676 4685
rect 4644 4635 4676 4636
rect 4644 4605 4645 4635
rect 4645 4605 4675 4635
rect 4675 4605 4676 4635
rect 4644 4604 4676 4605
rect 4644 4524 4676 4556
rect 4644 4475 4676 4476
rect 4644 4445 4645 4475
rect 4645 4445 4675 4475
rect 4675 4445 4676 4475
rect 4644 4444 4676 4445
rect 4724 5515 4756 5516
rect 4724 5485 4725 5515
rect 4725 5485 4755 5515
rect 4755 5485 4756 5515
rect 4724 5484 4756 5485
rect 4724 5435 4756 5436
rect 4724 5405 4725 5435
rect 4725 5405 4755 5435
rect 4755 5405 4756 5435
rect 4724 5404 4756 5405
rect 4724 5324 4756 5356
rect 4724 5275 4756 5276
rect 4724 5245 4725 5275
rect 4725 5245 4755 5275
rect 4755 5245 4756 5275
rect 4724 5244 4756 5245
rect 4724 5195 4756 5196
rect 4724 5165 4725 5195
rect 4725 5165 4755 5195
rect 4755 5165 4756 5195
rect 4724 5164 4756 5165
rect 4724 5115 4756 5116
rect 4724 5085 4725 5115
rect 4725 5085 4755 5115
rect 4755 5085 4756 5115
rect 4724 5084 4756 5085
rect 4724 5035 4756 5036
rect 4724 5005 4725 5035
rect 4725 5005 4755 5035
rect 4755 5005 4756 5035
rect 4724 5004 4756 5005
rect 4724 4924 4756 4956
rect 4724 4875 4756 4876
rect 4724 4845 4725 4875
rect 4725 4845 4755 4875
rect 4755 4845 4756 4875
rect 4724 4844 4756 4845
rect 4724 4764 4756 4796
rect 4724 4715 4756 4716
rect 4724 4685 4725 4715
rect 4725 4685 4755 4715
rect 4755 4685 4756 4715
rect 4724 4684 4756 4685
rect 4724 4635 4756 4636
rect 4724 4605 4725 4635
rect 4725 4605 4755 4635
rect 4755 4605 4756 4635
rect 4724 4604 4756 4605
rect 4724 4524 4756 4556
rect 4724 4475 4756 4476
rect 4724 4445 4725 4475
rect 4725 4445 4755 4475
rect 4755 4445 4756 4475
rect 4724 4444 4756 4445
rect 4804 5515 4836 5516
rect 4804 5485 4805 5515
rect 4805 5485 4835 5515
rect 4835 5485 4836 5515
rect 4804 5484 4836 5485
rect 4804 5435 4836 5436
rect 4804 5405 4805 5435
rect 4805 5405 4835 5435
rect 4835 5405 4836 5435
rect 4804 5404 4836 5405
rect 4804 5324 4836 5356
rect 4804 5275 4836 5276
rect 4804 5245 4805 5275
rect 4805 5245 4835 5275
rect 4835 5245 4836 5275
rect 4804 5244 4836 5245
rect 4804 5195 4836 5196
rect 4804 5165 4805 5195
rect 4805 5165 4835 5195
rect 4835 5165 4836 5195
rect 4804 5164 4836 5165
rect 4804 5115 4836 5116
rect 4804 5085 4805 5115
rect 4805 5085 4835 5115
rect 4835 5085 4836 5115
rect 4804 5084 4836 5085
rect 4804 5035 4836 5036
rect 4804 5005 4805 5035
rect 4805 5005 4835 5035
rect 4835 5005 4836 5035
rect 4804 5004 4836 5005
rect 4804 4924 4836 4956
rect 4804 4875 4836 4876
rect 4804 4845 4805 4875
rect 4805 4845 4835 4875
rect 4835 4845 4836 4875
rect 4804 4844 4836 4845
rect 4804 4764 4836 4796
rect 4804 4715 4836 4716
rect 4804 4685 4805 4715
rect 4805 4685 4835 4715
rect 4835 4685 4836 4715
rect 4804 4684 4836 4685
rect 4804 4635 4836 4636
rect 4804 4605 4805 4635
rect 4805 4605 4835 4635
rect 4835 4605 4836 4635
rect 4804 4604 4836 4605
rect 4804 4524 4836 4556
rect 4804 4475 4836 4476
rect 4804 4445 4805 4475
rect 4805 4445 4835 4475
rect 4835 4445 4836 4475
rect 4804 4444 4836 4445
rect 4884 5515 4916 5516
rect 4884 5485 4885 5515
rect 4885 5485 4915 5515
rect 4915 5485 4916 5515
rect 4884 5484 4916 5485
rect 4884 5435 4916 5436
rect 4884 5405 4885 5435
rect 4885 5405 4915 5435
rect 4915 5405 4916 5435
rect 4884 5404 4916 5405
rect 4884 5355 4916 5356
rect 4884 5325 4885 5355
rect 4885 5325 4915 5355
rect 4915 5325 4916 5355
rect 4884 5324 4916 5325
rect 4884 5275 4916 5276
rect 4884 5245 4885 5275
rect 4885 5245 4915 5275
rect 4915 5245 4916 5275
rect 4884 5244 4916 5245
rect 4884 5195 4916 5196
rect 4884 5165 4885 5195
rect 4885 5165 4915 5195
rect 4915 5165 4916 5195
rect 4884 5164 4916 5165
rect 4884 5115 4916 5116
rect 4884 5085 4885 5115
rect 4885 5085 4915 5115
rect 4915 5085 4916 5115
rect 4884 5084 4916 5085
rect 4884 5035 4916 5036
rect 4884 5005 4885 5035
rect 4885 5005 4915 5035
rect 4915 5005 4916 5035
rect 4884 5004 4916 5005
rect 4884 4955 4916 4956
rect 4884 4925 4885 4955
rect 4885 4925 4915 4955
rect 4915 4925 4916 4955
rect 4884 4924 4916 4925
rect 4884 4875 4916 4876
rect 4884 4845 4885 4875
rect 4885 4845 4915 4875
rect 4915 4845 4916 4875
rect 4884 4844 4916 4845
rect 4884 4795 4916 4796
rect 4884 4765 4885 4795
rect 4885 4765 4915 4795
rect 4915 4765 4916 4795
rect 4884 4764 4916 4765
rect 4884 4715 4916 4716
rect 4884 4685 4885 4715
rect 4885 4685 4915 4715
rect 4915 4685 4916 4715
rect 4884 4684 4916 4685
rect 4884 4635 4916 4636
rect 4884 4605 4885 4635
rect 4885 4605 4915 4635
rect 4915 4605 4916 4635
rect 4884 4604 4916 4605
rect 4884 4555 4916 4556
rect 4884 4525 4885 4555
rect 4885 4525 4915 4555
rect 4915 4525 4916 4555
rect 4884 4524 4916 4525
rect 4884 4475 4916 4476
rect 4884 4445 4885 4475
rect 4885 4445 4915 4475
rect 4915 4445 4916 4475
rect 4884 4444 4916 4445
rect -876 4395 -844 4396
rect -876 4365 -875 4395
rect -875 4365 -845 4395
rect -845 4365 -844 4395
rect -876 4364 -844 4365
rect -876 4315 -844 4316
rect -876 4285 -875 4315
rect -875 4285 -845 4315
rect -845 4285 -844 4315
rect -876 4284 -844 4285
rect -876 4235 -844 4236
rect -876 4205 -875 4235
rect -875 4205 -845 4235
rect -845 4205 -844 4235
rect -876 4204 -844 4205
rect -876 4155 -844 4156
rect -876 4125 -875 4155
rect -875 4125 -845 4155
rect -845 4125 -844 4155
rect -876 4124 -844 4125
rect -876 4075 -844 4076
rect -876 4045 -875 4075
rect -875 4045 -845 4075
rect -845 4045 -844 4075
rect -876 4044 -844 4045
rect -876 3995 -844 3996
rect -876 3965 -875 3995
rect -875 3965 -845 3995
rect -845 3965 -844 3995
rect -876 3964 -844 3965
rect -876 3915 -844 3916
rect -876 3885 -875 3915
rect -875 3885 -845 3915
rect -845 3885 -844 3915
rect -876 3884 -844 3885
rect -876 3835 -844 3836
rect -876 3805 -875 3835
rect -875 3805 -845 3835
rect -845 3805 -844 3835
rect -876 3804 -844 3805
rect -876 3755 -844 3756
rect -876 3725 -875 3755
rect -875 3725 -845 3755
rect -845 3725 -844 3755
rect -876 3724 -844 3725
rect -876 3675 -844 3676
rect -876 3645 -875 3675
rect -875 3645 -845 3675
rect -845 3645 -844 3675
rect -876 3644 -844 3645
rect -796 4395 -764 4396
rect -796 4365 -795 4395
rect -795 4365 -765 4395
rect -765 4365 -764 4395
rect -796 4364 -764 4365
rect -796 4284 -764 4316
rect -796 4235 -764 4236
rect -796 4205 -795 4235
rect -795 4205 -765 4235
rect -765 4205 -764 4235
rect -796 4204 -764 4205
rect -796 4124 -764 4156
rect -796 4075 -764 4076
rect -796 4045 -795 4075
rect -795 4045 -765 4075
rect -765 4045 -764 4075
rect -796 4044 -764 4045
rect -796 3995 -764 3996
rect -796 3965 -795 3995
rect -795 3965 -765 3995
rect -765 3965 -764 3995
rect -796 3964 -764 3965
rect -796 3915 -764 3916
rect -796 3885 -795 3915
rect -795 3885 -765 3915
rect -765 3885 -764 3915
rect -796 3884 -764 3885
rect -796 3835 -764 3836
rect -796 3805 -795 3835
rect -795 3805 -765 3835
rect -765 3805 -764 3835
rect -796 3804 -764 3805
rect -796 3755 -764 3756
rect -796 3725 -795 3755
rect -795 3725 -765 3755
rect -765 3725 -764 3755
rect -796 3724 -764 3725
rect -796 3675 -764 3676
rect -796 3645 -795 3675
rect -795 3645 -765 3675
rect -765 3645 -764 3675
rect -796 3644 -764 3645
rect -716 4395 -684 4396
rect -716 4365 -715 4395
rect -715 4365 -685 4395
rect -685 4365 -684 4395
rect -716 4364 -684 4365
rect -716 4284 -684 4316
rect -716 4235 -684 4236
rect -716 4205 -715 4235
rect -715 4205 -685 4235
rect -685 4205 -684 4235
rect -716 4204 -684 4205
rect -716 4124 -684 4156
rect -716 4075 -684 4076
rect -716 4045 -715 4075
rect -715 4045 -685 4075
rect -685 4045 -684 4075
rect -716 4044 -684 4045
rect -716 3995 -684 3996
rect -716 3965 -715 3995
rect -715 3965 -685 3995
rect -685 3965 -684 3995
rect -716 3964 -684 3965
rect -716 3915 -684 3916
rect -716 3885 -715 3915
rect -715 3885 -685 3915
rect -685 3885 -684 3915
rect -716 3884 -684 3885
rect -716 3835 -684 3836
rect -716 3805 -715 3835
rect -715 3805 -685 3835
rect -685 3805 -684 3835
rect -716 3804 -684 3805
rect -716 3755 -684 3756
rect -716 3725 -715 3755
rect -715 3725 -685 3755
rect -685 3725 -684 3755
rect -716 3724 -684 3725
rect -716 3675 -684 3676
rect -716 3645 -715 3675
rect -715 3645 -685 3675
rect -685 3645 -684 3675
rect -716 3644 -684 3645
rect -636 4395 -604 4396
rect -636 4365 -635 4395
rect -635 4365 -605 4395
rect -605 4365 -604 4395
rect -636 4364 -604 4365
rect -636 4284 -604 4316
rect -636 4235 -604 4236
rect -636 4205 -635 4235
rect -635 4205 -605 4235
rect -605 4205 -604 4235
rect -636 4204 -604 4205
rect -636 4124 -604 4156
rect -636 4075 -604 4076
rect -636 4045 -635 4075
rect -635 4045 -605 4075
rect -605 4045 -604 4075
rect -636 4044 -604 4045
rect -636 3995 -604 3996
rect -636 3965 -635 3995
rect -635 3965 -605 3995
rect -605 3965 -604 3995
rect -636 3964 -604 3965
rect -636 3915 -604 3916
rect -636 3885 -635 3915
rect -635 3885 -605 3915
rect -605 3885 -604 3915
rect -636 3884 -604 3885
rect -636 3835 -604 3836
rect -636 3805 -635 3835
rect -635 3805 -605 3835
rect -605 3805 -604 3835
rect -636 3804 -604 3805
rect -636 3755 -604 3756
rect -636 3725 -635 3755
rect -635 3725 -605 3755
rect -605 3725 -604 3755
rect -636 3724 -604 3725
rect -636 3675 -604 3676
rect -636 3645 -635 3675
rect -635 3645 -605 3675
rect -605 3645 -604 3675
rect -636 3644 -604 3645
rect -556 4395 -524 4396
rect -556 4365 -555 4395
rect -555 4365 -525 4395
rect -525 4365 -524 4395
rect -556 4364 -524 4365
rect -556 4284 -524 4316
rect -556 4235 -524 4236
rect -556 4205 -555 4235
rect -555 4205 -525 4235
rect -525 4205 -524 4235
rect -556 4204 -524 4205
rect -556 4124 -524 4156
rect -556 4075 -524 4076
rect -556 4045 -555 4075
rect -555 4045 -525 4075
rect -525 4045 -524 4075
rect -556 4044 -524 4045
rect -556 3995 -524 3996
rect -556 3965 -555 3995
rect -555 3965 -525 3995
rect -525 3965 -524 3995
rect -556 3964 -524 3965
rect -556 3915 -524 3916
rect -556 3885 -555 3915
rect -555 3885 -525 3915
rect -525 3885 -524 3915
rect -556 3884 -524 3885
rect -556 3835 -524 3836
rect -556 3805 -555 3835
rect -555 3805 -525 3835
rect -525 3805 -524 3835
rect -556 3804 -524 3805
rect -556 3755 -524 3756
rect -556 3725 -555 3755
rect -555 3725 -525 3755
rect -525 3725 -524 3755
rect -556 3724 -524 3725
rect -556 3675 -524 3676
rect -556 3645 -555 3675
rect -555 3645 -525 3675
rect -525 3645 -524 3675
rect -556 3644 -524 3645
rect -476 4395 -444 4396
rect -476 4365 -475 4395
rect -475 4365 -445 4395
rect -445 4365 -444 4395
rect -476 4364 -444 4365
rect -476 4284 -444 4316
rect -476 4235 -444 4236
rect -476 4205 -475 4235
rect -475 4205 -445 4235
rect -445 4205 -444 4235
rect -476 4204 -444 4205
rect -476 4124 -444 4156
rect -476 4075 -444 4076
rect -476 4045 -475 4075
rect -475 4045 -445 4075
rect -445 4045 -444 4075
rect -476 4044 -444 4045
rect -476 3995 -444 3996
rect -476 3965 -475 3995
rect -475 3965 -445 3995
rect -445 3965 -444 3995
rect -476 3964 -444 3965
rect -476 3915 -444 3916
rect -476 3885 -475 3915
rect -475 3885 -445 3915
rect -445 3885 -444 3915
rect -476 3884 -444 3885
rect -476 3835 -444 3836
rect -476 3805 -475 3835
rect -475 3805 -445 3835
rect -445 3805 -444 3835
rect -476 3804 -444 3805
rect -476 3755 -444 3756
rect -476 3725 -475 3755
rect -475 3725 -445 3755
rect -445 3725 -444 3755
rect -476 3724 -444 3725
rect -476 3675 -444 3676
rect -476 3645 -475 3675
rect -475 3645 -445 3675
rect -445 3645 -444 3675
rect -476 3644 -444 3645
rect -396 4395 -364 4396
rect -396 4365 -395 4395
rect -395 4365 -365 4395
rect -365 4365 -364 4395
rect -396 4364 -364 4365
rect -396 4284 -364 4316
rect -396 4235 -364 4236
rect -396 4205 -395 4235
rect -395 4205 -365 4235
rect -365 4205 -364 4235
rect -396 4204 -364 4205
rect -396 4124 -364 4156
rect -396 4075 -364 4076
rect -396 4045 -395 4075
rect -395 4045 -365 4075
rect -365 4045 -364 4075
rect -396 4044 -364 4045
rect -396 3995 -364 3996
rect -396 3965 -395 3995
rect -395 3965 -365 3995
rect -365 3965 -364 3995
rect -396 3964 -364 3965
rect -396 3915 -364 3916
rect -396 3885 -395 3915
rect -395 3885 -365 3915
rect -365 3885 -364 3915
rect -396 3884 -364 3885
rect -396 3835 -364 3836
rect -396 3805 -395 3835
rect -395 3805 -365 3835
rect -365 3805 -364 3835
rect -396 3804 -364 3805
rect -396 3755 -364 3756
rect -396 3725 -395 3755
rect -395 3725 -365 3755
rect -365 3725 -364 3755
rect -396 3724 -364 3725
rect -396 3675 -364 3676
rect -396 3645 -395 3675
rect -395 3645 -365 3675
rect -365 3645 -364 3675
rect -396 3644 -364 3645
rect -316 4395 -284 4396
rect -316 4365 -315 4395
rect -315 4365 -285 4395
rect -285 4365 -284 4395
rect -316 4364 -284 4365
rect -316 4284 -284 4316
rect -316 4235 -284 4236
rect -316 4205 -315 4235
rect -315 4205 -285 4235
rect -285 4205 -284 4235
rect -316 4204 -284 4205
rect -316 4124 -284 4156
rect -316 4075 -284 4076
rect -316 4045 -315 4075
rect -315 4045 -285 4075
rect -285 4045 -284 4075
rect -316 4044 -284 4045
rect -316 3995 -284 3996
rect -316 3965 -315 3995
rect -315 3965 -285 3995
rect -285 3965 -284 3995
rect -316 3964 -284 3965
rect -316 3915 -284 3916
rect -316 3885 -315 3915
rect -315 3885 -285 3915
rect -285 3885 -284 3915
rect -316 3884 -284 3885
rect -316 3835 -284 3836
rect -316 3805 -315 3835
rect -315 3805 -285 3835
rect -285 3805 -284 3835
rect -316 3804 -284 3805
rect -316 3755 -284 3756
rect -316 3725 -315 3755
rect -315 3725 -285 3755
rect -285 3725 -284 3755
rect -316 3724 -284 3725
rect -316 3675 -284 3676
rect -316 3645 -315 3675
rect -315 3645 -285 3675
rect -285 3645 -284 3675
rect -316 3644 -284 3645
rect -236 4395 -204 4396
rect -236 4365 -235 4395
rect -235 4365 -205 4395
rect -205 4365 -204 4395
rect -236 4364 -204 4365
rect -236 4284 -204 4316
rect -236 4235 -204 4236
rect -236 4205 -235 4235
rect -235 4205 -205 4235
rect -205 4205 -204 4235
rect -236 4204 -204 4205
rect -236 4124 -204 4156
rect -236 4075 -204 4076
rect -236 4045 -235 4075
rect -235 4045 -205 4075
rect -205 4045 -204 4075
rect -236 4044 -204 4045
rect -236 3995 -204 3996
rect -236 3965 -235 3995
rect -235 3965 -205 3995
rect -205 3965 -204 3995
rect -236 3964 -204 3965
rect -236 3915 -204 3916
rect -236 3885 -235 3915
rect -235 3885 -205 3915
rect -205 3885 -204 3915
rect -236 3884 -204 3885
rect -236 3835 -204 3836
rect -236 3805 -235 3835
rect -235 3805 -205 3835
rect -205 3805 -204 3835
rect -236 3804 -204 3805
rect -236 3755 -204 3756
rect -236 3725 -235 3755
rect -235 3725 -205 3755
rect -205 3725 -204 3755
rect -236 3724 -204 3725
rect -236 3675 -204 3676
rect -236 3645 -235 3675
rect -235 3645 -205 3675
rect -205 3645 -204 3675
rect -236 3644 -204 3645
rect -156 4395 -124 4396
rect -156 4365 -155 4395
rect -155 4365 -125 4395
rect -125 4365 -124 4395
rect -156 4364 -124 4365
rect -156 4284 -124 4316
rect -156 4235 -124 4236
rect -156 4205 -155 4235
rect -155 4205 -125 4235
rect -125 4205 -124 4235
rect -156 4204 -124 4205
rect -156 4124 -124 4156
rect -156 4075 -124 4076
rect -156 4045 -155 4075
rect -155 4045 -125 4075
rect -125 4045 -124 4075
rect -156 4044 -124 4045
rect -156 3995 -124 3996
rect -156 3965 -155 3995
rect -155 3965 -125 3995
rect -125 3965 -124 3995
rect -156 3964 -124 3965
rect -156 3915 -124 3916
rect -156 3885 -155 3915
rect -155 3885 -125 3915
rect -125 3885 -124 3915
rect -156 3884 -124 3885
rect -156 3835 -124 3836
rect -156 3805 -155 3835
rect -155 3805 -125 3835
rect -125 3805 -124 3835
rect -156 3804 -124 3805
rect -156 3755 -124 3756
rect -156 3725 -155 3755
rect -155 3725 -125 3755
rect -125 3725 -124 3755
rect -156 3724 -124 3725
rect -156 3675 -124 3676
rect -156 3645 -155 3675
rect -155 3645 -125 3675
rect -125 3645 -124 3675
rect -156 3644 -124 3645
rect -76 4395 -44 4396
rect -76 4365 -75 4395
rect -75 4365 -45 4395
rect -45 4365 -44 4395
rect -76 4364 -44 4365
rect -76 4284 -44 4316
rect -76 4235 -44 4236
rect -76 4205 -75 4235
rect -75 4205 -45 4235
rect -45 4205 -44 4235
rect -76 4204 -44 4205
rect -76 4124 -44 4156
rect -76 4075 -44 4076
rect -76 4045 -75 4075
rect -75 4045 -45 4075
rect -45 4045 -44 4075
rect -76 4044 -44 4045
rect -76 3995 -44 3996
rect -76 3965 -75 3995
rect -75 3965 -45 3995
rect -45 3965 -44 3995
rect -76 3964 -44 3965
rect -76 3915 -44 3916
rect -76 3885 -75 3915
rect -75 3885 -45 3915
rect -45 3885 -44 3915
rect -76 3884 -44 3885
rect -76 3835 -44 3836
rect -76 3805 -75 3835
rect -75 3805 -45 3835
rect -45 3805 -44 3835
rect -76 3804 -44 3805
rect -76 3755 -44 3756
rect -76 3725 -75 3755
rect -75 3725 -45 3755
rect -45 3725 -44 3755
rect -76 3724 -44 3725
rect -76 3675 -44 3676
rect -76 3645 -75 3675
rect -75 3645 -45 3675
rect -45 3645 -44 3675
rect -76 3644 -44 3645
rect 4 4395 36 4396
rect 4 4365 5 4395
rect 5 4365 35 4395
rect 35 4365 36 4395
rect 4 4364 36 4365
rect 4 4284 36 4316
rect 4 4235 36 4236
rect 4 4205 5 4235
rect 5 4205 35 4235
rect 35 4205 36 4235
rect 4 4204 36 4205
rect 4 4124 36 4156
rect 4 4075 36 4076
rect 4 4045 5 4075
rect 5 4045 35 4075
rect 35 4045 36 4075
rect 4 4044 36 4045
rect 4 3995 36 3996
rect 4 3965 5 3995
rect 5 3965 35 3995
rect 35 3965 36 3995
rect 4 3964 36 3965
rect 4 3915 36 3916
rect 4 3885 5 3915
rect 5 3885 35 3915
rect 35 3885 36 3915
rect 4 3884 36 3885
rect 4 3835 36 3836
rect 4 3805 5 3835
rect 5 3805 35 3835
rect 35 3805 36 3835
rect 4 3804 36 3805
rect 4 3755 36 3756
rect 4 3725 5 3755
rect 5 3725 35 3755
rect 35 3725 36 3755
rect 4 3724 36 3725
rect 4 3675 36 3676
rect 4 3645 5 3675
rect 5 3645 35 3675
rect 35 3645 36 3675
rect 4 3644 36 3645
rect 84 4395 116 4396
rect 84 4365 85 4395
rect 85 4365 115 4395
rect 115 4365 116 4395
rect 84 4364 116 4365
rect 84 4284 116 4316
rect 84 4235 116 4236
rect 84 4205 85 4235
rect 85 4205 115 4235
rect 115 4205 116 4235
rect 84 4204 116 4205
rect 84 4124 116 4156
rect 84 4075 116 4076
rect 84 4045 85 4075
rect 85 4045 115 4075
rect 115 4045 116 4075
rect 84 4044 116 4045
rect 84 3995 116 3996
rect 84 3965 85 3995
rect 85 3965 115 3995
rect 115 3965 116 3995
rect 84 3964 116 3965
rect 84 3915 116 3916
rect 84 3885 85 3915
rect 85 3885 115 3915
rect 115 3885 116 3915
rect 84 3884 116 3885
rect 84 3835 116 3836
rect 84 3805 85 3835
rect 85 3805 115 3835
rect 115 3805 116 3835
rect 84 3804 116 3805
rect 84 3755 116 3756
rect 84 3725 85 3755
rect 85 3725 115 3755
rect 115 3725 116 3755
rect 84 3724 116 3725
rect 84 3675 116 3676
rect 84 3645 85 3675
rect 85 3645 115 3675
rect 115 3645 116 3675
rect 84 3644 116 3645
rect 164 4395 196 4396
rect 164 4365 165 4395
rect 165 4365 195 4395
rect 195 4365 196 4395
rect 164 4364 196 4365
rect 164 4284 196 4316
rect 164 4235 196 4236
rect 164 4205 165 4235
rect 165 4205 195 4235
rect 195 4205 196 4235
rect 164 4204 196 4205
rect 164 4124 196 4156
rect 164 4075 196 4076
rect 164 4045 165 4075
rect 165 4045 195 4075
rect 195 4045 196 4075
rect 164 4044 196 4045
rect 164 3995 196 3996
rect 164 3965 165 3995
rect 165 3965 195 3995
rect 195 3965 196 3995
rect 164 3964 196 3965
rect 164 3915 196 3916
rect 164 3885 165 3915
rect 165 3885 195 3915
rect 195 3885 196 3915
rect 164 3884 196 3885
rect 164 3835 196 3836
rect 164 3805 165 3835
rect 165 3805 195 3835
rect 195 3805 196 3835
rect 164 3804 196 3805
rect 164 3755 196 3756
rect 164 3725 165 3755
rect 165 3725 195 3755
rect 195 3725 196 3755
rect 164 3724 196 3725
rect 164 3675 196 3676
rect 164 3645 165 3675
rect 165 3645 195 3675
rect 195 3645 196 3675
rect 164 3644 196 3645
rect 244 4395 276 4396
rect 244 4365 245 4395
rect 245 4365 275 4395
rect 275 4365 276 4395
rect 244 4364 276 4365
rect 244 4284 276 4316
rect 244 4235 276 4236
rect 244 4205 245 4235
rect 245 4205 275 4235
rect 275 4205 276 4235
rect 244 4204 276 4205
rect 244 4124 276 4156
rect 244 4075 276 4076
rect 244 4045 245 4075
rect 245 4045 275 4075
rect 275 4045 276 4075
rect 244 4044 276 4045
rect 244 3995 276 3996
rect 244 3965 245 3995
rect 245 3965 275 3995
rect 275 3965 276 3995
rect 244 3964 276 3965
rect 244 3915 276 3916
rect 244 3885 245 3915
rect 245 3885 275 3915
rect 275 3885 276 3915
rect 244 3884 276 3885
rect 244 3835 276 3836
rect 244 3805 245 3835
rect 245 3805 275 3835
rect 275 3805 276 3835
rect 244 3804 276 3805
rect 244 3755 276 3756
rect 244 3725 245 3755
rect 245 3725 275 3755
rect 275 3725 276 3755
rect 244 3724 276 3725
rect 244 3675 276 3676
rect 244 3645 245 3675
rect 245 3645 275 3675
rect 275 3645 276 3675
rect 244 3644 276 3645
rect 324 4395 356 4396
rect 324 4365 325 4395
rect 325 4365 355 4395
rect 355 4365 356 4395
rect 324 4364 356 4365
rect 324 4284 356 4316
rect 324 4235 356 4236
rect 324 4205 325 4235
rect 325 4205 355 4235
rect 355 4205 356 4235
rect 324 4204 356 4205
rect 324 4124 356 4156
rect 324 4075 356 4076
rect 324 4045 325 4075
rect 325 4045 355 4075
rect 355 4045 356 4075
rect 324 4044 356 4045
rect 324 3995 356 3996
rect 324 3965 325 3995
rect 325 3965 355 3995
rect 355 3965 356 3995
rect 324 3964 356 3965
rect 324 3915 356 3916
rect 324 3885 325 3915
rect 325 3885 355 3915
rect 355 3885 356 3915
rect 324 3884 356 3885
rect 324 3835 356 3836
rect 324 3805 325 3835
rect 325 3805 355 3835
rect 355 3805 356 3835
rect 324 3804 356 3805
rect 324 3755 356 3756
rect 324 3725 325 3755
rect 325 3725 355 3755
rect 355 3725 356 3755
rect 324 3724 356 3725
rect 324 3675 356 3676
rect 324 3645 325 3675
rect 325 3645 355 3675
rect 355 3645 356 3675
rect 324 3644 356 3645
rect 404 4395 436 4396
rect 404 4365 405 4395
rect 405 4365 435 4395
rect 435 4365 436 4395
rect 404 4364 436 4365
rect 404 4284 436 4316
rect 404 4235 436 4236
rect 404 4205 405 4235
rect 405 4205 435 4235
rect 435 4205 436 4235
rect 404 4204 436 4205
rect 404 4124 436 4156
rect 404 4075 436 4076
rect 404 4045 405 4075
rect 405 4045 435 4075
rect 435 4045 436 4075
rect 404 4044 436 4045
rect 404 3995 436 3996
rect 404 3965 405 3995
rect 405 3965 435 3995
rect 435 3965 436 3995
rect 404 3964 436 3965
rect 404 3915 436 3916
rect 404 3885 405 3915
rect 405 3885 435 3915
rect 435 3885 436 3915
rect 404 3884 436 3885
rect 404 3835 436 3836
rect 404 3805 405 3835
rect 405 3805 435 3835
rect 435 3805 436 3835
rect 404 3804 436 3805
rect 404 3755 436 3756
rect 404 3725 405 3755
rect 405 3725 435 3755
rect 435 3725 436 3755
rect 404 3724 436 3725
rect 404 3675 436 3676
rect 404 3645 405 3675
rect 405 3645 435 3675
rect 435 3645 436 3675
rect 404 3644 436 3645
rect 484 4395 516 4396
rect 484 4365 485 4395
rect 485 4365 515 4395
rect 515 4365 516 4395
rect 484 4364 516 4365
rect 484 4284 516 4316
rect 484 4235 516 4236
rect 484 4205 485 4235
rect 485 4205 515 4235
rect 515 4205 516 4235
rect 484 4204 516 4205
rect 484 4124 516 4156
rect 484 4075 516 4076
rect 484 4045 485 4075
rect 485 4045 515 4075
rect 515 4045 516 4075
rect 484 4044 516 4045
rect 484 3995 516 3996
rect 484 3965 485 3995
rect 485 3965 515 3995
rect 515 3965 516 3995
rect 484 3964 516 3965
rect 484 3915 516 3916
rect 484 3885 485 3915
rect 485 3885 515 3915
rect 515 3885 516 3915
rect 484 3884 516 3885
rect 484 3835 516 3836
rect 484 3805 485 3835
rect 485 3805 515 3835
rect 515 3805 516 3835
rect 484 3804 516 3805
rect 484 3755 516 3756
rect 484 3725 485 3755
rect 485 3725 515 3755
rect 515 3725 516 3755
rect 484 3724 516 3725
rect 484 3675 516 3676
rect 484 3645 485 3675
rect 485 3645 515 3675
rect 515 3645 516 3675
rect 484 3644 516 3645
rect 564 4395 596 4396
rect 564 4365 565 4395
rect 565 4365 595 4395
rect 595 4365 596 4395
rect 564 4364 596 4365
rect 564 4284 596 4316
rect 564 4235 596 4236
rect 564 4205 565 4235
rect 565 4205 595 4235
rect 595 4205 596 4235
rect 564 4204 596 4205
rect 564 4124 596 4156
rect 564 4075 596 4076
rect 564 4045 565 4075
rect 565 4045 595 4075
rect 595 4045 596 4075
rect 564 4044 596 4045
rect 564 3995 596 3996
rect 564 3965 565 3995
rect 565 3965 595 3995
rect 595 3965 596 3995
rect 564 3964 596 3965
rect 564 3915 596 3916
rect 564 3885 565 3915
rect 565 3885 595 3915
rect 595 3885 596 3915
rect 564 3884 596 3885
rect 564 3835 596 3836
rect 564 3805 565 3835
rect 565 3805 595 3835
rect 595 3805 596 3835
rect 564 3804 596 3805
rect 564 3755 596 3756
rect 564 3725 565 3755
rect 565 3725 595 3755
rect 595 3725 596 3755
rect 564 3724 596 3725
rect 564 3675 596 3676
rect 564 3645 565 3675
rect 565 3645 595 3675
rect 595 3645 596 3675
rect 564 3644 596 3645
rect 644 4395 676 4396
rect 644 4365 645 4395
rect 645 4365 675 4395
rect 675 4365 676 4395
rect 644 4364 676 4365
rect 644 4284 676 4316
rect 644 4235 676 4236
rect 644 4205 645 4235
rect 645 4205 675 4235
rect 675 4205 676 4235
rect 644 4204 676 4205
rect 644 4124 676 4156
rect 644 4075 676 4076
rect 644 4045 645 4075
rect 645 4045 675 4075
rect 675 4045 676 4075
rect 644 4044 676 4045
rect 644 3995 676 3996
rect 644 3965 645 3995
rect 645 3965 675 3995
rect 675 3965 676 3995
rect 644 3964 676 3965
rect 644 3915 676 3916
rect 644 3885 645 3915
rect 645 3885 675 3915
rect 675 3885 676 3915
rect 644 3884 676 3885
rect 644 3835 676 3836
rect 644 3805 645 3835
rect 645 3805 675 3835
rect 675 3805 676 3835
rect 644 3804 676 3805
rect 644 3755 676 3756
rect 644 3725 645 3755
rect 645 3725 675 3755
rect 675 3725 676 3755
rect 644 3724 676 3725
rect 644 3675 676 3676
rect 644 3645 645 3675
rect 645 3645 675 3675
rect 675 3645 676 3675
rect 644 3644 676 3645
rect 724 4395 756 4396
rect 724 4365 725 4395
rect 725 4365 755 4395
rect 755 4365 756 4395
rect 724 4364 756 4365
rect 724 4284 756 4316
rect 724 4235 756 4236
rect 724 4205 725 4235
rect 725 4205 755 4235
rect 755 4205 756 4235
rect 724 4204 756 4205
rect 724 4124 756 4156
rect 724 4075 756 4076
rect 724 4045 725 4075
rect 725 4045 755 4075
rect 755 4045 756 4075
rect 724 4044 756 4045
rect 724 3995 756 3996
rect 724 3965 725 3995
rect 725 3965 755 3995
rect 755 3965 756 3995
rect 724 3964 756 3965
rect 724 3915 756 3916
rect 724 3885 725 3915
rect 725 3885 755 3915
rect 755 3885 756 3915
rect 724 3884 756 3885
rect 724 3835 756 3836
rect 724 3805 725 3835
rect 725 3805 755 3835
rect 755 3805 756 3835
rect 724 3804 756 3805
rect 724 3755 756 3756
rect 724 3725 725 3755
rect 725 3725 755 3755
rect 755 3725 756 3755
rect 724 3724 756 3725
rect 724 3675 756 3676
rect 724 3645 725 3675
rect 725 3645 755 3675
rect 755 3645 756 3675
rect 724 3644 756 3645
rect 804 4395 836 4396
rect 804 4365 805 4395
rect 805 4365 835 4395
rect 835 4365 836 4395
rect 804 4364 836 4365
rect 804 4284 836 4316
rect 804 4235 836 4236
rect 804 4205 805 4235
rect 805 4205 835 4235
rect 835 4205 836 4235
rect 804 4204 836 4205
rect 804 4124 836 4156
rect 804 4075 836 4076
rect 804 4045 805 4075
rect 805 4045 835 4075
rect 835 4045 836 4075
rect 804 4044 836 4045
rect 804 3995 836 3996
rect 804 3965 805 3995
rect 805 3965 835 3995
rect 835 3965 836 3995
rect 804 3964 836 3965
rect 804 3915 836 3916
rect 804 3885 805 3915
rect 805 3885 835 3915
rect 835 3885 836 3915
rect 804 3884 836 3885
rect 804 3835 836 3836
rect 804 3805 805 3835
rect 805 3805 835 3835
rect 835 3805 836 3835
rect 804 3804 836 3805
rect 804 3755 836 3756
rect 804 3725 805 3755
rect 805 3725 835 3755
rect 835 3725 836 3755
rect 804 3724 836 3725
rect 804 3675 836 3676
rect 804 3645 805 3675
rect 805 3645 835 3675
rect 835 3645 836 3675
rect 804 3644 836 3645
rect 884 4395 916 4396
rect 884 4365 885 4395
rect 885 4365 915 4395
rect 915 4365 916 4395
rect 884 4364 916 4365
rect 884 4284 916 4316
rect 884 4235 916 4236
rect 884 4205 885 4235
rect 885 4205 915 4235
rect 915 4205 916 4235
rect 884 4204 916 4205
rect 884 4124 916 4156
rect 884 4075 916 4076
rect 884 4045 885 4075
rect 885 4045 915 4075
rect 915 4045 916 4075
rect 884 4044 916 4045
rect 884 3995 916 3996
rect 884 3965 885 3995
rect 885 3965 915 3995
rect 915 3965 916 3995
rect 884 3964 916 3965
rect 884 3915 916 3916
rect 884 3885 885 3915
rect 885 3885 915 3915
rect 915 3885 916 3915
rect 884 3884 916 3885
rect 884 3835 916 3836
rect 884 3805 885 3835
rect 885 3805 915 3835
rect 915 3805 916 3835
rect 884 3804 916 3805
rect 884 3755 916 3756
rect 884 3725 885 3755
rect 885 3725 915 3755
rect 915 3725 916 3755
rect 884 3724 916 3725
rect 884 3675 916 3676
rect 884 3645 885 3675
rect 885 3645 915 3675
rect 915 3645 916 3675
rect 884 3644 916 3645
rect 964 4395 996 4396
rect 964 4365 965 4395
rect 965 4365 995 4395
rect 995 4365 996 4395
rect 964 4364 996 4365
rect 964 4284 996 4316
rect 964 4235 996 4236
rect 964 4205 965 4235
rect 965 4205 995 4235
rect 995 4205 996 4235
rect 964 4204 996 4205
rect 964 4124 996 4156
rect 964 4075 996 4076
rect 964 4045 965 4075
rect 965 4045 995 4075
rect 995 4045 996 4075
rect 964 4044 996 4045
rect 964 3995 996 3996
rect 964 3965 965 3995
rect 965 3965 995 3995
rect 995 3965 996 3995
rect 964 3964 996 3965
rect 964 3915 996 3916
rect 964 3885 965 3915
rect 965 3885 995 3915
rect 995 3885 996 3915
rect 964 3884 996 3885
rect 964 3835 996 3836
rect 964 3805 965 3835
rect 965 3805 995 3835
rect 995 3805 996 3835
rect 964 3804 996 3805
rect 964 3755 996 3756
rect 964 3725 965 3755
rect 965 3725 995 3755
rect 995 3725 996 3755
rect 964 3724 996 3725
rect 964 3675 996 3676
rect 964 3645 965 3675
rect 965 3645 995 3675
rect 995 3645 996 3675
rect 964 3644 996 3645
rect 1044 4395 1076 4396
rect 1044 4365 1045 4395
rect 1045 4365 1075 4395
rect 1075 4365 1076 4395
rect 1044 4364 1076 4365
rect 1044 4284 1076 4316
rect 1044 4235 1076 4236
rect 1044 4205 1045 4235
rect 1045 4205 1075 4235
rect 1075 4205 1076 4235
rect 1044 4204 1076 4205
rect 1044 4124 1076 4156
rect 1044 4075 1076 4076
rect 1044 4045 1045 4075
rect 1045 4045 1075 4075
rect 1075 4045 1076 4075
rect 1044 4044 1076 4045
rect 1044 3995 1076 3996
rect 1044 3965 1045 3995
rect 1045 3965 1075 3995
rect 1075 3965 1076 3995
rect 1044 3964 1076 3965
rect 1044 3915 1076 3916
rect 1044 3885 1045 3915
rect 1045 3885 1075 3915
rect 1075 3885 1076 3915
rect 1044 3884 1076 3885
rect 1044 3835 1076 3836
rect 1044 3805 1045 3835
rect 1045 3805 1075 3835
rect 1075 3805 1076 3835
rect 1044 3804 1076 3805
rect 1044 3755 1076 3756
rect 1044 3725 1045 3755
rect 1045 3725 1075 3755
rect 1075 3725 1076 3755
rect 1044 3724 1076 3725
rect 1044 3675 1076 3676
rect 1044 3645 1045 3675
rect 1045 3645 1075 3675
rect 1075 3645 1076 3675
rect 1044 3644 1076 3645
rect 1124 4395 1156 4396
rect 1124 4365 1125 4395
rect 1125 4365 1155 4395
rect 1155 4365 1156 4395
rect 1124 4364 1156 4365
rect 1124 4284 1156 4316
rect 1124 4235 1156 4236
rect 1124 4205 1125 4235
rect 1125 4205 1155 4235
rect 1155 4205 1156 4235
rect 1124 4204 1156 4205
rect 1124 4124 1156 4156
rect 1124 4075 1156 4076
rect 1124 4045 1125 4075
rect 1125 4045 1155 4075
rect 1155 4045 1156 4075
rect 1124 4044 1156 4045
rect 1124 3995 1156 3996
rect 1124 3965 1125 3995
rect 1125 3965 1155 3995
rect 1155 3965 1156 3995
rect 1124 3964 1156 3965
rect 1124 3915 1156 3916
rect 1124 3885 1125 3915
rect 1125 3885 1155 3915
rect 1155 3885 1156 3915
rect 1124 3884 1156 3885
rect 1124 3835 1156 3836
rect 1124 3805 1125 3835
rect 1125 3805 1155 3835
rect 1155 3805 1156 3835
rect 1124 3804 1156 3805
rect 1124 3755 1156 3756
rect 1124 3725 1125 3755
rect 1125 3725 1155 3755
rect 1155 3725 1156 3755
rect 1124 3724 1156 3725
rect 1124 3675 1156 3676
rect 1124 3645 1125 3675
rect 1125 3645 1155 3675
rect 1155 3645 1156 3675
rect 1124 3644 1156 3645
rect 1204 4395 1236 4396
rect 1204 4365 1205 4395
rect 1205 4365 1235 4395
rect 1235 4365 1236 4395
rect 1204 4364 1236 4365
rect 1204 4284 1236 4316
rect 1204 4235 1236 4236
rect 1204 4205 1205 4235
rect 1205 4205 1235 4235
rect 1235 4205 1236 4235
rect 1204 4204 1236 4205
rect 1204 4124 1236 4156
rect 1204 4075 1236 4076
rect 1204 4045 1205 4075
rect 1205 4045 1235 4075
rect 1235 4045 1236 4075
rect 1204 4044 1236 4045
rect 1204 3995 1236 3996
rect 1204 3965 1205 3995
rect 1205 3965 1235 3995
rect 1235 3965 1236 3995
rect 1204 3964 1236 3965
rect 1204 3915 1236 3916
rect 1204 3885 1205 3915
rect 1205 3885 1235 3915
rect 1235 3885 1236 3915
rect 1204 3884 1236 3885
rect 1204 3835 1236 3836
rect 1204 3805 1205 3835
rect 1205 3805 1235 3835
rect 1235 3805 1236 3835
rect 1204 3804 1236 3805
rect 1204 3755 1236 3756
rect 1204 3725 1205 3755
rect 1205 3725 1235 3755
rect 1235 3725 1236 3755
rect 1204 3724 1236 3725
rect 1204 3675 1236 3676
rect 1204 3645 1205 3675
rect 1205 3645 1235 3675
rect 1235 3645 1236 3675
rect 1204 3644 1236 3645
rect 1284 4395 1316 4396
rect 1284 4365 1285 4395
rect 1285 4365 1315 4395
rect 1315 4365 1316 4395
rect 1284 4364 1316 4365
rect 1284 4284 1316 4316
rect 1284 4235 1316 4236
rect 1284 4205 1285 4235
rect 1285 4205 1315 4235
rect 1315 4205 1316 4235
rect 1284 4204 1316 4205
rect 1284 4124 1316 4156
rect 1284 4075 1316 4076
rect 1284 4045 1285 4075
rect 1285 4045 1315 4075
rect 1315 4045 1316 4075
rect 1284 4044 1316 4045
rect 1284 3995 1316 3996
rect 1284 3965 1285 3995
rect 1285 3965 1315 3995
rect 1315 3965 1316 3995
rect 1284 3964 1316 3965
rect 1284 3915 1316 3916
rect 1284 3885 1285 3915
rect 1285 3885 1315 3915
rect 1315 3885 1316 3915
rect 1284 3884 1316 3885
rect 1284 3835 1316 3836
rect 1284 3805 1285 3835
rect 1285 3805 1315 3835
rect 1315 3805 1316 3835
rect 1284 3804 1316 3805
rect 1284 3755 1316 3756
rect 1284 3725 1285 3755
rect 1285 3725 1315 3755
rect 1315 3725 1316 3755
rect 1284 3724 1316 3725
rect 1284 3675 1316 3676
rect 1284 3645 1285 3675
rect 1285 3645 1315 3675
rect 1315 3645 1316 3675
rect 1284 3644 1316 3645
rect 1364 4395 1396 4396
rect 1364 4365 1365 4395
rect 1365 4365 1395 4395
rect 1395 4365 1396 4395
rect 1364 4364 1396 4365
rect 1364 4284 1396 4316
rect 1364 4235 1396 4236
rect 1364 4205 1365 4235
rect 1365 4205 1395 4235
rect 1395 4205 1396 4235
rect 1364 4204 1396 4205
rect 1364 4124 1396 4156
rect 1364 4075 1396 4076
rect 1364 4045 1365 4075
rect 1365 4045 1395 4075
rect 1395 4045 1396 4075
rect 1364 4044 1396 4045
rect 1364 3995 1396 3996
rect 1364 3965 1365 3995
rect 1365 3965 1395 3995
rect 1395 3965 1396 3995
rect 1364 3964 1396 3965
rect 1364 3915 1396 3916
rect 1364 3885 1365 3915
rect 1365 3885 1395 3915
rect 1395 3885 1396 3915
rect 1364 3884 1396 3885
rect 1364 3835 1396 3836
rect 1364 3805 1365 3835
rect 1365 3805 1395 3835
rect 1395 3805 1396 3835
rect 1364 3804 1396 3805
rect 1364 3755 1396 3756
rect 1364 3725 1365 3755
rect 1365 3725 1395 3755
rect 1395 3725 1396 3755
rect 1364 3724 1396 3725
rect 1364 3675 1396 3676
rect 1364 3645 1365 3675
rect 1365 3645 1395 3675
rect 1395 3645 1396 3675
rect 1364 3644 1396 3645
rect 1444 4395 1476 4396
rect 1444 4365 1445 4395
rect 1445 4365 1475 4395
rect 1475 4365 1476 4395
rect 1444 4364 1476 4365
rect 1444 4284 1476 4316
rect 1444 4235 1476 4236
rect 1444 4205 1445 4235
rect 1445 4205 1475 4235
rect 1475 4205 1476 4235
rect 1444 4204 1476 4205
rect 1444 4124 1476 4156
rect 1444 4075 1476 4076
rect 1444 4045 1445 4075
rect 1445 4045 1475 4075
rect 1475 4045 1476 4075
rect 1444 4044 1476 4045
rect 1444 3995 1476 3996
rect 1444 3965 1445 3995
rect 1445 3965 1475 3995
rect 1475 3965 1476 3995
rect 1444 3964 1476 3965
rect 1444 3915 1476 3916
rect 1444 3885 1445 3915
rect 1445 3885 1475 3915
rect 1475 3885 1476 3915
rect 1444 3884 1476 3885
rect 1444 3835 1476 3836
rect 1444 3805 1445 3835
rect 1445 3805 1475 3835
rect 1475 3805 1476 3835
rect 1444 3804 1476 3805
rect 1444 3755 1476 3756
rect 1444 3725 1445 3755
rect 1445 3725 1475 3755
rect 1475 3725 1476 3755
rect 1444 3724 1476 3725
rect 1444 3675 1476 3676
rect 1444 3645 1445 3675
rect 1445 3645 1475 3675
rect 1475 3645 1476 3675
rect 1444 3644 1476 3645
rect 1524 4395 1556 4396
rect 1524 4365 1525 4395
rect 1525 4365 1555 4395
rect 1555 4365 1556 4395
rect 1524 4364 1556 4365
rect 1524 4284 1556 4316
rect 1524 4235 1556 4236
rect 1524 4205 1525 4235
rect 1525 4205 1555 4235
rect 1555 4205 1556 4235
rect 1524 4204 1556 4205
rect 1524 4124 1556 4156
rect 1524 4075 1556 4076
rect 1524 4045 1525 4075
rect 1525 4045 1555 4075
rect 1555 4045 1556 4075
rect 1524 4044 1556 4045
rect 1524 3995 1556 3996
rect 1524 3965 1525 3995
rect 1525 3965 1555 3995
rect 1555 3965 1556 3995
rect 1524 3964 1556 3965
rect 1524 3915 1556 3916
rect 1524 3885 1525 3915
rect 1525 3885 1555 3915
rect 1555 3885 1556 3915
rect 1524 3884 1556 3885
rect 1524 3835 1556 3836
rect 1524 3805 1525 3835
rect 1525 3805 1555 3835
rect 1555 3805 1556 3835
rect 1524 3804 1556 3805
rect 1524 3755 1556 3756
rect 1524 3725 1525 3755
rect 1525 3725 1555 3755
rect 1555 3725 1556 3755
rect 1524 3724 1556 3725
rect 1524 3675 1556 3676
rect 1524 3645 1525 3675
rect 1525 3645 1555 3675
rect 1555 3645 1556 3675
rect 1524 3644 1556 3645
rect 1604 4395 1636 4396
rect 1604 4365 1605 4395
rect 1605 4365 1635 4395
rect 1635 4365 1636 4395
rect 1604 4364 1636 4365
rect 1604 4284 1636 4316
rect 1604 4235 1636 4236
rect 1604 4205 1605 4235
rect 1605 4205 1635 4235
rect 1635 4205 1636 4235
rect 1604 4204 1636 4205
rect 1604 4124 1636 4156
rect 1604 4075 1636 4076
rect 1604 4045 1605 4075
rect 1605 4045 1635 4075
rect 1635 4045 1636 4075
rect 1604 4044 1636 4045
rect 1604 3995 1636 3996
rect 1604 3965 1605 3995
rect 1605 3965 1635 3995
rect 1635 3965 1636 3995
rect 1604 3964 1636 3965
rect 1604 3915 1636 3916
rect 1604 3885 1605 3915
rect 1605 3885 1635 3915
rect 1635 3885 1636 3915
rect 1604 3884 1636 3885
rect 1604 3835 1636 3836
rect 1604 3805 1605 3835
rect 1605 3805 1635 3835
rect 1635 3805 1636 3835
rect 1604 3804 1636 3805
rect 1604 3755 1636 3756
rect 1604 3725 1605 3755
rect 1605 3725 1635 3755
rect 1635 3725 1636 3755
rect 1604 3724 1636 3725
rect 1604 3675 1636 3676
rect 1604 3645 1605 3675
rect 1605 3645 1635 3675
rect 1635 3645 1636 3675
rect 1604 3644 1636 3645
rect 1684 4395 1716 4396
rect 1684 4365 1685 4395
rect 1685 4365 1715 4395
rect 1715 4365 1716 4395
rect 1684 4364 1716 4365
rect 1684 4284 1716 4316
rect 1684 4235 1716 4236
rect 1684 4205 1685 4235
rect 1685 4205 1715 4235
rect 1715 4205 1716 4235
rect 1684 4204 1716 4205
rect 1684 4124 1716 4156
rect 1684 4075 1716 4076
rect 1684 4045 1685 4075
rect 1685 4045 1715 4075
rect 1715 4045 1716 4075
rect 1684 4044 1716 4045
rect 1684 3995 1716 3996
rect 1684 3965 1685 3995
rect 1685 3965 1715 3995
rect 1715 3965 1716 3995
rect 1684 3964 1716 3965
rect 1684 3915 1716 3916
rect 1684 3885 1685 3915
rect 1685 3885 1715 3915
rect 1715 3885 1716 3915
rect 1684 3884 1716 3885
rect 1684 3835 1716 3836
rect 1684 3805 1685 3835
rect 1685 3805 1715 3835
rect 1715 3805 1716 3835
rect 1684 3804 1716 3805
rect 1684 3755 1716 3756
rect 1684 3725 1685 3755
rect 1685 3725 1715 3755
rect 1715 3725 1716 3755
rect 1684 3724 1716 3725
rect 1684 3675 1716 3676
rect 1684 3645 1685 3675
rect 1685 3645 1715 3675
rect 1715 3645 1716 3675
rect 1684 3644 1716 3645
rect 1764 4395 1796 4396
rect 1764 4365 1765 4395
rect 1765 4365 1795 4395
rect 1795 4365 1796 4395
rect 1764 4364 1796 4365
rect 1764 4284 1796 4316
rect 1764 4235 1796 4236
rect 1764 4205 1765 4235
rect 1765 4205 1795 4235
rect 1795 4205 1796 4235
rect 1764 4204 1796 4205
rect 1764 4124 1796 4156
rect 1764 4075 1796 4076
rect 1764 4045 1765 4075
rect 1765 4045 1795 4075
rect 1795 4045 1796 4075
rect 1764 4044 1796 4045
rect 1764 3995 1796 3996
rect 1764 3965 1765 3995
rect 1765 3965 1795 3995
rect 1795 3965 1796 3995
rect 1764 3964 1796 3965
rect 1764 3915 1796 3916
rect 1764 3885 1765 3915
rect 1765 3885 1795 3915
rect 1795 3885 1796 3915
rect 1764 3884 1796 3885
rect 1764 3835 1796 3836
rect 1764 3805 1765 3835
rect 1765 3805 1795 3835
rect 1795 3805 1796 3835
rect 1764 3804 1796 3805
rect 1764 3755 1796 3756
rect 1764 3725 1765 3755
rect 1765 3725 1795 3755
rect 1795 3725 1796 3755
rect 1764 3724 1796 3725
rect 1764 3675 1796 3676
rect 1764 3645 1765 3675
rect 1765 3645 1795 3675
rect 1795 3645 1796 3675
rect 1764 3644 1796 3645
rect 1844 4395 1876 4396
rect 1844 4365 1845 4395
rect 1845 4365 1875 4395
rect 1875 4365 1876 4395
rect 1844 4364 1876 4365
rect 1844 4284 1876 4316
rect 1844 4235 1876 4236
rect 1844 4205 1845 4235
rect 1845 4205 1875 4235
rect 1875 4205 1876 4235
rect 1844 4204 1876 4205
rect 1844 4124 1876 4156
rect 1844 4075 1876 4076
rect 1844 4045 1845 4075
rect 1845 4045 1875 4075
rect 1875 4045 1876 4075
rect 1844 4044 1876 4045
rect 1844 3995 1876 3996
rect 1844 3965 1845 3995
rect 1845 3965 1875 3995
rect 1875 3965 1876 3995
rect 1844 3964 1876 3965
rect 1844 3915 1876 3916
rect 1844 3885 1845 3915
rect 1845 3885 1875 3915
rect 1875 3885 1876 3915
rect 1844 3884 1876 3885
rect 1844 3835 1876 3836
rect 1844 3805 1845 3835
rect 1845 3805 1875 3835
rect 1875 3805 1876 3835
rect 1844 3804 1876 3805
rect 1844 3755 1876 3756
rect 1844 3725 1845 3755
rect 1845 3725 1875 3755
rect 1875 3725 1876 3755
rect 1844 3724 1876 3725
rect 1844 3675 1876 3676
rect 1844 3645 1845 3675
rect 1845 3645 1875 3675
rect 1875 3645 1876 3675
rect 1844 3644 1876 3645
rect 1924 4395 1956 4396
rect 1924 4365 1925 4395
rect 1925 4365 1955 4395
rect 1955 4365 1956 4395
rect 1924 4364 1956 4365
rect 1924 4284 1956 4316
rect 1924 4235 1956 4236
rect 1924 4205 1925 4235
rect 1925 4205 1955 4235
rect 1955 4205 1956 4235
rect 1924 4204 1956 4205
rect 1924 4124 1956 4156
rect 1924 4075 1956 4076
rect 1924 4045 1925 4075
rect 1925 4045 1955 4075
rect 1955 4045 1956 4075
rect 1924 4044 1956 4045
rect 1924 3995 1956 3996
rect 1924 3965 1925 3995
rect 1925 3965 1955 3995
rect 1955 3965 1956 3995
rect 1924 3964 1956 3965
rect 1924 3915 1956 3916
rect 1924 3885 1925 3915
rect 1925 3885 1955 3915
rect 1955 3885 1956 3915
rect 1924 3884 1956 3885
rect 1924 3835 1956 3836
rect 1924 3805 1925 3835
rect 1925 3805 1955 3835
rect 1955 3805 1956 3835
rect 1924 3804 1956 3805
rect 1924 3755 1956 3756
rect 1924 3725 1925 3755
rect 1925 3725 1955 3755
rect 1955 3725 1956 3755
rect 1924 3724 1956 3725
rect 1924 3675 1956 3676
rect 1924 3645 1925 3675
rect 1925 3645 1955 3675
rect 1955 3645 1956 3675
rect 1924 3644 1956 3645
rect 2004 4395 2036 4396
rect 2004 4365 2005 4395
rect 2005 4365 2035 4395
rect 2035 4365 2036 4395
rect 2004 4364 2036 4365
rect 2004 4284 2036 4316
rect 2004 4235 2036 4236
rect 2004 4205 2005 4235
rect 2005 4205 2035 4235
rect 2035 4205 2036 4235
rect 2004 4204 2036 4205
rect 2004 4124 2036 4156
rect 2004 4075 2036 4076
rect 2004 4045 2005 4075
rect 2005 4045 2035 4075
rect 2035 4045 2036 4075
rect 2004 4044 2036 4045
rect 2004 3995 2036 3996
rect 2004 3965 2005 3995
rect 2005 3965 2035 3995
rect 2035 3965 2036 3995
rect 2004 3964 2036 3965
rect 2004 3915 2036 3916
rect 2004 3885 2005 3915
rect 2005 3885 2035 3915
rect 2035 3885 2036 3915
rect 2004 3884 2036 3885
rect 2004 3835 2036 3836
rect 2004 3805 2005 3835
rect 2005 3805 2035 3835
rect 2035 3805 2036 3835
rect 2004 3804 2036 3805
rect 2004 3755 2036 3756
rect 2004 3725 2005 3755
rect 2005 3725 2035 3755
rect 2035 3725 2036 3755
rect 2004 3724 2036 3725
rect 2004 3675 2036 3676
rect 2004 3645 2005 3675
rect 2005 3645 2035 3675
rect 2035 3645 2036 3675
rect 2004 3644 2036 3645
rect 2084 4395 2116 4396
rect 2084 4365 2085 4395
rect 2085 4365 2115 4395
rect 2115 4365 2116 4395
rect 2084 4364 2116 4365
rect 2084 4284 2116 4316
rect 2084 4235 2116 4236
rect 2084 4205 2085 4235
rect 2085 4205 2115 4235
rect 2115 4205 2116 4235
rect 2084 4204 2116 4205
rect 2084 4124 2116 4156
rect 2084 4075 2116 4076
rect 2084 4045 2085 4075
rect 2085 4045 2115 4075
rect 2115 4045 2116 4075
rect 2084 4044 2116 4045
rect 2084 3995 2116 3996
rect 2084 3965 2085 3995
rect 2085 3965 2115 3995
rect 2115 3965 2116 3995
rect 2084 3964 2116 3965
rect 2084 3915 2116 3916
rect 2084 3885 2085 3915
rect 2085 3885 2115 3915
rect 2115 3885 2116 3915
rect 2084 3884 2116 3885
rect 2084 3835 2116 3836
rect 2084 3805 2085 3835
rect 2085 3805 2115 3835
rect 2115 3805 2116 3835
rect 2084 3804 2116 3805
rect 2084 3755 2116 3756
rect 2084 3725 2085 3755
rect 2085 3725 2115 3755
rect 2115 3725 2116 3755
rect 2084 3724 2116 3725
rect 2084 3675 2116 3676
rect 2084 3645 2085 3675
rect 2085 3645 2115 3675
rect 2115 3645 2116 3675
rect 2084 3644 2116 3645
rect 2164 4395 2196 4396
rect 2164 4365 2165 4395
rect 2165 4365 2195 4395
rect 2195 4365 2196 4395
rect 2164 4364 2196 4365
rect 2164 4284 2196 4316
rect 2164 4235 2196 4236
rect 2164 4205 2165 4235
rect 2165 4205 2195 4235
rect 2195 4205 2196 4235
rect 2164 4204 2196 4205
rect 2164 4124 2196 4156
rect 2164 4075 2196 4076
rect 2164 4045 2165 4075
rect 2165 4045 2195 4075
rect 2195 4045 2196 4075
rect 2164 4044 2196 4045
rect 2164 3995 2196 3996
rect 2164 3965 2165 3995
rect 2165 3965 2195 3995
rect 2195 3965 2196 3995
rect 2164 3964 2196 3965
rect 2164 3915 2196 3916
rect 2164 3885 2165 3915
rect 2165 3885 2195 3915
rect 2195 3885 2196 3915
rect 2164 3884 2196 3885
rect 2164 3835 2196 3836
rect 2164 3805 2165 3835
rect 2165 3805 2195 3835
rect 2195 3805 2196 3835
rect 2164 3804 2196 3805
rect 2164 3755 2196 3756
rect 2164 3725 2165 3755
rect 2165 3725 2195 3755
rect 2195 3725 2196 3755
rect 2164 3724 2196 3725
rect 2164 3675 2196 3676
rect 2164 3645 2165 3675
rect 2165 3645 2195 3675
rect 2195 3645 2196 3675
rect 2164 3644 2196 3645
rect 2244 4395 2276 4396
rect 2244 4365 2245 4395
rect 2245 4365 2275 4395
rect 2275 4365 2276 4395
rect 2244 4364 2276 4365
rect 2244 4284 2276 4316
rect 2244 4235 2276 4236
rect 2244 4205 2245 4235
rect 2245 4205 2275 4235
rect 2275 4205 2276 4235
rect 2244 4204 2276 4205
rect 2244 4124 2276 4156
rect 2244 4075 2276 4076
rect 2244 4045 2245 4075
rect 2245 4045 2275 4075
rect 2275 4045 2276 4075
rect 2244 4044 2276 4045
rect 2244 3995 2276 3996
rect 2244 3965 2245 3995
rect 2245 3965 2275 3995
rect 2275 3965 2276 3995
rect 2244 3964 2276 3965
rect 2244 3915 2276 3916
rect 2244 3885 2245 3915
rect 2245 3885 2275 3915
rect 2275 3885 2276 3915
rect 2244 3884 2276 3885
rect 2244 3835 2276 3836
rect 2244 3805 2245 3835
rect 2245 3805 2275 3835
rect 2275 3805 2276 3835
rect 2244 3804 2276 3805
rect 2244 3755 2276 3756
rect 2244 3725 2245 3755
rect 2245 3725 2275 3755
rect 2275 3725 2276 3755
rect 2244 3724 2276 3725
rect 2244 3675 2276 3676
rect 2244 3645 2245 3675
rect 2245 3645 2275 3675
rect 2275 3645 2276 3675
rect 2244 3644 2276 3645
rect 2324 4395 2356 4396
rect 2324 4365 2325 4395
rect 2325 4365 2355 4395
rect 2355 4365 2356 4395
rect 2324 4364 2356 4365
rect 2324 4284 2356 4316
rect 2324 4235 2356 4236
rect 2324 4205 2325 4235
rect 2325 4205 2355 4235
rect 2355 4205 2356 4235
rect 2324 4204 2356 4205
rect 2324 4124 2356 4156
rect 2324 4075 2356 4076
rect 2324 4045 2325 4075
rect 2325 4045 2355 4075
rect 2355 4045 2356 4075
rect 2324 4044 2356 4045
rect 2324 3995 2356 3996
rect 2324 3965 2325 3995
rect 2325 3965 2355 3995
rect 2355 3965 2356 3995
rect 2324 3964 2356 3965
rect 2324 3915 2356 3916
rect 2324 3885 2325 3915
rect 2325 3885 2355 3915
rect 2355 3885 2356 3915
rect 2324 3884 2356 3885
rect 2324 3835 2356 3836
rect 2324 3805 2325 3835
rect 2325 3805 2355 3835
rect 2355 3805 2356 3835
rect 2324 3804 2356 3805
rect 2324 3755 2356 3756
rect 2324 3725 2325 3755
rect 2325 3725 2355 3755
rect 2355 3725 2356 3755
rect 2324 3724 2356 3725
rect 2324 3675 2356 3676
rect 2324 3645 2325 3675
rect 2325 3645 2355 3675
rect 2355 3645 2356 3675
rect 2324 3644 2356 3645
rect 2404 4395 2436 4396
rect 2404 4365 2405 4395
rect 2405 4365 2435 4395
rect 2435 4365 2436 4395
rect 2404 4364 2436 4365
rect 2404 4284 2436 4316
rect 2404 4235 2436 4236
rect 2404 4205 2405 4235
rect 2405 4205 2435 4235
rect 2435 4205 2436 4235
rect 2404 4204 2436 4205
rect 2404 4124 2436 4156
rect 2404 4075 2436 4076
rect 2404 4045 2405 4075
rect 2405 4045 2435 4075
rect 2435 4045 2436 4075
rect 2404 4044 2436 4045
rect 2404 3995 2436 3996
rect 2404 3965 2405 3995
rect 2405 3965 2435 3995
rect 2435 3965 2436 3995
rect 2404 3964 2436 3965
rect 2404 3915 2436 3916
rect 2404 3885 2405 3915
rect 2405 3885 2435 3915
rect 2435 3885 2436 3915
rect 2404 3884 2436 3885
rect 2404 3835 2436 3836
rect 2404 3805 2405 3835
rect 2405 3805 2435 3835
rect 2435 3805 2436 3835
rect 2404 3804 2436 3805
rect 2404 3755 2436 3756
rect 2404 3725 2405 3755
rect 2405 3725 2435 3755
rect 2435 3725 2436 3755
rect 2404 3724 2436 3725
rect 2404 3675 2436 3676
rect 2404 3645 2405 3675
rect 2405 3645 2435 3675
rect 2435 3645 2436 3675
rect 2404 3644 2436 3645
rect 2484 4395 2516 4396
rect 2484 4365 2485 4395
rect 2485 4365 2515 4395
rect 2515 4365 2516 4395
rect 2484 4364 2516 4365
rect 2484 4284 2516 4316
rect 2484 4235 2516 4236
rect 2484 4205 2485 4235
rect 2485 4205 2515 4235
rect 2515 4205 2516 4235
rect 2484 4204 2516 4205
rect 2484 4124 2516 4156
rect 2484 4075 2516 4076
rect 2484 4045 2485 4075
rect 2485 4045 2515 4075
rect 2515 4045 2516 4075
rect 2484 4044 2516 4045
rect 2484 3995 2516 3996
rect 2484 3965 2485 3995
rect 2485 3965 2515 3995
rect 2515 3965 2516 3995
rect 2484 3964 2516 3965
rect 2484 3915 2516 3916
rect 2484 3885 2485 3915
rect 2485 3885 2515 3915
rect 2515 3885 2516 3915
rect 2484 3884 2516 3885
rect 2484 3835 2516 3836
rect 2484 3805 2485 3835
rect 2485 3805 2515 3835
rect 2515 3805 2516 3835
rect 2484 3804 2516 3805
rect 2484 3755 2516 3756
rect 2484 3725 2485 3755
rect 2485 3725 2515 3755
rect 2515 3725 2516 3755
rect 2484 3724 2516 3725
rect 2484 3675 2516 3676
rect 2484 3645 2485 3675
rect 2485 3645 2515 3675
rect 2515 3645 2516 3675
rect 2484 3644 2516 3645
rect 2564 4395 2596 4396
rect 2564 4365 2565 4395
rect 2565 4365 2595 4395
rect 2595 4365 2596 4395
rect 2564 4364 2596 4365
rect 2564 4284 2596 4316
rect 2564 4235 2596 4236
rect 2564 4205 2565 4235
rect 2565 4205 2595 4235
rect 2595 4205 2596 4235
rect 2564 4204 2596 4205
rect 2564 4124 2596 4156
rect 2564 4075 2596 4076
rect 2564 4045 2565 4075
rect 2565 4045 2595 4075
rect 2595 4045 2596 4075
rect 2564 4044 2596 4045
rect 2564 3995 2596 3996
rect 2564 3965 2565 3995
rect 2565 3965 2595 3995
rect 2595 3965 2596 3995
rect 2564 3964 2596 3965
rect 2564 3915 2596 3916
rect 2564 3885 2565 3915
rect 2565 3885 2595 3915
rect 2595 3885 2596 3915
rect 2564 3884 2596 3885
rect 2564 3835 2596 3836
rect 2564 3805 2565 3835
rect 2565 3805 2595 3835
rect 2595 3805 2596 3835
rect 2564 3804 2596 3805
rect 2564 3755 2596 3756
rect 2564 3725 2565 3755
rect 2565 3725 2595 3755
rect 2595 3725 2596 3755
rect 2564 3724 2596 3725
rect 2564 3675 2596 3676
rect 2564 3645 2565 3675
rect 2565 3645 2595 3675
rect 2595 3645 2596 3675
rect 2564 3644 2596 3645
rect 2644 4395 2676 4396
rect 2644 4365 2645 4395
rect 2645 4365 2675 4395
rect 2675 4365 2676 4395
rect 2644 4364 2676 4365
rect 2644 4284 2676 4316
rect 2644 4235 2676 4236
rect 2644 4205 2645 4235
rect 2645 4205 2675 4235
rect 2675 4205 2676 4235
rect 2644 4204 2676 4205
rect 2644 4124 2676 4156
rect 2644 4075 2676 4076
rect 2644 4045 2645 4075
rect 2645 4045 2675 4075
rect 2675 4045 2676 4075
rect 2644 4044 2676 4045
rect 2644 3995 2676 3996
rect 2644 3965 2645 3995
rect 2645 3965 2675 3995
rect 2675 3965 2676 3995
rect 2644 3964 2676 3965
rect 2644 3915 2676 3916
rect 2644 3885 2645 3915
rect 2645 3885 2675 3915
rect 2675 3885 2676 3915
rect 2644 3884 2676 3885
rect 2644 3835 2676 3836
rect 2644 3805 2645 3835
rect 2645 3805 2675 3835
rect 2675 3805 2676 3835
rect 2644 3804 2676 3805
rect 2644 3755 2676 3756
rect 2644 3725 2645 3755
rect 2645 3725 2675 3755
rect 2675 3725 2676 3755
rect 2644 3724 2676 3725
rect 2644 3675 2676 3676
rect 2644 3645 2645 3675
rect 2645 3645 2675 3675
rect 2675 3645 2676 3675
rect 2644 3644 2676 3645
rect 2724 4395 2756 4396
rect 2724 4365 2725 4395
rect 2725 4365 2755 4395
rect 2755 4365 2756 4395
rect 2724 4364 2756 4365
rect 2724 4284 2756 4316
rect 2724 4235 2756 4236
rect 2724 4205 2725 4235
rect 2725 4205 2755 4235
rect 2755 4205 2756 4235
rect 2724 4204 2756 4205
rect 2724 4124 2756 4156
rect 2724 4075 2756 4076
rect 2724 4045 2725 4075
rect 2725 4045 2755 4075
rect 2755 4045 2756 4075
rect 2724 4044 2756 4045
rect 2724 3995 2756 3996
rect 2724 3965 2725 3995
rect 2725 3965 2755 3995
rect 2755 3965 2756 3995
rect 2724 3964 2756 3965
rect 2724 3915 2756 3916
rect 2724 3885 2725 3915
rect 2725 3885 2755 3915
rect 2755 3885 2756 3915
rect 2724 3884 2756 3885
rect 2724 3835 2756 3836
rect 2724 3805 2725 3835
rect 2725 3805 2755 3835
rect 2755 3805 2756 3835
rect 2724 3804 2756 3805
rect 2724 3755 2756 3756
rect 2724 3725 2725 3755
rect 2725 3725 2755 3755
rect 2755 3725 2756 3755
rect 2724 3724 2756 3725
rect 2724 3675 2756 3676
rect 2724 3645 2725 3675
rect 2725 3645 2755 3675
rect 2755 3645 2756 3675
rect 2724 3644 2756 3645
rect 2804 4395 2836 4396
rect 2804 4365 2805 4395
rect 2805 4365 2835 4395
rect 2835 4365 2836 4395
rect 2804 4364 2836 4365
rect 2804 4284 2836 4316
rect 2804 4235 2836 4236
rect 2804 4205 2805 4235
rect 2805 4205 2835 4235
rect 2835 4205 2836 4235
rect 2804 4204 2836 4205
rect 2804 4124 2836 4156
rect 2804 4075 2836 4076
rect 2804 4045 2805 4075
rect 2805 4045 2835 4075
rect 2835 4045 2836 4075
rect 2804 4044 2836 4045
rect 2804 3995 2836 3996
rect 2804 3965 2805 3995
rect 2805 3965 2835 3995
rect 2835 3965 2836 3995
rect 2804 3964 2836 3965
rect 2804 3915 2836 3916
rect 2804 3885 2805 3915
rect 2805 3885 2835 3915
rect 2835 3885 2836 3915
rect 2804 3884 2836 3885
rect 2804 3835 2836 3836
rect 2804 3805 2805 3835
rect 2805 3805 2835 3835
rect 2835 3805 2836 3835
rect 2804 3804 2836 3805
rect 2804 3755 2836 3756
rect 2804 3725 2805 3755
rect 2805 3725 2835 3755
rect 2835 3725 2836 3755
rect 2804 3724 2836 3725
rect 2804 3675 2836 3676
rect 2804 3645 2805 3675
rect 2805 3645 2835 3675
rect 2835 3645 2836 3675
rect 2804 3644 2836 3645
rect 2884 4395 2916 4396
rect 2884 4365 2885 4395
rect 2885 4365 2915 4395
rect 2915 4365 2916 4395
rect 2884 4364 2916 4365
rect 2884 4284 2916 4316
rect 2884 4235 2916 4236
rect 2884 4205 2885 4235
rect 2885 4205 2915 4235
rect 2915 4205 2916 4235
rect 2884 4204 2916 4205
rect 2884 4124 2916 4156
rect 2884 4075 2916 4076
rect 2884 4045 2885 4075
rect 2885 4045 2915 4075
rect 2915 4045 2916 4075
rect 2884 4044 2916 4045
rect 2884 3995 2916 3996
rect 2884 3965 2885 3995
rect 2885 3965 2915 3995
rect 2915 3965 2916 3995
rect 2884 3964 2916 3965
rect 2884 3915 2916 3916
rect 2884 3885 2885 3915
rect 2885 3885 2915 3915
rect 2915 3885 2916 3915
rect 2884 3884 2916 3885
rect 2884 3835 2916 3836
rect 2884 3805 2885 3835
rect 2885 3805 2915 3835
rect 2915 3805 2916 3835
rect 2884 3804 2916 3805
rect 2884 3755 2916 3756
rect 2884 3725 2885 3755
rect 2885 3725 2915 3755
rect 2915 3725 2916 3755
rect 2884 3724 2916 3725
rect 2884 3675 2916 3676
rect 2884 3645 2885 3675
rect 2885 3645 2915 3675
rect 2915 3645 2916 3675
rect 2884 3644 2916 3645
rect 2964 4395 2996 4396
rect 2964 4365 2965 4395
rect 2965 4365 2995 4395
rect 2995 4365 2996 4395
rect 2964 4364 2996 4365
rect 2964 4284 2996 4316
rect 2964 4235 2996 4236
rect 2964 4205 2965 4235
rect 2965 4205 2995 4235
rect 2995 4205 2996 4235
rect 2964 4204 2996 4205
rect 2964 4124 2996 4156
rect 2964 4075 2996 4076
rect 2964 4045 2965 4075
rect 2965 4045 2995 4075
rect 2995 4045 2996 4075
rect 2964 4044 2996 4045
rect 2964 3995 2996 3996
rect 2964 3965 2965 3995
rect 2965 3965 2995 3995
rect 2995 3965 2996 3995
rect 2964 3964 2996 3965
rect 2964 3915 2996 3916
rect 2964 3885 2965 3915
rect 2965 3885 2995 3915
rect 2995 3885 2996 3915
rect 2964 3884 2996 3885
rect 2964 3835 2996 3836
rect 2964 3805 2965 3835
rect 2965 3805 2995 3835
rect 2995 3805 2996 3835
rect 2964 3804 2996 3805
rect 2964 3755 2996 3756
rect 2964 3725 2965 3755
rect 2965 3725 2995 3755
rect 2995 3725 2996 3755
rect 2964 3724 2996 3725
rect 2964 3675 2996 3676
rect 2964 3645 2965 3675
rect 2965 3645 2995 3675
rect 2995 3645 2996 3675
rect 2964 3644 2996 3645
rect 3044 4395 3076 4396
rect 3044 4365 3045 4395
rect 3045 4365 3075 4395
rect 3075 4365 3076 4395
rect 3044 4364 3076 4365
rect 3044 4284 3076 4316
rect 3044 4235 3076 4236
rect 3044 4205 3045 4235
rect 3045 4205 3075 4235
rect 3075 4205 3076 4235
rect 3044 4204 3076 4205
rect 3044 4124 3076 4156
rect 3044 4075 3076 4076
rect 3044 4045 3045 4075
rect 3045 4045 3075 4075
rect 3075 4045 3076 4075
rect 3044 4044 3076 4045
rect 3044 3995 3076 3996
rect 3044 3965 3045 3995
rect 3045 3965 3075 3995
rect 3075 3965 3076 3995
rect 3044 3964 3076 3965
rect 3044 3915 3076 3916
rect 3044 3885 3045 3915
rect 3045 3885 3075 3915
rect 3075 3885 3076 3915
rect 3044 3884 3076 3885
rect 3044 3835 3076 3836
rect 3044 3805 3045 3835
rect 3045 3805 3075 3835
rect 3075 3805 3076 3835
rect 3044 3804 3076 3805
rect 3044 3755 3076 3756
rect 3044 3725 3045 3755
rect 3045 3725 3075 3755
rect 3075 3725 3076 3755
rect 3044 3724 3076 3725
rect 3044 3675 3076 3676
rect 3044 3645 3045 3675
rect 3045 3645 3075 3675
rect 3075 3645 3076 3675
rect 3044 3644 3076 3645
rect 3124 4395 3156 4396
rect 3124 4365 3125 4395
rect 3125 4365 3155 4395
rect 3155 4365 3156 4395
rect 3124 4364 3156 4365
rect 3124 4284 3156 4316
rect 3124 4235 3156 4236
rect 3124 4205 3125 4235
rect 3125 4205 3155 4235
rect 3155 4205 3156 4235
rect 3124 4204 3156 4205
rect 3124 4124 3156 4156
rect 3124 4075 3156 4076
rect 3124 4045 3125 4075
rect 3125 4045 3155 4075
rect 3155 4045 3156 4075
rect 3124 4044 3156 4045
rect 3124 3995 3156 3996
rect 3124 3965 3125 3995
rect 3125 3965 3155 3995
rect 3155 3965 3156 3995
rect 3124 3964 3156 3965
rect 3124 3915 3156 3916
rect 3124 3885 3125 3915
rect 3125 3885 3155 3915
rect 3155 3885 3156 3915
rect 3124 3884 3156 3885
rect 3124 3835 3156 3836
rect 3124 3805 3125 3835
rect 3125 3805 3155 3835
rect 3155 3805 3156 3835
rect 3124 3804 3156 3805
rect 3124 3755 3156 3756
rect 3124 3725 3125 3755
rect 3125 3725 3155 3755
rect 3155 3725 3156 3755
rect 3124 3724 3156 3725
rect 3124 3675 3156 3676
rect 3124 3645 3125 3675
rect 3125 3645 3155 3675
rect 3155 3645 3156 3675
rect 3124 3644 3156 3645
rect 3204 4395 3236 4396
rect 3204 4365 3205 4395
rect 3205 4365 3235 4395
rect 3235 4365 3236 4395
rect 3204 4364 3236 4365
rect 3204 4284 3236 4316
rect 3204 4235 3236 4236
rect 3204 4205 3205 4235
rect 3205 4205 3235 4235
rect 3235 4205 3236 4235
rect 3204 4204 3236 4205
rect 3204 4124 3236 4156
rect 3204 4075 3236 4076
rect 3204 4045 3205 4075
rect 3205 4045 3235 4075
rect 3235 4045 3236 4075
rect 3204 4044 3236 4045
rect 3204 3995 3236 3996
rect 3204 3965 3205 3995
rect 3205 3965 3235 3995
rect 3235 3965 3236 3995
rect 3204 3964 3236 3965
rect 3204 3915 3236 3916
rect 3204 3885 3205 3915
rect 3205 3885 3235 3915
rect 3235 3885 3236 3915
rect 3204 3884 3236 3885
rect 3204 3835 3236 3836
rect 3204 3805 3205 3835
rect 3205 3805 3235 3835
rect 3235 3805 3236 3835
rect 3204 3804 3236 3805
rect 3204 3755 3236 3756
rect 3204 3725 3205 3755
rect 3205 3725 3235 3755
rect 3235 3725 3236 3755
rect 3204 3724 3236 3725
rect 3204 3675 3236 3676
rect 3204 3645 3205 3675
rect 3205 3645 3235 3675
rect 3235 3645 3236 3675
rect 3204 3644 3236 3645
rect 3284 4395 3316 4396
rect 3284 4365 3285 4395
rect 3285 4365 3315 4395
rect 3315 4365 3316 4395
rect 3284 4364 3316 4365
rect 3284 4284 3316 4316
rect 3284 4235 3316 4236
rect 3284 4205 3285 4235
rect 3285 4205 3315 4235
rect 3315 4205 3316 4235
rect 3284 4204 3316 4205
rect 3284 4124 3316 4156
rect 3284 4075 3316 4076
rect 3284 4045 3285 4075
rect 3285 4045 3315 4075
rect 3315 4045 3316 4075
rect 3284 4044 3316 4045
rect 3284 3995 3316 3996
rect 3284 3965 3285 3995
rect 3285 3965 3315 3995
rect 3315 3965 3316 3995
rect 3284 3964 3316 3965
rect 3284 3915 3316 3916
rect 3284 3885 3285 3915
rect 3285 3885 3315 3915
rect 3315 3885 3316 3915
rect 3284 3884 3316 3885
rect 3284 3835 3316 3836
rect 3284 3805 3285 3835
rect 3285 3805 3315 3835
rect 3315 3805 3316 3835
rect 3284 3804 3316 3805
rect 3284 3755 3316 3756
rect 3284 3725 3285 3755
rect 3285 3725 3315 3755
rect 3315 3725 3316 3755
rect 3284 3724 3316 3725
rect 3284 3675 3316 3676
rect 3284 3645 3285 3675
rect 3285 3645 3315 3675
rect 3315 3645 3316 3675
rect 3284 3644 3316 3645
rect 3364 4395 3396 4396
rect 3364 4365 3365 4395
rect 3365 4365 3395 4395
rect 3395 4365 3396 4395
rect 3364 4364 3396 4365
rect 3364 4284 3396 4316
rect 3364 4235 3396 4236
rect 3364 4205 3365 4235
rect 3365 4205 3395 4235
rect 3395 4205 3396 4235
rect 3364 4204 3396 4205
rect 3364 4124 3396 4156
rect 3364 4075 3396 4076
rect 3364 4045 3365 4075
rect 3365 4045 3395 4075
rect 3395 4045 3396 4075
rect 3364 4044 3396 4045
rect 3364 3995 3396 3996
rect 3364 3965 3365 3995
rect 3365 3965 3395 3995
rect 3395 3965 3396 3995
rect 3364 3964 3396 3965
rect 3364 3915 3396 3916
rect 3364 3885 3365 3915
rect 3365 3885 3395 3915
rect 3395 3885 3396 3915
rect 3364 3884 3396 3885
rect 3364 3835 3396 3836
rect 3364 3805 3365 3835
rect 3365 3805 3395 3835
rect 3395 3805 3396 3835
rect 3364 3804 3396 3805
rect 3364 3755 3396 3756
rect 3364 3725 3365 3755
rect 3365 3725 3395 3755
rect 3395 3725 3396 3755
rect 3364 3724 3396 3725
rect 3364 3675 3396 3676
rect 3364 3645 3365 3675
rect 3365 3645 3395 3675
rect 3395 3645 3396 3675
rect 3364 3644 3396 3645
rect 3444 4395 3476 4396
rect 3444 4365 3445 4395
rect 3445 4365 3475 4395
rect 3475 4365 3476 4395
rect 3444 4364 3476 4365
rect 3444 4284 3476 4316
rect 3444 4235 3476 4236
rect 3444 4205 3445 4235
rect 3445 4205 3475 4235
rect 3475 4205 3476 4235
rect 3444 4204 3476 4205
rect 3444 4124 3476 4156
rect 3444 4075 3476 4076
rect 3444 4045 3445 4075
rect 3445 4045 3475 4075
rect 3475 4045 3476 4075
rect 3444 4044 3476 4045
rect 3444 3995 3476 3996
rect 3444 3965 3445 3995
rect 3445 3965 3475 3995
rect 3475 3965 3476 3995
rect 3444 3964 3476 3965
rect 3444 3915 3476 3916
rect 3444 3885 3445 3915
rect 3445 3885 3475 3915
rect 3475 3885 3476 3915
rect 3444 3884 3476 3885
rect 3444 3835 3476 3836
rect 3444 3805 3445 3835
rect 3445 3805 3475 3835
rect 3475 3805 3476 3835
rect 3444 3804 3476 3805
rect 3444 3755 3476 3756
rect 3444 3725 3445 3755
rect 3445 3725 3475 3755
rect 3475 3725 3476 3755
rect 3444 3724 3476 3725
rect 3444 3675 3476 3676
rect 3444 3645 3445 3675
rect 3445 3645 3475 3675
rect 3475 3645 3476 3675
rect 3444 3644 3476 3645
rect 3524 4395 3556 4396
rect 3524 4365 3525 4395
rect 3525 4365 3555 4395
rect 3555 4365 3556 4395
rect 3524 4364 3556 4365
rect 3524 4284 3556 4316
rect 3524 4235 3556 4236
rect 3524 4205 3525 4235
rect 3525 4205 3555 4235
rect 3555 4205 3556 4235
rect 3524 4204 3556 4205
rect 3524 4124 3556 4156
rect 3524 4075 3556 4076
rect 3524 4045 3525 4075
rect 3525 4045 3555 4075
rect 3555 4045 3556 4075
rect 3524 4044 3556 4045
rect 3524 3995 3556 3996
rect 3524 3965 3525 3995
rect 3525 3965 3555 3995
rect 3555 3965 3556 3995
rect 3524 3964 3556 3965
rect 3524 3915 3556 3916
rect 3524 3885 3525 3915
rect 3525 3885 3555 3915
rect 3555 3885 3556 3915
rect 3524 3884 3556 3885
rect 3524 3835 3556 3836
rect 3524 3805 3525 3835
rect 3525 3805 3555 3835
rect 3555 3805 3556 3835
rect 3524 3804 3556 3805
rect 3524 3755 3556 3756
rect 3524 3725 3525 3755
rect 3525 3725 3555 3755
rect 3555 3725 3556 3755
rect 3524 3724 3556 3725
rect 3524 3675 3556 3676
rect 3524 3645 3525 3675
rect 3525 3645 3555 3675
rect 3555 3645 3556 3675
rect 3524 3644 3556 3645
rect 3604 4395 3636 4396
rect 3604 4365 3605 4395
rect 3605 4365 3635 4395
rect 3635 4365 3636 4395
rect 3604 4364 3636 4365
rect 3604 4284 3636 4316
rect 3604 4235 3636 4236
rect 3604 4205 3605 4235
rect 3605 4205 3635 4235
rect 3635 4205 3636 4235
rect 3604 4204 3636 4205
rect 3604 4124 3636 4156
rect 3604 4075 3636 4076
rect 3604 4045 3605 4075
rect 3605 4045 3635 4075
rect 3635 4045 3636 4075
rect 3604 4044 3636 4045
rect 3604 3995 3636 3996
rect 3604 3965 3605 3995
rect 3605 3965 3635 3995
rect 3635 3965 3636 3995
rect 3604 3964 3636 3965
rect 3604 3915 3636 3916
rect 3604 3885 3605 3915
rect 3605 3885 3635 3915
rect 3635 3885 3636 3915
rect 3604 3884 3636 3885
rect 3604 3835 3636 3836
rect 3604 3805 3605 3835
rect 3605 3805 3635 3835
rect 3635 3805 3636 3835
rect 3604 3804 3636 3805
rect 3604 3755 3636 3756
rect 3604 3725 3605 3755
rect 3605 3725 3635 3755
rect 3635 3725 3636 3755
rect 3604 3724 3636 3725
rect 3604 3675 3636 3676
rect 3604 3645 3605 3675
rect 3605 3645 3635 3675
rect 3635 3645 3636 3675
rect 3604 3644 3636 3645
rect 3684 4395 3716 4396
rect 3684 4365 3685 4395
rect 3685 4365 3715 4395
rect 3715 4365 3716 4395
rect 3684 4364 3716 4365
rect 3684 4284 3716 4316
rect 3684 4235 3716 4236
rect 3684 4205 3685 4235
rect 3685 4205 3715 4235
rect 3715 4205 3716 4235
rect 3684 4204 3716 4205
rect 3684 4124 3716 4156
rect 3684 4075 3716 4076
rect 3684 4045 3685 4075
rect 3685 4045 3715 4075
rect 3715 4045 3716 4075
rect 3684 4044 3716 4045
rect 3684 3995 3716 3996
rect 3684 3965 3685 3995
rect 3685 3965 3715 3995
rect 3715 3965 3716 3995
rect 3684 3964 3716 3965
rect 3684 3915 3716 3916
rect 3684 3885 3685 3915
rect 3685 3885 3715 3915
rect 3715 3885 3716 3915
rect 3684 3884 3716 3885
rect 3684 3835 3716 3836
rect 3684 3805 3685 3835
rect 3685 3805 3715 3835
rect 3715 3805 3716 3835
rect 3684 3804 3716 3805
rect 3684 3755 3716 3756
rect 3684 3725 3685 3755
rect 3685 3725 3715 3755
rect 3715 3725 3716 3755
rect 3684 3724 3716 3725
rect 3684 3675 3716 3676
rect 3684 3645 3685 3675
rect 3685 3645 3715 3675
rect 3715 3645 3716 3675
rect 3684 3644 3716 3645
rect 3764 4395 3796 4396
rect 3764 4365 3765 4395
rect 3765 4365 3795 4395
rect 3795 4365 3796 4395
rect 3764 4364 3796 4365
rect 3764 4284 3796 4316
rect 3764 4235 3796 4236
rect 3764 4205 3765 4235
rect 3765 4205 3795 4235
rect 3795 4205 3796 4235
rect 3764 4204 3796 4205
rect 3764 4124 3796 4156
rect 3764 4075 3796 4076
rect 3764 4045 3765 4075
rect 3765 4045 3795 4075
rect 3795 4045 3796 4075
rect 3764 4044 3796 4045
rect 3764 3995 3796 3996
rect 3764 3965 3765 3995
rect 3765 3965 3795 3995
rect 3795 3965 3796 3995
rect 3764 3964 3796 3965
rect 3764 3915 3796 3916
rect 3764 3885 3765 3915
rect 3765 3885 3795 3915
rect 3795 3885 3796 3915
rect 3764 3884 3796 3885
rect 3764 3835 3796 3836
rect 3764 3805 3765 3835
rect 3765 3805 3795 3835
rect 3795 3805 3796 3835
rect 3764 3804 3796 3805
rect 3764 3755 3796 3756
rect 3764 3725 3765 3755
rect 3765 3725 3795 3755
rect 3795 3725 3796 3755
rect 3764 3724 3796 3725
rect 3764 3675 3796 3676
rect 3764 3645 3765 3675
rect 3765 3645 3795 3675
rect 3795 3645 3796 3675
rect 3764 3644 3796 3645
rect 3844 4395 3876 4396
rect 3844 4365 3845 4395
rect 3845 4365 3875 4395
rect 3875 4365 3876 4395
rect 3844 4364 3876 4365
rect 3844 4284 3876 4316
rect 3844 4235 3876 4236
rect 3844 4205 3845 4235
rect 3845 4205 3875 4235
rect 3875 4205 3876 4235
rect 3844 4204 3876 4205
rect 3844 4124 3876 4156
rect 3844 4075 3876 4076
rect 3844 4045 3845 4075
rect 3845 4045 3875 4075
rect 3875 4045 3876 4075
rect 3844 4044 3876 4045
rect 3844 3995 3876 3996
rect 3844 3965 3845 3995
rect 3845 3965 3875 3995
rect 3875 3965 3876 3995
rect 3844 3964 3876 3965
rect 3844 3915 3876 3916
rect 3844 3885 3845 3915
rect 3845 3885 3875 3915
rect 3875 3885 3876 3915
rect 3844 3884 3876 3885
rect 3844 3835 3876 3836
rect 3844 3805 3845 3835
rect 3845 3805 3875 3835
rect 3875 3805 3876 3835
rect 3844 3804 3876 3805
rect 3844 3755 3876 3756
rect 3844 3725 3845 3755
rect 3845 3725 3875 3755
rect 3875 3725 3876 3755
rect 3844 3724 3876 3725
rect 3844 3675 3876 3676
rect 3844 3645 3845 3675
rect 3845 3645 3875 3675
rect 3875 3645 3876 3675
rect 3844 3644 3876 3645
rect 3924 4395 3956 4396
rect 3924 4365 3925 4395
rect 3925 4365 3955 4395
rect 3955 4365 3956 4395
rect 3924 4364 3956 4365
rect 3924 4284 3956 4316
rect 3924 4235 3956 4236
rect 3924 4205 3925 4235
rect 3925 4205 3955 4235
rect 3955 4205 3956 4235
rect 3924 4204 3956 4205
rect 3924 4124 3956 4156
rect 3924 4075 3956 4076
rect 3924 4045 3925 4075
rect 3925 4045 3955 4075
rect 3955 4045 3956 4075
rect 3924 4044 3956 4045
rect 3924 3995 3956 3996
rect 3924 3965 3925 3995
rect 3925 3965 3955 3995
rect 3955 3965 3956 3995
rect 3924 3964 3956 3965
rect 3924 3915 3956 3916
rect 3924 3885 3925 3915
rect 3925 3885 3955 3915
rect 3955 3885 3956 3915
rect 3924 3884 3956 3885
rect 3924 3835 3956 3836
rect 3924 3805 3925 3835
rect 3925 3805 3955 3835
rect 3955 3805 3956 3835
rect 3924 3804 3956 3805
rect 3924 3755 3956 3756
rect 3924 3725 3925 3755
rect 3925 3725 3955 3755
rect 3955 3725 3956 3755
rect 3924 3724 3956 3725
rect 3924 3675 3956 3676
rect 3924 3645 3925 3675
rect 3925 3645 3955 3675
rect 3955 3645 3956 3675
rect 3924 3644 3956 3645
rect 4004 4395 4036 4396
rect 4004 4365 4005 4395
rect 4005 4365 4035 4395
rect 4035 4365 4036 4395
rect 4004 4364 4036 4365
rect 4004 4284 4036 4316
rect 4004 4235 4036 4236
rect 4004 4205 4005 4235
rect 4005 4205 4035 4235
rect 4035 4205 4036 4235
rect 4004 4204 4036 4205
rect 4004 4124 4036 4156
rect 4004 4075 4036 4076
rect 4004 4045 4005 4075
rect 4005 4045 4035 4075
rect 4035 4045 4036 4075
rect 4004 4044 4036 4045
rect 4004 3995 4036 3996
rect 4004 3965 4005 3995
rect 4005 3965 4035 3995
rect 4035 3965 4036 3995
rect 4004 3964 4036 3965
rect 4004 3915 4036 3916
rect 4004 3885 4005 3915
rect 4005 3885 4035 3915
rect 4035 3885 4036 3915
rect 4004 3884 4036 3885
rect 4004 3835 4036 3836
rect 4004 3805 4005 3835
rect 4005 3805 4035 3835
rect 4035 3805 4036 3835
rect 4004 3804 4036 3805
rect 4004 3755 4036 3756
rect 4004 3725 4005 3755
rect 4005 3725 4035 3755
rect 4035 3725 4036 3755
rect 4004 3724 4036 3725
rect 4004 3675 4036 3676
rect 4004 3645 4005 3675
rect 4005 3645 4035 3675
rect 4035 3645 4036 3675
rect 4004 3644 4036 3645
rect 4084 4395 4116 4396
rect 4084 4365 4085 4395
rect 4085 4365 4115 4395
rect 4115 4365 4116 4395
rect 4084 4364 4116 4365
rect 4084 4284 4116 4316
rect 4084 4235 4116 4236
rect 4084 4205 4085 4235
rect 4085 4205 4115 4235
rect 4115 4205 4116 4235
rect 4084 4204 4116 4205
rect 4084 4124 4116 4156
rect 4084 4075 4116 4076
rect 4084 4045 4085 4075
rect 4085 4045 4115 4075
rect 4115 4045 4116 4075
rect 4084 4044 4116 4045
rect 4084 3995 4116 3996
rect 4084 3965 4085 3995
rect 4085 3965 4115 3995
rect 4115 3965 4116 3995
rect 4084 3964 4116 3965
rect 4084 3915 4116 3916
rect 4084 3885 4085 3915
rect 4085 3885 4115 3915
rect 4115 3885 4116 3915
rect 4084 3884 4116 3885
rect 4084 3835 4116 3836
rect 4084 3805 4085 3835
rect 4085 3805 4115 3835
rect 4115 3805 4116 3835
rect 4084 3804 4116 3805
rect 4084 3755 4116 3756
rect 4084 3725 4085 3755
rect 4085 3725 4115 3755
rect 4115 3725 4116 3755
rect 4084 3724 4116 3725
rect 4084 3675 4116 3676
rect 4084 3645 4085 3675
rect 4085 3645 4115 3675
rect 4115 3645 4116 3675
rect 4084 3644 4116 3645
rect 4164 4395 4196 4396
rect 4164 4365 4165 4395
rect 4165 4365 4195 4395
rect 4195 4365 4196 4395
rect 4164 4364 4196 4365
rect 4164 4284 4196 4316
rect 4164 4235 4196 4236
rect 4164 4205 4165 4235
rect 4165 4205 4195 4235
rect 4195 4205 4196 4235
rect 4164 4204 4196 4205
rect 4164 4124 4196 4156
rect 4164 4075 4196 4076
rect 4164 4045 4165 4075
rect 4165 4045 4195 4075
rect 4195 4045 4196 4075
rect 4164 4044 4196 4045
rect 4164 3995 4196 3996
rect 4164 3965 4165 3995
rect 4165 3965 4195 3995
rect 4195 3965 4196 3995
rect 4164 3964 4196 3965
rect 4164 3915 4196 3916
rect 4164 3885 4165 3915
rect 4165 3885 4195 3915
rect 4195 3885 4196 3915
rect 4164 3884 4196 3885
rect 4164 3835 4196 3836
rect 4164 3805 4165 3835
rect 4165 3805 4195 3835
rect 4195 3805 4196 3835
rect 4164 3804 4196 3805
rect 4164 3755 4196 3756
rect 4164 3725 4165 3755
rect 4165 3725 4195 3755
rect 4195 3725 4196 3755
rect 4164 3724 4196 3725
rect 4164 3675 4196 3676
rect 4164 3645 4165 3675
rect 4165 3645 4195 3675
rect 4195 3645 4196 3675
rect 4164 3644 4196 3645
rect 4244 4395 4276 4396
rect 4244 4365 4245 4395
rect 4245 4365 4275 4395
rect 4275 4365 4276 4395
rect 4244 4364 4276 4365
rect 4244 4284 4276 4316
rect 4244 4235 4276 4236
rect 4244 4205 4245 4235
rect 4245 4205 4275 4235
rect 4275 4205 4276 4235
rect 4244 4204 4276 4205
rect 4244 4124 4276 4156
rect 4244 4075 4276 4076
rect 4244 4045 4245 4075
rect 4245 4045 4275 4075
rect 4275 4045 4276 4075
rect 4244 4044 4276 4045
rect 4244 3995 4276 3996
rect 4244 3965 4245 3995
rect 4245 3965 4275 3995
rect 4275 3965 4276 3995
rect 4244 3964 4276 3965
rect 4244 3915 4276 3916
rect 4244 3885 4245 3915
rect 4245 3885 4275 3915
rect 4275 3885 4276 3915
rect 4244 3884 4276 3885
rect 4244 3835 4276 3836
rect 4244 3805 4245 3835
rect 4245 3805 4275 3835
rect 4275 3805 4276 3835
rect 4244 3804 4276 3805
rect 4244 3755 4276 3756
rect 4244 3725 4245 3755
rect 4245 3725 4275 3755
rect 4275 3725 4276 3755
rect 4244 3724 4276 3725
rect 4244 3675 4276 3676
rect 4244 3645 4245 3675
rect 4245 3645 4275 3675
rect 4275 3645 4276 3675
rect 4244 3644 4276 3645
rect 4324 4395 4356 4396
rect 4324 4365 4325 4395
rect 4325 4365 4355 4395
rect 4355 4365 4356 4395
rect 4324 4364 4356 4365
rect 4324 4284 4356 4316
rect 4324 4235 4356 4236
rect 4324 4205 4325 4235
rect 4325 4205 4355 4235
rect 4355 4205 4356 4235
rect 4324 4204 4356 4205
rect 4324 4124 4356 4156
rect 4324 4075 4356 4076
rect 4324 4045 4325 4075
rect 4325 4045 4355 4075
rect 4355 4045 4356 4075
rect 4324 4044 4356 4045
rect 4324 3995 4356 3996
rect 4324 3965 4325 3995
rect 4325 3965 4355 3995
rect 4355 3965 4356 3995
rect 4324 3964 4356 3965
rect 4324 3915 4356 3916
rect 4324 3885 4325 3915
rect 4325 3885 4355 3915
rect 4355 3885 4356 3915
rect 4324 3884 4356 3885
rect 4324 3835 4356 3836
rect 4324 3805 4325 3835
rect 4325 3805 4355 3835
rect 4355 3805 4356 3835
rect 4324 3804 4356 3805
rect 4324 3755 4356 3756
rect 4324 3725 4325 3755
rect 4325 3725 4355 3755
rect 4355 3725 4356 3755
rect 4324 3724 4356 3725
rect 4324 3675 4356 3676
rect 4324 3645 4325 3675
rect 4325 3645 4355 3675
rect 4355 3645 4356 3675
rect 4324 3644 4356 3645
rect 4404 4395 4436 4396
rect 4404 4365 4405 4395
rect 4405 4365 4435 4395
rect 4435 4365 4436 4395
rect 4404 4364 4436 4365
rect 4404 4284 4436 4316
rect 4404 4235 4436 4236
rect 4404 4205 4405 4235
rect 4405 4205 4435 4235
rect 4435 4205 4436 4235
rect 4404 4204 4436 4205
rect 4404 4124 4436 4156
rect 4404 4075 4436 4076
rect 4404 4045 4405 4075
rect 4405 4045 4435 4075
rect 4435 4045 4436 4075
rect 4404 4044 4436 4045
rect 4404 3995 4436 3996
rect 4404 3965 4405 3995
rect 4405 3965 4435 3995
rect 4435 3965 4436 3995
rect 4404 3964 4436 3965
rect 4404 3915 4436 3916
rect 4404 3885 4405 3915
rect 4405 3885 4435 3915
rect 4435 3885 4436 3915
rect 4404 3884 4436 3885
rect 4404 3835 4436 3836
rect 4404 3805 4405 3835
rect 4405 3805 4435 3835
rect 4435 3805 4436 3835
rect 4404 3804 4436 3805
rect 4404 3755 4436 3756
rect 4404 3725 4405 3755
rect 4405 3725 4435 3755
rect 4435 3725 4436 3755
rect 4404 3724 4436 3725
rect 4404 3675 4436 3676
rect 4404 3645 4405 3675
rect 4405 3645 4435 3675
rect 4435 3645 4436 3675
rect 4404 3644 4436 3645
rect 4484 4395 4516 4396
rect 4484 4365 4485 4395
rect 4485 4365 4515 4395
rect 4515 4365 4516 4395
rect 4484 4364 4516 4365
rect 4484 4284 4516 4316
rect 4484 4235 4516 4236
rect 4484 4205 4485 4235
rect 4485 4205 4515 4235
rect 4515 4205 4516 4235
rect 4484 4204 4516 4205
rect 4484 4124 4516 4156
rect 4484 4075 4516 4076
rect 4484 4045 4485 4075
rect 4485 4045 4515 4075
rect 4515 4045 4516 4075
rect 4484 4044 4516 4045
rect 4484 3995 4516 3996
rect 4484 3965 4485 3995
rect 4485 3965 4515 3995
rect 4515 3965 4516 3995
rect 4484 3964 4516 3965
rect 4484 3915 4516 3916
rect 4484 3885 4485 3915
rect 4485 3885 4515 3915
rect 4515 3885 4516 3915
rect 4484 3884 4516 3885
rect 4484 3835 4516 3836
rect 4484 3805 4485 3835
rect 4485 3805 4515 3835
rect 4515 3805 4516 3835
rect 4484 3804 4516 3805
rect 4484 3755 4516 3756
rect 4484 3725 4485 3755
rect 4485 3725 4515 3755
rect 4515 3725 4516 3755
rect 4484 3724 4516 3725
rect 4484 3675 4516 3676
rect 4484 3645 4485 3675
rect 4485 3645 4515 3675
rect 4515 3645 4516 3675
rect 4484 3644 4516 3645
rect 4564 4395 4596 4396
rect 4564 4365 4565 4395
rect 4565 4365 4595 4395
rect 4595 4365 4596 4395
rect 4564 4364 4596 4365
rect 4564 4284 4596 4316
rect 4564 4235 4596 4236
rect 4564 4205 4565 4235
rect 4565 4205 4595 4235
rect 4595 4205 4596 4235
rect 4564 4204 4596 4205
rect 4564 4124 4596 4156
rect 4564 4075 4596 4076
rect 4564 4045 4565 4075
rect 4565 4045 4595 4075
rect 4595 4045 4596 4075
rect 4564 4044 4596 4045
rect 4564 3995 4596 3996
rect 4564 3965 4565 3995
rect 4565 3965 4595 3995
rect 4595 3965 4596 3995
rect 4564 3964 4596 3965
rect 4564 3915 4596 3916
rect 4564 3885 4565 3915
rect 4565 3885 4595 3915
rect 4595 3885 4596 3915
rect 4564 3884 4596 3885
rect 4564 3835 4596 3836
rect 4564 3805 4565 3835
rect 4565 3805 4595 3835
rect 4595 3805 4596 3835
rect 4564 3804 4596 3805
rect 4564 3755 4596 3756
rect 4564 3725 4565 3755
rect 4565 3725 4595 3755
rect 4595 3725 4596 3755
rect 4564 3724 4596 3725
rect 4564 3675 4596 3676
rect 4564 3645 4565 3675
rect 4565 3645 4595 3675
rect 4595 3645 4596 3675
rect 4564 3644 4596 3645
rect 4644 4395 4676 4396
rect 4644 4365 4645 4395
rect 4645 4365 4675 4395
rect 4675 4365 4676 4395
rect 4644 4364 4676 4365
rect 4644 4284 4676 4316
rect 4644 4235 4676 4236
rect 4644 4205 4645 4235
rect 4645 4205 4675 4235
rect 4675 4205 4676 4235
rect 4644 4204 4676 4205
rect 4644 4124 4676 4156
rect 4644 4075 4676 4076
rect 4644 4045 4645 4075
rect 4645 4045 4675 4075
rect 4675 4045 4676 4075
rect 4644 4044 4676 4045
rect 4644 3995 4676 3996
rect 4644 3965 4645 3995
rect 4645 3965 4675 3995
rect 4675 3965 4676 3995
rect 4644 3964 4676 3965
rect 4644 3915 4676 3916
rect 4644 3885 4645 3915
rect 4645 3885 4675 3915
rect 4675 3885 4676 3915
rect 4644 3884 4676 3885
rect 4644 3835 4676 3836
rect 4644 3805 4645 3835
rect 4645 3805 4675 3835
rect 4675 3805 4676 3835
rect 4644 3804 4676 3805
rect 4644 3755 4676 3756
rect 4644 3725 4645 3755
rect 4645 3725 4675 3755
rect 4675 3725 4676 3755
rect 4644 3724 4676 3725
rect 4644 3675 4676 3676
rect 4644 3645 4645 3675
rect 4645 3645 4675 3675
rect 4675 3645 4676 3675
rect 4644 3644 4676 3645
rect 4724 4395 4756 4396
rect 4724 4365 4725 4395
rect 4725 4365 4755 4395
rect 4755 4365 4756 4395
rect 4724 4364 4756 4365
rect 4724 4284 4756 4316
rect 4724 4235 4756 4236
rect 4724 4205 4725 4235
rect 4725 4205 4755 4235
rect 4755 4205 4756 4235
rect 4724 4204 4756 4205
rect 4724 4124 4756 4156
rect 4724 4075 4756 4076
rect 4724 4045 4725 4075
rect 4725 4045 4755 4075
rect 4755 4045 4756 4075
rect 4724 4044 4756 4045
rect 4724 3995 4756 3996
rect 4724 3965 4725 3995
rect 4725 3965 4755 3995
rect 4755 3965 4756 3995
rect 4724 3964 4756 3965
rect 4724 3915 4756 3916
rect 4724 3885 4725 3915
rect 4725 3885 4755 3915
rect 4755 3885 4756 3915
rect 4724 3884 4756 3885
rect 4724 3835 4756 3836
rect 4724 3805 4725 3835
rect 4725 3805 4755 3835
rect 4755 3805 4756 3835
rect 4724 3804 4756 3805
rect 4724 3755 4756 3756
rect 4724 3725 4725 3755
rect 4725 3725 4755 3755
rect 4755 3725 4756 3755
rect 4724 3724 4756 3725
rect 4724 3675 4756 3676
rect 4724 3645 4725 3675
rect 4725 3645 4755 3675
rect 4755 3645 4756 3675
rect 4724 3644 4756 3645
rect 4804 4395 4836 4396
rect 4804 4365 4805 4395
rect 4805 4365 4835 4395
rect 4835 4365 4836 4395
rect 4804 4364 4836 4365
rect 4804 4284 4836 4316
rect 4804 4235 4836 4236
rect 4804 4205 4805 4235
rect 4805 4205 4835 4235
rect 4835 4205 4836 4235
rect 4804 4204 4836 4205
rect 4804 4124 4836 4156
rect 4804 4075 4836 4076
rect 4804 4045 4805 4075
rect 4805 4045 4835 4075
rect 4835 4045 4836 4075
rect 4804 4044 4836 4045
rect 4804 3995 4836 3996
rect 4804 3965 4805 3995
rect 4805 3965 4835 3995
rect 4835 3965 4836 3995
rect 4804 3964 4836 3965
rect 4804 3915 4836 3916
rect 4804 3885 4805 3915
rect 4805 3885 4835 3915
rect 4835 3885 4836 3915
rect 4804 3884 4836 3885
rect 4804 3835 4836 3836
rect 4804 3805 4805 3835
rect 4805 3805 4835 3835
rect 4835 3805 4836 3835
rect 4804 3804 4836 3805
rect 4804 3755 4836 3756
rect 4804 3725 4805 3755
rect 4805 3725 4835 3755
rect 4835 3725 4836 3755
rect 4804 3724 4836 3725
rect 4804 3675 4836 3676
rect 4804 3645 4805 3675
rect 4805 3645 4835 3675
rect 4835 3645 4836 3675
rect 4804 3644 4836 3645
rect 4884 4395 4916 4396
rect 4884 4365 4885 4395
rect 4885 4365 4915 4395
rect 4915 4365 4916 4395
rect 4884 4364 4916 4365
rect 4884 4284 4916 4316
rect 4884 4235 4916 4236
rect 4884 4205 4885 4235
rect 4885 4205 4915 4235
rect 4915 4205 4916 4235
rect 4884 4204 4916 4205
rect 4884 4124 4916 4156
rect 4884 4075 4916 4076
rect 4884 4045 4885 4075
rect 4885 4045 4915 4075
rect 4915 4045 4916 4075
rect 4884 4044 4916 4045
rect 4884 3995 4916 3996
rect 4884 3965 4885 3995
rect 4885 3965 4915 3995
rect 4915 3965 4916 3995
rect 4884 3964 4916 3965
rect 4884 3915 4916 3916
rect 4884 3885 4885 3915
rect 4885 3885 4915 3915
rect 4915 3885 4916 3915
rect 4884 3884 4916 3885
rect 4884 3835 4916 3836
rect 4884 3805 4885 3835
rect 4885 3805 4915 3835
rect 4915 3805 4916 3835
rect 4884 3804 4916 3805
rect 4884 3755 4916 3756
rect 4884 3725 4885 3755
rect 4885 3725 4915 3755
rect 4915 3725 4916 3755
rect 4884 3724 4916 3725
rect 4884 3675 4916 3676
rect 4884 3645 4885 3675
rect 4885 3645 4915 3675
rect 4915 3645 4916 3675
rect 4884 3644 4916 3645
rect -876 3595 -844 3596
rect -876 3565 -875 3595
rect -875 3565 -845 3595
rect -845 3565 -844 3595
rect -876 3564 -844 3565
rect -876 3515 -844 3516
rect -876 3485 -875 3515
rect -875 3485 -845 3515
rect -845 3485 -844 3515
rect -876 3484 -844 3485
rect -876 3404 -844 3436
rect -876 3355 -844 3356
rect -876 3325 -875 3355
rect -875 3325 -845 3355
rect -845 3325 -844 3355
rect -876 3324 -844 3325
rect -876 3275 -844 3276
rect -876 3245 -875 3275
rect -875 3245 -845 3275
rect -845 3245 -844 3275
rect -876 3244 -844 3245
rect -876 3195 -844 3196
rect -876 3165 -875 3195
rect -875 3165 -845 3195
rect -845 3165 -844 3195
rect -876 3164 -844 3165
rect -876 3115 -844 3116
rect -876 3085 -875 3115
rect -875 3085 -845 3115
rect -845 3085 -844 3115
rect -876 3084 -844 3085
rect -876 3004 -844 3036
rect -876 2955 -844 2956
rect -876 2925 -875 2955
rect -875 2925 -845 2955
rect -845 2925 -844 2955
rect -876 2924 -844 2925
rect -876 2844 -844 2876
rect -876 2795 -844 2796
rect -876 2765 -875 2795
rect -875 2765 -845 2795
rect -845 2765 -844 2795
rect -876 2764 -844 2765
rect -876 2715 -844 2716
rect -876 2685 -875 2715
rect -875 2685 -845 2715
rect -845 2685 -844 2715
rect -876 2684 -844 2685
rect -876 2604 -844 2636
rect -876 2555 -844 2556
rect -876 2525 -875 2555
rect -875 2525 -845 2555
rect -845 2525 -844 2555
rect -876 2524 -844 2525
rect -796 3595 -764 3596
rect -796 3565 -795 3595
rect -795 3565 -765 3595
rect -765 3565 -764 3595
rect -796 3564 -764 3565
rect -796 3515 -764 3516
rect -796 3485 -795 3515
rect -795 3485 -765 3515
rect -765 3485 -764 3515
rect -796 3484 -764 3485
rect -796 3404 -764 3436
rect -796 3355 -764 3356
rect -796 3325 -795 3355
rect -795 3325 -765 3355
rect -765 3325 -764 3355
rect -796 3324 -764 3325
rect -796 3275 -764 3276
rect -796 3245 -795 3275
rect -795 3245 -765 3275
rect -765 3245 -764 3275
rect -796 3244 -764 3245
rect -796 3195 -764 3196
rect -796 3165 -795 3195
rect -795 3165 -765 3195
rect -765 3165 -764 3195
rect -796 3164 -764 3165
rect -796 3115 -764 3116
rect -796 3085 -795 3115
rect -795 3085 -765 3115
rect -765 3085 -764 3115
rect -796 3084 -764 3085
rect -796 3004 -764 3036
rect -796 2955 -764 2956
rect -796 2925 -795 2955
rect -795 2925 -765 2955
rect -765 2925 -764 2955
rect -796 2924 -764 2925
rect -796 2844 -764 2876
rect -796 2795 -764 2796
rect -796 2765 -795 2795
rect -795 2765 -765 2795
rect -765 2765 -764 2795
rect -796 2764 -764 2765
rect -796 2715 -764 2716
rect -796 2685 -795 2715
rect -795 2685 -765 2715
rect -765 2685 -764 2715
rect -796 2684 -764 2685
rect -796 2604 -764 2636
rect -796 2555 -764 2556
rect -796 2525 -795 2555
rect -795 2525 -765 2555
rect -765 2525 -764 2555
rect -796 2524 -764 2525
rect -716 3595 -684 3596
rect -716 3565 -715 3595
rect -715 3565 -685 3595
rect -685 3565 -684 3595
rect -716 3564 -684 3565
rect -716 3515 -684 3516
rect -716 3485 -715 3515
rect -715 3485 -685 3515
rect -685 3485 -684 3515
rect -716 3484 -684 3485
rect -716 3404 -684 3436
rect -716 3355 -684 3356
rect -716 3325 -715 3355
rect -715 3325 -685 3355
rect -685 3325 -684 3355
rect -716 3324 -684 3325
rect -716 3275 -684 3276
rect -716 3245 -715 3275
rect -715 3245 -685 3275
rect -685 3245 -684 3275
rect -716 3244 -684 3245
rect -716 3195 -684 3196
rect -716 3165 -715 3195
rect -715 3165 -685 3195
rect -685 3165 -684 3195
rect -716 3164 -684 3165
rect -716 3115 -684 3116
rect -716 3085 -715 3115
rect -715 3085 -685 3115
rect -685 3085 -684 3115
rect -716 3084 -684 3085
rect -716 3004 -684 3036
rect -716 2955 -684 2956
rect -716 2925 -715 2955
rect -715 2925 -685 2955
rect -685 2925 -684 2955
rect -716 2924 -684 2925
rect -716 2844 -684 2876
rect -716 2795 -684 2796
rect -716 2765 -715 2795
rect -715 2765 -685 2795
rect -685 2765 -684 2795
rect -716 2764 -684 2765
rect -716 2715 -684 2716
rect -716 2685 -715 2715
rect -715 2685 -685 2715
rect -685 2685 -684 2715
rect -716 2684 -684 2685
rect -716 2604 -684 2636
rect -716 2555 -684 2556
rect -716 2525 -715 2555
rect -715 2525 -685 2555
rect -685 2525 -684 2555
rect -716 2524 -684 2525
rect -636 3595 -604 3596
rect -636 3565 -635 3595
rect -635 3565 -605 3595
rect -605 3565 -604 3595
rect -636 3564 -604 3565
rect -636 3515 -604 3516
rect -636 3485 -635 3515
rect -635 3485 -605 3515
rect -605 3485 -604 3515
rect -636 3484 -604 3485
rect -636 3404 -604 3436
rect -636 3355 -604 3356
rect -636 3325 -635 3355
rect -635 3325 -605 3355
rect -605 3325 -604 3355
rect -636 3324 -604 3325
rect -636 3275 -604 3276
rect -636 3245 -635 3275
rect -635 3245 -605 3275
rect -605 3245 -604 3275
rect -636 3244 -604 3245
rect -636 3195 -604 3196
rect -636 3165 -635 3195
rect -635 3165 -605 3195
rect -605 3165 -604 3195
rect -636 3164 -604 3165
rect -636 3115 -604 3116
rect -636 3085 -635 3115
rect -635 3085 -605 3115
rect -605 3085 -604 3115
rect -636 3084 -604 3085
rect -636 3004 -604 3036
rect -636 2955 -604 2956
rect -636 2925 -635 2955
rect -635 2925 -605 2955
rect -605 2925 -604 2955
rect -636 2924 -604 2925
rect -636 2844 -604 2876
rect -636 2795 -604 2796
rect -636 2765 -635 2795
rect -635 2765 -605 2795
rect -605 2765 -604 2795
rect -636 2764 -604 2765
rect -636 2715 -604 2716
rect -636 2685 -635 2715
rect -635 2685 -605 2715
rect -605 2685 -604 2715
rect -636 2684 -604 2685
rect -636 2604 -604 2636
rect -636 2555 -604 2556
rect -636 2525 -635 2555
rect -635 2525 -605 2555
rect -605 2525 -604 2555
rect -636 2524 -604 2525
rect -556 3595 -524 3596
rect -556 3565 -555 3595
rect -555 3565 -525 3595
rect -525 3565 -524 3595
rect -556 3564 -524 3565
rect -556 3515 -524 3516
rect -556 3485 -555 3515
rect -555 3485 -525 3515
rect -525 3485 -524 3515
rect -556 3484 -524 3485
rect -556 3404 -524 3436
rect -556 3355 -524 3356
rect -556 3325 -555 3355
rect -555 3325 -525 3355
rect -525 3325 -524 3355
rect -556 3324 -524 3325
rect -556 3275 -524 3276
rect -556 3245 -555 3275
rect -555 3245 -525 3275
rect -525 3245 -524 3275
rect -556 3244 -524 3245
rect -556 3195 -524 3196
rect -556 3165 -555 3195
rect -555 3165 -525 3195
rect -525 3165 -524 3195
rect -556 3164 -524 3165
rect -556 3115 -524 3116
rect -556 3085 -555 3115
rect -555 3085 -525 3115
rect -525 3085 -524 3115
rect -556 3084 -524 3085
rect -556 3004 -524 3036
rect -556 2955 -524 2956
rect -556 2925 -555 2955
rect -555 2925 -525 2955
rect -525 2925 -524 2955
rect -556 2924 -524 2925
rect -556 2844 -524 2876
rect -556 2795 -524 2796
rect -556 2765 -555 2795
rect -555 2765 -525 2795
rect -525 2765 -524 2795
rect -556 2764 -524 2765
rect -556 2715 -524 2716
rect -556 2685 -555 2715
rect -555 2685 -525 2715
rect -525 2685 -524 2715
rect -556 2684 -524 2685
rect -556 2604 -524 2636
rect -556 2555 -524 2556
rect -556 2525 -555 2555
rect -555 2525 -525 2555
rect -525 2525 -524 2555
rect -556 2524 -524 2525
rect -476 3595 -444 3596
rect -476 3565 -475 3595
rect -475 3565 -445 3595
rect -445 3565 -444 3595
rect -476 3564 -444 3565
rect -476 3515 -444 3516
rect -476 3485 -475 3515
rect -475 3485 -445 3515
rect -445 3485 -444 3515
rect -476 3484 -444 3485
rect -476 3404 -444 3436
rect -476 3355 -444 3356
rect -476 3325 -475 3355
rect -475 3325 -445 3355
rect -445 3325 -444 3355
rect -476 3324 -444 3325
rect -476 3275 -444 3276
rect -476 3245 -475 3275
rect -475 3245 -445 3275
rect -445 3245 -444 3275
rect -476 3244 -444 3245
rect -476 3195 -444 3196
rect -476 3165 -475 3195
rect -475 3165 -445 3195
rect -445 3165 -444 3195
rect -476 3164 -444 3165
rect -476 3115 -444 3116
rect -476 3085 -475 3115
rect -475 3085 -445 3115
rect -445 3085 -444 3115
rect -476 3084 -444 3085
rect -476 3004 -444 3036
rect -476 2955 -444 2956
rect -476 2925 -475 2955
rect -475 2925 -445 2955
rect -445 2925 -444 2955
rect -476 2924 -444 2925
rect -476 2844 -444 2876
rect -476 2795 -444 2796
rect -476 2765 -475 2795
rect -475 2765 -445 2795
rect -445 2765 -444 2795
rect -476 2764 -444 2765
rect -476 2715 -444 2716
rect -476 2685 -475 2715
rect -475 2685 -445 2715
rect -445 2685 -444 2715
rect -476 2684 -444 2685
rect -476 2604 -444 2636
rect -476 2555 -444 2556
rect -476 2525 -475 2555
rect -475 2525 -445 2555
rect -445 2525 -444 2555
rect -476 2524 -444 2525
rect -396 3595 -364 3596
rect -396 3565 -395 3595
rect -395 3565 -365 3595
rect -365 3565 -364 3595
rect -396 3564 -364 3565
rect -396 3515 -364 3516
rect -396 3485 -395 3515
rect -395 3485 -365 3515
rect -365 3485 -364 3515
rect -396 3484 -364 3485
rect -396 3404 -364 3436
rect -396 3355 -364 3356
rect -396 3325 -395 3355
rect -395 3325 -365 3355
rect -365 3325 -364 3355
rect -396 3324 -364 3325
rect -396 3275 -364 3276
rect -396 3245 -395 3275
rect -395 3245 -365 3275
rect -365 3245 -364 3275
rect -396 3244 -364 3245
rect -396 3195 -364 3196
rect -396 3165 -395 3195
rect -395 3165 -365 3195
rect -365 3165 -364 3195
rect -396 3164 -364 3165
rect -396 3115 -364 3116
rect -396 3085 -395 3115
rect -395 3085 -365 3115
rect -365 3085 -364 3115
rect -396 3084 -364 3085
rect -396 3004 -364 3036
rect -396 2955 -364 2956
rect -396 2925 -395 2955
rect -395 2925 -365 2955
rect -365 2925 -364 2955
rect -396 2924 -364 2925
rect -396 2844 -364 2876
rect -396 2795 -364 2796
rect -396 2765 -395 2795
rect -395 2765 -365 2795
rect -365 2765 -364 2795
rect -396 2764 -364 2765
rect -396 2715 -364 2716
rect -396 2685 -395 2715
rect -395 2685 -365 2715
rect -365 2685 -364 2715
rect -396 2684 -364 2685
rect -396 2604 -364 2636
rect -396 2555 -364 2556
rect -396 2525 -395 2555
rect -395 2525 -365 2555
rect -365 2525 -364 2555
rect -396 2524 -364 2525
rect -316 3595 -284 3596
rect -316 3565 -315 3595
rect -315 3565 -285 3595
rect -285 3565 -284 3595
rect -316 3564 -284 3565
rect -316 3515 -284 3516
rect -316 3485 -315 3515
rect -315 3485 -285 3515
rect -285 3485 -284 3515
rect -316 3484 -284 3485
rect -316 3404 -284 3436
rect -316 3355 -284 3356
rect -316 3325 -315 3355
rect -315 3325 -285 3355
rect -285 3325 -284 3355
rect -316 3324 -284 3325
rect -316 3275 -284 3276
rect -316 3245 -315 3275
rect -315 3245 -285 3275
rect -285 3245 -284 3275
rect -316 3244 -284 3245
rect -316 3195 -284 3196
rect -316 3165 -315 3195
rect -315 3165 -285 3195
rect -285 3165 -284 3195
rect -316 3164 -284 3165
rect -316 3115 -284 3116
rect -316 3085 -315 3115
rect -315 3085 -285 3115
rect -285 3085 -284 3115
rect -316 3084 -284 3085
rect -316 3004 -284 3036
rect -316 2955 -284 2956
rect -316 2925 -315 2955
rect -315 2925 -285 2955
rect -285 2925 -284 2955
rect -316 2924 -284 2925
rect -316 2844 -284 2876
rect -316 2795 -284 2796
rect -316 2765 -315 2795
rect -315 2765 -285 2795
rect -285 2765 -284 2795
rect -316 2764 -284 2765
rect -316 2715 -284 2716
rect -316 2685 -315 2715
rect -315 2685 -285 2715
rect -285 2685 -284 2715
rect -316 2684 -284 2685
rect -316 2604 -284 2636
rect -316 2555 -284 2556
rect -316 2525 -315 2555
rect -315 2525 -285 2555
rect -285 2525 -284 2555
rect -316 2524 -284 2525
rect -236 3595 -204 3596
rect -236 3565 -235 3595
rect -235 3565 -205 3595
rect -205 3565 -204 3595
rect -236 3564 -204 3565
rect -236 3515 -204 3516
rect -236 3485 -235 3515
rect -235 3485 -205 3515
rect -205 3485 -204 3515
rect -236 3484 -204 3485
rect -236 3404 -204 3436
rect -236 3355 -204 3356
rect -236 3325 -235 3355
rect -235 3325 -205 3355
rect -205 3325 -204 3355
rect -236 3324 -204 3325
rect -236 3275 -204 3276
rect -236 3245 -235 3275
rect -235 3245 -205 3275
rect -205 3245 -204 3275
rect -236 3244 -204 3245
rect -236 3195 -204 3196
rect -236 3165 -235 3195
rect -235 3165 -205 3195
rect -205 3165 -204 3195
rect -236 3164 -204 3165
rect -236 3115 -204 3116
rect -236 3085 -235 3115
rect -235 3085 -205 3115
rect -205 3085 -204 3115
rect -236 3084 -204 3085
rect -236 3004 -204 3036
rect -236 2955 -204 2956
rect -236 2925 -235 2955
rect -235 2925 -205 2955
rect -205 2925 -204 2955
rect -236 2924 -204 2925
rect -236 2844 -204 2876
rect -236 2795 -204 2796
rect -236 2765 -235 2795
rect -235 2765 -205 2795
rect -205 2765 -204 2795
rect -236 2764 -204 2765
rect -236 2715 -204 2716
rect -236 2685 -235 2715
rect -235 2685 -205 2715
rect -205 2685 -204 2715
rect -236 2684 -204 2685
rect -236 2604 -204 2636
rect -236 2555 -204 2556
rect -236 2525 -235 2555
rect -235 2525 -205 2555
rect -205 2525 -204 2555
rect -236 2524 -204 2525
rect -156 3595 -124 3596
rect -156 3565 -155 3595
rect -155 3565 -125 3595
rect -125 3565 -124 3595
rect -156 3564 -124 3565
rect -156 3515 -124 3516
rect -156 3485 -155 3515
rect -155 3485 -125 3515
rect -125 3485 -124 3515
rect -156 3484 -124 3485
rect -156 3404 -124 3436
rect -156 3355 -124 3356
rect -156 3325 -155 3355
rect -155 3325 -125 3355
rect -125 3325 -124 3355
rect -156 3324 -124 3325
rect -156 3275 -124 3276
rect -156 3245 -155 3275
rect -155 3245 -125 3275
rect -125 3245 -124 3275
rect -156 3244 -124 3245
rect -156 3195 -124 3196
rect -156 3165 -155 3195
rect -155 3165 -125 3195
rect -125 3165 -124 3195
rect -156 3164 -124 3165
rect -156 3115 -124 3116
rect -156 3085 -155 3115
rect -155 3085 -125 3115
rect -125 3085 -124 3115
rect -156 3084 -124 3085
rect -156 3004 -124 3036
rect -156 2955 -124 2956
rect -156 2925 -155 2955
rect -155 2925 -125 2955
rect -125 2925 -124 2955
rect -156 2924 -124 2925
rect -156 2844 -124 2876
rect -156 2795 -124 2796
rect -156 2765 -155 2795
rect -155 2765 -125 2795
rect -125 2765 -124 2795
rect -156 2764 -124 2765
rect -156 2715 -124 2716
rect -156 2685 -155 2715
rect -155 2685 -125 2715
rect -125 2685 -124 2715
rect -156 2684 -124 2685
rect -156 2604 -124 2636
rect -156 2555 -124 2556
rect -156 2525 -155 2555
rect -155 2525 -125 2555
rect -125 2525 -124 2555
rect -156 2524 -124 2525
rect -76 3595 -44 3596
rect -76 3565 -75 3595
rect -75 3565 -45 3595
rect -45 3565 -44 3595
rect -76 3564 -44 3565
rect -76 3515 -44 3516
rect -76 3485 -75 3515
rect -75 3485 -45 3515
rect -45 3485 -44 3515
rect -76 3484 -44 3485
rect -76 3404 -44 3436
rect -76 3355 -44 3356
rect -76 3325 -75 3355
rect -75 3325 -45 3355
rect -45 3325 -44 3355
rect -76 3324 -44 3325
rect -76 3275 -44 3276
rect -76 3245 -75 3275
rect -75 3245 -45 3275
rect -45 3245 -44 3275
rect -76 3244 -44 3245
rect -76 3195 -44 3196
rect -76 3165 -75 3195
rect -75 3165 -45 3195
rect -45 3165 -44 3195
rect -76 3164 -44 3165
rect -76 3115 -44 3116
rect -76 3085 -75 3115
rect -75 3085 -45 3115
rect -45 3085 -44 3115
rect -76 3084 -44 3085
rect -76 3004 -44 3036
rect -76 2955 -44 2956
rect -76 2925 -75 2955
rect -75 2925 -45 2955
rect -45 2925 -44 2955
rect -76 2924 -44 2925
rect -76 2844 -44 2876
rect -76 2795 -44 2796
rect -76 2765 -75 2795
rect -75 2765 -45 2795
rect -45 2765 -44 2795
rect -76 2764 -44 2765
rect -76 2715 -44 2716
rect -76 2685 -75 2715
rect -75 2685 -45 2715
rect -45 2685 -44 2715
rect -76 2684 -44 2685
rect -76 2604 -44 2636
rect -76 2555 -44 2556
rect -76 2525 -75 2555
rect -75 2525 -45 2555
rect -45 2525 -44 2555
rect -76 2524 -44 2525
rect 4 3595 36 3596
rect 4 3565 5 3595
rect 5 3565 35 3595
rect 35 3565 36 3595
rect 4 3564 36 3565
rect 4 3515 36 3516
rect 4 3485 5 3515
rect 5 3485 35 3515
rect 35 3485 36 3515
rect 4 3484 36 3485
rect 4 3404 36 3436
rect 4 3355 36 3356
rect 4 3325 5 3355
rect 5 3325 35 3355
rect 35 3325 36 3355
rect 4 3324 36 3325
rect 4 3275 36 3276
rect 4 3245 5 3275
rect 5 3245 35 3275
rect 35 3245 36 3275
rect 4 3244 36 3245
rect 4 3195 36 3196
rect 4 3165 5 3195
rect 5 3165 35 3195
rect 35 3165 36 3195
rect 4 3164 36 3165
rect 4 3115 36 3116
rect 4 3085 5 3115
rect 5 3085 35 3115
rect 35 3085 36 3115
rect 4 3084 36 3085
rect 4 3004 36 3036
rect 4 2955 36 2956
rect 4 2925 5 2955
rect 5 2925 35 2955
rect 35 2925 36 2955
rect 4 2924 36 2925
rect 4 2844 36 2876
rect 4 2795 36 2796
rect 4 2765 5 2795
rect 5 2765 35 2795
rect 35 2765 36 2795
rect 4 2764 36 2765
rect 4 2715 36 2716
rect 4 2685 5 2715
rect 5 2685 35 2715
rect 35 2685 36 2715
rect 4 2684 36 2685
rect 4 2604 36 2636
rect 4 2555 36 2556
rect 4 2525 5 2555
rect 5 2525 35 2555
rect 35 2525 36 2555
rect 4 2524 36 2525
rect 84 3595 116 3596
rect 84 3565 85 3595
rect 85 3565 115 3595
rect 115 3565 116 3595
rect 84 3564 116 3565
rect 84 3515 116 3516
rect 84 3485 85 3515
rect 85 3485 115 3515
rect 115 3485 116 3515
rect 84 3484 116 3485
rect 84 3404 116 3436
rect 84 3355 116 3356
rect 84 3325 85 3355
rect 85 3325 115 3355
rect 115 3325 116 3355
rect 84 3324 116 3325
rect 84 3275 116 3276
rect 84 3245 85 3275
rect 85 3245 115 3275
rect 115 3245 116 3275
rect 84 3244 116 3245
rect 84 3195 116 3196
rect 84 3165 85 3195
rect 85 3165 115 3195
rect 115 3165 116 3195
rect 84 3164 116 3165
rect 84 3115 116 3116
rect 84 3085 85 3115
rect 85 3085 115 3115
rect 115 3085 116 3115
rect 84 3084 116 3085
rect 84 3004 116 3036
rect 84 2955 116 2956
rect 84 2925 85 2955
rect 85 2925 115 2955
rect 115 2925 116 2955
rect 84 2924 116 2925
rect 84 2844 116 2876
rect 84 2795 116 2796
rect 84 2765 85 2795
rect 85 2765 115 2795
rect 115 2765 116 2795
rect 84 2764 116 2765
rect 84 2715 116 2716
rect 84 2685 85 2715
rect 85 2685 115 2715
rect 115 2685 116 2715
rect 84 2684 116 2685
rect 84 2604 116 2636
rect 84 2555 116 2556
rect 84 2525 85 2555
rect 85 2525 115 2555
rect 115 2525 116 2555
rect 84 2524 116 2525
rect 164 3595 196 3596
rect 164 3565 165 3595
rect 165 3565 195 3595
rect 195 3565 196 3595
rect 164 3564 196 3565
rect 164 3515 196 3516
rect 164 3485 165 3515
rect 165 3485 195 3515
rect 195 3485 196 3515
rect 164 3484 196 3485
rect 164 3404 196 3436
rect 164 3355 196 3356
rect 164 3325 165 3355
rect 165 3325 195 3355
rect 195 3325 196 3355
rect 164 3324 196 3325
rect 164 3275 196 3276
rect 164 3245 165 3275
rect 165 3245 195 3275
rect 195 3245 196 3275
rect 164 3244 196 3245
rect 164 3195 196 3196
rect 164 3165 165 3195
rect 165 3165 195 3195
rect 195 3165 196 3195
rect 164 3164 196 3165
rect 164 3115 196 3116
rect 164 3085 165 3115
rect 165 3085 195 3115
rect 195 3085 196 3115
rect 164 3084 196 3085
rect 164 3004 196 3036
rect 164 2955 196 2956
rect 164 2925 165 2955
rect 165 2925 195 2955
rect 195 2925 196 2955
rect 164 2924 196 2925
rect 164 2844 196 2876
rect 164 2795 196 2796
rect 164 2765 165 2795
rect 165 2765 195 2795
rect 195 2765 196 2795
rect 164 2764 196 2765
rect 164 2715 196 2716
rect 164 2685 165 2715
rect 165 2685 195 2715
rect 195 2685 196 2715
rect 164 2684 196 2685
rect 164 2604 196 2636
rect 164 2555 196 2556
rect 164 2525 165 2555
rect 165 2525 195 2555
rect 195 2525 196 2555
rect 164 2524 196 2525
rect 244 3595 276 3596
rect 244 3565 245 3595
rect 245 3565 275 3595
rect 275 3565 276 3595
rect 244 3564 276 3565
rect 244 3515 276 3516
rect 244 3485 245 3515
rect 245 3485 275 3515
rect 275 3485 276 3515
rect 244 3484 276 3485
rect 244 3404 276 3436
rect 244 3355 276 3356
rect 244 3325 245 3355
rect 245 3325 275 3355
rect 275 3325 276 3355
rect 244 3324 276 3325
rect 244 3275 276 3276
rect 244 3245 245 3275
rect 245 3245 275 3275
rect 275 3245 276 3275
rect 244 3244 276 3245
rect 244 3195 276 3196
rect 244 3165 245 3195
rect 245 3165 275 3195
rect 275 3165 276 3195
rect 244 3164 276 3165
rect 244 3115 276 3116
rect 244 3085 245 3115
rect 245 3085 275 3115
rect 275 3085 276 3115
rect 244 3084 276 3085
rect 244 3004 276 3036
rect 244 2955 276 2956
rect 244 2925 245 2955
rect 245 2925 275 2955
rect 275 2925 276 2955
rect 244 2924 276 2925
rect 244 2844 276 2876
rect 244 2795 276 2796
rect 244 2765 245 2795
rect 245 2765 275 2795
rect 275 2765 276 2795
rect 244 2764 276 2765
rect 244 2715 276 2716
rect 244 2685 245 2715
rect 245 2685 275 2715
rect 275 2685 276 2715
rect 244 2684 276 2685
rect 244 2604 276 2636
rect 244 2555 276 2556
rect 244 2525 245 2555
rect 245 2525 275 2555
rect 275 2525 276 2555
rect 244 2524 276 2525
rect 324 3595 356 3596
rect 324 3565 325 3595
rect 325 3565 355 3595
rect 355 3565 356 3595
rect 324 3564 356 3565
rect 324 3515 356 3516
rect 324 3485 325 3515
rect 325 3485 355 3515
rect 355 3485 356 3515
rect 324 3484 356 3485
rect 324 3404 356 3436
rect 324 3355 356 3356
rect 324 3325 325 3355
rect 325 3325 355 3355
rect 355 3325 356 3355
rect 324 3324 356 3325
rect 324 3275 356 3276
rect 324 3245 325 3275
rect 325 3245 355 3275
rect 355 3245 356 3275
rect 324 3244 356 3245
rect 324 3195 356 3196
rect 324 3165 325 3195
rect 325 3165 355 3195
rect 355 3165 356 3195
rect 324 3164 356 3165
rect 324 3115 356 3116
rect 324 3085 325 3115
rect 325 3085 355 3115
rect 355 3085 356 3115
rect 324 3084 356 3085
rect 324 3004 356 3036
rect 324 2955 356 2956
rect 324 2925 325 2955
rect 325 2925 355 2955
rect 355 2925 356 2955
rect 324 2924 356 2925
rect 324 2844 356 2876
rect 324 2795 356 2796
rect 324 2765 325 2795
rect 325 2765 355 2795
rect 355 2765 356 2795
rect 324 2764 356 2765
rect 324 2715 356 2716
rect 324 2685 325 2715
rect 325 2685 355 2715
rect 355 2685 356 2715
rect 324 2684 356 2685
rect 324 2604 356 2636
rect 324 2555 356 2556
rect 324 2525 325 2555
rect 325 2525 355 2555
rect 355 2525 356 2555
rect 324 2524 356 2525
rect 404 3595 436 3596
rect 404 3565 405 3595
rect 405 3565 435 3595
rect 435 3565 436 3595
rect 404 3564 436 3565
rect 404 3515 436 3516
rect 404 3485 405 3515
rect 405 3485 435 3515
rect 435 3485 436 3515
rect 404 3484 436 3485
rect 404 3404 436 3436
rect 404 3355 436 3356
rect 404 3325 405 3355
rect 405 3325 435 3355
rect 435 3325 436 3355
rect 404 3324 436 3325
rect 404 3275 436 3276
rect 404 3245 405 3275
rect 405 3245 435 3275
rect 435 3245 436 3275
rect 404 3244 436 3245
rect 404 3195 436 3196
rect 404 3165 405 3195
rect 405 3165 435 3195
rect 435 3165 436 3195
rect 404 3164 436 3165
rect 404 3115 436 3116
rect 404 3085 405 3115
rect 405 3085 435 3115
rect 435 3085 436 3115
rect 404 3084 436 3085
rect 404 3004 436 3036
rect 404 2955 436 2956
rect 404 2925 405 2955
rect 405 2925 435 2955
rect 435 2925 436 2955
rect 404 2924 436 2925
rect 404 2844 436 2876
rect 404 2795 436 2796
rect 404 2765 405 2795
rect 405 2765 435 2795
rect 435 2765 436 2795
rect 404 2764 436 2765
rect 404 2715 436 2716
rect 404 2685 405 2715
rect 405 2685 435 2715
rect 435 2685 436 2715
rect 404 2684 436 2685
rect 404 2604 436 2636
rect 404 2555 436 2556
rect 404 2525 405 2555
rect 405 2525 435 2555
rect 435 2525 436 2555
rect 404 2524 436 2525
rect 484 3595 516 3596
rect 484 3565 485 3595
rect 485 3565 515 3595
rect 515 3565 516 3595
rect 484 3564 516 3565
rect 484 3515 516 3516
rect 484 3485 485 3515
rect 485 3485 515 3515
rect 515 3485 516 3515
rect 484 3484 516 3485
rect 484 3404 516 3436
rect 484 3355 516 3356
rect 484 3325 485 3355
rect 485 3325 515 3355
rect 515 3325 516 3355
rect 484 3324 516 3325
rect 484 3275 516 3276
rect 484 3245 485 3275
rect 485 3245 515 3275
rect 515 3245 516 3275
rect 484 3244 516 3245
rect 484 3195 516 3196
rect 484 3165 485 3195
rect 485 3165 515 3195
rect 515 3165 516 3195
rect 484 3164 516 3165
rect 484 3115 516 3116
rect 484 3085 485 3115
rect 485 3085 515 3115
rect 515 3085 516 3115
rect 484 3084 516 3085
rect 484 3004 516 3036
rect 484 2955 516 2956
rect 484 2925 485 2955
rect 485 2925 515 2955
rect 515 2925 516 2955
rect 484 2924 516 2925
rect 484 2844 516 2876
rect 484 2795 516 2796
rect 484 2765 485 2795
rect 485 2765 515 2795
rect 515 2765 516 2795
rect 484 2764 516 2765
rect 484 2715 516 2716
rect 484 2685 485 2715
rect 485 2685 515 2715
rect 515 2685 516 2715
rect 484 2684 516 2685
rect 484 2604 516 2636
rect 484 2555 516 2556
rect 484 2525 485 2555
rect 485 2525 515 2555
rect 515 2525 516 2555
rect 484 2524 516 2525
rect 564 3595 596 3596
rect 564 3565 565 3595
rect 565 3565 595 3595
rect 595 3565 596 3595
rect 564 3564 596 3565
rect 564 3515 596 3516
rect 564 3485 565 3515
rect 565 3485 595 3515
rect 595 3485 596 3515
rect 564 3484 596 3485
rect 564 3404 596 3436
rect 564 3355 596 3356
rect 564 3325 565 3355
rect 565 3325 595 3355
rect 595 3325 596 3355
rect 564 3324 596 3325
rect 564 3275 596 3276
rect 564 3245 565 3275
rect 565 3245 595 3275
rect 595 3245 596 3275
rect 564 3244 596 3245
rect 564 3195 596 3196
rect 564 3165 565 3195
rect 565 3165 595 3195
rect 595 3165 596 3195
rect 564 3164 596 3165
rect 564 3115 596 3116
rect 564 3085 565 3115
rect 565 3085 595 3115
rect 595 3085 596 3115
rect 564 3084 596 3085
rect 564 3004 596 3036
rect 564 2955 596 2956
rect 564 2925 565 2955
rect 565 2925 595 2955
rect 595 2925 596 2955
rect 564 2924 596 2925
rect 564 2844 596 2876
rect 564 2795 596 2796
rect 564 2765 565 2795
rect 565 2765 595 2795
rect 595 2765 596 2795
rect 564 2764 596 2765
rect 564 2715 596 2716
rect 564 2685 565 2715
rect 565 2685 595 2715
rect 595 2685 596 2715
rect 564 2684 596 2685
rect 564 2604 596 2636
rect 564 2555 596 2556
rect 564 2525 565 2555
rect 565 2525 595 2555
rect 595 2525 596 2555
rect 564 2524 596 2525
rect 644 3595 676 3596
rect 644 3565 645 3595
rect 645 3565 675 3595
rect 675 3565 676 3595
rect 644 3564 676 3565
rect 644 3515 676 3516
rect 644 3485 645 3515
rect 645 3485 675 3515
rect 675 3485 676 3515
rect 644 3484 676 3485
rect 644 3404 676 3436
rect 644 3355 676 3356
rect 644 3325 645 3355
rect 645 3325 675 3355
rect 675 3325 676 3355
rect 644 3324 676 3325
rect 644 3275 676 3276
rect 644 3245 645 3275
rect 645 3245 675 3275
rect 675 3245 676 3275
rect 644 3244 676 3245
rect 644 3195 676 3196
rect 644 3165 645 3195
rect 645 3165 675 3195
rect 675 3165 676 3195
rect 644 3164 676 3165
rect 644 3115 676 3116
rect 644 3085 645 3115
rect 645 3085 675 3115
rect 675 3085 676 3115
rect 644 3084 676 3085
rect 644 3004 676 3036
rect 644 2955 676 2956
rect 644 2925 645 2955
rect 645 2925 675 2955
rect 675 2925 676 2955
rect 644 2924 676 2925
rect 644 2844 676 2876
rect 644 2795 676 2796
rect 644 2765 645 2795
rect 645 2765 675 2795
rect 675 2765 676 2795
rect 644 2764 676 2765
rect 644 2715 676 2716
rect 644 2685 645 2715
rect 645 2685 675 2715
rect 675 2685 676 2715
rect 644 2684 676 2685
rect 644 2604 676 2636
rect 644 2555 676 2556
rect 644 2525 645 2555
rect 645 2525 675 2555
rect 675 2525 676 2555
rect 644 2524 676 2525
rect 724 3595 756 3596
rect 724 3565 725 3595
rect 725 3565 755 3595
rect 755 3565 756 3595
rect 724 3564 756 3565
rect 724 3515 756 3516
rect 724 3485 725 3515
rect 725 3485 755 3515
rect 755 3485 756 3515
rect 724 3484 756 3485
rect 724 3404 756 3436
rect 724 3355 756 3356
rect 724 3325 725 3355
rect 725 3325 755 3355
rect 755 3325 756 3355
rect 724 3324 756 3325
rect 724 3275 756 3276
rect 724 3245 725 3275
rect 725 3245 755 3275
rect 755 3245 756 3275
rect 724 3244 756 3245
rect 724 3195 756 3196
rect 724 3165 725 3195
rect 725 3165 755 3195
rect 755 3165 756 3195
rect 724 3164 756 3165
rect 724 3115 756 3116
rect 724 3085 725 3115
rect 725 3085 755 3115
rect 755 3085 756 3115
rect 724 3084 756 3085
rect 724 3004 756 3036
rect 724 2955 756 2956
rect 724 2925 725 2955
rect 725 2925 755 2955
rect 755 2925 756 2955
rect 724 2924 756 2925
rect 724 2844 756 2876
rect 724 2795 756 2796
rect 724 2765 725 2795
rect 725 2765 755 2795
rect 755 2765 756 2795
rect 724 2764 756 2765
rect 724 2715 756 2716
rect 724 2685 725 2715
rect 725 2685 755 2715
rect 755 2685 756 2715
rect 724 2684 756 2685
rect 724 2604 756 2636
rect 724 2555 756 2556
rect 724 2525 725 2555
rect 725 2525 755 2555
rect 755 2525 756 2555
rect 724 2524 756 2525
rect 804 3595 836 3596
rect 804 3565 805 3595
rect 805 3565 835 3595
rect 835 3565 836 3595
rect 804 3564 836 3565
rect 804 3515 836 3516
rect 804 3485 805 3515
rect 805 3485 835 3515
rect 835 3485 836 3515
rect 804 3484 836 3485
rect 804 3404 836 3436
rect 804 3355 836 3356
rect 804 3325 805 3355
rect 805 3325 835 3355
rect 835 3325 836 3355
rect 804 3324 836 3325
rect 804 3275 836 3276
rect 804 3245 805 3275
rect 805 3245 835 3275
rect 835 3245 836 3275
rect 804 3244 836 3245
rect 804 3195 836 3196
rect 804 3165 805 3195
rect 805 3165 835 3195
rect 835 3165 836 3195
rect 804 3164 836 3165
rect 804 3115 836 3116
rect 804 3085 805 3115
rect 805 3085 835 3115
rect 835 3085 836 3115
rect 804 3084 836 3085
rect 804 3004 836 3036
rect 804 2955 836 2956
rect 804 2925 805 2955
rect 805 2925 835 2955
rect 835 2925 836 2955
rect 804 2924 836 2925
rect 804 2844 836 2876
rect 804 2795 836 2796
rect 804 2765 805 2795
rect 805 2765 835 2795
rect 835 2765 836 2795
rect 804 2764 836 2765
rect 804 2715 836 2716
rect 804 2685 805 2715
rect 805 2685 835 2715
rect 835 2685 836 2715
rect 804 2684 836 2685
rect 804 2604 836 2636
rect 804 2555 836 2556
rect 804 2525 805 2555
rect 805 2525 835 2555
rect 835 2525 836 2555
rect 804 2524 836 2525
rect 884 3595 916 3596
rect 884 3565 885 3595
rect 885 3565 915 3595
rect 915 3565 916 3595
rect 884 3564 916 3565
rect 884 3515 916 3516
rect 884 3485 885 3515
rect 885 3485 915 3515
rect 915 3485 916 3515
rect 884 3484 916 3485
rect 884 3404 916 3436
rect 884 3355 916 3356
rect 884 3325 885 3355
rect 885 3325 915 3355
rect 915 3325 916 3355
rect 884 3324 916 3325
rect 884 3275 916 3276
rect 884 3245 885 3275
rect 885 3245 915 3275
rect 915 3245 916 3275
rect 884 3244 916 3245
rect 884 3195 916 3196
rect 884 3165 885 3195
rect 885 3165 915 3195
rect 915 3165 916 3195
rect 884 3164 916 3165
rect 884 3115 916 3116
rect 884 3085 885 3115
rect 885 3085 915 3115
rect 915 3085 916 3115
rect 884 3084 916 3085
rect 884 3004 916 3036
rect 884 2955 916 2956
rect 884 2925 885 2955
rect 885 2925 915 2955
rect 915 2925 916 2955
rect 884 2924 916 2925
rect 884 2844 916 2876
rect 884 2795 916 2796
rect 884 2765 885 2795
rect 885 2765 915 2795
rect 915 2765 916 2795
rect 884 2764 916 2765
rect 884 2715 916 2716
rect 884 2685 885 2715
rect 885 2685 915 2715
rect 915 2685 916 2715
rect 884 2684 916 2685
rect 884 2604 916 2636
rect 884 2555 916 2556
rect 884 2525 885 2555
rect 885 2525 915 2555
rect 915 2525 916 2555
rect 884 2524 916 2525
rect 964 3595 996 3596
rect 964 3565 965 3595
rect 965 3565 995 3595
rect 995 3565 996 3595
rect 964 3564 996 3565
rect 964 3515 996 3516
rect 964 3485 965 3515
rect 965 3485 995 3515
rect 995 3485 996 3515
rect 964 3484 996 3485
rect 964 3404 996 3436
rect 964 3355 996 3356
rect 964 3325 965 3355
rect 965 3325 995 3355
rect 995 3325 996 3355
rect 964 3324 996 3325
rect 964 3275 996 3276
rect 964 3245 965 3275
rect 965 3245 995 3275
rect 995 3245 996 3275
rect 964 3244 996 3245
rect 964 3195 996 3196
rect 964 3165 965 3195
rect 965 3165 995 3195
rect 995 3165 996 3195
rect 964 3164 996 3165
rect 964 3115 996 3116
rect 964 3085 965 3115
rect 965 3085 995 3115
rect 995 3085 996 3115
rect 964 3084 996 3085
rect 964 3004 996 3036
rect 964 2955 996 2956
rect 964 2925 965 2955
rect 965 2925 995 2955
rect 995 2925 996 2955
rect 964 2924 996 2925
rect 964 2844 996 2876
rect 964 2795 996 2796
rect 964 2765 965 2795
rect 965 2765 995 2795
rect 995 2765 996 2795
rect 964 2764 996 2765
rect 964 2715 996 2716
rect 964 2685 965 2715
rect 965 2685 995 2715
rect 995 2685 996 2715
rect 964 2684 996 2685
rect 964 2604 996 2636
rect 964 2555 996 2556
rect 964 2525 965 2555
rect 965 2525 995 2555
rect 995 2525 996 2555
rect 964 2524 996 2525
rect 1044 3595 1076 3596
rect 1044 3565 1045 3595
rect 1045 3565 1075 3595
rect 1075 3565 1076 3595
rect 1044 3564 1076 3565
rect 1044 3515 1076 3516
rect 1044 3485 1045 3515
rect 1045 3485 1075 3515
rect 1075 3485 1076 3515
rect 1044 3484 1076 3485
rect 1044 3404 1076 3436
rect 1044 3355 1076 3356
rect 1044 3325 1045 3355
rect 1045 3325 1075 3355
rect 1075 3325 1076 3355
rect 1044 3324 1076 3325
rect 1044 3275 1076 3276
rect 1044 3245 1045 3275
rect 1045 3245 1075 3275
rect 1075 3245 1076 3275
rect 1044 3244 1076 3245
rect 1044 3195 1076 3196
rect 1044 3165 1045 3195
rect 1045 3165 1075 3195
rect 1075 3165 1076 3195
rect 1044 3164 1076 3165
rect 1044 3115 1076 3116
rect 1044 3085 1045 3115
rect 1045 3085 1075 3115
rect 1075 3085 1076 3115
rect 1044 3084 1076 3085
rect 1044 3004 1076 3036
rect 1044 2955 1076 2956
rect 1044 2925 1045 2955
rect 1045 2925 1075 2955
rect 1075 2925 1076 2955
rect 1044 2924 1076 2925
rect 1044 2844 1076 2876
rect 1044 2795 1076 2796
rect 1044 2765 1045 2795
rect 1045 2765 1075 2795
rect 1075 2765 1076 2795
rect 1044 2764 1076 2765
rect 1044 2715 1076 2716
rect 1044 2685 1045 2715
rect 1045 2685 1075 2715
rect 1075 2685 1076 2715
rect 1044 2684 1076 2685
rect 1044 2604 1076 2636
rect 1044 2555 1076 2556
rect 1044 2525 1045 2555
rect 1045 2525 1075 2555
rect 1075 2525 1076 2555
rect 1044 2524 1076 2525
rect 1124 3595 1156 3596
rect 1124 3565 1125 3595
rect 1125 3565 1155 3595
rect 1155 3565 1156 3595
rect 1124 3564 1156 3565
rect 1124 3515 1156 3516
rect 1124 3485 1125 3515
rect 1125 3485 1155 3515
rect 1155 3485 1156 3515
rect 1124 3484 1156 3485
rect 1124 3404 1156 3436
rect 1124 3355 1156 3356
rect 1124 3325 1125 3355
rect 1125 3325 1155 3355
rect 1155 3325 1156 3355
rect 1124 3324 1156 3325
rect 1124 3275 1156 3276
rect 1124 3245 1125 3275
rect 1125 3245 1155 3275
rect 1155 3245 1156 3275
rect 1124 3244 1156 3245
rect 1124 3195 1156 3196
rect 1124 3165 1125 3195
rect 1125 3165 1155 3195
rect 1155 3165 1156 3195
rect 1124 3164 1156 3165
rect 1124 3115 1156 3116
rect 1124 3085 1125 3115
rect 1125 3085 1155 3115
rect 1155 3085 1156 3115
rect 1124 3084 1156 3085
rect 1124 3004 1156 3036
rect 1124 2955 1156 2956
rect 1124 2925 1125 2955
rect 1125 2925 1155 2955
rect 1155 2925 1156 2955
rect 1124 2924 1156 2925
rect 1124 2844 1156 2876
rect 1124 2795 1156 2796
rect 1124 2765 1125 2795
rect 1125 2765 1155 2795
rect 1155 2765 1156 2795
rect 1124 2764 1156 2765
rect 1124 2715 1156 2716
rect 1124 2685 1125 2715
rect 1125 2685 1155 2715
rect 1155 2685 1156 2715
rect 1124 2684 1156 2685
rect 1124 2604 1156 2636
rect 1124 2555 1156 2556
rect 1124 2525 1125 2555
rect 1125 2525 1155 2555
rect 1155 2525 1156 2555
rect 1124 2524 1156 2525
rect 1204 3595 1236 3596
rect 1204 3565 1205 3595
rect 1205 3565 1235 3595
rect 1235 3565 1236 3595
rect 1204 3564 1236 3565
rect 1204 3515 1236 3516
rect 1204 3485 1205 3515
rect 1205 3485 1235 3515
rect 1235 3485 1236 3515
rect 1204 3484 1236 3485
rect 1204 3404 1236 3436
rect 1204 3355 1236 3356
rect 1204 3325 1205 3355
rect 1205 3325 1235 3355
rect 1235 3325 1236 3355
rect 1204 3324 1236 3325
rect 1204 3275 1236 3276
rect 1204 3245 1205 3275
rect 1205 3245 1235 3275
rect 1235 3245 1236 3275
rect 1204 3244 1236 3245
rect 1204 3195 1236 3196
rect 1204 3165 1205 3195
rect 1205 3165 1235 3195
rect 1235 3165 1236 3195
rect 1204 3164 1236 3165
rect 1204 3115 1236 3116
rect 1204 3085 1205 3115
rect 1205 3085 1235 3115
rect 1235 3085 1236 3115
rect 1204 3084 1236 3085
rect 1204 3004 1236 3036
rect 1204 2955 1236 2956
rect 1204 2925 1205 2955
rect 1205 2925 1235 2955
rect 1235 2925 1236 2955
rect 1204 2924 1236 2925
rect 1204 2844 1236 2876
rect 1204 2795 1236 2796
rect 1204 2765 1205 2795
rect 1205 2765 1235 2795
rect 1235 2765 1236 2795
rect 1204 2764 1236 2765
rect 1204 2715 1236 2716
rect 1204 2685 1205 2715
rect 1205 2685 1235 2715
rect 1235 2685 1236 2715
rect 1204 2684 1236 2685
rect 1204 2604 1236 2636
rect 1204 2555 1236 2556
rect 1204 2525 1205 2555
rect 1205 2525 1235 2555
rect 1235 2525 1236 2555
rect 1204 2524 1236 2525
rect 1284 3595 1316 3596
rect 1284 3565 1285 3595
rect 1285 3565 1315 3595
rect 1315 3565 1316 3595
rect 1284 3564 1316 3565
rect 1284 3515 1316 3516
rect 1284 3485 1285 3515
rect 1285 3485 1315 3515
rect 1315 3485 1316 3515
rect 1284 3484 1316 3485
rect 1284 3404 1316 3436
rect 1284 3355 1316 3356
rect 1284 3325 1285 3355
rect 1285 3325 1315 3355
rect 1315 3325 1316 3355
rect 1284 3324 1316 3325
rect 1284 3275 1316 3276
rect 1284 3245 1285 3275
rect 1285 3245 1315 3275
rect 1315 3245 1316 3275
rect 1284 3244 1316 3245
rect 1284 3195 1316 3196
rect 1284 3165 1285 3195
rect 1285 3165 1315 3195
rect 1315 3165 1316 3195
rect 1284 3164 1316 3165
rect 1284 3115 1316 3116
rect 1284 3085 1285 3115
rect 1285 3085 1315 3115
rect 1315 3085 1316 3115
rect 1284 3084 1316 3085
rect 1284 3004 1316 3036
rect 1284 2955 1316 2956
rect 1284 2925 1285 2955
rect 1285 2925 1315 2955
rect 1315 2925 1316 2955
rect 1284 2924 1316 2925
rect 1284 2844 1316 2876
rect 1284 2795 1316 2796
rect 1284 2765 1285 2795
rect 1285 2765 1315 2795
rect 1315 2765 1316 2795
rect 1284 2764 1316 2765
rect 1284 2715 1316 2716
rect 1284 2685 1285 2715
rect 1285 2685 1315 2715
rect 1315 2685 1316 2715
rect 1284 2684 1316 2685
rect 1284 2604 1316 2636
rect 1284 2555 1316 2556
rect 1284 2525 1285 2555
rect 1285 2525 1315 2555
rect 1315 2525 1316 2555
rect 1284 2524 1316 2525
rect 1364 3595 1396 3596
rect 1364 3565 1365 3595
rect 1365 3565 1395 3595
rect 1395 3565 1396 3595
rect 1364 3564 1396 3565
rect 1364 3515 1396 3516
rect 1364 3485 1365 3515
rect 1365 3485 1395 3515
rect 1395 3485 1396 3515
rect 1364 3484 1396 3485
rect 1364 3404 1396 3436
rect 1364 3355 1396 3356
rect 1364 3325 1365 3355
rect 1365 3325 1395 3355
rect 1395 3325 1396 3355
rect 1364 3324 1396 3325
rect 1364 3275 1396 3276
rect 1364 3245 1365 3275
rect 1365 3245 1395 3275
rect 1395 3245 1396 3275
rect 1364 3244 1396 3245
rect 1364 3195 1396 3196
rect 1364 3165 1365 3195
rect 1365 3165 1395 3195
rect 1395 3165 1396 3195
rect 1364 3164 1396 3165
rect 1364 3115 1396 3116
rect 1364 3085 1365 3115
rect 1365 3085 1395 3115
rect 1395 3085 1396 3115
rect 1364 3084 1396 3085
rect 1364 3004 1396 3036
rect 1364 2955 1396 2956
rect 1364 2925 1365 2955
rect 1365 2925 1395 2955
rect 1395 2925 1396 2955
rect 1364 2924 1396 2925
rect 1364 2844 1396 2876
rect 1364 2795 1396 2796
rect 1364 2765 1365 2795
rect 1365 2765 1395 2795
rect 1395 2765 1396 2795
rect 1364 2764 1396 2765
rect 1364 2715 1396 2716
rect 1364 2685 1365 2715
rect 1365 2685 1395 2715
rect 1395 2685 1396 2715
rect 1364 2684 1396 2685
rect 1364 2604 1396 2636
rect 1364 2555 1396 2556
rect 1364 2525 1365 2555
rect 1365 2525 1395 2555
rect 1395 2525 1396 2555
rect 1364 2524 1396 2525
rect 1444 3595 1476 3596
rect 1444 3565 1445 3595
rect 1445 3565 1475 3595
rect 1475 3565 1476 3595
rect 1444 3564 1476 3565
rect 1444 3515 1476 3516
rect 1444 3485 1445 3515
rect 1445 3485 1475 3515
rect 1475 3485 1476 3515
rect 1444 3484 1476 3485
rect 1444 3404 1476 3436
rect 1444 3355 1476 3356
rect 1444 3325 1445 3355
rect 1445 3325 1475 3355
rect 1475 3325 1476 3355
rect 1444 3324 1476 3325
rect 1444 3275 1476 3276
rect 1444 3245 1445 3275
rect 1445 3245 1475 3275
rect 1475 3245 1476 3275
rect 1444 3244 1476 3245
rect 1444 3195 1476 3196
rect 1444 3165 1445 3195
rect 1445 3165 1475 3195
rect 1475 3165 1476 3195
rect 1444 3164 1476 3165
rect 1444 3115 1476 3116
rect 1444 3085 1445 3115
rect 1445 3085 1475 3115
rect 1475 3085 1476 3115
rect 1444 3084 1476 3085
rect 1444 3004 1476 3036
rect 1444 2955 1476 2956
rect 1444 2925 1445 2955
rect 1445 2925 1475 2955
rect 1475 2925 1476 2955
rect 1444 2924 1476 2925
rect 1444 2844 1476 2876
rect 1444 2795 1476 2796
rect 1444 2765 1445 2795
rect 1445 2765 1475 2795
rect 1475 2765 1476 2795
rect 1444 2764 1476 2765
rect 1444 2715 1476 2716
rect 1444 2685 1445 2715
rect 1445 2685 1475 2715
rect 1475 2685 1476 2715
rect 1444 2684 1476 2685
rect 1444 2604 1476 2636
rect 1444 2555 1476 2556
rect 1444 2525 1445 2555
rect 1445 2525 1475 2555
rect 1475 2525 1476 2555
rect 1444 2524 1476 2525
rect 1524 3595 1556 3596
rect 1524 3565 1525 3595
rect 1525 3565 1555 3595
rect 1555 3565 1556 3595
rect 1524 3564 1556 3565
rect 1524 3515 1556 3516
rect 1524 3485 1525 3515
rect 1525 3485 1555 3515
rect 1555 3485 1556 3515
rect 1524 3484 1556 3485
rect 1524 3404 1556 3436
rect 1524 3355 1556 3356
rect 1524 3325 1525 3355
rect 1525 3325 1555 3355
rect 1555 3325 1556 3355
rect 1524 3324 1556 3325
rect 1524 3275 1556 3276
rect 1524 3245 1525 3275
rect 1525 3245 1555 3275
rect 1555 3245 1556 3275
rect 1524 3244 1556 3245
rect 1524 3195 1556 3196
rect 1524 3165 1525 3195
rect 1525 3165 1555 3195
rect 1555 3165 1556 3195
rect 1524 3164 1556 3165
rect 1524 3115 1556 3116
rect 1524 3085 1525 3115
rect 1525 3085 1555 3115
rect 1555 3085 1556 3115
rect 1524 3084 1556 3085
rect 1524 3004 1556 3036
rect 1524 2955 1556 2956
rect 1524 2925 1525 2955
rect 1525 2925 1555 2955
rect 1555 2925 1556 2955
rect 1524 2924 1556 2925
rect 1524 2844 1556 2876
rect 1524 2795 1556 2796
rect 1524 2765 1525 2795
rect 1525 2765 1555 2795
rect 1555 2765 1556 2795
rect 1524 2764 1556 2765
rect 1524 2715 1556 2716
rect 1524 2685 1525 2715
rect 1525 2685 1555 2715
rect 1555 2685 1556 2715
rect 1524 2684 1556 2685
rect 1524 2604 1556 2636
rect 1524 2555 1556 2556
rect 1524 2525 1525 2555
rect 1525 2525 1555 2555
rect 1555 2525 1556 2555
rect 1524 2524 1556 2525
rect 1604 3595 1636 3596
rect 1604 3565 1605 3595
rect 1605 3565 1635 3595
rect 1635 3565 1636 3595
rect 1604 3564 1636 3565
rect 1604 3515 1636 3516
rect 1604 3485 1605 3515
rect 1605 3485 1635 3515
rect 1635 3485 1636 3515
rect 1604 3484 1636 3485
rect 1604 3404 1636 3436
rect 1604 3355 1636 3356
rect 1604 3325 1605 3355
rect 1605 3325 1635 3355
rect 1635 3325 1636 3355
rect 1604 3324 1636 3325
rect 1604 3275 1636 3276
rect 1604 3245 1605 3275
rect 1605 3245 1635 3275
rect 1635 3245 1636 3275
rect 1604 3244 1636 3245
rect 1604 3195 1636 3196
rect 1604 3165 1605 3195
rect 1605 3165 1635 3195
rect 1635 3165 1636 3195
rect 1604 3164 1636 3165
rect 1604 3115 1636 3116
rect 1604 3085 1605 3115
rect 1605 3085 1635 3115
rect 1635 3085 1636 3115
rect 1604 3084 1636 3085
rect 1604 3004 1636 3036
rect 1604 2955 1636 2956
rect 1604 2925 1605 2955
rect 1605 2925 1635 2955
rect 1635 2925 1636 2955
rect 1604 2924 1636 2925
rect 1604 2844 1636 2876
rect 1604 2795 1636 2796
rect 1604 2765 1605 2795
rect 1605 2765 1635 2795
rect 1635 2765 1636 2795
rect 1604 2764 1636 2765
rect 1604 2715 1636 2716
rect 1604 2685 1605 2715
rect 1605 2685 1635 2715
rect 1635 2685 1636 2715
rect 1604 2684 1636 2685
rect 1604 2604 1636 2636
rect 1604 2555 1636 2556
rect 1604 2525 1605 2555
rect 1605 2525 1635 2555
rect 1635 2525 1636 2555
rect 1604 2524 1636 2525
rect 1684 3595 1716 3596
rect 1684 3565 1685 3595
rect 1685 3565 1715 3595
rect 1715 3565 1716 3595
rect 1684 3564 1716 3565
rect 1684 3515 1716 3516
rect 1684 3485 1685 3515
rect 1685 3485 1715 3515
rect 1715 3485 1716 3515
rect 1684 3484 1716 3485
rect 1684 3404 1716 3436
rect 1684 3355 1716 3356
rect 1684 3325 1685 3355
rect 1685 3325 1715 3355
rect 1715 3325 1716 3355
rect 1684 3324 1716 3325
rect 1684 3275 1716 3276
rect 1684 3245 1685 3275
rect 1685 3245 1715 3275
rect 1715 3245 1716 3275
rect 1684 3244 1716 3245
rect 1684 3195 1716 3196
rect 1684 3165 1685 3195
rect 1685 3165 1715 3195
rect 1715 3165 1716 3195
rect 1684 3164 1716 3165
rect 1684 3115 1716 3116
rect 1684 3085 1685 3115
rect 1685 3085 1715 3115
rect 1715 3085 1716 3115
rect 1684 3084 1716 3085
rect 1684 3004 1716 3036
rect 1684 2955 1716 2956
rect 1684 2925 1685 2955
rect 1685 2925 1715 2955
rect 1715 2925 1716 2955
rect 1684 2924 1716 2925
rect 1684 2844 1716 2876
rect 1684 2795 1716 2796
rect 1684 2765 1685 2795
rect 1685 2765 1715 2795
rect 1715 2765 1716 2795
rect 1684 2764 1716 2765
rect 1684 2715 1716 2716
rect 1684 2685 1685 2715
rect 1685 2685 1715 2715
rect 1715 2685 1716 2715
rect 1684 2684 1716 2685
rect 1684 2604 1716 2636
rect 1684 2555 1716 2556
rect 1684 2525 1685 2555
rect 1685 2525 1715 2555
rect 1715 2525 1716 2555
rect 1684 2524 1716 2525
rect 1764 3595 1796 3596
rect 1764 3565 1765 3595
rect 1765 3565 1795 3595
rect 1795 3565 1796 3595
rect 1764 3564 1796 3565
rect 1764 3515 1796 3516
rect 1764 3485 1765 3515
rect 1765 3485 1795 3515
rect 1795 3485 1796 3515
rect 1764 3484 1796 3485
rect 1764 3404 1796 3436
rect 1764 3355 1796 3356
rect 1764 3325 1765 3355
rect 1765 3325 1795 3355
rect 1795 3325 1796 3355
rect 1764 3324 1796 3325
rect 1764 3275 1796 3276
rect 1764 3245 1765 3275
rect 1765 3245 1795 3275
rect 1795 3245 1796 3275
rect 1764 3244 1796 3245
rect 1764 3195 1796 3196
rect 1764 3165 1765 3195
rect 1765 3165 1795 3195
rect 1795 3165 1796 3195
rect 1764 3164 1796 3165
rect 1764 3115 1796 3116
rect 1764 3085 1765 3115
rect 1765 3085 1795 3115
rect 1795 3085 1796 3115
rect 1764 3084 1796 3085
rect 1764 3004 1796 3036
rect 1764 2955 1796 2956
rect 1764 2925 1765 2955
rect 1765 2925 1795 2955
rect 1795 2925 1796 2955
rect 1764 2924 1796 2925
rect 1764 2844 1796 2876
rect 1764 2795 1796 2796
rect 1764 2765 1765 2795
rect 1765 2765 1795 2795
rect 1795 2765 1796 2795
rect 1764 2764 1796 2765
rect 1764 2715 1796 2716
rect 1764 2685 1765 2715
rect 1765 2685 1795 2715
rect 1795 2685 1796 2715
rect 1764 2684 1796 2685
rect 1764 2604 1796 2636
rect 1764 2555 1796 2556
rect 1764 2525 1765 2555
rect 1765 2525 1795 2555
rect 1795 2525 1796 2555
rect 1764 2524 1796 2525
rect 1844 3595 1876 3596
rect 1844 3565 1845 3595
rect 1845 3565 1875 3595
rect 1875 3565 1876 3595
rect 1844 3564 1876 3565
rect 1844 3515 1876 3516
rect 1844 3485 1845 3515
rect 1845 3485 1875 3515
rect 1875 3485 1876 3515
rect 1844 3484 1876 3485
rect 1844 3404 1876 3436
rect 1844 3355 1876 3356
rect 1844 3325 1845 3355
rect 1845 3325 1875 3355
rect 1875 3325 1876 3355
rect 1844 3324 1876 3325
rect 1844 3275 1876 3276
rect 1844 3245 1845 3275
rect 1845 3245 1875 3275
rect 1875 3245 1876 3275
rect 1844 3244 1876 3245
rect 1844 3195 1876 3196
rect 1844 3165 1845 3195
rect 1845 3165 1875 3195
rect 1875 3165 1876 3195
rect 1844 3164 1876 3165
rect 1844 3115 1876 3116
rect 1844 3085 1845 3115
rect 1845 3085 1875 3115
rect 1875 3085 1876 3115
rect 1844 3084 1876 3085
rect 1844 3004 1876 3036
rect 1844 2955 1876 2956
rect 1844 2925 1845 2955
rect 1845 2925 1875 2955
rect 1875 2925 1876 2955
rect 1844 2924 1876 2925
rect 1844 2844 1876 2876
rect 1844 2795 1876 2796
rect 1844 2765 1845 2795
rect 1845 2765 1875 2795
rect 1875 2765 1876 2795
rect 1844 2764 1876 2765
rect 1844 2715 1876 2716
rect 1844 2685 1845 2715
rect 1845 2685 1875 2715
rect 1875 2685 1876 2715
rect 1844 2684 1876 2685
rect 1844 2604 1876 2636
rect 1844 2555 1876 2556
rect 1844 2525 1845 2555
rect 1845 2525 1875 2555
rect 1875 2525 1876 2555
rect 1844 2524 1876 2525
rect 1924 3595 1956 3596
rect 1924 3565 1925 3595
rect 1925 3565 1955 3595
rect 1955 3565 1956 3595
rect 1924 3564 1956 3565
rect 1924 3515 1956 3516
rect 1924 3485 1925 3515
rect 1925 3485 1955 3515
rect 1955 3485 1956 3515
rect 1924 3484 1956 3485
rect 1924 3404 1956 3436
rect 1924 3355 1956 3356
rect 1924 3325 1925 3355
rect 1925 3325 1955 3355
rect 1955 3325 1956 3355
rect 1924 3324 1956 3325
rect 1924 3275 1956 3276
rect 1924 3245 1925 3275
rect 1925 3245 1955 3275
rect 1955 3245 1956 3275
rect 1924 3244 1956 3245
rect 1924 3195 1956 3196
rect 1924 3165 1925 3195
rect 1925 3165 1955 3195
rect 1955 3165 1956 3195
rect 1924 3164 1956 3165
rect 1924 3115 1956 3116
rect 1924 3085 1925 3115
rect 1925 3085 1955 3115
rect 1955 3085 1956 3115
rect 1924 3084 1956 3085
rect 1924 3004 1956 3036
rect 1924 2955 1956 2956
rect 1924 2925 1925 2955
rect 1925 2925 1955 2955
rect 1955 2925 1956 2955
rect 1924 2924 1956 2925
rect 1924 2844 1956 2876
rect 1924 2795 1956 2796
rect 1924 2765 1925 2795
rect 1925 2765 1955 2795
rect 1955 2765 1956 2795
rect 1924 2764 1956 2765
rect 1924 2715 1956 2716
rect 1924 2685 1925 2715
rect 1925 2685 1955 2715
rect 1955 2685 1956 2715
rect 1924 2684 1956 2685
rect 1924 2604 1956 2636
rect 1924 2555 1956 2556
rect 1924 2525 1925 2555
rect 1925 2525 1955 2555
rect 1955 2525 1956 2555
rect 1924 2524 1956 2525
rect 2004 3595 2036 3596
rect 2004 3565 2005 3595
rect 2005 3565 2035 3595
rect 2035 3565 2036 3595
rect 2004 3564 2036 3565
rect 2004 3515 2036 3516
rect 2004 3485 2005 3515
rect 2005 3485 2035 3515
rect 2035 3485 2036 3515
rect 2004 3484 2036 3485
rect 2004 3404 2036 3436
rect 2004 3355 2036 3356
rect 2004 3325 2005 3355
rect 2005 3325 2035 3355
rect 2035 3325 2036 3355
rect 2004 3324 2036 3325
rect 2004 3275 2036 3276
rect 2004 3245 2005 3275
rect 2005 3245 2035 3275
rect 2035 3245 2036 3275
rect 2004 3244 2036 3245
rect 2004 3195 2036 3196
rect 2004 3165 2005 3195
rect 2005 3165 2035 3195
rect 2035 3165 2036 3195
rect 2004 3164 2036 3165
rect 2004 3115 2036 3116
rect 2004 3085 2005 3115
rect 2005 3085 2035 3115
rect 2035 3085 2036 3115
rect 2004 3084 2036 3085
rect 2004 3004 2036 3036
rect 2004 2955 2036 2956
rect 2004 2925 2005 2955
rect 2005 2925 2035 2955
rect 2035 2925 2036 2955
rect 2004 2924 2036 2925
rect 2004 2844 2036 2876
rect 2004 2795 2036 2796
rect 2004 2765 2005 2795
rect 2005 2765 2035 2795
rect 2035 2765 2036 2795
rect 2004 2764 2036 2765
rect 2004 2715 2036 2716
rect 2004 2685 2005 2715
rect 2005 2685 2035 2715
rect 2035 2685 2036 2715
rect 2004 2684 2036 2685
rect 2004 2604 2036 2636
rect 2004 2555 2036 2556
rect 2004 2525 2005 2555
rect 2005 2525 2035 2555
rect 2035 2525 2036 2555
rect 2004 2524 2036 2525
rect 2084 3595 2116 3596
rect 2084 3565 2085 3595
rect 2085 3565 2115 3595
rect 2115 3565 2116 3595
rect 2084 3564 2116 3565
rect 2084 3515 2116 3516
rect 2084 3485 2085 3515
rect 2085 3485 2115 3515
rect 2115 3485 2116 3515
rect 2084 3484 2116 3485
rect 2084 3404 2116 3436
rect 2084 3355 2116 3356
rect 2084 3325 2085 3355
rect 2085 3325 2115 3355
rect 2115 3325 2116 3355
rect 2084 3324 2116 3325
rect 2084 3275 2116 3276
rect 2084 3245 2085 3275
rect 2085 3245 2115 3275
rect 2115 3245 2116 3275
rect 2084 3244 2116 3245
rect 2084 3195 2116 3196
rect 2084 3165 2085 3195
rect 2085 3165 2115 3195
rect 2115 3165 2116 3195
rect 2084 3164 2116 3165
rect 2084 3115 2116 3116
rect 2084 3085 2085 3115
rect 2085 3085 2115 3115
rect 2115 3085 2116 3115
rect 2084 3084 2116 3085
rect 2084 3004 2116 3036
rect 2084 2955 2116 2956
rect 2084 2925 2085 2955
rect 2085 2925 2115 2955
rect 2115 2925 2116 2955
rect 2084 2924 2116 2925
rect 2084 2844 2116 2876
rect 2084 2795 2116 2796
rect 2084 2765 2085 2795
rect 2085 2765 2115 2795
rect 2115 2765 2116 2795
rect 2084 2764 2116 2765
rect 2084 2715 2116 2716
rect 2084 2685 2085 2715
rect 2085 2685 2115 2715
rect 2115 2685 2116 2715
rect 2084 2684 2116 2685
rect 2084 2604 2116 2636
rect 2084 2555 2116 2556
rect 2084 2525 2085 2555
rect 2085 2525 2115 2555
rect 2115 2525 2116 2555
rect 2084 2524 2116 2525
rect 2164 3595 2196 3596
rect 2164 3565 2165 3595
rect 2165 3565 2195 3595
rect 2195 3565 2196 3595
rect 2164 3564 2196 3565
rect 2164 3515 2196 3516
rect 2164 3485 2165 3515
rect 2165 3485 2195 3515
rect 2195 3485 2196 3515
rect 2164 3484 2196 3485
rect 2164 3404 2196 3436
rect 2164 3355 2196 3356
rect 2164 3325 2165 3355
rect 2165 3325 2195 3355
rect 2195 3325 2196 3355
rect 2164 3324 2196 3325
rect 2164 3275 2196 3276
rect 2164 3245 2165 3275
rect 2165 3245 2195 3275
rect 2195 3245 2196 3275
rect 2164 3244 2196 3245
rect 2164 3195 2196 3196
rect 2164 3165 2165 3195
rect 2165 3165 2195 3195
rect 2195 3165 2196 3195
rect 2164 3164 2196 3165
rect 2164 3115 2196 3116
rect 2164 3085 2165 3115
rect 2165 3085 2195 3115
rect 2195 3085 2196 3115
rect 2164 3084 2196 3085
rect 2164 3004 2196 3036
rect 2164 2955 2196 2956
rect 2164 2925 2165 2955
rect 2165 2925 2195 2955
rect 2195 2925 2196 2955
rect 2164 2924 2196 2925
rect 2164 2844 2196 2876
rect 2164 2795 2196 2796
rect 2164 2765 2165 2795
rect 2165 2765 2195 2795
rect 2195 2765 2196 2795
rect 2164 2764 2196 2765
rect 2164 2715 2196 2716
rect 2164 2685 2165 2715
rect 2165 2685 2195 2715
rect 2195 2685 2196 2715
rect 2164 2684 2196 2685
rect 2164 2604 2196 2636
rect 2164 2555 2196 2556
rect 2164 2525 2165 2555
rect 2165 2525 2195 2555
rect 2195 2525 2196 2555
rect 2164 2524 2196 2525
rect 2244 3595 2276 3596
rect 2244 3565 2245 3595
rect 2245 3565 2275 3595
rect 2275 3565 2276 3595
rect 2244 3564 2276 3565
rect 2244 3515 2276 3516
rect 2244 3485 2245 3515
rect 2245 3485 2275 3515
rect 2275 3485 2276 3515
rect 2244 3484 2276 3485
rect 2244 3404 2276 3436
rect 2244 3355 2276 3356
rect 2244 3325 2245 3355
rect 2245 3325 2275 3355
rect 2275 3325 2276 3355
rect 2244 3324 2276 3325
rect 2244 3275 2276 3276
rect 2244 3245 2245 3275
rect 2245 3245 2275 3275
rect 2275 3245 2276 3275
rect 2244 3244 2276 3245
rect 2244 3195 2276 3196
rect 2244 3165 2245 3195
rect 2245 3165 2275 3195
rect 2275 3165 2276 3195
rect 2244 3164 2276 3165
rect 2244 3115 2276 3116
rect 2244 3085 2245 3115
rect 2245 3085 2275 3115
rect 2275 3085 2276 3115
rect 2244 3084 2276 3085
rect 2244 3004 2276 3036
rect 2244 2955 2276 2956
rect 2244 2925 2245 2955
rect 2245 2925 2275 2955
rect 2275 2925 2276 2955
rect 2244 2924 2276 2925
rect 2244 2844 2276 2876
rect 2244 2795 2276 2796
rect 2244 2765 2245 2795
rect 2245 2765 2275 2795
rect 2275 2765 2276 2795
rect 2244 2764 2276 2765
rect 2244 2715 2276 2716
rect 2244 2685 2245 2715
rect 2245 2685 2275 2715
rect 2275 2685 2276 2715
rect 2244 2684 2276 2685
rect 2244 2604 2276 2636
rect 2244 2555 2276 2556
rect 2244 2525 2245 2555
rect 2245 2525 2275 2555
rect 2275 2525 2276 2555
rect 2244 2524 2276 2525
rect 2324 3595 2356 3596
rect 2324 3565 2325 3595
rect 2325 3565 2355 3595
rect 2355 3565 2356 3595
rect 2324 3564 2356 3565
rect 2324 3515 2356 3516
rect 2324 3485 2325 3515
rect 2325 3485 2355 3515
rect 2355 3485 2356 3515
rect 2324 3484 2356 3485
rect 2324 3404 2356 3436
rect 2324 3355 2356 3356
rect 2324 3325 2325 3355
rect 2325 3325 2355 3355
rect 2355 3325 2356 3355
rect 2324 3324 2356 3325
rect 2324 3275 2356 3276
rect 2324 3245 2325 3275
rect 2325 3245 2355 3275
rect 2355 3245 2356 3275
rect 2324 3244 2356 3245
rect 2324 3195 2356 3196
rect 2324 3165 2325 3195
rect 2325 3165 2355 3195
rect 2355 3165 2356 3195
rect 2324 3164 2356 3165
rect 2324 3115 2356 3116
rect 2324 3085 2325 3115
rect 2325 3085 2355 3115
rect 2355 3085 2356 3115
rect 2324 3084 2356 3085
rect 2324 3004 2356 3036
rect 2324 2955 2356 2956
rect 2324 2925 2325 2955
rect 2325 2925 2355 2955
rect 2355 2925 2356 2955
rect 2324 2924 2356 2925
rect 2324 2844 2356 2876
rect 2324 2795 2356 2796
rect 2324 2765 2325 2795
rect 2325 2765 2355 2795
rect 2355 2765 2356 2795
rect 2324 2764 2356 2765
rect 2324 2715 2356 2716
rect 2324 2685 2325 2715
rect 2325 2685 2355 2715
rect 2355 2685 2356 2715
rect 2324 2684 2356 2685
rect 2324 2604 2356 2636
rect 2324 2555 2356 2556
rect 2324 2525 2325 2555
rect 2325 2525 2355 2555
rect 2355 2525 2356 2555
rect 2324 2524 2356 2525
rect 2404 3595 2436 3596
rect 2404 3565 2405 3595
rect 2405 3565 2435 3595
rect 2435 3565 2436 3595
rect 2404 3564 2436 3565
rect 2404 3515 2436 3516
rect 2404 3485 2405 3515
rect 2405 3485 2435 3515
rect 2435 3485 2436 3515
rect 2404 3484 2436 3485
rect 2404 3404 2436 3436
rect 2404 3355 2436 3356
rect 2404 3325 2405 3355
rect 2405 3325 2435 3355
rect 2435 3325 2436 3355
rect 2404 3324 2436 3325
rect 2404 3275 2436 3276
rect 2404 3245 2405 3275
rect 2405 3245 2435 3275
rect 2435 3245 2436 3275
rect 2404 3244 2436 3245
rect 2404 3195 2436 3196
rect 2404 3165 2405 3195
rect 2405 3165 2435 3195
rect 2435 3165 2436 3195
rect 2404 3164 2436 3165
rect 2404 3115 2436 3116
rect 2404 3085 2405 3115
rect 2405 3085 2435 3115
rect 2435 3085 2436 3115
rect 2404 3084 2436 3085
rect 2404 3004 2436 3036
rect 2404 2955 2436 2956
rect 2404 2925 2405 2955
rect 2405 2925 2435 2955
rect 2435 2925 2436 2955
rect 2404 2924 2436 2925
rect 2404 2844 2436 2876
rect 2404 2795 2436 2796
rect 2404 2765 2405 2795
rect 2405 2765 2435 2795
rect 2435 2765 2436 2795
rect 2404 2764 2436 2765
rect 2404 2715 2436 2716
rect 2404 2685 2405 2715
rect 2405 2685 2435 2715
rect 2435 2685 2436 2715
rect 2404 2684 2436 2685
rect 2404 2604 2436 2636
rect 2404 2555 2436 2556
rect 2404 2525 2405 2555
rect 2405 2525 2435 2555
rect 2435 2525 2436 2555
rect 2404 2524 2436 2525
rect 2484 3595 2516 3596
rect 2484 3565 2485 3595
rect 2485 3565 2515 3595
rect 2515 3565 2516 3595
rect 2484 3564 2516 3565
rect 2484 3515 2516 3516
rect 2484 3485 2485 3515
rect 2485 3485 2515 3515
rect 2515 3485 2516 3515
rect 2484 3484 2516 3485
rect 2484 3404 2516 3436
rect 2484 3355 2516 3356
rect 2484 3325 2485 3355
rect 2485 3325 2515 3355
rect 2515 3325 2516 3355
rect 2484 3324 2516 3325
rect 2484 3275 2516 3276
rect 2484 3245 2485 3275
rect 2485 3245 2515 3275
rect 2515 3245 2516 3275
rect 2484 3244 2516 3245
rect 2484 3195 2516 3196
rect 2484 3165 2485 3195
rect 2485 3165 2515 3195
rect 2515 3165 2516 3195
rect 2484 3164 2516 3165
rect 2484 3115 2516 3116
rect 2484 3085 2485 3115
rect 2485 3085 2515 3115
rect 2515 3085 2516 3115
rect 2484 3084 2516 3085
rect 2484 3004 2516 3036
rect 2484 2955 2516 2956
rect 2484 2925 2485 2955
rect 2485 2925 2515 2955
rect 2515 2925 2516 2955
rect 2484 2924 2516 2925
rect 2484 2844 2516 2876
rect 2484 2795 2516 2796
rect 2484 2765 2485 2795
rect 2485 2765 2515 2795
rect 2515 2765 2516 2795
rect 2484 2764 2516 2765
rect 2484 2715 2516 2716
rect 2484 2685 2485 2715
rect 2485 2685 2515 2715
rect 2515 2685 2516 2715
rect 2484 2684 2516 2685
rect 2484 2604 2516 2636
rect 2484 2555 2516 2556
rect 2484 2525 2485 2555
rect 2485 2525 2515 2555
rect 2515 2525 2516 2555
rect 2484 2524 2516 2525
rect 2564 3595 2596 3596
rect 2564 3565 2565 3595
rect 2565 3565 2595 3595
rect 2595 3565 2596 3595
rect 2564 3564 2596 3565
rect 2564 3515 2596 3516
rect 2564 3485 2565 3515
rect 2565 3485 2595 3515
rect 2595 3485 2596 3515
rect 2564 3484 2596 3485
rect 2564 3404 2596 3436
rect 2564 3355 2596 3356
rect 2564 3325 2565 3355
rect 2565 3325 2595 3355
rect 2595 3325 2596 3355
rect 2564 3324 2596 3325
rect 2564 3275 2596 3276
rect 2564 3245 2565 3275
rect 2565 3245 2595 3275
rect 2595 3245 2596 3275
rect 2564 3244 2596 3245
rect 2564 3195 2596 3196
rect 2564 3165 2565 3195
rect 2565 3165 2595 3195
rect 2595 3165 2596 3195
rect 2564 3164 2596 3165
rect 2564 3115 2596 3116
rect 2564 3085 2565 3115
rect 2565 3085 2595 3115
rect 2595 3085 2596 3115
rect 2564 3084 2596 3085
rect 2564 3004 2596 3036
rect 2564 2955 2596 2956
rect 2564 2925 2565 2955
rect 2565 2925 2595 2955
rect 2595 2925 2596 2955
rect 2564 2924 2596 2925
rect 2564 2844 2596 2876
rect 2564 2795 2596 2796
rect 2564 2765 2565 2795
rect 2565 2765 2595 2795
rect 2595 2765 2596 2795
rect 2564 2764 2596 2765
rect 2564 2715 2596 2716
rect 2564 2685 2565 2715
rect 2565 2685 2595 2715
rect 2595 2685 2596 2715
rect 2564 2684 2596 2685
rect 2564 2604 2596 2636
rect 2564 2555 2596 2556
rect 2564 2525 2565 2555
rect 2565 2525 2595 2555
rect 2595 2525 2596 2555
rect 2564 2524 2596 2525
rect 2644 3595 2676 3596
rect 2644 3565 2645 3595
rect 2645 3565 2675 3595
rect 2675 3565 2676 3595
rect 2644 3564 2676 3565
rect 2644 3515 2676 3516
rect 2644 3485 2645 3515
rect 2645 3485 2675 3515
rect 2675 3485 2676 3515
rect 2644 3484 2676 3485
rect 2644 3404 2676 3436
rect 2644 3355 2676 3356
rect 2644 3325 2645 3355
rect 2645 3325 2675 3355
rect 2675 3325 2676 3355
rect 2644 3324 2676 3325
rect 2644 3275 2676 3276
rect 2644 3245 2645 3275
rect 2645 3245 2675 3275
rect 2675 3245 2676 3275
rect 2644 3244 2676 3245
rect 2644 3195 2676 3196
rect 2644 3165 2645 3195
rect 2645 3165 2675 3195
rect 2675 3165 2676 3195
rect 2644 3164 2676 3165
rect 2644 3115 2676 3116
rect 2644 3085 2645 3115
rect 2645 3085 2675 3115
rect 2675 3085 2676 3115
rect 2644 3084 2676 3085
rect 2644 3004 2676 3036
rect 2644 2955 2676 2956
rect 2644 2925 2645 2955
rect 2645 2925 2675 2955
rect 2675 2925 2676 2955
rect 2644 2924 2676 2925
rect 2644 2844 2676 2876
rect 2644 2795 2676 2796
rect 2644 2765 2645 2795
rect 2645 2765 2675 2795
rect 2675 2765 2676 2795
rect 2644 2764 2676 2765
rect 2644 2715 2676 2716
rect 2644 2685 2645 2715
rect 2645 2685 2675 2715
rect 2675 2685 2676 2715
rect 2644 2684 2676 2685
rect 2644 2604 2676 2636
rect 2644 2555 2676 2556
rect 2644 2525 2645 2555
rect 2645 2525 2675 2555
rect 2675 2525 2676 2555
rect 2644 2524 2676 2525
rect 2724 3595 2756 3596
rect 2724 3565 2725 3595
rect 2725 3565 2755 3595
rect 2755 3565 2756 3595
rect 2724 3564 2756 3565
rect 2724 3515 2756 3516
rect 2724 3485 2725 3515
rect 2725 3485 2755 3515
rect 2755 3485 2756 3515
rect 2724 3484 2756 3485
rect 2724 3404 2756 3436
rect 2724 3355 2756 3356
rect 2724 3325 2725 3355
rect 2725 3325 2755 3355
rect 2755 3325 2756 3355
rect 2724 3324 2756 3325
rect 2724 3275 2756 3276
rect 2724 3245 2725 3275
rect 2725 3245 2755 3275
rect 2755 3245 2756 3275
rect 2724 3244 2756 3245
rect 2724 3195 2756 3196
rect 2724 3165 2725 3195
rect 2725 3165 2755 3195
rect 2755 3165 2756 3195
rect 2724 3164 2756 3165
rect 2724 3115 2756 3116
rect 2724 3085 2725 3115
rect 2725 3085 2755 3115
rect 2755 3085 2756 3115
rect 2724 3084 2756 3085
rect 2724 3004 2756 3036
rect 2724 2955 2756 2956
rect 2724 2925 2725 2955
rect 2725 2925 2755 2955
rect 2755 2925 2756 2955
rect 2724 2924 2756 2925
rect 2724 2844 2756 2876
rect 2724 2795 2756 2796
rect 2724 2765 2725 2795
rect 2725 2765 2755 2795
rect 2755 2765 2756 2795
rect 2724 2764 2756 2765
rect 2724 2715 2756 2716
rect 2724 2685 2725 2715
rect 2725 2685 2755 2715
rect 2755 2685 2756 2715
rect 2724 2684 2756 2685
rect 2724 2604 2756 2636
rect 2724 2555 2756 2556
rect 2724 2525 2725 2555
rect 2725 2525 2755 2555
rect 2755 2525 2756 2555
rect 2724 2524 2756 2525
rect 2804 3595 2836 3596
rect 2804 3565 2805 3595
rect 2805 3565 2835 3595
rect 2835 3565 2836 3595
rect 2804 3564 2836 3565
rect 2804 3515 2836 3516
rect 2804 3485 2805 3515
rect 2805 3485 2835 3515
rect 2835 3485 2836 3515
rect 2804 3484 2836 3485
rect 2804 3404 2836 3436
rect 2804 3355 2836 3356
rect 2804 3325 2805 3355
rect 2805 3325 2835 3355
rect 2835 3325 2836 3355
rect 2804 3324 2836 3325
rect 2804 3275 2836 3276
rect 2804 3245 2805 3275
rect 2805 3245 2835 3275
rect 2835 3245 2836 3275
rect 2804 3244 2836 3245
rect 2804 3195 2836 3196
rect 2804 3165 2805 3195
rect 2805 3165 2835 3195
rect 2835 3165 2836 3195
rect 2804 3164 2836 3165
rect 2804 3115 2836 3116
rect 2804 3085 2805 3115
rect 2805 3085 2835 3115
rect 2835 3085 2836 3115
rect 2804 3084 2836 3085
rect 2804 3004 2836 3036
rect 2804 2955 2836 2956
rect 2804 2925 2805 2955
rect 2805 2925 2835 2955
rect 2835 2925 2836 2955
rect 2804 2924 2836 2925
rect 2804 2844 2836 2876
rect 2804 2795 2836 2796
rect 2804 2765 2805 2795
rect 2805 2765 2835 2795
rect 2835 2765 2836 2795
rect 2804 2764 2836 2765
rect 2804 2715 2836 2716
rect 2804 2685 2805 2715
rect 2805 2685 2835 2715
rect 2835 2685 2836 2715
rect 2804 2684 2836 2685
rect 2804 2604 2836 2636
rect 2804 2555 2836 2556
rect 2804 2525 2805 2555
rect 2805 2525 2835 2555
rect 2835 2525 2836 2555
rect 2804 2524 2836 2525
rect 2884 3595 2916 3596
rect 2884 3565 2885 3595
rect 2885 3565 2915 3595
rect 2915 3565 2916 3595
rect 2884 3564 2916 3565
rect 2884 3515 2916 3516
rect 2884 3485 2885 3515
rect 2885 3485 2915 3515
rect 2915 3485 2916 3515
rect 2884 3484 2916 3485
rect 2884 3404 2916 3436
rect 2884 3355 2916 3356
rect 2884 3325 2885 3355
rect 2885 3325 2915 3355
rect 2915 3325 2916 3355
rect 2884 3324 2916 3325
rect 2884 3275 2916 3276
rect 2884 3245 2885 3275
rect 2885 3245 2915 3275
rect 2915 3245 2916 3275
rect 2884 3244 2916 3245
rect 2884 3195 2916 3196
rect 2884 3165 2885 3195
rect 2885 3165 2915 3195
rect 2915 3165 2916 3195
rect 2884 3164 2916 3165
rect 2884 3115 2916 3116
rect 2884 3085 2885 3115
rect 2885 3085 2915 3115
rect 2915 3085 2916 3115
rect 2884 3084 2916 3085
rect 2884 3004 2916 3036
rect 2884 2955 2916 2956
rect 2884 2925 2885 2955
rect 2885 2925 2915 2955
rect 2915 2925 2916 2955
rect 2884 2924 2916 2925
rect 2884 2844 2916 2876
rect 2884 2795 2916 2796
rect 2884 2765 2885 2795
rect 2885 2765 2915 2795
rect 2915 2765 2916 2795
rect 2884 2764 2916 2765
rect 2884 2715 2916 2716
rect 2884 2685 2885 2715
rect 2885 2685 2915 2715
rect 2915 2685 2916 2715
rect 2884 2684 2916 2685
rect 2884 2604 2916 2636
rect 2884 2555 2916 2556
rect 2884 2525 2885 2555
rect 2885 2525 2915 2555
rect 2915 2525 2916 2555
rect 2884 2524 2916 2525
rect 2964 3595 2996 3596
rect 2964 3565 2965 3595
rect 2965 3565 2995 3595
rect 2995 3565 2996 3595
rect 2964 3564 2996 3565
rect 2964 3515 2996 3516
rect 2964 3485 2965 3515
rect 2965 3485 2995 3515
rect 2995 3485 2996 3515
rect 2964 3484 2996 3485
rect 2964 3404 2996 3436
rect 2964 3355 2996 3356
rect 2964 3325 2965 3355
rect 2965 3325 2995 3355
rect 2995 3325 2996 3355
rect 2964 3324 2996 3325
rect 2964 3275 2996 3276
rect 2964 3245 2965 3275
rect 2965 3245 2995 3275
rect 2995 3245 2996 3275
rect 2964 3244 2996 3245
rect 2964 3195 2996 3196
rect 2964 3165 2965 3195
rect 2965 3165 2995 3195
rect 2995 3165 2996 3195
rect 2964 3164 2996 3165
rect 2964 3115 2996 3116
rect 2964 3085 2965 3115
rect 2965 3085 2995 3115
rect 2995 3085 2996 3115
rect 2964 3084 2996 3085
rect 2964 3004 2996 3036
rect 2964 2955 2996 2956
rect 2964 2925 2965 2955
rect 2965 2925 2995 2955
rect 2995 2925 2996 2955
rect 2964 2924 2996 2925
rect 2964 2844 2996 2876
rect 2964 2795 2996 2796
rect 2964 2765 2965 2795
rect 2965 2765 2995 2795
rect 2995 2765 2996 2795
rect 2964 2764 2996 2765
rect 2964 2715 2996 2716
rect 2964 2685 2965 2715
rect 2965 2685 2995 2715
rect 2995 2685 2996 2715
rect 2964 2684 2996 2685
rect 2964 2604 2996 2636
rect 2964 2555 2996 2556
rect 2964 2525 2965 2555
rect 2965 2525 2995 2555
rect 2995 2525 2996 2555
rect 2964 2524 2996 2525
rect 3044 3595 3076 3596
rect 3044 3565 3045 3595
rect 3045 3565 3075 3595
rect 3075 3565 3076 3595
rect 3044 3564 3076 3565
rect 3044 3515 3076 3516
rect 3044 3485 3045 3515
rect 3045 3485 3075 3515
rect 3075 3485 3076 3515
rect 3044 3484 3076 3485
rect 3044 3404 3076 3436
rect 3044 3355 3076 3356
rect 3044 3325 3045 3355
rect 3045 3325 3075 3355
rect 3075 3325 3076 3355
rect 3044 3324 3076 3325
rect 3044 3275 3076 3276
rect 3044 3245 3045 3275
rect 3045 3245 3075 3275
rect 3075 3245 3076 3275
rect 3044 3244 3076 3245
rect 3044 3195 3076 3196
rect 3044 3165 3045 3195
rect 3045 3165 3075 3195
rect 3075 3165 3076 3195
rect 3044 3164 3076 3165
rect 3044 3115 3076 3116
rect 3044 3085 3045 3115
rect 3045 3085 3075 3115
rect 3075 3085 3076 3115
rect 3044 3084 3076 3085
rect 3044 3004 3076 3036
rect 3044 2955 3076 2956
rect 3044 2925 3045 2955
rect 3045 2925 3075 2955
rect 3075 2925 3076 2955
rect 3044 2924 3076 2925
rect 3044 2844 3076 2876
rect 3044 2795 3076 2796
rect 3044 2765 3045 2795
rect 3045 2765 3075 2795
rect 3075 2765 3076 2795
rect 3044 2764 3076 2765
rect 3044 2715 3076 2716
rect 3044 2685 3045 2715
rect 3045 2685 3075 2715
rect 3075 2685 3076 2715
rect 3044 2684 3076 2685
rect 3044 2604 3076 2636
rect 3044 2555 3076 2556
rect 3044 2525 3045 2555
rect 3045 2525 3075 2555
rect 3075 2525 3076 2555
rect 3044 2524 3076 2525
rect 3124 3595 3156 3596
rect 3124 3565 3125 3595
rect 3125 3565 3155 3595
rect 3155 3565 3156 3595
rect 3124 3564 3156 3565
rect 3124 3515 3156 3516
rect 3124 3485 3125 3515
rect 3125 3485 3155 3515
rect 3155 3485 3156 3515
rect 3124 3484 3156 3485
rect 3124 3404 3156 3436
rect 3124 3355 3156 3356
rect 3124 3325 3125 3355
rect 3125 3325 3155 3355
rect 3155 3325 3156 3355
rect 3124 3324 3156 3325
rect 3124 3275 3156 3276
rect 3124 3245 3125 3275
rect 3125 3245 3155 3275
rect 3155 3245 3156 3275
rect 3124 3244 3156 3245
rect 3124 3195 3156 3196
rect 3124 3165 3125 3195
rect 3125 3165 3155 3195
rect 3155 3165 3156 3195
rect 3124 3164 3156 3165
rect 3124 3115 3156 3116
rect 3124 3085 3125 3115
rect 3125 3085 3155 3115
rect 3155 3085 3156 3115
rect 3124 3084 3156 3085
rect 3124 3004 3156 3036
rect 3124 2955 3156 2956
rect 3124 2925 3125 2955
rect 3125 2925 3155 2955
rect 3155 2925 3156 2955
rect 3124 2924 3156 2925
rect 3124 2844 3156 2876
rect 3124 2795 3156 2796
rect 3124 2765 3125 2795
rect 3125 2765 3155 2795
rect 3155 2765 3156 2795
rect 3124 2764 3156 2765
rect 3124 2715 3156 2716
rect 3124 2685 3125 2715
rect 3125 2685 3155 2715
rect 3155 2685 3156 2715
rect 3124 2684 3156 2685
rect 3124 2604 3156 2636
rect 3124 2555 3156 2556
rect 3124 2525 3125 2555
rect 3125 2525 3155 2555
rect 3155 2525 3156 2555
rect 3124 2524 3156 2525
rect 3204 3595 3236 3596
rect 3204 3565 3205 3595
rect 3205 3565 3235 3595
rect 3235 3565 3236 3595
rect 3204 3564 3236 3565
rect 3204 3515 3236 3516
rect 3204 3485 3205 3515
rect 3205 3485 3235 3515
rect 3235 3485 3236 3515
rect 3204 3484 3236 3485
rect 3204 3404 3236 3436
rect 3204 3355 3236 3356
rect 3204 3325 3205 3355
rect 3205 3325 3235 3355
rect 3235 3325 3236 3355
rect 3204 3324 3236 3325
rect 3204 3275 3236 3276
rect 3204 3245 3205 3275
rect 3205 3245 3235 3275
rect 3235 3245 3236 3275
rect 3204 3244 3236 3245
rect 3204 3195 3236 3196
rect 3204 3165 3205 3195
rect 3205 3165 3235 3195
rect 3235 3165 3236 3195
rect 3204 3164 3236 3165
rect 3204 3115 3236 3116
rect 3204 3085 3205 3115
rect 3205 3085 3235 3115
rect 3235 3085 3236 3115
rect 3204 3084 3236 3085
rect 3204 3004 3236 3036
rect 3204 2955 3236 2956
rect 3204 2925 3205 2955
rect 3205 2925 3235 2955
rect 3235 2925 3236 2955
rect 3204 2924 3236 2925
rect 3204 2844 3236 2876
rect 3204 2795 3236 2796
rect 3204 2765 3205 2795
rect 3205 2765 3235 2795
rect 3235 2765 3236 2795
rect 3204 2764 3236 2765
rect 3204 2715 3236 2716
rect 3204 2685 3205 2715
rect 3205 2685 3235 2715
rect 3235 2685 3236 2715
rect 3204 2684 3236 2685
rect 3204 2604 3236 2636
rect 3204 2555 3236 2556
rect 3204 2525 3205 2555
rect 3205 2525 3235 2555
rect 3235 2525 3236 2555
rect 3204 2524 3236 2525
rect 3284 3595 3316 3596
rect 3284 3565 3285 3595
rect 3285 3565 3315 3595
rect 3315 3565 3316 3595
rect 3284 3564 3316 3565
rect 3284 3515 3316 3516
rect 3284 3485 3285 3515
rect 3285 3485 3315 3515
rect 3315 3485 3316 3515
rect 3284 3484 3316 3485
rect 3284 3404 3316 3436
rect 3284 3355 3316 3356
rect 3284 3325 3285 3355
rect 3285 3325 3315 3355
rect 3315 3325 3316 3355
rect 3284 3324 3316 3325
rect 3284 3275 3316 3276
rect 3284 3245 3285 3275
rect 3285 3245 3315 3275
rect 3315 3245 3316 3275
rect 3284 3244 3316 3245
rect 3284 3195 3316 3196
rect 3284 3165 3285 3195
rect 3285 3165 3315 3195
rect 3315 3165 3316 3195
rect 3284 3164 3316 3165
rect 3284 3115 3316 3116
rect 3284 3085 3285 3115
rect 3285 3085 3315 3115
rect 3315 3085 3316 3115
rect 3284 3084 3316 3085
rect 3284 3004 3316 3036
rect 3284 2955 3316 2956
rect 3284 2925 3285 2955
rect 3285 2925 3315 2955
rect 3315 2925 3316 2955
rect 3284 2924 3316 2925
rect 3284 2844 3316 2876
rect 3284 2795 3316 2796
rect 3284 2765 3285 2795
rect 3285 2765 3315 2795
rect 3315 2765 3316 2795
rect 3284 2764 3316 2765
rect 3284 2715 3316 2716
rect 3284 2685 3285 2715
rect 3285 2685 3315 2715
rect 3315 2685 3316 2715
rect 3284 2684 3316 2685
rect 3284 2604 3316 2636
rect 3284 2555 3316 2556
rect 3284 2525 3285 2555
rect 3285 2525 3315 2555
rect 3315 2525 3316 2555
rect 3284 2524 3316 2525
rect 3364 3595 3396 3596
rect 3364 3565 3365 3595
rect 3365 3565 3395 3595
rect 3395 3565 3396 3595
rect 3364 3564 3396 3565
rect 3364 3515 3396 3516
rect 3364 3485 3365 3515
rect 3365 3485 3395 3515
rect 3395 3485 3396 3515
rect 3364 3484 3396 3485
rect 3364 3404 3396 3436
rect 3364 3355 3396 3356
rect 3364 3325 3365 3355
rect 3365 3325 3395 3355
rect 3395 3325 3396 3355
rect 3364 3324 3396 3325
rect 3364 3275 3396 3276
rect 3364 3245 3365 3275
rect 3365 3245 3395 3275
rect 3395 3245 3396 3275
rect 3364 3244 3396 3245
rect 3364 3195 3396 3196
rect 3364 3165 3365 3195
rect 3365 3165 3395 3195
rect 3395 3165 3396 3195
rect 3364 3164 3396 3165
rect 3364 3115 3396 3116
rect 3364 3085 3365 3115
rect 3365 3085 3395 3115
rect 3395 3085 3396 3115
rect 3364 3084 3396 3085
rect 3364 3004 3396 3036
rect 3364 2955 3396 2956
rect 3364 2925 3365 2955
rect 3365 2925 3395 2955
rect 3395 2925 3396 2955
rect 3364 2924 3396 2925
rect 3364 2844 3396 2876
rect 3364 2795 3396 2796
rect 3364 2765 3365 2795
rect 3365 2765 3395 2795
rect 3395 2765 3396 2795
rect 3364 2764 3396 2765
rect 3364 2715 3396 2716
rect 3364 2685 3365 2715
rect 3365 2685 3395 2715
rect 3395 2685 3396 2715
rect 3364 2684 3396 2685
rect 3364 2604 3396 2636
rect 3364 2555 3396 2556
rect 3364 2525 3365 2555
rect 3365 2525 3395 2555
rect 3395 2525 3396 2555
rect 3364 2524 3396 2525
rect 3444 3595 3476 3596
rect 3444 3565 3445 3595
rect 3445 3565 3475 3595
rect 3475 3565 3476 3595
rect 3444 3564 3476 3565
rect 3444 3515 3476 3516
rect 3444 3485 3445 3515
rect 3445 3485 3475 3515
rect 3475 3485 3476 3515
rect 3444 3484 3476 3485
rect 3444 3404 3476 3436
rect 3444 3355 3476 3356
rect 3444 3325 3445 3355
rect 3445 3325 3475 3355
rect 3475 3325 3476 3355
rect 3444 3324 3476 3325
rect 3444 3275 3476 3276
rect 3444 3245 3445 3275
rect 3445 3245 3475 3275
rect 3475 3245 3476 3275
rect 3444 3244 3476 3245
rect 3444 3195 3476 3196
rect 3444 3165 3445 3195
rect 3445 3165 3475 3195
rect 3475 3165 3476 3195
rect 3444 3164 3476 3165
rect 3444 3115 3476 3116
rect 3444 3085 3445 3115
rect 3445 3085 3475 3115
rect 3475 3085 3476 3115
rect 3444 3084 3476 3085
rect 3444 3004 3476 3036
rect 3444 2955 3476 2956
rect 3444 2925 3445 2955
rect 3445 2925 3475 2955
rect 3475 2925 3476 2955
rect 3444 2924 3476 2925
rect 3444 2844 3476 2876
rect 3444 2795 3476 2796
rect 3444 2765 3445 2795
rect 3445 2765 3475 2795
rect 3475 2765 3476 2795
rect 3444 2764 3476 2765
rect 3444 2715 3476 2716
rect 3444 2685 3445 2715
rect 3445 2685 3475 2715
rect 3475 2685 3476 2715
rect 3444 2684 3476 2685
rect 3444 2604 3476 2636
rect 3444 2555 3476 2556
rect 3444 2525 3445 2555
rect 3445 2525 3475 2555
rect 3475 2525 3476 2555
rect 3444 2524 3476 2525
rect 3524 3595 3556 3596
rect 3524 3565 3525 3595
rect 3525 3565 3555 3595
rect 3555 3565 3556 3595
rect 3524 3564 3556 3565
rect 3524 3515 3556 3516
rect 3524 3485 3525 3515
rect 3525 3485 3555 3515
rect 3555 3485 3556 3515
rect 3524 3484 3556 3485
rect 3524 3404 3556 3436
rect 3524 3355 3556 3356
rect 3524 3325 3525 3355
rect 3525 3325 3555 3355
rect 3555 3325 3556 3355
rect 3524 3324 3556 3325
rect 3524 3275 3556 3276
rect 3524 3245 3525 3275
rect 3525 3245 3555 3275
rect 3555 3245 3556 3275
rect 3524 3244 3556 3245
rect 3524 3195 3556 3196
rect 3524 3165 3525 3195
rect 3525 3165 3555 3195
rect 3555 3165 3556 3195
rect 3524 3164 3556 3165
rect 3524 3115 3556 3116
rect 3524 3085 3525 3115
rect 3525 3085 3555 3115
rect 3555 3085 3556 3115
rect 3524 3084 3556 3085
rect 3524 3004 3556 3036
rect 3524 2955 3556 2956
rect 3524 2925 3525 2955
rect 3525 2925 3555 2955
rect 3555 2925 3556 2955
rect 3524 2924 3556 2925
rect 3524 2844 3556 2876
rect 3524 2795 3556 2796
rect 3524 2765 3525 2795
rect 3525 2765 3555 2795
rect 3555 2765 3556 2795
rect 3524 2764 3556 2765
rect 3524 2715 3556 2716
rect 3524 2685 3525 2715
rect 3525 2685 3555 2715
rect 3555 2685 3556 2715
rect 3524 2684 3556 2685
rect 3524 2604 3556 2636
rect 3524 2555 3556 2556
rect 3524 2525 3525 2555
rect 3525 2525 3555 2555
rect 3555 2525 3556 2555
rect 3524 2524 3556 2525
rect 3604 3595 3636 3596
rect 3604 3565 3605 3595
rect 3605 3565 3635 3595
rect 3635 3565 3636 3595
rect 3604 3564 3636 3565
rect 3604 3515 3636 3516
rect 3604 3485 3605 3515
rect 3605 3485 3635 3515
rect 3635 3485 3636 3515
rect 3604 3484 3636 3485
rect 3604 3404 3636 3436
rect 3604 3355 3636 3356
rect 3604 3325 3605 3355
rect 3605 3325 3635 3355
rect 3635 3325 3636 3355
rect 3604 3324 3636 3325
rect 3604 3275 3636 3276
rect 3604 3245 3605 3275
rect 3605 3245 3635 3275
rect 3635 3245 3636 3275
rect 3604 3244 3636 3245
rect 3604 3195 3636 3196
rect 3604 3165 3605 3195
rect 3605 3165 3635 3195
rect 3635 3165 3636 3195
rect 3604 3164 3636 3165
rect 3604 3115 3636 3116
rect 3604 3085 3605 3115
rect 3605 3085 3635 3115
rect 3635 3085 3636 3115
rect 3604 3084 3636 3085
rect 3604 3004 3636 3036
rect 3604 2955 3636 2956
rect 3604 2925 3605 2955
rect 3605 2925 3635 2955
rect 3635 2925 3636 2955
rect 3604 2924 3636 2925
rect 3604 2844 3636 2876
rect 3604 2795 3636 2796
rect 3604 2765 3605 2795
rect 3605 2765 3635 2795
rect 3635 2765 3636 2795
rect 3604 2764 3636 2765
rect 3604 2715 3636 2716
rect 3604 2685 3605 2715
rect 3605 2685 3635 2715
rect 3635 2685 3636 2715
rect 3604 2684 3636 2685
rect 3604 2604 3636 2636
rect 3604 2555 3636 2556
rect 3604 2525 3605 2555
rect 3605 2525 3635 2555
rect 3635 2525 3636 2555
rect 3604 2524 3636 2525
rect 3684 3595 3716 3596
rect 3684 3565 3685 3595
rect 3685 3565 3715 3595
rect 3715 3565 3716 3595
rect 3684 3564 3716 3565
rect 3684 3515 3716 3516
rect 3684 3485 3685 3515
rect 3685 3485 3715 3515
rect 3715 3485 3716 3515
rect 3684 3484 3716 3485
rect 3684 3404 3716 3436
rect 3684 3355 3716 3356
rect 3684 3325 3685 3355
rect 3685 3325 3715 3355
rect 3715 3325 3716 3355
rect 3684 3324 3716 3325
rect 3684 3275 3716 3276
rect 3684 3245 3685 3275
rect 3685 3245 3715 3275
rect 3715 3245 3716 3275
rect 3684 3244 3716 3245
rect 3684 3195 3716 3196
rect 3684 3165 3685 3195
rect 3685 3165 3715 3195
rect 3715 3165 3716 3195
rect 3684 3164 3716 3165
rect 3684 3115 3716 3116
rect 3684 3085 3685 3115
rect 3685 3085 3715 3115
rect 3715 3085 3716 3115
rect 3684 3084 3716 3085
rect 3684 3004 3716 3036
rect 3684 2955 3716 2956
rect 3684 2925 3685 2955
rect 3685 2925 3715 2955
rect 3715 2925 3716 2955
rect 3684 2924 3716 2925
rect 3684 2844 3716 2876
rect 3684 2795 3716 2796
rect 3684 2765 3685 2795
rect 3685 2765 3715 2795
rect 3715 2765 3716 2795
rect 3684 2764 3716 2765
rect 3684 2715 3716 2716
rect 3684 2685 3685 2715
rect 3685 2685 3715 2715
rect 3715 2685 3716 2715
rect 3684 2684 3716 2685
rect 3684 2604 3716 2636
rect 3684 2555 3716 2556
rect 3684 2525 3685 2555
rect 3685 2525 3715 2555
rect 3715 2525 3716 2555
rect 3684 2524 3716 2525
rect 3764 3595 3796 3596
rect 3764 3565 3765 3595
rect 3765 3565 3795 3595
rect 3795 3565 3796 3595
rect 3764 3564 3796 3565
rect 3764 3515 3796 3516
rect 3764 3485 3765 3515
rect 3765 3485 3795 3515
rect 3795 3485 3796 3515
rect 3764 3484 3796 3485
rect 3764 3404 3796 3436
rect 3764 3355 3796 3356
rect 3764 3325 3765 3355
rect 3765 3325 3795 3355
rect 3795 3325 3796 3355
rect 3764 3324 3796 3325
rect 3764 3275 3796 3276
rect 3764 3245 3765 3275
rect 3765 3245 3795 3275
rect 3795 3245 3796 3275
rect 3764 3244 3796 3245
rect 3764 3195 3796 3196
rect 3764 3165 3765 3195
rect 3765 3165 3795 3195
rect 3795 3165 3796 3195
rect 3764 3164 3796 3165
rect 3764 3115 3796 3116
rect 3764 3085 3765 3115
rect 3765 3085 3795 3115
rect 3795 3085 3796 3115
rect 3764 3084 3796 3085
rect 3764 3004 3796 3036
rect 3764 2955 3796 2956
rect 3764 2925 3765 2955
rect 3765 2925 3795 2955
rect 3795 2925 3796 2955
rect 3764 2924 3796 2925
rect 3764 2844 3796 2876
rect 3764 2795 3796 2796
rect 3764 2765 3765 2795
rect 3765 2765 3795 2795
rect 3795 2765 3796 2795
rect 3764 2764 3796 2765
rect 3764 2715 3796 2716
rect 3764 2685 3765 2715
rect 3765 2685 3795 2715
rect 3795 2685 3796 2715
rect 3764 2684 3796 2685
rect 3764 2604 3796 2636
rect 3764 2555 3796 2556
rect 3764 2525 3765 2555
rect 3765 2525 3795 2555
rect 3795 2525 3796 2555
rect 3764 2524 3796 2525
rect 3844 3595 3876 3596
rect 3844 3565 3845 3595
rect 3845 3565 3875 3595
rect 3875 3565 3876 3595
rect 3844 3564 3876 3565
rect 3844 3515 3876 3516
rect 3844 3485 3845 3515
rect 3845 3485 3875 3515
rect 3875 3485 3876 3515
rect 3844 3484 3876 3485
rect 3844 3404 3876 3436
rect 3844 3355 3876 3356
rect 3844 3325 3845 3355
rect 3845 3325 3875 3355
rect 3875 3325 3876 3355
rect 3844 3324 3876 3325
rect 3844 3275 3876 3276
rect 3844 3245 3845 3275
rect 3845 3245 3875 3275
rect 3875 3245 3876 3275
rect 3844 3244 3876 3245
rect 3844 3195 3876 3196
rect 3844 3165 3845 3195
rect 3845 3165 3875 3195
rect 3875 3165 3876 3195
rect 3844 3164 3876 3165
rect 3844 3115 3876 3116
rect 3844 3085 3845 3115
rect 3845 3085 3875 3115
rect 3875 3085 3876 3115
rect 3844 3084 3876 3085
rect 3844 3004 3876 3036
rect 3844 2955 3876 2956
rect 3844 2925 3845 2955
rect 3845 2925 3875 2955
rect 3875 2925 3876 2955
rect 3844 2924 3876 2925
rect 3844 2844 3876 2876
rect 3844 2795 3876 2796
rect 3844 2765 3845 2795
rect 3845 2765 3875 2795
rect 3875 2765 3876 2795
rect 3844 2764 3876 2765
rect 3844 2715 3876 2716
rect 3844 2685 3845 2715
rect 3845 2685 3875 2715
rect 3875 2685 3876 2715
rect 3844 2684 3876 2685
rect 3844 2604 3876 2636
rect 3844 2555 3876 2556
rect 3844 2525 3845 2555
rect 3845 2525 3875 2555
rect 3875 2525 3876 2555
rect 3844 2524 3876 2525
rect 3924 3595 3956 3596
rect 3924 3565 3925 3595
rect 3925 3565 3955 3595
rect 3955 3565 3956 3595
rect 3924 3564 3956 3565
rect 3924 3515 3956 3516
rect 3924 3485 3925 3515
rect 3925 3485 3955 3515
rect 3955 3485 3956 3515
rect 3924 3484 3956 3485
rect 3924 3404 3956 3436
rect 3924 3355 3956 3356
rect 3924 3325 3925 3355
rect 3925 3325 3955 3355
rect 3955 3325 3956 3355
rect 3924 3324 3956 3325
rect 3924 3275 3956 3276
rect 3924 3245 3925 3275
rect 3925 3245 3955 3275
rect 3955 3245 3956 3275
rect 3924 3244 3956 3245
rect 3924 3195 3956 3196
rect 3924 3165 3925 3195
rect 3925 3165 3955 3195
rect 3955 3165 3956 3195
rect 3924 3164 3956 3165
rect 3924 3115 3956 3116
rect 3924 3085 3925 3115
rect 3925 3085 3955 3115
rect 3955 3085 3956 3115
rect 3924 3084 3956 3085
rect 3924 3004 3956 3036
rect 3924 2955 3956 2956
rect 3924 2925 3925 2955
rect 3925 2925 3955 2955
rect 3955 2925 3956 2955
rect 3924 2924 3956 2925
rect 3924 2844 3956 2876
rect 3924 2795 3956 2796
rect 3924 2765 3925 2795
rect 3925 2765 3955 2795
rect 3955 2765 3956 2795
rect 3924 2764 3956 2765
rect 3924 2715 3956 2716
rect 3924 2685 3925 2715
rect 3925 2685 3955 2715
rect 3955 2685 3956 2715
rect 3924 2684 3956 2685
rect 3924 2604 3956 2636
rect 3924 2555 3956 2556
rect 3924 2525 3925 2555
rect 3925 2525 3955 2555
rect 3955 2525 3956 2555
rect 3924 2524 3956 2525
rect 4004 3595 4036 3596
rect 4004 3565 4005 3595
rect 4005 3565 4035 3595
rect 4035 3565 4036 3595
rect 4004 3564 4036 3565
rect 4004 3515 4036 3516
rect 4004 3485 4005 3515
rect 4005 3485 4035 3515
rect 4035 3485 4036 3515
rect 4004 3484 4036 3485
rect 4004 3404 4036 3436
rect 4004 3355 4036 3356
rect 4004 3325 4005 3355
rect 4005 3325 4035 3355
rect 4035 3325 4036 3355
rect 4004 3324 4036 3325
rect 4004 3275 4036 3276
rect 4004 3245 4005 3275
rect 4005 3245 4035 3275
rect 4035 3245 4036 3275
rect 4004 3244 4036 3245
rect 4004 3195 4036 3196
rect 4004 3165 4005 3195
rect 4005 3165 4035 3195
rect 4035 3165 4036 3195
rect 4004 3164 4036 3165
rect 4004 3115 4036 3116
rect 4004 3085 4005 3115
rect 4005 3085 4035 3115
rect 4035 3085 4036 3115
rect 4004 3084 4036 3085
rect 4004 3004 4036 3036
rect 4004 2955 4036 2956
rect 4004 2925 4005 2955
rect 4005 2925 4035 2955
rect 4035 2925 4036 2955
rect 4004 2924 4036 2925
rect 4004 2844 4036 2876
rect 4004 2795 4036 2796
rect 4004 2765 4005 2795
rect 4005 2765 4035 2795
rect 4035 2765 4036 2795
rect 4004 2764 4036 2765
rect 4004 2715 4036 2716
rect 4004 2685 4005 2715
rect 4005 2685 4035 2715
rect 4035 2685 4036 2715
rect 4004 2684 4036 2685
rect 4004 2604 4036 2636
rect 4004 2555 4036 2556
rect 4004 2525 4005 2555
rect 4005 2525 4035 2555
rect 4035 2525 4036 2555
rect 4004 2524 4036 2525
rect 4084 3595 4116 3596
rect 4084 3565 4085 3595
rect 4085 3565 4115 3595
rect 4115 3565 4116 3595
rect 4084 3564 4116 3565
rect 4084 3515 4116 3516
rect 4084 3485 4085 3515
rect 4085 3485 4115 3515
rect 4115 3485 4116 3515
rect 4084 3484 4116 3485
rect 4084 3404 4116 3436
rect 4084 3355 4116 3356
rect 4084 3325 4085 3355
rect 4085 3325 4115 3355
rect 4115 3325 4116 3355
rect 4084 3324 4116 3325
rect 4084 3275 4116 3276
rect 4084 3245 4085 3275
rect 4085 3245 4115 3275
rect 4115 3245 4116 3275
rect 4084 3244 4116 3245
rect 4084 3195 4116 3196
rect 4084 3165 4085 3195
rect 4085 3165 4115 3195
rect 4115 3165 4116 3195
rect 4084 3164 4116 3165
rect 4084 3115 4116 3116
rect 4084 3085 4085 3115
rect 4085 3085 4115 3115
rect 4115 3085 4116 3115
rect 4084 3084 4116 3085
rect 4084 3004 4116 3036
rect 4084 2955 4116 2956
rect 4084 2925 4085 2955
rect 4085 2925 4115 2955
rect 4115 2925 4116 2955
rect 4084 2924 4116 2925
rect 4084 2844 4116 2876
rect 4084 2795 4116 2796
rect 4084 2765 4085 2795
rect 4085 2765 4115 2795
rect 4115 2765 4116 2795
rect 4084 2764 4116 2765
rect 4084 2715 4116 2716
rect 4084 2685 4085 2715
rect 4085 2685 4115 2715
rect 4115 2685 4116 2715
rect 4084 2684 4116 2685
rect 4084 2604 4116 2636
rect 4084 2555 4116 2556
rect 4084 2525 4085 2555
rect 4085 2525 4115 2555
rect 4115 2525 4116 2555
rect 4084 2524 4116 2525
rect 4164 3595 4196 3596
rect 4164 3565 4165 3595
rect 4165 3565 4195 3595
rect 4195 3565 4196 3595
rect 4164 3564 4196 3565
rect 4164 3515 4196 3516
rect 4164 3485 4165 3515
rect 4165 3485 4195 3515
rect 4195 3485 4196 3515
rect 4164 3484 4196 3485
rect 4164 3404 4196 3436
rect 4164 3355 4196 3356
rect 4164 3325 4165 3355
rect 4165 3325 4195 3355
rect 4195 3325 4196 3355
rect 4164 3324 4196 3325
rect 4164 3275 4196 3276
rect 4164 3245 4165 3275
rect 4165 3245 4195 3275
rect 4195 3245 4196 3275
rect 4164 3244 4196 3245
rect 4164 3195 4196 3196
rect 4164 3165 4165 3195
rect 4165 3165 4195 3195
rect 4195 3165 4196 3195
rect 4164 3164 4196 3165
rect 4164 3115 4196 3116
rect 4164 3085 4165 3115
rect 4165 3085 4195 3115
rect 4195 3085 4196 3115
rect 4164 3084 4196 3085
rect 4164 3004 4196 3036
rect 4164 2955 4196 2956
rect 4164 2925 4165 2955
rect 4165 2925 4195 2955
rect 4195 2925 4196 2955
rect 4164 2924 4196 2925
rect 4164 2844 4196 2876
rect 4164 2795 4196 2796
rect 4164 2765 4165 2795
rect 4165 2765 4195 2795
rect 4195 2765 4196 2795
rect 4164 2764 4196 2765
rect 4164 2715 4196 2716
rect 4164 2685 4165 2715
rect 4165 2685 4195 2715
rect 4195 2685 4196 2715
rect 4164 2684 4196 2685
rect 4164 2604 4196 2636
rect 4164 2555 4196 2556
rect 4164 2525 4165 2555
rect 4165 2525 4195 2555
rect 4195 2525 4196 2555
rect 4164 2524 4196 2525
rect 4244 3595 4276 3596
rect 4244 3565 4245 3595
rect 4245 3565 4275 3595
rect 4275 3565 4276 3595
rect 4244 3564 4276 3565
rect 4244 3515 4276 3516
rect 4244 3485 4245 3515
rect 4245 3485 4275 3515
rect 4275 3485 4276 3515
rect 4244 3484 4276 3485
rect 4244 3404 4276 3436
rect 4244 3355 4276 3356
rect 4244 3325 4245 3355
rect 4245 3325 4275 3355
rect 4275 3325 4276 3355
rect 4244 3324 4276 3325
rect 4244 3275 4276 3276
rect 4244 3245 4245 3275
rect 4245 3245 4275 3275
rect 4275 3245 4276 3275
rect 4244 3244 4276 3245
rect 4244 3195 4276 3196
rect 4244 3165 4245 3195
rect 4245 3165 4275 3195
rect 4275 3165 4276 3195
rect 4244 3164 4276 3165
rect 4244 3115 4276 3116
rect 4244 3085 4245 3115
rect 4245 3085 4275 3115
rect 4275 3085 4276 3115
rect 4244 3084 4276 3085
rect 4244 3004 4276 3036
rect 4244 2955 4276 2956
rect 4244 2925 4245 2955
rect 4245 2925 4275 2955
rect 4275 2925 4276 2955
rect 4244 2924 4276 2925
rect 4244 2844 4276 2876
rect 4244 2795 4276 2796
rect 4244 2765 4245 2795
rect 4245 2765 4275 2795
rect 4275 2765 4276 2795
rect 4244 2764 4276 2765
rect 4244 2715 4276 2716
rect 4244 2685 4245 2715
rect 4245 2685 4275 2715
rect 4275 2685 4276 2715
rect 4244 2684 4276 2685
rect 4244 2604 4276 2636
rect 4244 2555 4276 2556
rect 4244 2525 4245 2555
rect 4245 2525 4275 2555
rect 4275 2525 4276 2555
rect 4244 2524 4276 2525
rect 4324 3595 4356 3596
rect 4324 3565 4325 3595
rect 4325 3565 4355 3595
rect 4355 3565 4356 3595
rect 4324 3564 4356 3565
rect 4324 3515 4356 3516
rect 4324 3485 4325 3515
rect 4325 3485 4355 3515
rect 4355 3485 4356 3515
rect 4324 3484 4356 3485
rect 4324 3404 4356 3436
rect 4324 3355 4356 3356
rect 4324 3325 4325 3355
rect 4325 3325 4355 3355
rect 4355 3325 4356 3355
rect 4324 3324 4356 3325
rect 4324 3275 4356 3276
rect 4324 3245 4325 3275
rect 4325 3245 4355 3275
rect 4355 3245 4356 3275
rect 4324 3244 4356 3245
rect 4324 3195 4356 3196
rect 4324 3165 4325 3195
rect 4325 3165 4355 3195
rect 4355 3165 4356 3195
rect 4324 3164 4356 3165
rect 4324 3115 4356 3116
rect 4324 3085 4325 3115
rect 4325 3085 4355 3115
rect 4355 3085 4356 3115
rect 4324 3084 4356 3085
rect 4324 3004 4356 3036
rect 4324 2955 4356 2956
rect 4324 2925 4325 2955
rect 4325 2925 4355 2955
rect 4355 2925 4356 2955
rect 4324 2924 4356 2925
rect 4324 2844 4356 2876
rect 4324 2795 4356 2796
rect 4324 2765 4325 2795
rect 4325 2765 4355 2795
rect 4355 2765 4356 2795
rect 4324 2764 4356 2765
rect 4324 2715 4356 2716
rect 4324 2685 4325 2715
rect 4325 2685 4355 2715
rect 4355 2685 4356 2715
rect 4324 2684 4356 2685
rect 4324 2604 4356 2636
rect 4324 2555 4356 2556
rect 4324 2525 4325 2555
rect 4325 2525 4355 2555
rect 4355 2525 4356 2555
rect 4324 2524 4356 2525
rect 4404 3595 4436 3596
rect 4404 3565 4405 3595
rect 4405 3565 4435 3595
rect 4435 3565 4436 3595
rect 4404 3564 4436 3565
rect 4404 3515 4436 3516
rect 4404 3485 4405 3515
rect 4405 3485 4435 3515
rect 4435 3485 4436 3515
rect 4404 3484 4436 3485
rect 4404 3404 4436 3436
rect 4404 3355 4436 3356
rect 4404 3325 4405 3355
rect 4405 3325 4435 3355
rect 4435 3325 4436 3355
rect 4404 3324 4436 3325
rect 4404 3275 4436 3276
rect 4404 3245 4405 3275
rect 4405 3245 4435 3275
rect 4435 3245 4436 3275
rect 4404 3244 4436 3245
rect 4404 3195 4436 3196
rect 4404 3165 4405 3195
rect 4405 3165 4435 3195
rect 4435 3165 4436 3195
rect 4404 3164 4436 3165
rect 4404 3115 4436 3116
rect 4404 3085 4405 3115
rect 4405 3085 4435 3115
rect 4435 3085 4436 3115
rect 4404 3084 4436 3085
rect 4404 3004 4436 3036
rect 4404 2955 4436 2956
rect 4404 2925 4405 2955
rect 4405 2925 4435 2955
rect 4435 2925 4436 2955
rect 4404 2924 4436 2925
rect 4404 2844 4436 2876
rect 4404 2795 4436 2796
rect 4404 2765 4405 2795
rect 4405 2765 4435 2795
rect 4435 2765 4436 2795
rect 4404 2764 4436 2765
rect 4404 2715 4436 2716
rect 4404 2685 4405 2715
rect 4405 2685 4435 2715
rect 4435 2685 4436 2715
rect 4404 2684 4436 2685
rect 4404 2604 4436 2636
rect 4404 2555 4436 2556
rect 4404 2525 4405 2555
rect 4405 2525 4435 2555
rect 4435 2525 4436 2555
rect 4404 2524 4436 2525
rect 4484 3595 4516 3596
rect 4484 3565 4485 3595
rect 4485 3565 4515 3595
rect 4515 3565 4516 3595
rect 4484 3564 4516 3565
rect 4484 3515 4516 3516
rect 4484 3485 4485 3515
rect 4485 3485 4515 3515
rect 4515 3485 4516 3515
rect 4484 3484 4516 3485
rect 4484 3404 4516 3436
rect 4484 3355 4516 3356
rect 4484 3325 4485 3355
rect 4485 3325 4515 3355
rect 4515 3325 4516 3355
rect 4484 3324 4516 3325
rect 4484 3275 4516 3276
rect 4484 3245 4485 3275
rect 4485 3245 4515 3275
rect 4515 3245 4516 3275
rect 4484 3244 4516 3245
rect 4484 3195 4516 3196
rect 4484 3165 4485 3195
rect 4485 3165 4515 3195
rect 4515 3165 4516 3195
rect 4484 3164 4516 3165
rect 4484 3115 4516 3116
rect 4484 3085 4485 3115
rect 4485 3085 4515 3115
rect 4515 3085 4516 3115
rect 4484 3084 4516 3085
rect 4484 3004 4516 3036
rect 4484 2955 4516 2956
rect 4484 2925 4485 2955
rect 4485 2925 4515 2955
rect 4515 2925 4516 2955
rect 4484 2924 4516 2925
rect 4484 2844 4516 2876
rect 4484 2795 4516 2796
rect 4484 2765 4485 2795
rect 4485 2765 4515 2795
rect 4515 2765 4516 2795
rect 4484 2764 4516 2765
rect 4484 2715 4516 2716
rect 4484 2685 4485 2715
rect 4485 2685 4515 2715
rect 4515 2685 4516 2715
rect 4484 2684 4516 2685
rect 4484 2604 4516 2636
rect 4484 2555 4516 2556
rect 4484 2525 4485 2555
rect 4485 2525 4515 2555
rect 4515 2525 4516 2555
rect 4484 2524 4516 2525
rect 4564 3595 4596 3596
rect 4564 3565 4565 3595
rect 4565 3565 4595 3595
rect 4595 3565 4596 3595
rect 4564 3564 4596 3565
rect 4564 3515 4596 3516
rect 4564 3485 4565 3515
rect 4565 3485 4595 3515
rect 4595 3485 4596 3515
rect 4564 3484 4596 3485
rect 4564 3404 4596 3436
rect 4564 3355 4596 3356
rect 4564 3325 4565 3355
rect 4565 3325 4595 3355
rect 4595 3325 4596 3355
rect 4564 3324 4596 3325
rect 4564 3275 4596 3276
rect 4564 3245 4565 3275
rect 4565 3245 4595 3275
rect 4595 3245 4596 3275
rect 4564 3244 4596 3245
rect 4564 3195 4596 3196
rect 4564 3165 4565 3195
rect 4565 3165 4595 3195
rect 4595 3165 4596 3195
rect 4564 3164 4596 3165
rect 4564 3115 4596 3116
rect 4564 3085 4565 3115
rect 4565 3085 4595 3115
rect 4595 3085 4596 3115
rect 4564 3084 4596 3085
rect 4564 3004 4596 3036
rect 4564 2955 4596 2956
rect 4564 2925 4565 2955
rect 4565 2925 4595 2955
rect 4595 2925 4596 2955
rect 4564 2924 4596 2925
rect 4564 2844 4596 2876
rect 4564 2795 4596 2796
rect 4564 2765 4565 2795
rect 4565 2765 4595 2795
rect 4595 2765 4596 2795
rect 4564 2764 4596 2765
rect 4564 2715 4596 2716
rect 4564 2685 4565 2715
rect 4565 2685 4595 2715
rect 4595 2685 4596 2715
rect 4564 2684 4596 2685
rect 4564 2604 4596 2636
rect 4564 2555 4596 2556
rect 4564 2525 4565 2555
rect 4565 2525 4595 2555
rect 4595 2525 4596 2555
rect 4564 2524 4596 2525
rect 4644 3595 4676 3596
rect 4644 3565 4645 3595
rect 4645 3565 4675 3595
rect 4675 3565 4676 3595
rect 4644 3564 4676 3565
rect 4644 3515 4676 3516
rect 4644 3485 4645 3515
rect 4645 3485 4675 3515
rect 4675 3485 4676 3515
rect 4644 3484 4676 3485
rect 4644 3404 4676 3436
rect 4644 3355 4676 3356
rect 4644 3325 4645 3355
rect 4645 3325 4675 3355
rect 4675 3325 4676 3355
rect 4644 3324 4676 3325
rect 4644 3275 4676 3276
rect 4644 3245 4645 3275
rect 4645 3245 4675 3275
rect 4675 3245 4676 3275
rect 4644 3244 4676 3245
rect 4644 3195 4676 3196
rect 4644 3165 4645 3195
rect 4645 3165 4675 3195
rect 4675 3165 4676 3195
rect 4644 3164 4676 3165
rect 4644 3115 4676 3116
rect 4644 3085 4645 3115
rect 4645 3085 4675 3115
rect 4675 3085 4676 3115
rect 4644 3084 4676 3085
rect 4644 3004 4676 3036
rect 4644 2955 4676 2956
rect 4644 2925 4645 2955
rect 4645 2925 4675 2955
rect 4675 2925 4676 2955
rect 4644 2924 4676 2925
rect 4644 2844 4676 2876
rect 4644 2795 4676 2796
rect 4644 2765 4645 2795
rect 4645 2765 4675 2795
rect 4675 2765 4676 2795
rect 4644 2764 4676 2765
rect 4644 2715 4676 2716
rect 4644 2685 4645 2715
rect 4645 2685 4675 2715
rect 4675 2685 4676 2715
rect 4644 2684 4676 2685
rect 4644 2604 4676 2636
rect 4644 2555 4676 2556
rect 4644 2525 4645 2555
rect 4645 2525 4675 2555
rect 4675 2525 4676 2555
rect 4644 2524 4676 2525
rect 4724 3595 4756 3596
rect 4724 3565 4725 3595
rect 4725 3565 4755 3595
rect 4755 3565 4756 3595
rect 4724 3564 4756 3565
rect 4724 3515 4756 3516
rect 4724 3485 4725 3515
rect 4725 3485 4755 3515
rect 4755 3485 4756 3515
rect 4724 3484 4756 3485
rect 4724 3404 4756 3436
rect 4724 3355 4756 3356
rect 4724 3325 4725 3355
rect 4725 3325 4755 3355
rect 4755 3325 4756 3355
rect 4724 3324 4756 3325
rect 4724 3275 4756 3276
rect 4724 3245 4725 3275
rect 4725 3245 4755 3275
rect 4755 3245 4756 3275
rect 4724 3244 4756 3245
rect 4724 3195 4756 3196
rect 4724 3165 4725 3195
rect 4725 3165 4755 3195
rect 4755 3165 4756 3195
rect 4724 3164 4756 3165
rect 4724 3115 4756 3116
rect 4724 3085 4725 3115
rect 4725 3085 4755 3115
rect 4755 3085 4756 3115
rect 4724 3084 4756 3085
rect 4724 3004 4756 3036
rect 4724 2955 4756 2956
rect 4724 2925 4725 2955
rect 4725 2925 4755 2955
rect 4755 2925 4756 2955
rect 4724 2924 4756 2925
rect 4724 2844 4756 2876
rect 4724 2795 4756 2796
rect 4724 2765 4725 2795
rect 4725 2765 4755 2795
rect 4755 2765 4756 2795
rect 4724 2764 4756 2765
rect 4724 2715 4756 2716
rect 4724 2685 4725 2715
rect 4725 2685 4755 2715
rect 4755 2685 4756 2715
rect 4724 2684 4756 2685
rect 4724 2604 4756 2636
rect 4724 2555 4756 2556
rect 4724 2525 4725 2555
rect 4725 2525 4755 2555
rect 4755 2525 4756 2555
rect 4724 2524 4756 2525
rect 4804 3595 4836 3596
rect 4804 3565 4805 3595
rect 4805 3565 4835 3595
rect 4835 3565 4836 3595
rect 4804 3564 4836 3565
rect 4804 3515 4836 3516
rect 4804 3485 4805 3515
rect 4805 3485 4835 3515
rect 4835 3485 4836 3515
rect 4804 3484 4836 3485
rect 4804 3404 4836 3436
rect 4804 3355 4836 3356
rect 4804 3325 4805 3355
rect 4805 3325 4835 3355
rect 4835 3325 4836 3355
rect 4804 3324 4836 3325
rect 4804 3275 4836 3276
rect 4804 3245 4805 3275
rect 4805 3245 4835 3275
rect 4835 3245 4836 3275
rect 4804 3244 4836 3245
rect 4804 3195 4836 3196
rect 4804 3165 4805 3195
rect 4805 3165 4835 3195
rect 4835 3165 4836 3195
rect 4804 3164 4836 3165
rect 4804 3115 4836 3116
rect 4804 3085 4805 3115
rect 4805 3085 4835 3115
rect 4835 3085 4836 3115
rect 4804 3084 4836 3085
rect 4804 3004 4836 3036
rect 4804 2955 4836 2956
rect 4804 2925 4805 2955
rect 4805 2925 4835 2955
rect 4835 2925 4836 2955
rect 4804 2924 4836 2925
rect 4804 2844 4836 2876
rect 4804 2795 4836 2796
rect 4804 2765 4805 2795
rect 4805 2765 4835 2795
rect 4835 2765 4836 2795
rect 4804 2764 4836 2765
rect 4804 2715 4836 2716
rect 4804 2685 4805 2715
rect 4805 2685 4835 2715
rect 4835 2685 4836 2715
rect 4804 2684 4836 2685
rect 4804 2604 4836 2636
rect 4804 2555 4836 2556
rect 4804 2525 4805 2555
rect 4805 2525 4835 2555
rect 4835 2525 4836 2555
rect 4804 2524 4836 2525
rect 4884 3595 4916 3596
rect 4884 3565 4885 3595
rect 4885 3565 4915 3595
rect 4915 3565 4916 3595
rect 4884 3564 4916 3565
rect 4884 3515 4916 3516
rect 4884 3485 4885 3515
rect 4885 3485 4915 3515
rect 4915 3485 4916 3515
rect 4884 3484 4916 3485
rect 4884 3435 4916 3436
rect 4884 3405 4885 3435
rect 4885 3405 4915 3435
rect 4915 3405 4916 3435
rect 4884 3404 4916 3405
rect 4884 3355 4916 3356
rect 4884 3325 4885 3355
rect 4885 3325 4915 3355
rect 4915 3325 4916 3355
rect 4884 3324 4916 3325
rect 4884 3275 4916 3276
rect 4884 3245 4885 3275
rect 4885 3245 4915 3275
rect 4915 3245 4916 3275
rect 4884 3244 4916 3245
rect 4884 3195 4916 3196
rect 4884 3165 4885 3195
rect 4885 3165 4915 3195
rect 4915 3165 4916 3195
rect 4884 3164 4916 3165
rect 4884 3115 4916 3116
rect 4884 3085 4885 3115
rect 4885 3085 4915 3115
rect 4915 3085 4916 3115
rect 4884 3084 4916 3085
rect 4884 3035 4916 3036
rect 4884 3005 4885 3035
rect 4885 3005 4915 3035
rect 4915 3005 4916 3035
rect 4884 3004 4916 3005
rect 4884 2955 4916 2956
rect 4884 2925 4885 2955
rect 4885 2925 4915 2955
rect 4915 2925 4916 2955
rect 4884 2924 4916 2925
rect 4884 2875 4916 2876
rect 4884 2845 4885 2875
rect 4885 2845 4915 2875
rect 4915 2845 4916 2875
rect 4884 2844 4916 2845
rect 4884 2795 4916 2796
rect 4884 2765 4885 2795
rect 4885 2765 4915 2795
rect 4915 2765 4916 2795
rect 4884 2764 4916 2765
rect 4884 2715 4916 2716
rect 4884 2685 4885 2715
rect 4885 2685 4915 2715
rect 4915 2685 4916 2715
rect 4884 2684 4916 2685
rect 4884 2635 4916 2636
rect 4884 2605 4885 2635
rect 4885 2605 4915 2635
rect 4915 2605 4916 2635
rect 4884 2604 4916 2605
rect 4884 2555 4916 2556
rect 4884 2525 4885 2555
rect 4885 2525 4915 2555
rect 4915 2525 4916 2555
rect 4884 2524 4916 2525
rect -876 2475 -844 2476
rect -876 2445 -875 2475
rect -875 2445 -845 2475
rect -845 2445 -844 2475
rect -876 2444 -844 2445
rect -876 2395 -844 2396
rect -876 2365 -875 2395
rect -875 2365 -845 2395
rect -845 2365 -844 2395
rect -876 2364 -844 2365
rect -876 2315 -844 2316
rect -876 2285 -875 2315
rect -875 2285 -845 2315
rect -845 2285 -844 2315
rect -876 2284 -844 2285
rect -876 2235 -844 2236
rect -876 2205 -875 2235
rect -875 2205 -845 2235
rect -845 2205 -844 2235
rect -876 2204 -844 2205
rect -876 2155 -844 2156
rect -876 2125 -875 2155
rect -875 2125 -845 2155
rect -845 2125 -844 2155
rect -876 2124 -844 2125
rect -876 2075 -844 2076
rect -876 2045 -875 2075
rect -875 2045 -845 2075
rect -845 2045 -844 2075
rect -876 2044 -844 2045
rect -876 1995 -844 1996
rect -876 1965 -875 1995
rect -875 1965 -845 1995
rect -845 1965 -844 1995
rect -876 1964 -844 1965
rect -876 1915 -844 1916
rect -876 1885 -875 1915
rect -875 1885 -845 1915
rect -845 1885 -844 1915
rect -876 1884 -844 1885
rect -876 1835 -844 1836
rect -876 1805 -875 1835
rect -875 1805 -845 1835
rect -845 1805 -844 1835
rect -876 1804 -844 1805
rect -876 1755 -844 1756
rect -876 1725 -875 1755
rect -875 1725 -845 1755
rect -845 1725 -844 1755
rect -876 1724 -844 1725
rect -796 2475 -764 2476
rect -796 2445 -795 2475
rect -795 2445 -765 2475
rect -765 2445 -764 2475
rect -796 2444 -764 2445
rect -796 2364 -764 2396
rect -796 2315 -764 2316
rect -796 2285 -795 2315
rect -795 2285 -765 2315
rect -765 2285 -764 2315
rect -796 2284 -764 2285
rect -796 2204 -764 2236
rect -796 2155 -764 2156
rect -796 2125 -795 2155
rect -795 2125 -765 2155
rect -765 2125 -764 2155
rect -796 2124 -764 2125
rect -796 2075 -764 2076
rect -796 2045 -795 2075
rect -795 2045 -765 2075
rect -765 2045 -764 2075
rect -796 2044 -764 2045
rect -796 1995 -764 1996
rect -796 1965 -795 1995
rect -795 1965 -765 1995
rect -765 1965 -764 1995
rect -796 1964 -764 1965
rect -796 1915 -764 1916
rect -796 1885 -795 1915
rect -795 1885 -765 1915
rect -765 1885 -764 1915
rect -796 1884 -764 1885
rect -796 1835 -764 1836
rect -796 1805 -795 1835
rect -795 1805 -765 1835
rect -765 1805 -764 1835
rect -796 1804 -764 1805
rect -796 1755 -764 1756
rect -796 1725 -795 1755
rect -795 1725 -765 1755
rect -765 1725 -764 1755
rect -796 1724 -764 1725
rect -716 2475 -684 2476
rect -716 2445 -715 2475
rect -715 2445 -685 2475
rect -685 2445 -684 2475
rect -716 2444 -684 2445
rect -716 2364 -684 2396
rect -716 2315 -684 2316
rect -716 2285 -715 2315
rect -715 2285 -685 2315
rect -685 2285 -684 2315
rect -716 2284 -684 2285
rect -716 2204 -684 2236
rect -716 2155 -684 2156
rect -716 2125 -715 2155
rect -715 2125 -685 2155
rect -685 2125 -684 2155
rect -716 2124 -684 2125
rect -716 2075 -684 2076
rect -716 2045 -715 2075
rect -715 2045 -685 2075
rect -685 2045 -684 2075
rect -716 2044 -684 2045
rect -716 1995 -684 1996
rect -716 1965 -715 1995
rect -715 1965 -685 1995
rect -685 1965 -684 1995
rect -716 1964 -684 1965
rect -716 1915 -684 1916
rect -716 1885 -715 1915
rect -715 1885 -685 1915
rect -685 1885 -684 1915
rect -716 1884 -684 1885
rect -716 1835 -684 1836
rect -716 1805 -715 1835
rect -715 1805 -685 1835
rect -685 1805 -684 1835
rect -716 1804 -684 1805
rect -716 1755 -684 1756
rect -716 1725 -715 1755
rect -715 1725 -685 1755
rect -685 1725 -684 1755
rect -716 1724 -684 1725
rect -636 2475 -604 2476
rect -636 2445 -635 2475
rect -635 2445 -605 2475
rect -605 2445 -604 2475
rect -636 2444 -604 2445
rect -636 2364 -604 2396
rect -636 2315 -604 2316
rect -636 2285 -635 2315
rect -635 2285 -605 2315
rect -605 2285 -604 2315
rect -636 2284 -604 2285
rect -636 2204 -604 2236
rect -636 2155 -604 2156
rect -636 2125 -635 2155
rect -635 2125 -605 2155
rect -605 2125 -604 2155
rect -636 2124 -604 2125
rect -636 2075 -604 2076
rect -636 2045 -635 2075
rect -635 2045 -605 2075
rect -605 2045 -604 2075
rect -636 2044 -604 2045
rect -636 1995 -604 1996
rect -636 1965 -635 1995
rect -635 1965 -605 1995
rect -605 1965 -604 1995
rect -636 1964 -604 1965
rect -636 1915 -604 1916
rect -636 1885 -635 1915
rect -635 1885 -605 1915
rect -605 1885 -604 1915
rect -636 1884 -604 1885
rect -636 1835 -604 1836
rect -636 1805 -635 1835
rect -635 1805 -605 1835
rect -605 1805 -604 1835
rect -636 1804 -604 1805
rect -636 1755 -604 1756
rect -636 1725 -635 1755
rect -635 1725 -605 1755
rect -605 1725 -604 1755
rect -636 1724 -604 1725
rect -556 2475 -524 2476
rect -556 2445 -555 2475
rect -555 2445 -525 2475
rect -525 2445 -524 2475
rect -556 2444 -524 2445
rect -556 2364 -524 2396
rect -556 2315 -524 2316
rect -556 2285 -555 2315
rect -555 2285 -525 2315
rect -525 2285 -524 2315
rect -556 2284 -524 2285
rect -556 2204 -524 2236
rect -556 2155 -524 2156
rect -556 2125 -555 2155
rect -555 2125 -525 2155
rect -525 2125 -524 2155
rect -556 2124 -524 2125
rect -556 2075 -524 2076
rect -556 2045 -555 2075
rect -555 2045 -525 2075
rect -525 2045 -524 2075
rect -556 2044 -524 2045
rect -556 1995 -524 1996
rect -556 1965 -555 1995
rect -555 1965 -525 1995
rect -525 1965 -524 1995
rect -556 1964 -524 1965
rect -556 1915 -524 1916
rect -556 1885 -555 1915
rect -555 1885 -525 1915
rect -525 1885 -524 1915
rect -556 1884 -524 1885
rect -556 1835 -524 1836
rect -556 1805 -555 1835
rect -555 1805 -525 1835
rect -525 1805 -524 1835
rect -556 1804 -524 1805
rect -556 1755 -524 1756
rect -556 1725 -555 1755
rect -555 1725 -525 1755
rect -525 1725 -524 1755
rect -556 1724 -524 1725
rect -476 2475 -444 2476
rect -476 2445 -475 2475
rect -475 2445 -445 2475
rect -445 2445 -444 2475
rect -476 2444 -444 2445
rect -476 2364 -444 2396
rect -476 2315 -444 2316
rect -476 2285 -475 2315
rect -475 2285 -445 2315
rect -445 2285 -444 2315
rect -476 2284 -444 2285
rect -476 2204 -444 2236
rect -476 2155 -444 2156
rect -476 2125 -475 2155
rect -475 2125 -445 2155
rect -445 2125 -444 2155
rect -476 2124 -444 2125
rect -476 2075 -444 2076
rect -476 2045 -475 2075
rect -475 2045 -445 2075
rect -445 2045 -444 2075
rect -476 2044 -444 2045
rect -476 1995 -444 1996
rect -476 1965 -475 1995
rect -475 1965 -445 1995
rect -445 1965 -444 1995
rect -476 1964 -444 1965
rect -476 1915 -444 1916
rect -476 1885 -475 1915
rect -475 1885 -445 1915
rect -445 1885 -444 1915
rect -476 1884 -444 1885
rect -476 1835 -444 1836
rect -476 1805 -475 1835
rect -475 1805 -445 1835
rect -445 1805 -444 1835
rect -476 1804 -444 1805
rect -476 1755 -444 1756
rect -476 1725 -475 1755
rect -475 1725 -445 1755
rect -445 1725 -444 1755
rect -476 1724 -444 1725
rect -396 2475 -364 2476
rect -396 2445 -395 2475
rect -395 2445 -365 2475
rect -365 2445 -364 2475
rect -396 2444 -364 2445
rect -396 2364 -364 2396
rect -396 2315 -364 2316
rect -396 2285 -395 2315
rect -395 2285 -365 2315
rect -365 2285 -364 2315
rect -396 2284 -364 2285
rect -396 2204 -364 2236
rect -396 2155 -364 2156
rect -396 2125 -395 2155
rect -395 2125 -365 2155
rect -365 2125 -364 2155
rect -396 2124 -364 2125
rect -396 2075 -364 2076
rect -396 2045 -395 2075
rect -395 2045 -365 2075
rect -365 2045 -364 2075
rect -396 2044 -364 2045
rect -396 1995 -364 1996
rect -396 1965 -395 1995
rect -395 1965 -365 1995
rect -365 1965 -364 1995
rect -396 1964 -364 1965
rect -396 1915 -364 1916
rect -396 1885 -395 1915
rect -395 1885 -365 1915
rect -365 1885 -364 1915
rect -396 1884 -364 1885
rect -396 1835 -364 1836
rect -396 1805 -395 1835
rect -395 1805 -365 1835
rect -365 1805 -364 1835
rect -396 1804 -364 1805
rect -396 1755 -364 1756
rect -396 1725 -395 1755
rect -395 1725 -365 1755
rect -365 1725 -364 1755
rect -396 1724 -364 1725
rect -316 2475 -284 2476
rect -316 2445 -315 2475
rect -315 2445 -285 2475
rect -285 2445 -284 2475
rect -316 2444 -284 2445
rect -316 2364 -284 2396
rect -316 2315 -284 2316
rect -316 2285 -315 2315
rect -315 2285 -285 2315
rect -285 2285 -284 2315
rect -316 2284 -284 2285
rect -316 2204 -284 2236
rect -316 2155 -284 2156
rect -316 2125 -315 2155
rect -315 2125 -285 2155
rect -285 2125 -284 2155
rect -316 2124 -284 2125
rect -316 2075 -284 2076
rect -316 2045 -315 2075
rect -315 2045 -285 2075
rect -285 2045 -284 2075
rect -316 2044 -284 2045
rect -316 1995 -284 1996
rect -316 1965 -315 1995
rect -315 1965 -285 1995
rect -285 1965 -284 1995
rect -316 1964 -284 1965
rect -316 1915 -284 1916
rect -316 1885 -315 1915
rect -315 1885 -285 1915
rect -285 1885 -284 1915
rect -316 1884 -284 1885
rect -316 1835 -284 1836
rect -316 1805 -315 1835
rect -315 1805 -285 1835
rect -285 1805 -284 1835
rect -316 1804 -284 1805
rect -316 1755 -284 1756
rect -316 1725 -315 1755
rect -315 1725 -285 1755
rect -285 1725 -284 1755
rect -316 1724 -284 1725
rect -236 2475 -204 2476
rect -236 2445 -235 2475
rect -235 2445 -205 2475
rect -205 2445 -204 2475
rect -236 2444 -204 2445
rect -236 2364 -204 2396
rect -236 2315 -204 2316
rect -236 2285 -235 2315
rect -235 2285 -205 2315
rect -205 2285 -204 2315
rect -236 2284 -204 2285
rect -236 2204 -204 2236
rect -236 2155 -204 2156
rect -236 2125 -235 2155
rect -235 2125 -205 2155
rect -205 2125 -204 2155
rect -236 2124 -204 2125
rect -236 2075 -204 2076
rect -236 2045 -235 2075
rect -235 2045 -205 2075
rect -205 2045 -204 2075
rect -236 2044 -204 2045
rect -236 1995 -204 1996
rect -236 1965 -235 1995
rect -235 1965 -205 1995
rect -205 1965 -204 1995
rect -236 1964 -204 1965
rect -236 1915 -204 1916
rect -236 1885 -235 1915
rect -235 1885 -205 1915
rect -205 1885 -204 1915
rect -236 1884 -204 1885
rect -236 1835 -204 1836
rect -236 1805 -235 1835
rect -235 1805 -205 1835
rect -205 1805 -204 1835
rect -236 1804 -204 1805
rect -236 1755 -204 1756
rect -236 1725 -235 1755
rect -235 1725 -205 1755
rect -205 1725 -204 1755
rect -236 1724 -204 1725
rect -156 2475 -124 2476
rect -156 2445 -155 2475
rect -155 2445 -125 2475
rect -125 2445 -124 2475
rect -156 2444 -124 2445
rect -156 2364 -124 2396
rect -156 2315 -124 2316
rect -156 2285 -155 2315
rect -155 2285 -125 2315
rect -125 2285 -124 2315
rect -156 2284 -124 2285
rect -156 2204 -124 2236
rect -156 2155 -124 2156
rect -156 2125 -155 2155
rect -155 2125 -125 2155
rect -125 2125 -124 2155
rect -156 2124 -124 2125
rect -156 2075 -124 2076
rect -156 2045 -155 2075
rect -155 2045 -125 2075
rect -125 2045 -124 2075
rect -156 2044 -124 2045
rect -156 1995 -124 1996
rect -156 1965 -155 1995
rect -155 1965 -125 1995
rect -125 1965 -124 1995
rect -156 1964 -124 1965
rect -156 1915 -124 1916
rect -156 1885 -155 1915
rect -155 1885 -125 1915
rect -125 1885 -124 1915
rect -156 1884 -124 1885
rect -156 1835 -124 1836
rect -156 1805 -155 1835
rect -155 1805 -125 1835
rect -125 1805 -124 1835
rect -156 1804 -124 1805
rect -156 1755 -124 1756
rect -156 1725 -155 1755
rect -155 1725 -125 1755
rect -125 1725 -124 1755
rect -156 1724 -124 1725
rect -76 2475 -44 2476
rect -76 2445 -75 2475
rect -75 2445 -45 2475
rect -45 2445 -44 2475
rect -76 2444 -44 2445
rect -76 2364 -44 2396
rect -76 2315 -44 2316
rect -76 2285 -75 2315
rect -75 2285 -45 2315
rect -45 2285 -44 2315
rect -76 2284 -44 2285
rect -76 2204 -44 2236
rect -76 2155 -44 2156
rect -76 2125 -75 2155
rect -75 2125 -45 2155
rect -45 2125 -44 2155
rect -76 2124 -44 2125
rect -76 2075 -44 2076
rect -76 2045 -75 2075
rect -75 2045 -45 2075
rect -45 2045 -44 2075
rect -76 2044 -44 2045
rect -76 1995 -44 1996
rect -76 1965 -75 1995
rect -75 1965 -45 1995
rect -45 1965 -44 1995
rect -76 1964 -44 1965
rect -76 1915 -44 1916
rect -76 1885 -75 1915
rect -75 1885 -45 1915
rect -45 1885 -44 1915
rect -76 1884 -44 1885
rect -76 1835 -44 1836
rect -76 1805 -75 1835
rect -75 1805 -45 1835
rect -45 1805 -44 1835
rect -76 1804 -44 1805
rect -76 1755 -44 1756
rect -76 1725 -75 1755
rect -75 1725 -45 1755
rect -45 1725 -44 1755
rect -76 1724 -44 1725
rect 4 2475 36 2476
rect 4 2445 5 2475
rect 5 2445 35 2475
rect 35 2445 36 2475
rect 4 2444 36 2445
rect 4 2364 36 2396
rect 4 2315 36 2316
rect 4 2285 5 2315
rect 5 2285 35 2315
rect 35 2285 36 2315
rect 4 2284 36 2285
rect 4 2204 36 2236
rect 4 2155 36 2156
rect 4 2125 5 2155
rect 5 2125 35 2155
rect 35 2125 36 2155
rect 4 2124 36 2125
rect 4 2075 36 2076
rect 4 2045 5 2075
rect 5 2045 35 2075
rect 35 2045 36 2075
rect 4 2044 36 2045
rect 4 1995 36 1996
rect 4 1965 5 1995
rect 5 1965 35 1995
rect 35 1965 36 1995
rect 4 1964 36 1965
rect 4 1915 36 1916
rect 4 1885 5 1915
rect 5 1885 35 1915
rect 35 1885 36 1915
rect 4 1884 36 1885
rect 4 1835 36 1836
rect 4 1805 5 1835
rect 5 1805 35 1835
rect 35 1805 36 1835
rect 4 1804 36 1805
rect 4 1755 36 1756
rect 4 1725 5 1755
rect 5 1725 35 1755
rect 35 1725 36 1755
rect 4 1724 36 1725
rect 84 2475 116 2476
rect 84 2445 85 2475
rect 85 2445 115 2475
rect 115 2445 116 2475
rect 84 2444 116 2445
rect 84 2364 116 2396
rect 84 2315 116 2316
rect 84 2285 85 2315
rect 85 2285 115 2315
rect 115 2285 116 2315
rect 84 2284 116 2285
rect 84 2204 116 2236
rect 84 2155 116 2156
rect 84 2125 85 2155
rect 85 2125 115 2155
rect 115 2125 116 2155
rect 84 2124 116 2125
rect 84 2075 116 2076
rect 84 2045 85 2075
rect 85 2045 115 2075
rect 115 2045 116 2075
rect 84 2044 116 2045
rect 84 1995 116 1996
rect 84 1965 85 1995
rect 85 1965 115 1995
rect 115 1965 116 1995
rect 84 1964 116 1965
rect 84 1915 116 1916
rect 84 1885 85 1915
rect 85 1885 115 1915
rect 115 1885 116 1915
rect 84 1884 116 1885
rect 84 1835 116 1836
rect 84 1805 85 1835
rect 85 1805 115 1835
rect 115 1805 116 1835
rect 84 1804 116 1805
rect 84 1755 116 1756
rect 84 1725 85 1755
rect 85 1725 115 1755
rect 115 1725 116 1755
rect 84 1724 116 1725
rect 164 2475 196 2476
rect 164 2445 165 2475
rect 165 2445 195 2475
rect 195 2445 196 2475
rect 164 2444 196 2445
rect 164 2364 196 2396
rect 164 2315 196 2316
rect 164 2285 165 2315
rect 165 2285 195 2315
rect 195 2285 196 2315
rect 164 2284 196 2285
rect 164 2204 196 2236
rect 164 2155 196 2156
rect 164 2125 165 2155
rect 165 2125 195 2155
rect 195 2125 196 2155
rect 164 2124 196 2125
rect 164 2075 196 2076
rect 164 2045 165 2075
rect 165 2045 195 2075
rect 195 2045 196 2075
rect 164 2044 196 2045
rect 164 1995 196 1996
rect 164 1965 165 1995
rect 165 1965 195 1995
rect 195 1965 196 1995
rect 164 1964 196 1965
rect 164 1915 196 1916
rect 164 1885 165 1915
rect 165 1885 195 1915
rect 195 1885 196 1915
rect 164 1884 196 1885
rect 164 1835 196 1836
rect 164 1805 165 1835
rect 165 1805 195 1835
rect 195 1805 196 1835
rect 164 1804 196 1805
rect 164 1755 196 1756
rect 164 1725 165 1755
rect 165 1725 195 1755
rect 195 1725 196 1755
rect 164 1724 196 1725
rect 244 2475 276 2476
rect 244 2445 245 2475
rect 245 2445 275 2475
rect 275 2445 276 2475
rect 244 2444 276 2445
rect 244 2364 276 2396
rect 244 2315 276 2316
rect 244 2285 245 2315
rect 245 2285 275 2315
rect 275 2285 276 2315
rect 244 2284 276 2285
rect 244 2204 276 2236
rect 244 2155 276 2156
rect 244 2125 245 2155
rect 245 2125 275 2155
rect 275 2125 276 2155
rect 244 2124 276 2125
rect 244 2075 276 2076
rect 244 2045 245 2075
rect 245 2045 275 2075
rect 275 2045 276 2075
rect 244 2044 276 2045
rect 244 1995 276 1996
rect 244 1965 245 1995
rect 245 1965 275 1995
rect 275 1965 276 1995
rect 244 1964 276 1965
rect 244 1915 276 1916
rect 244 1885 245 1915
rect 245 1885 275 1915
rect 275 1885 276 1915
rect 244 1884 276 1885
rect 244 1835 276 1836
rect 244 1805 245 1835
rect 245 1805 275 1835
rect 275 1805 276 1835
rect 244 1804 276 1805
rect 244 1755 276 1756
rect 244 1725 245 1755
rect 245 1725 275 1755
rect 275 1725 276 1755
rect 244 1724 276 1725
rect 324 2475 356 2476
rect 324 2445 325 2475
rect 325 2445 355 2475
rect 355 2445 356 2475
rect 324 2444 356 2445
rect 324 2364 356 2396
rect 324 2315 356 2316
rect 324 2285 325 2315
rect 325 2285 355 2315
rect 355 2285 356 2315
rect 324 2284 356 2285
rect 324 2204 356 2236
rect 324 2155 356 2156
rect 324 2125 325 2155
rect 325 2125 355 2155
rect 355 2125 356 2155
rect 324 2124 356 2125
rect 324 2075 356 2076
rect 324 2045 325 2075
rect 325 2045 355 2075
rect 355 2045 356 2075
rect 324 2044 356 2045
rect 324 1995 356 1996
rect 324 1965 325 1995
rect 325 1965 355 1995
rect 355 1965 356 1995
rect 324 1964 356 1965
rect 324 1915 356 1916
rect 324 1885 325 1915
rect 325 1885 355 1915
rect 355 1885 356 1915
rect 324 1884 356 1885
rect 324 1835 356 1836
rect 324 1805 325 1835
rect 325 1805 355 1835
rect 355 1805 356 1835
rect 324 1804 356 1805
rect 324 1755 356 1756
rect 324 1725 325 1755
rect 325 1725 355 1755
rect 355 1725 356 1755
rect 324 1724 356 1725
rect 404 2475 436 2476
rect 404 2445 405 2475
rect 405 2445 435 2475
rect 435 2445 436 2475
rect 404 2444 436 2445
rect 404 2364 436 2396
rect 404 2315 436 2316
rect 404 2285 405 2315
rect 405 2285 435 2315
rect 435 2285 436 2315
rect 404 2284 436 2285
rect 404 2204 436 2236
rect 404 2155 436 2156
rect 404 2125 405 2155
rect 405 2125 435 2155
rect 435 2125 436 2155
rect 404 2124 436 2125
rect 404 2075 436 2076
rect 404 2045 405 2075
rect 405 2045 435 2075
rect 435 2045 436 2075
rect 404 2044 436 2045
rect 404 1995 436 1996
rect 404 1965 405 1995
rect 405 1965 435 1995
rect 435 1965 436 1995
rect 404 1964 436 1965
rect 404 1915 436 1916
rect 404 1885 405 1915
rect 405 1885 435 1915
rect 435 1885 436 1915
rect 404 1884 436 1885
rect 404 1835 436 1836
rect 404 1805 405 1835
rect 405 1805 435 1835
rect 435 1805 436 1835
rect 404 1804 436 1805
rect 404 1755 436 1756
rect 404 1725 405 1755
rect 405 1725 435 1755
rect 435 1725 436 1755
rect 404 1724 436 1725
rect 484 2475 516 2476
rect 484 2445 485 2475
rect 485 2445 515 2475
rect 515 2445 516 2475
rect 484 2444 516 2445
rect 484 2364 516 2396
rect 484 2315 516 2316
rect 484 2285 485 2315
rect 485 2285 515 2315
rect 515 2285 516 2315
rect 484 2284 516 2285
rect 484 2204 516 2236
rect 484 2155 516 2156
rect 484 2125 485 2155
rect 485 2125 515 2155
rect 515 2125 516 2155
rect 484 2124 516 2125
rect 484 2075 516 2076
rect 484 2045 485 2075
rect 485 2045 515 2075
rect 515 2045 516 2075
rect 484 2044 516 2045
rect 484 1995 516 1996
rect 484 1965 485 1995
rect 485 1965 515 1995
rect 515 1965 516 1995
rect 484 1964 516 1965
rect 484 1915 516 1916
rect 484 1885 485 1915
rect 485 1885 515 1915
rect 515 1885 516 1915
rect 484 1884 516 1885
rect 484 1835 516 1836
rect 484 1805 485 1835
rect 485 1805 515 1835
rect 515 1805 516 1835
rect 484 1804 516 1805
rect 484 1755 516 1756
rect 484 1725 485 1755
rect 485 1725 515 1755
rect 515 1725 516 1755
rect 484 1724 516 1725
rect 564 2475 596 2476
rect 564 2445 565 2475
rect 565 2445 595 2475
rect 595 2445 596 2475
rect 564 2444 596 2445
rect 564 2364 596 2396
rect 564 2315 596 2316
rect 564 2285 565 2315
rect 565 2285 595 2315
rect 595 2285 596 2315
rect 564 2284 596 2285
rect 564 2204 596 2236
rect 564 2155 596 2156
rect 564 2125 565 2155
rect 565 2125 595 2155
rect 595 2125 596 2155
rect 564 2124 596 2125
rect 564 2075 596 2076
rect 564 2045 565 2075
rect 565 2045 595 2075
rect 595 2045 596 2075
rect 564 2044 596 2045
rect 564 1995 596 1996
rect 564 1965 565 1995
rect 565 1965 595 1995
rect 595 1965 596 1995
rect 564 1964 596 1965
rect 564 1915 596 1916
rect 564 1885 565 1915
rect 565 1885 595 1915
rect 595 1885 596 1915
rect 564 1884 596 1885
rect 564 1835 596 1836
rect 564 1805 565 1835
rect 565 1805 595 1835
rect 595 1805 596 1835
rect 564 1804 596 1805
rect 564 1755 596 1756
rect 564 1725 565 1755
rect 565 1725 595 1755
rect 595 1725 596 1755
rect 564 1724 596 1725
rect 644 2475 676 2476
rect 644 2445 645 2475
rect 645 2445 675 2475
rect 675 2445 676 2475
rect 644 2444 676 2445
rect 644 2364 676 2396
rect 644 2315 676 2316
rect 644 2285 645 2315
rect 645 2285 675 2315
rect 675 2285 676 2315
rect 644 2284 676 2285
rect 644 2204 676 2236
rect 644 2155 676 2156
rect 644 2125 645 2155
rect 645 2125 675 2155
rect 675 2125 676 2155
rect 644 2124 676 2125
rect 644 2075 676 2076
rect 644 2045 645 2075
rect 645 2045 675 2075
rect 675 2045 676 2075
rect 644 2044 676 2045
rect 644 1995 676 1996
rect 644 1965 645 1995
rect 645 1965 675 1995
rect 675 1965 676 1995
rect 644 1964 676 1965
rect 644 1915 676 1916
rect 644 1885 645 1915
rect 645 1885 675 1915
rect 675 1885 676 1915
rect 644 1884 676 1885
rect 644 1835 676 1836
rect 644 1805 645 1835
rect 645 1805 675 1835
rect 675 1805 676 1835
rect 644 1804 676 1805
rect 644 1755 676 1756
rect 644 1725 645 1755
rect 645 1725 675 1755
rect 675 1725 676 1755
rect 644 1724 676 1725
rect 724 2475 756 2476
rect 724 2445 725 2475
rect 725 2445 755 2475
rect 755 2445 756 2475
rect 724 2444 756 2445
rect 724 2364 756 2396
rect 724 2315 756 2316
rect 724 2285 725 2315
rect 725 2285 755 2315
rect 755 2285 756 2315
rect 724 2284 756 2285
rect 724 2204 756 2236
rect 724 2155 756 2156
rect 724 2125 725 2155
rect 725 2125 755 2155
rect 755 2125 756 2155
rect 724 2124 756 2125
rect 724 2075 756 2076
rect 724 2045 725 2075
rect 725 2045 755 2075
rect 755 2045 756 2075
rect 724 2044 756 2045
rect 724 1995 756 1996
rect 724 1965 725 1995
rect 725 1965 755 1995
rect 755 1965 756 1995
rect 724 1964 756 1965
rect 724 1915 756 1916
rect 724 1885 725 1915
rect 725 1885 755 1915
rect 755 1885 756 1915
rect 724 1884 756 1885
rect 724 1835 756 1836
rect 724 1805 725 1835
rect 725 1805 755 1835
rect 755 1805 756 1835
rect 724 1804 756 1805
rect 724 1755 756 1756
rect 724 1725 725 1755
rect 725 1725 755 1755
rect 755 1725 756 1755
rect 724 1724 756 1725
rect 804 2475 836 2476
rect 804 2445 805 2475
rect 805 2445 835 2475
rect 835 2445 836 2475
rect 804 2444 836 2445
rect 804 2364 836 2396
rect 804 2315 836 2316
rect 804 2285 805 2315
rect 805 2285 835 2315
rect 835 2285 836 2315
rect 804 2284 836 2285
rect 804 2204 836 2236
rect 804 2155 836 2156
rect 804 2125 805 2155
rect 805 2125 835 2155
rect 835 2125 836 2155
rect 804 2124 836 2125
rect 804 2075 836 2076
rect 804 2045 805 2075
rect 805 2045 835 2075
rect 835 2045 836 2075
rect 804 2044 836 2045
rect 804 1995 836 1996
rect 804 1965 805 1995
rect 805 1965 835 1995
rect 835 1965 836 1995
rect 804 1964 836 1965
rect 804 1915 836 1916
rect 804 1885 805 1915
rect 805 1885 835 1915
rect 835 1885 836 1915
rect 804 1884 836 1885
rect 804 1835 836 1836
rect 804 1805 805 1835
rect 805 1805 835 1835
rect 835 1805 836 1835
rect 804 1804 836 1805
rect 804 1755 836 1756
rect 804 1725 805 1755
rect 805 1725 835 1755
rect 835 1725 836 1755
rect 804 1724 836 1725
rect 884 2475 916 2476
rect 884 2445 885 2475
rect 885 2445 915 2475
rect 915 2445 916 2475
rect 884 2444 916 2445
rect 884 2364 916 2396
rect 884 2315 916 2316
rect 884 2285 885 2315
rect 885 2285 915 2315
rect 915 2285 916 2315
rect 884 2284 916 2285
rect 884 2204 916 2236
rect 884 2155 916 2156
rect 884 2125 885 2155
rect 885 2125 915 2155
rect 915 2125 916 2155
rect 884 2124 916 2125
rect 884 2075 916 2076
rect 884 2045 885 2075
rect 885 2045 915 2075
rect 915 2045 916 2075
rect 884 2044 916 2045
rect 884 1995 916 1996
rect 884 1965 885 1995
rect 885 1965 915 1995
rect 915 1965 916 1995
rect 884 1964 916 1965
rect 884 1915 916 1916
rect 884 1885 885 1915
rect 885 1885 915 1915
rect 915 1885 916 1915
rect 884 1884 916 1885
rect 884 1835 916 1836
rect 884 1805 885 1835
rect 885 1805 915 1835
rect 915 1805 916 1835
rect 884 1804 916 1805
rect 884 1755 916 1756
rect 884 1725 885 1755
rect 885 1725 915 1755
rect 915 1725 916 1755
rect 884 1724 916 1725
rect 964 2475 996 2476
rect 964 2445 965 2475
rect 965 2445 995 2475
rect 995 2445 996 2475
rect 964 2444 996 2445
rect 964 2364 996 2396
rect 964 2315 996 2316
rect 964 2285 965 2315
rect 965 2285 995 2315
rect 995 2285 996 2315
rect 964 2284 996 2285
rect 964 2204 996 2236
rect 964 2155 996 2156
rect 964 2125 965 2155
rect 965 2125 995 2155
rect 995 2125 996 2155
rect 964 2124 996 2125
rect 964 2075 996 2076
rect 964 2045 965 2075
rect 965 2045 995 2075
rect 995 2045 996 2075
rect 964 2044 996 2045
rect 964 1995 996 1996
rect 964 1965 965 1995
rect 965 1965 995 1995
rect 995 1965 996 1995
rect 964 1964 996 1965
rect 964 1915 996 1916
rect 964 1885 965 1915
rect 965 1885 995 1915
rect 995 1885 996 1915
rect 964 1884 996 1885
rect 964 1835 996 1836
rect 964 1805 965 1835
rect 965 1805 995 1835
rect 995 1805 996 1835
rect 964 1804 996 1805
rect 964 1755 996 1756
rect 964 1725 965 1755
rect 965 1725 995 1755
rect 995 1725 996 1755
rect 964 1724 996 1725
rect 1044 2475 1076 2476
rect 1044 2445 1045 2475
rect 1045 2445 1075 2475
rect 1075 2445 1076 2475
rect 1044 2444 1076 2445
rect 1044 2364 1076 2396
rect 1044 2315 1076 2316
rect 1044 2285 1045 2315
rect 1045 2285 1075 2315
rect 1075 2285 1076 2315
rect 1044 2284 1076 2285
rect 1044 2204 1076 2236
rect 1044 2155 1076 2156
rect 1044 2125 1045 2155
rect 1045 2125 1075 2155
rect 1075 2125 1076 2155
rect 1044 2124 1076 2125
rect 1044 2075 1076 2076
rect 1044 2045 1045 2075
rect 1045 2045 1075 2075
rect 1075 2045 1076 2075
rect 1044 2044 1076 2045
rect 1044 1995 1076 1996
rect 1044 1965 1045 1995
rect 1045 1965 1075 1995
rect 1075 1965 1076 1995
rect 1044 1964 1076 1965
rect 1044 1915 1076 1916
rect 1044 1885 1045 1915
rect 1045 1885 1075 1915
rect 1075 1885 1076 1915
rect 1044 1884 1076 1885
rect 1044 1835 1076 1836
rect 1044 1805 1045 1835
rect 1045 1805 1075 1835
rect 1075 1805 1076 1835
rect 1044 1804 1076 1805
rect 1044 1755 1076 1756
rect 1044 1725 1045 1755
rect 1045 1725 1075 1755
rect 1075 1725 1076 1755
rect 1044 1724 1076 1725
rect 1124 2475 1156 2476
rect 1124 2445 1125 2475
rect 1125 2445 1155 2475
rect 1155 2445 1156 2475
rect 1124 2444 1156 2445
rect 1124 2364 1156 2396
rect 1124 2315 1156 2316
rect 1124 2285 1125 2315
rect 1125 2285 1155 2315
rect 1155 2285 1156 2315
rect 1124 2284 1156 2285
rect 1124 2204 1156 2236
rect 1124 2155 1156 2156
rect 1124 2125 1125 2155
rect 1125 2125 1155 2155
rect 1155 2125 1156 2155
rect 1124 2124 1156 2125
rect 1124 2075 1156 2076
rect 1124 2045 1125 2075
rect 1125 2045 1155 2075
rect 1155 2045 1156 2075
rect 1124 2044 1156 2045
rect 1124 1995 1156 1996
rect 1124 1965 1125 1995
rect 1125 1965 1155 1995
rect 1155 1965 1156 1995
rect 1124 1964 1156 1965
rect 1124 1915 1156 1916
rect 1124 1885 1125 1915
rect 1125 1885 1155 1915
rect 1155 1885 1156 1915
rect 1124 1884 1156 1885
rect 1124 1835 1156 1836
rect 1124 1805 1125 1835
rect 1125 1805 1155 1835
rect 1155 1805 1156 1835
rect 1124 1804 1156 1805
rect 1124 1755 1156 1756
rect 1124 1725 1125 1755
rect 1125 1725 1155 1755
rect 1155 1725 1156 1755
rect 1124 1724 1156 1725
rect 1204 2475 1236 2476
rect 1204 2445 1205 2475
rect 1205 2445 1235 2475
rect 1235 2445 1236 2475
rect 1204 2444 1236 2445
rect 1204 2364 1236 2396
rect 1204 2315 1236 2316
rect 1204 2285 1205 2315
rect 1205 2285 1235 2315
rect 1235 2285 1236 2315
rect 1204 2284 1236 2285
rect 1204 2204 1236 2236
rect 1204 2155 1236 2156
rect 1204 2125 1205 2155
rect 1205 2125 1235 2155
rect 1235 2125 1236 2155
rect 1204 2124 1236 2125
rect 1204 2075 1236 2076
rect 1204 2045 1205 2075
rect 1205 2045 1235 2075
rect 1235 2045 1236 2075
rect 1204 2044 1236 2045
rect 1204 1995 1236 1996
rect 1204 1965 1205 1995
rect 1205 1965 1235 1995
rect 1235 1965 1236 1995
rect 1204 1964 1236 1965
rect 1204 1915 1236 1916
rect 1204 1885 1205 1915
rect 1205 1885 1235 1915
rect 1235 1885 1236 1915
rect 1204 1884 1236 1885
rect 1204 1835 1236 1836
rect 1204 1805 1205 1835
rect 1205 1805 1235 1835
rect 1235 1805 1236 1835
rect 1204 1804 1236 1805
rect 1204 1755 1236 1756
rect 1204 1725 1205 1755
rect 1205 1725 1235 1755
rect 1235 1725 1236 1755
rect 1204 1724 1236 1725
rect 1284 2475 1316 2476
rect 1284 2445 1285 2475
rect 1285 2445 1315 2475
rect 1315 2445 1316 2475
rect 1284 2444 1316 2445
rect 1284 2364 1316 2396
rect 1284 2315 1316 2316
rect 1284 2285 1285 2315
rect 1285 2285 1315 2315
rect 1315 2285 1316 2315
rect 1284 2284 1316 2285
rect 1284 2204 1316 2236
rect 1284 2155 1316 2156
rect 1284 2125 1285 2155
rect 1285 2125 1315 2155
rect 1315 2125 1316 2155
rect 1284 2124 1316 2125
rect 1284 2075 1316 2076
rect 1284 2045 1285 2075
rect 1285 2045 1315 2075
rect 1315 2045 1316 2075
rect 1284 2044 1316 2045
rect 1284 1995 1316 1996
rect 1284 1965 1285 1995
rect 1285 1965 1315 1995
rect 1315 1965 1316 1995
rect 1284 1964 1316 1965
rect 1284 1915 1316 1916
rect 1284 1885 1285 1915
rect 1285 1885 1315 1915
rect 1315 1885 1316 1915
rect 1284 1884 1316 1885
rect 1284 1835 1316 1836
rect 1284 1805 1285 1835
rect 1285 1805 1315 1835
rect 1315 1805 1316 1835
rect 1284 1804 1316 1805
rect 1284 1755 1316 1756
rect 1284 1725 1285 1755
rect 1285 1725 1315 1755
rect 1315 1725 1316 1755
rect 1284 1724 1316 1725
rect 1364 2475 1396 2476
rect 1364 2445 1365 2475
rect 1365 2445 1395 2475
rect 1395 2445 1396 2475
rect 1364 2444 1396 2445
rect 1364 2364 1396 2396
rect 1364 2315 1396 2316
rect 1364 2285 1365 2315
rect 1365 2285 1395 2315
rect 1395 2285 1396 2315
rect 1364 2284 1396 2285
rect 1364 2204 1396 2236
rect 1364 2155 1396 2156
rect 1364 2125 1365 2155
rect 1365 2125 1395 2155
rect 1395 2125 1396 2155
rect 1364 2124 1396 2125
rect 1364 2075 1396 2076
rect 1364 2045 1365 2075
rect 1365 2045 1395 2075
rect 1395 2045 1396 2075
rect 1364 2044 1396 2045
rect 1364 1995 1396 1996
rect 1364 1965 1365 1995
rect 1365 1965 1395 1995
rect 1395 1965 1396 1995
rect 1364 1964 1396 1965
rect 1364 1915 1396 1916
rect 1364 1885 1365 1915
rect 1365 1885 1395 1915
rect 1395 1885 1396 1915
rect 1364 1884 1396 1885
rect 1364 1835 1396 1836
rect 1364 1805 1365 1835
rect 1365 1805 1395 1835
rect 1395 1805 1396 1835
rect 1364 1804 1396 1805
rect 1364 1755 1396 1756
rect 1364 1725 1365 1755
rect 1365 1725 1395 1755
rect 1395 1725 1396 1755
rect 1364 1724 1396 1725
rect 1444 2475 1476 2476
rect 1444 2445 1445 2475
rect 1445 2445 1475 2475
rect 1475 2445 1476 2475
rect 1444 2444 1476 2445
rect 1444 2364 1476 2396
rect 1444 2315 1476 2316
rect 1444 2285 1445 2315
rect 1445 2285 1475 2315
rect 1475 2285 1476 2315
rect 1444 2284 1476 2285
rect 1444 2204 1476 2236
rect 1444 2155 1476 2156
rect 1444 2125 1445 2155
rect 1445 2125 1475 2155
rect 1475 2125 1476 2155
rect 1444 2124 1476 2125
rect 1444 2075 1476 2076
rect 1444 2045 1445 2075
rect 1445 2045 1475 2075
rect 1475 2045 1476 2075
rect 1444 2044 1476 2045
rect 1444 1995 1476 1996
rect 1444 1965 1445 1995
rect 1445 1965 1475 1995
rect 1475 1965 1476 1995
rect 1444 1964 1476 1965
rect 1444 1915 1476 1916
rect 1444 1885 1445 1915
rect 1445 1885 1475 1915
rect 1475 1885 1476 1915
rect 1444 1884 1476 1885
rect 1444 1835 1476 1836
rect 1444 1805 1445 1835
rect 1445 1805 1475 1835
rect 1475 1805 1476 1835
rect 1444 1804 1476 1805
rect 1444 1755 1476 1756
rect 1444 1725 1445 1755
rect 1445 1725 1475 1755
rect 1475 1725 1476 1755
rect 1444 1724 1476 1725
rect 1524 2475 1556 2476
rect 1524 2445 1525 2475
rect 1525 2445 1555 2475
rect 1555 2445 1556 2475
rect 1524 2444 1556 2445
rect 1524 2364 1556 2396
rect 1524 2315 1556 2316
rect 1524 2285 1525 2315
rect 1525 2285 1555 2315
rect 1555 2285 1556 2315
rect 1524 2284 1556 2285
rect 1524 2204 1556 2236
rect 1524 2155 1556 2156
rect 1524 2125 1525 2155
rect 1525 2125 1555 2155
rect 1555 2125 1556 2155
rect 1524 2124 1556 2125
rect 1524 2075 1556 2076
rect 1524 2045 1525 2075
rect 1525 2045 1555 2075
rect 1555 2045 1556 2075
rect 1524 2044 1556 2045
rect 1524 1995 1556 1996
rect 1524 1965 1525 1995
rect 1525 1965 1555 1995
rect 1555 1965 1556 1995
rect 1524 1964 1556 1965
rect 1524 1915 1556 1916
rect 1524 1885 1525 1915
rect 1525 1885 1555 1915
rect 1555 1885 1556 1915
rect 1524 1884 1556 1885
rect 1524 1835 1556 1836
rect 1524 1805 1525 1835
rect 1525 1805 1555 1835
rect 1555 1805 1556 1835
rect 1524 1804 1556 1805
rect 1524 1755 1556 1756
rect 1524 1725 1525 1755
rect 1525 1725 1555 1755
rect 1555 1725 1556 1755
rect 1524 1724 1556 1725
rect 1604 2475 1636 2476
rect 1604 2445 1605 2475
rect 1605 2445 1635 2475
rect 1635 2445 1636 2475
rect 1604 2444 1636 2445
rect 1604 2364 1636 2396
rect 1604 2315 1636 2316
rect 1604 2285 1605 2315
rect 1605 2285 1635 2315
rect 1635 2285 1636 2315
rect 1604 2284 1636 2285
rect 1604 2204 1636 2236
rect 1604 2155 1636 2156
rect 1604 2125 1605 2155
rect 1605 2125 1635 2155
rect 1635 2125 1636 2155
rect 1604 2124 1636 2125
rect 1604 2075 1636 2076
rect 1604 2045 1605 2075
rect 1605 2045 1635 2075
rect 1635 2045 1636 2075
rect 1604 2044 1636 2045
rect 1604 1995 1636 1996
rect 1604 1965 1605 1995
rect 1605 1965 1635 1995
rect 1635 1965 1636 1995
rect 1604 1964 1636 1965
rect 1604 1915 1636 1916
rect 1604 1885 1605 1915
rect 1605 1885 1635 1915
rect 1635 1885 1636 1915
rect 1604 1884 1636 1885
rect 1604 1835 1636 1836
rect 1604 1805 1605 1835
rect 1605 1805 1635 1835
rect 1635 1805 1636 1835
rect 1604 1804 1636 1805
rect 1604 1755 1636 1756
rect 1604 1725 1605 1755
rect 1605 1725 1635 1755
rect 1635 1725 1636 1755
rect 1604 1724 1636 1725
rect 1684 2475 1716 2476
rect 1684 2445 1685 2475
rect 1685 2445 1715 2475
rect 1715 2445 1716 2475
rect 1684 2444 1716 2445
rect 1684 2364 1716 2396
rect 1684 2315 1716 2316
rect 1684 2285 1685 2315
rect 1685 2285 1715 2315
rect 1715 2285 1716 2315
rect 1684 2284 1716 2285
rect 1684 2204 1716 2236
rect 1684 2155 1716 2156
rect 1684 2125 1685 2155
rect 1685 2125 1715 2155
rect 1715 2125 1716 2155
rect 1684 2124 1716 2125
rect 1684 2075 1716 2076
rect 1684 2045 1685 2075
rect 1685 2045 1715 2075
rect 1715 2045 1716 2075
rect 1684 2044 1716 2045
rect 1684 1995 1716 1996
rect 1684 1965 1685 1995
rect 1685 1965 1715 1995
rect 1715 1965 1716 1995
rect 1684 1964 1716 1965
rect 1684 1915 1716 1916
rect 1684 1885 1685 1915
rect 1685 1885 1715 1915
rect 1715 1885 1716 1915
rect 1684 1884 1716 1885
rect 1684 1835 1716 1836
rect 1684 1805 1685 1835
rect 1685 1805 1715 1835
rect 1715 1805 1716 1835
rect 1684 1804 1716 1805
rect 1684 1755 1716 1756
rect 1684 1725 1685 1755
rect 1685 1725 1715 1755
rect 1715 1725 1716 1755
rect 1684 1724 1716 1725
rect 1764 2475 1796 2476
rect 1764 2445 1765 2475
rect 1765 2445 1795 2475
rect 1795 2445 1796 2475
rect 1764 2444 1796 2445
rect 1764 2364 1796 2396
rect 1764 2315 1796 2316
rect 1764 2285 1765 2315
rect 1765 2285 1795 2315
rect 1795 2285 1796 2315
rect 1764 2284 1796 2285
rect 1764 2204 1796 2236
rect 1764 2155 1796 2156
rect 1764 2125 1765 2155
rect 1765 2125 1795 2155
rect 1795 2125 1796 2155
rect 1764 2124 1796 2125
rect 1764 2075 1796 2076
rect 1764 2045 1765 2075
rect 1765 2045 1795 2075
rect 1795 2045 1796 2075
rect 1764 2044 1796 2045
rect 1764 1995 1796 1996
rect 1764 1965 1765 1995
rect 1765 1965 1795 1995
rect 1795 1965 1796 1995
rect 1764 1964 1796 1965
rect 1764 1915 1796 1916
rect 1764 1885 1765 1915
rect 1765 1885 1795 1915
rect 1795 1885 1796 1915
rect 1764 1884 1796 1885
rect 1764 1835 1796 1836
rect 1764 1805 1765 1835
rect 1765 1805 1795 1835
rect 1795 1805 1796 1835
rect 1764 1804 1796 1805
rect 1764 1755 1796 1756
rect 1764 1725 1765 1755
rect 1765 1725 1795 1755
rect 1795 1725 1796 1755
rect 1764 1724 1796 1725
rect 1844 2475 1876 2476
rect 1844 2445 1845 2475
rect 1845 2445 1875 2475
rect 1875 2445 1876 2475
rect 1844 2444 1876 2445
rect 1844 2364 1876 2396
rect 1844 2315 1876 2316
rect 1844 2285 1845 2315
rect 1845 2285 1875 2315
rect 1875 2285 1876 2315
rect 1844 2284 1876 2285
rect 1844 2204 1876 2236
rect 1844 2155 1876 2156
rect 1844 2125 1845 2155
rect 1845 2125 1875 2155
rect 1875 2125 1876 2155
rect 1844 2124 1876 2125
rect 1844 2075 1876 2076
rect 1844 2045 1845 2075
rect 1845 2045 1875 2075
rect 1875 2045 1876 2075
rect 1844 2044 1876 2045
rect 1844 1995 1876 1996
rect 1844 1965 1845 1995
rect 1845 1965 1875 1995
rect 1875 1965 1876 1995
rect 1844 1964 1876 1965
rect 1844 1915 1876 1916
rect 1844 1885 1845 1915
rect 1845 1885 1875 1915
rect 1875 1885 1876 1915
rect 1844 1884 1876 1885
rect 1844 1835 1876 1836
rect 1844 1805 1845 1835
rect 1845 1805 1875 1835
rect 1875 1805 1876 1835
rect 1844 1804 1876 1805
rect 1844 1755 1876 1756
rect 1844 1725 1845 1755
rect 1845 1725 1875 1755
rect 1875 1725 1876 1755
rect 1844 1724 1876 1725
rect 1924 2475 1956 2476
rect 1924 2445 1925 2475
rect 1925 2445 1955 2475
rect 1955 2445 1956 2475
rect 1924 2444 1956 2445
rect 1924 2364 1956 2396
rect 1924 2315 1956 2316
rect 1924 2285 1925 2315
rect 1925 2285 1955 2315
rect 1955 2285 1956 2315
rect 1924 2284 1956 2285
rect 1924 2204 1956 2236
rect 1924 2155 1956 2156
rect 1924 2125 1925 2155
rect 1925 2125 1955 2155
rect 1955 2125 1956 2155
rect 1924 2124 1956 2125
rect 1924 2075 1956 2076
rect 1924 2045 1925 2075
rect 1925 2045 1955 2075
rect 1955 2045 1956 2075
rect 1924 2044 1956 2045
rect 1924 1995 1956 1996
rect 1924 1965 1925 1995
rect 1925 1965 1955 1995
rect 1955 1965 1956 1995
rect 1924 1964 1956 1965
rect 1924 1915 1956 1916
rect 1924 1885 1925 1915
rect 1925 1885 1955 1915
rect 1955 1885 1956 1915
rect 1924 1884 1956 1885
rect 1924 1835 1956 1836
rect 1924 1805 1925 1835
rect 1925 1805 1955 1835
rect 1955 1805 1956 1835
rect 1924 1804 1956 1805
rect 1924 1755 1956 1756
rect 1924 1725 1925 1755
rect 1925 1725 1955 1755
rect 1955 1725 1956 1755
rect 1924 1724 1956 1725
rect 2004 2475 2036 2476
rect 2004 2445 2005 2475
rect 2005 2445 2035 2475
rect 2035 2445 2036 2475
rect 2004 2444 2036 2445
rect 2004 2364 2036 2396
rect 2004 2315 2036 2316
rect 2004 2285 2005 2315
rect 2005 2285 2035 2315
rect 2035 2285 2036 2315
rect 2004 2284 2036 2285
rect 2004 2204 2036 2236
rect 2004 2155 2036 2156
rect 2004 2125 2005 2155
rect 2005 2125 2035 2155
rect 2035 2125 2036 2155
rect 2004 2124 2036 2125
rect 2004 2075 2036 2076
rect 2004 2045 2005 2075
rect 2005 2045 2035 2075
rect 2035 2045 2036 2075
rect 2004 2044 2036 2045
rect 2004 1995 2036 1996
rect 2004 1965 2005 1995
rect 2005 1965 2035 1995
rect 2035 1965 2036 1995
rect 2004 1964 2036 1965
rect 2004 1915 2036 1916
rect 2004 1885 2005 1915
rect 2005 1885 2035 1915
rect 2035 1885 2036 1915
rect 2004 1884 2036 1885
rect 2004 1835 2036 1836
rect 2004 1805 2005 1835
rect 2005 1805 2035 1835
rect 2035 1805 2036 1835
rect 2004 1804 2036 1805
rect 2004 1755 2036 1756
rect 2004 1725 2005 1755
rect 2005 1725 2035 1755
rect 2035 1725 2036 1755
rect 2004 1724 2036 1725
rect 2084 2475 2116 2476
rect 2084 2445 2085 2475
rect 2085 2445 2115 2475
rect 2115 2445 2116 2475
rect 2084 2444 2116 2445
rect 2084 2364 2116 2396
rect 2084 2315 2116 2316
rect 2084 2285 2085 2315
rect 2085 2285 2115 2315
rect 2115 2285 2116 2315
rect 2084 2284 2116 2285
rect 2084 2204 2116 2236
rect 2084 2155 2116 2156
rect 2084 2125 2085 2155
rect 2085 2125 2115 2155
rect 2115 2125 2116 2155
rect 2084 2124 2116 2125
rect 2084 2075 2116 2076
rect 2084 2045 2085 2075
rect 2085 2045 2115 2075
rect 2115 2045 2116 2075
rect 2084 2044 2116 2045
rect 2084 1995 2116 1996
rect 2084 1965 2085 1995
rect 2085 1965 2115 1995
rect 2115 1965 2116 1995
rect 2084 1964 2116 1965
rect 2084 1915 2116 1916
rect 2084 1885 2085 1915
rect 2085 1885 2115 1915
rect 2115 1885 2116 1915
rect 2084 1884 2116 1885
rect 2084 1835 2116 1836
rect 2084 1805 2085 1835
rect 2085 1805 2115 1835
rect 2115 1805 2116 1835
rect 2084 1804 2116 1805
rect 2084 1755 2116 1756
rect 2084 1725 2085 1755
rect 2085 1725 2115 1755
rect 2115 1725 2116 1755
rect 2084 1724 2116 1725
rect 2164 2475 2196 2476
rect 2164 2445 2165 2475
rect 2165 2445 2195 2475
rect 2195 2445 2196 2475
rect 2164 2444 2196 2445
rect 2164 2364 2196 2396
rect 2164 2315 2196 2316
rect 2164 2285 2165 2315
rect 2165 2285 2195 2315
rect 2195 2285 2196 2315
rect 2164 2284 2196 2285
rect 2164 2204 2196 2236
rect 2164 2155 2196 2156
rect 2164 2125 2165 2155
rect 2165 2125 2195 2155
rect 2195 2125 2196 2155
rect 2164 2124 2196 2125
rect 2164 2075 2196 2076
rect 2164 2045 2165 2075
rect 2165 2045 2195 2075
rect 2195 2045 2196 2075
rect 2164 2044 2196 2045
rect 2164 1995 2196 1996
rect 2164 1965 2165 1995
rect 2165 1965 2195 1995
rect 2195 1965 2196 1995
rect 2164 1964 2196 1965
rect 2164 1915 2196 1916
rect 2164 1885 2165 1915
rect 2165 1885 2195 1915
rect 2195 1885 2196 1915
rect 2164 1884 2196 1885
rect 2164 1835 2196 1836
rect 2164 1805 2165 1835
rect 2165 1805 2195 1835
rect 2195 1805 2196 1835
rect 2164 1804 2196 1805
rect 2164 1755 2196 1756
rect 2164 1725 2165 1755
rect 2165 1725 2195 1755
rect 2195 1725 2196 1755
rect 2164 1724 2196 1725
rect 2244 2475 2276 2476
rect 2244 2445 2245 2475
rect 2245 2445 2275 2475
rect 2275 2445 2276 2475
rect 2244 2444 2276 2445
rect 2244 2364 2276 2396
rect 2244 2315 2276 2316
rect 2244 2285 2245 2315
rect 2245 2285 2275 2315
rect 2275 2285 2276 2315
rect 2244 2284 2276 2285
rect 2244 2204 2276 2236
rect 2244 2155 2276 2156
rect 2244 2125 2245 2155
rect 2245 2125 2275 2155
rect 2275 2125 2276 2155
rect 2244 2124 2276 2125
rect 2244 2075 2276 2076
rect 2244 2045 2245 2075
rect 2245 2045 2275 2075
rect 2275 2045 2276 2075
rect 2244 2044 2276 2045
rect 2244 1995 2276 1996
rect 2244 1965 2245 1995
rect 2245 1965 2275 1995
rect 2275 1965 2276 1995
rect 2244 1964 2276 1965
rect 2244 1915 2276 1916
rect 2244 1885 2245 1915
rect 2245 1885 2275 1915
rect 2275 1885 2276 1915
rect 2244 1884 2276 1885
rect 2244 1835 2276 1836
rect 2244 1805 2245 1835
rect 2245 1805 2275 1835
rect 2275 1805 2276 1835
rect 2244 1804 2276 1805
rect 2244 1755 2276 1756
rect 2244 1725 2245 1755
rect 2245 1725 2275 1755
rect 2275 1725 2276 1755
rect 2244 1724 2276 1725
rect 2324 2475 2356 2476
rect 2324 2445 2325 2475
rect 2325 2445 2355 2475
rect 2355 2445 2356 2475
rect 2324 2444 2356 2445
rect 2324 2364 2356 2396
rect 2324 2315 2356 2316
rect 2324 2285 2325 2315
rect 2325 2285 2355 2315
rect 2355 2285 2356 2315
rect 2324 2284 2356 2285
rect 2324 2204 2356 2236
rect 2324 2155 2356 2156
rect 2324 2125 2325 2155
rect 2325 2125 2355 2155
rect 2355 2125 2356 2155
rect 2324 2124 2356 2125
rect 2324 2075 2356 2076
rect 2324 2045 2325 2075
rect 2325 2045 2355 2075
rect 2355 2045 2356 2075
rect 2324 2044 2356 2045
rect 2324 1995 2356 1996
rect 2324 1965 2325 1995
rect 2325 1965 2355 1995
rect 2355 1965 2356 1995
rect 2324 1964 2356 1965
rect 2324 1915 2356 1916
rect 2324 1885 2325 1915
rect 2325 1885 2355 1915
rect 2355 1885 2356 1915
rect 2324 1884 2356 1885
rect 2324 1835 2356 1836
rect 2324 1805 2325 1835
rect 2325 1805 2355 1835
rect 2355 1805 2356 1835
rect 2324 1804 2356 1805
rect 2324 1755 2356 1756
rect 2324 1725 2325 1755
rect 2325 1725 2355 1755
rect 2355 1725 2356 1755
rect 2324 1724 2356 1725
rect 2404 2475 2436 2476
rect 2404 2445 2405 2475
rect 2405 2445 2435 2475
rect 2435 2445 2436 2475
rect 2404 2444 2436 2445
rect 2404 2364 2436 2396
rect 2404 2315 2436 2316
rect 2404 2285 2405 2315
rect 2405 2285 2435 2315
rect 2435 2285 2436 2315
rect 2404 2284 2436 2285
rect 2404 2204 2436 2236
rect 2404 2155 2436 2156
rect 2404 2125 2405 2155
rect 2405 2125 2435 2155
rect 2435 2125 2436 2155
rect 2404 2124 2436 2125
rect 2404 2075 2436 2076
rect 2404 2045 2405 2075
rect 2405 2045 2435 2075
rect 2435 2045 2436 2075
rect 2404 2044 2436 2045
rect 2404 1995 2436 1996
rect 2404 1965 2405 1995
rect 2405 1965 2435 1995
rect 2435 1965 2436 1995
rect 2404 1964 2436 1965
rect 2404 1915 2436 1916
rect 2404 1885 2405 1915
rect 2405 1885 2435 1915
rect 2435 1885 2436 1915
rect 2404 1884 2436 1885
rect 2404 1835 2436 1836
rect 2404 1805 2405 1835
rect 2405 1805 2435 1835
rect 2435 1805 2436 1835
rect 2404 1804 2436 1805
rect 2404 1755 2436 1756
rect 2404 1725 2405 1755
rect 2405 1725 2435 1755
rect 2435 1725 2436 1755
rect 2404 1724 2436 1725
rect 2484 2475 2516 2476
rect 2484 2445 2485 2475
rect 2485 2445 2515 2475
rect 2515 2445 2516 2475
rect 2484 2444 2516 2445
rect 2484 2364 2516 2396
rect 2484 2315 2516 2316
rect 2484 2285 2485 2315
rect 2485 2285 2515 2315
rect 2515 2285 2516 2315
rect 2484 2284 2516 2285
rect 2484 2204 2516 2236
rect 2484 2155 2516 2156
rect 2484 2125 2485 2155
rect 2485 2125 2515 2155
rect 2515 2125 2516 2155
rect 2484 2124 2516 2125
rect 2484 2075 2516 2076
rect 2484 2045 2485 2075
rect 2485 2045 2515 2075
rect 2515 2045 2516 2075
rect 2484 2044 2516 2045
rect 2484 1995 2516 1996
rect 2484 1965 2485 1995
rect 2485 1965 2515 1995
rect 2515 1965 2516 1995
rect 2484 1964 2516 1965
rect 2484 1915 2516 1916
rect 2484 1885 2485 1915
rect 2485 1885 2515 1915
rect 2515 1885 2516 1915
rect 2484 1884 2516 1885
rect 2484 1835 2516 1836
rect 2484 1805 2485 1835
rect 2485 1805 2515 1835
rect 2515 1805 2516 1835
rect 2484 1804 2516 1805
rect 2484 1755 2516 1756
rect 2484 1725 2485 1755
rect 2485 1725 2515 1755
rect 2515 1725 2516 1755
rect 2484 1724 2516 1725
rect 2564 2475 2596 2476
rect 2564 2445 2565 2475
rect 2565 2445 2595 2475
rect 2595 2445 2596 2475
rect 2564 2444 2596 2445
rect 2564 2364 2596 2396
rect 2564 2315 2596 2316
rect 2564 2285 2565 2315
rect 2565 2285 2595 2315
rect 2595 2285 2596 2315
rect 2564 2284 2596 2285
rect 2564 2204 2596 2236
rect 2564 2155 2596 2156
rect 2564 2125 2565 2155
rect 2565 2125 2595 2155
rect 2595 2125 2596 2155
rect 2564 2124 2596 2125
rect 2564 2075 2596 2076
rect 2564 2045 2565 2075
rect 2565 2045 2595 2075
rect 2595 2045 2596 2075
rect 2564 2044 2596 2045
rect 2564 1995 2596 1996
rect 2564 1965 2565 1995
rect 2565 1965 2595 1995
rect 2595 1965 2596 1995
rect 2564 1964 2596 1965
rect 2564 1915 2596 1916
rect 2564 1885 2565 1915
rect 2565 1885 2595 1915
rect 2595 1885 2596 1915
rect 2564 1884 2596 1885
rect 2564 1835 2596 1836
rect 2564 1805 2565 1835
rect 2565 1805 2595 1835
rect 2595 1805 2596 1835
rect 2564 1804 2596 1805
rect 2564 1755 2596 1756
rect 2564 1725 2565 1755
rect 2565 1725 2595 1755
rect 2595 1725 2596 1755
rect 2564 1724 2596 1725
rect 2644 2475 2676 2476
rect 2644 2445 2645 2475
rect 2645 2445 2675 2475
rect 2675 2445 2676 2475
rect 2644 2444 2676 2445
rect 2644 2364 2676 2396
rect 2644 2315 2676 2316
rect 2644 2285 2645 2315
rect 2645 2285 2675 2315
rect 2675 2285 2676 2315
rect 2644 2284 2676 2285
rect 2644 2204 2676 2236
rect 2644 2155 2676 2156
rect 2644 2125 2645 2155
rect 2645 2125 2675 2155
rect 2675 2125 2676 2155
rect 2644 2124 2676 2125
rect 2644 2075 2676 2076
rect 2644 2045 2645 2075
rect 2645 2045 2675 2075
rect 2675 2045 2676 2075
rect 2644 2044 2676 2045
rect 2644 1995 2676 1996
rect 2644 1965 2645 1995
rect 2645 1965 2675 1995
rect 2675 1965 2676 1995
rect 2644 1964 2676 1965
rect 2644 1915 2676 1916
rect 2644 1885 2645 1915
rect 2645 1885 2675 1915
rect 2675 1885 2676 1915
rect 2644 1884 2676 1885
rect 2644 1835 2676 1836
rect 2644 1805 2645 1835
rect 2645 1805 2675 1835
rect 2675 1805 2676 1835
rect 2644 1804 2676 1805
rect 2644 1755 2676 1756
rect 2644 1725 2645 1755
rect 2645 1725 2675 1755
rect 2675 1725 2676 1755
rect 2644 1724 2676 1725
rect 2724 2475 2756 2476
rect 2724 2445 2725 2475
rect 2725 2445 2755 2475
rect 2755 2445 2756 2475
rect 2724 2444 2756 2445
rect 2724 2364 2756 2396
rect 2724 2315 2756 2316
rect 2724 2285 2725 2315
rect 2725 2285 2755 2315
rect 2755 2285 2756 2315
rect 2724 2284 2756 2285
rect 2724 2204 2756 2236
rect 2724 2155 2756 2156
rect 2724 2125 2725 2155
rect 2725 2125 2755 2155
rect 2755 2125 2756 2155
rect 2724 2124 2756 2125
rect 2724 2075 2756 2076
rect 2724 2045 2725 2075
rect 2725 2045 2755 2075
rect 2755 2045 2756 2075
rect 2724 2044 2756 2045
rect 2724 1995 2756 1996
rect 2724 1965 2725 1995
rect 2725 1965 2755 1995
rect 2755 1965 2756 1995
rect 2724 1964 2756 1965
rect 2724 1915 2756 1916
rect 2724 1885 2725 1915
rect 2725 1885 2755 1915
rect 2755 1885 2756 1915
rect 2724 1884 2756 1885
rect 2724 1835 2756 1836
rect 2724 1805 2725 1835
rect 2725 1805 2755 1835
rect 2755 1805 2756 1835
rect 2724 1804 2756 1805
rect 2724 1755 2756 1756
rect 2724 1725 2725 1755
rect 2725 1725 2755 1755
rect 2755 1725 2756 1755
rect 2724 1724 2756 1725
rect 2804 2475 2836 2476
rect 2804 2445 2805 2475
rect 2805 2445 2835 2475
rect 2835 2445 2836 2475
rect 2804 2444 2836 2445
rect 2804 2364 2836 2396
rect 2804 2315 2836 2316
rect 2804 2285 2805 2315
rect 2805 2285 2835 2315
rect 2835 2285 2836 2315
rect 2804 2284 2836 2285
rect 2804 2204 2836 2236
rect 2804 2155 2836 2156
rect 2804 2125 2805 2155
rect 2805 2125 2835 2155
rect 2835 2125 2836 2155
rect 2804 2124 2836 2125
rect 2804 2075 2836 2076
rect 2804 2045 2805 2075
rect 2805 2045 2835 2075
rect 2835 2045 2836 2075
rect 2804 2044 2836 2045
rect 2804 1995 2836 1996
rect 2804 1965 2805 1995
rect 2805 1965 2835 1995
rect 2835 1965 2836 1995
rect 2804 1964 2836 1965
rect 2804 1915 2836 1916
rect 2804 1885 2805 1915
rect 2805 1885 2835 1915
rect 2835 1885 2836 1915
rect 2804 1884 2836 1885
rect 2804 1835 2836 1836
rect 2804 1805 2805 1835
rect 2805 1805 2835 1835
rect 2835 1805 2836 1835
rect 2804 1804 2836 1805
rect 2804 1755 2836 1756
rect 2804 1725 2805 1755
rect 2805 1725 2835 1755
rect 2835 1725 2836 1755
rect 2804 1724 2836 1725
rect 2884 2475 2916 2476
rect 2884 2445 2885 2475
rect 2885 2445 2915 2475
rect 2915 2445 2916 2475
rect 2884 2444 2916 2445
rect 2884 2364 2916 2396
rect 2884 2315 2916 2316
rect 2884 2285 2885 2315
rect 2885 2285 2915 2315
rect 2915 2285 2916 2315
rect 2884 2284 2916 2285
rect 2884 2204 2916 2236
rect 2884 2155 2916 2156
rect 2884 2125 2885 2155
rect 2885 2125 2915 2155
rect 2915 2125 2916 2155
rect 2884 2124 2916 2125
rect 2884 2075 2916 2076
rect 2884 2045 2885 2075
rect 2885 2045 2915 2075
rect 2915 2045 2916 2075
rect 2884 2044 2916 2045
rect 2884 1995 2916 1996
rect 2884 1965 2885 1995
rect 2885 1965 2915 1995
rect 2915 1965 2916 1995
rect 2884 1964 2916 1965
rect 2884 1915 2916 1916
rect 2884 1885 2885 1915
rect 2885 1885 2915 1915
rect 2915 1885 2916 1915
rect 2884 1884 2916 1885
rect 2884 1835 2916 1836
rect 2884 1805 2885 1835
rect 2885 1805 2915 1835
rect 2915 1805 2916 1835
rect 2884 1804 2916 1805
rect 2884 1755 2916 1756
rect 2884 1725 2885 1755
rect 2885 1725 2915 1755
rect 2915 1725 2916 1755
rect 2884 1724 2916 1725
rect 2964 2475 2996 2476
rect 2964 2445 2965 2475
rect 2965 2445 2995 2475
rect 2995 2445 2996 2475
rect 2964 2444 2996 2445
rect 2964 2364 2996 2396
rect 2964 2315 2996 2316
rect 2964 2285 2965 2315
rect 2965 2285 2995 2315
rect 2995 2285 2996 2315
rect 2964 2284 2996 2285
rect 2964 2204 2996 2236
rect 2964 2155 2996 2156
rect 2964 2125 2965 2155
rect 2965 2125 2995 2155
rect 2995 2125 2996 2155
rect 2964 2124 2996 2125
rect 2964 2075 2996 2076
rect 2964 2045 2965 2075
rect 2965 2045 2995 2075
rect 2995 2045 2996 2075
rect 2964 2044 2996 2045
rect 2964 1995 2996 1996
rect 2964 1965 2965 1995
rect 2965 1965 2995 1995
rect 2995 1965 2996 1995
rect 2964 1964 2996 1965
rect 2964 1915 2996 1916
rect 2964 1885 2965 1915
rect 2965 1885 2995 1915
rect 2995 1885 2996 1915
rect 2964 1884 2996 1885
rect 2964 1835 2996 1836
rect 2964 1805 2965 1835
rect 2965 1805 2995 1835
rect 2995 1805 2996 1835
rect 2964 1804 2996 1805
rect 2964 1755 2996 1756
rect 2964 1725 2965 1755
rect 2965 1725 2995 1755
rect 2995 1725 2996 1755
rect 2964 1724 2996 1725
rect 3044 2475 3076 2476
rect 3044 2445 3045 2475
rect 3045 2445 3075 2475
rect 3075 2445 3076 2475
rect 3044 2444 3076 2445
rect 3044 2364 3076 2396
rect 3044 2315 3076 2316
rect 3044 2285 3045 2315
rect 3045 2285 3075 2315
rect 3075 2285 3076 2315
rect 3044 2284 3076 2285
rect 3044 2204 3076 2236
rect 3044 2155 3076 2156
rect 3044 2125 3045 2155
rect 3045 2125 3075 2155
rect 3075 2125 3076 2155
rect 3044 2124 3076 2125
rect 3044 2075 3076 2076
rect 3044 2045 3045 2075
rect 3045 2045 3075 2075
rect 3075 2045 3076 2075
rect 3044 2044 3076 2045
rect 3044 1995 3076 1996
rect 3044 1965 3045 1995
rect 3045 1965 3075 1995
rect 3075 1965 3076 1995
rect 3044 1964 3076 1965
rect 3044 1915 3076 1916
rect 3044 1885 3045 1915
rect 3045 1885 3075 1915
rect 3075 1885 3076 1915
rect 3044 1884 3076 1885
rect 3044 1835 3076 1836
rect 3044 1805 3045 1835
rect 3045 1805 3075 1835
rect 3075 1805 3076 1835
rect 3044 1804 3076 1805
rect 3044 1755 3076 1756
rect 3044 1725 3045 1755
rect 3045 1725 3075 1755
rect 3075 1725 3076 1755
rect 3044 1724 3076 1725
rect 3124 2475 3156 2476
rect 3124 2445 3125 2475
rect 3125 2445 3155 2475
rect 3155 2445 3156 2475
rect 3124 2444 3156 2445
rect 3124 2364 3156 2396
rect 3124 2315 3156 2316
rect 3124 2285 3125 2315
rect 3125 2285 3155 2315
rect 3155 2285 3156 2315
rect 3124 2284 3156 2285
rect 3124 2204 3156 2236
rect 3124 2155 3156 2156
rect 3124 2125 3125 2155
rect 3125 2125 3155 2155
rect 3155 2125 3156 2155
rect 3124 2124 3156 2125
rect 3124 2075 3156 2076
rect 3124 2045 3125 2075
rect 3125 2045 3155 2075
rect 3155 2045 3156 2075
rect 3124 2044 3156 2045
rect 3124 1995 3156 1996
rect 3124 1965 3125 1995
rect 3125 1965 3155 1995
rect 3155 1965 3156 1995
rect 3124 1964 3156 1965
rect 3124 1915 3156 1916
rect 3124 1885 3125 1915
rect 3125 1885 3155 1915
rect 3155 1885 3156 1915
rect 3124 1884 3156 1885
rect 3124 1835 3156 1836
rect 3124 1805 3125 1835
rect 3125 1805 3155 1835
rect 3155 1805 3156 1835
rect 3124 1804 3156 1805
rect 3124 1755 3156 1756
rect 3124 1725 3125 1755
rect 3125 1725 3155 1755
rect 3155 1725 3156 1755
rect 3124 1724 3156 1725
rect 3204 2475 3236 2476
rect 3204 2445 3205 2475
rect 3205 2445 3235 2475
rect 3235 2445 3236 2475
rect 3204 2444 3236 2445
rect 3204 2364 3236 2396
rect 3204 2315 3236 2316
rect 3204 2285 3205 2315
rect 3205 2285 3235 2315
rect 3235 2285 3236 2315
rect 3204 2284 3236 2285
rect 3204 2204 3236 2236
rect 3204 2155 3236 2156
rect 3204 2125 3205 2155
rect 3205 2125 3235 2155
rect 3235 2125 3236 2155
rect 3204 2124 3236 2125
rect 3204 2075 3236 2076
rect 3204 2045 3205 2075
rect 3205 2045 3235 2075
rect 3235 2045 3236 2075
rect 3204 2044 3236 2045
rect 3204 1995 3236 1996
rect 3204 1965 3205 1995
rect 3205 1965 3235 1995
rect 3235 1965 3236 1995
rect 3204 1964 3236 1965
rect 3204 1915 3236 1916
rect 3204 1885 3205 1915
rect 3205 1885 3235 1915
rect 3235 1885 3236 1915
rect 3204 1884 3236 1885
rect 3204 1835 3236 1836
rect 3204 1805 3205 1835
rect 3205 1805 3235 1835
rect 3235 1805 3236 1835
rect 3204 1804 3236 1805
rect 3204 1755 3236 1756
rect 3204 1725 3205 1755
rect 3205 1725 3235 1755
rect 3235 1725 3236 1755
rect 3204 1724 3236 1725
rect 3284 2475 3316 2476
rect 3284 2445 3285 2475
rect 3285 2445 3315 2475
rect 3315 2445 3316 2475
rect 3284 2444 3316 2445
rect 3284 2364 3316 2396
rect 3284 2315 3316 2316
rect 3284 2285 3285 2315
rect 3285 2285 3315 2315
rect 3315 2285 3316 2315
rect 3284 2284 3316 2285
rect 3284 2204 3316 2236
rect 3284 2155 3316 2156
rect 3284 2125 3285 2155
rect 3285 2125 3315 2155
rect 3315 2125 3316 2155
rect 3284 2124 3316 2125
rect 3284 2075 3316 2076
rect 3284 2045 3285 2075
rect 3285 2045 3315 2075
rect 3315 2045 3316 2075
rect 3284 2044 3316 2045
rect 3284 1995 3316 1996
rect 3284 1965 3285 1995
rect 3285 1965 3315 1995
rect 3315 1965 3316 1995
rect 3284 1964 3316 1965
rect 3284 1915 3316 1916
rect 3284 1885 3285 1915
rect 3285 1885 3315 1915
rect 3315 1885 3316 1915
rect 3284 1884 3316 1885
rect 3284 1835 3316 1836
rect 3284 1805 3285 1835
rect 3285 1805 3315 1835
rect 3315 1805 3316 1835
rect 3284 1804 3316 1805
rect 3284 1755 3316 1756
rect 3284 1725 3285 1755
rect 3285 1725 3315 1755
rect 3315 1725 3316 1755
rect 3284 1724 3316 1725
rect 3364 2475 3396 2476
rect 3364 2445 3365 2475
rect 3365 2445 3395 2475
rect 3395 2445 3396 2475
rect 3364 2444 3396 2445
rect 3364 2364 3396 2396
rect 3364 2315 3396 2316
rect 3364 2285 3365 2315
rect 3365 2285 3395 2315
rect 3395 2285 3396 2315
rect 3364 2284 3396 2285
rect 3364 2204 3396 2236
rect 3364 2155 3396 2156
rect 3364 2125 3365 2155
rect 3365 2125 3395 2155
rect 3395 2125 3396 2155
rect 3364 2124 3396 2125
rect 3364 2075 3396 2076
rect 3364 2045 3365 2075
rect 3365 2045 3395 2075
rect 3395 2045 3396 2075
rect 3364 2044 3396 2045
rect 3364 1995 3396 1996
rect 3364 1965 3365 1995
rect 3365 1965 3395 1995
rect 3395 1965 3396 1995
rect 3364 1964 3396 1965
rect 3364 1915 3396 1916
rect 3364 1885 3365 1915
rect 3365 1885 3395 1915
rect 3395 1885 3396 1915
rect 3364 1884 3396 1885
rect 3364 1835 3396 1836
rect 3364 1805 3365 1835
rect 3365 1805 3395 1835
rect 3395 1805 3396 1835
rect 3364 1804 3396 1805
rect 3364 1755 3396 1756
rect 3364 1725 3365 1755
rect 3365 1725 3395 1755
rect 3395 1725 3396 1755
rect 3364 1724 3396 1725
rect 3444 2475 3476 2476
rect 3444 2445 3445 2475
rect 3445 2445 3475 2475
rect 3475 2445 3476 2475
rect 3444 2444 3476 2445
rect 3444 2364 3476 2396
rect 3444 2315 3476 2316
rect 3444 2285 3445 2315
rect 3445 2285 3475 2315
rect 3475 2285 3476 2315
rect 3444 2284 3476 2285
rect 3444 2204 3476 2236
rect 3444 2155 3476 2156
rect 3444 2125 3445 2155
rect 3445 2125 3475 2155
rect 3475 2125 3476 2155
rect 3444 2124 3476 2125
rect 3444 2075 3476 2076
rect 3444 2045 3445 2075
rect 3445 2045 3475 2075
rect 3475 2045 3476 2075
rect 3444 2044 3476 2045
rect 3444 1995 3476 1996
rect 3444 1965 3445 1995
rect 3445 1965 3475 1995
rect 3475 1965 3476 1995
rect 3444 1964 3476 1965
rect 3444 1915 3476 1916
rect 3444 1885 3445 1915
rect 3445 1885 3475 1915
rect 3475 1885 3476 1915
rect 3444 1884 3476 1885
rect 3444 1835 3476 1836
rect 3444 1805 3445 1835
rect 3445 1805 3475 1835
rect 3475 1805 3476 1835
rect 3444 1804 3476 1805
rect 3444 1755 3476 1756
rect 3444 1725 3445 1755
rect 3445 1725 3475 1755
rect 3475 1725 3476 1755
rect 3444 1724 3476 1725
rect 3524 2475 3556 2476
rect 3524 2445 3525 2475
rect 3525 2445 3555 2475
rect 3555 2445 3556 2475
rect 3524 2444 3556 2445
rect 3524 2364 3556 2396
rect 3524 2315 3556 2316
rect 3524 2285 3525 2315
rect 3525 2285 3555 2315
rect 3555 2285 3556 2315
rect 3524 2284 3556 2285
rect 3524 2204 3556 2236
rect 3524 2155 3556 2156
rect 3524 2125 3525 2155
rect 3525 2125 3555 2155
rect 3555 2125 3556 2155
rect 3524 2124 3556 2125
rect 3524 2075 3556 2076
rect 3524 2045 3525 2075
rect 3525 2045 3555 2075
rect 3555 2045 3556 2075
rect 3524 2044 3556 2045
rect 3524 1995 3556 1996
rect 3524 1965 3525 1995
rect 3525 1965 3555 1995
rect 3555 1965 3556 1995
rect 3524 1964 3556 1965
rect 3524 1915 3556 1916
rect 3524 1885 3525 1915
rect 3525 1885 3555 1915
rect 3555 1885 3556 1915
rect 3524 1884 3556 1885
rect 3524 1835 3556 1836
rect 3524 1805 3525 1835
rect 3525 1805 3555 1835
rect 3555 1805 3556 1835
rect 3524 1804 3556 1805
rect 3524 1755 3556 1756
rect 3524 1725 3525 1755
rect 3525 1725 3555 1755
rect 3555 1725 3556 1755
rect 3524 1724 3556 1725
rect 3604 2475 3636 2476
rect 3604 2445 3605 2475
rect 3605 2445 3635 2475
rect 3635 2445 3636 2475
rect 3604 2444 3636 2445
rect 3604 2364 3636 2396
rect 3604 2315 3636 2316
rect 3604 2285 3605 2315
rect 3605 2285 3635 2315
rect 3635 2285 3636 2315
rect 3604 2284 3636 2285
rect 3604 2204 3636 2236
rect 3604 2155 3636 2156
rect 3604 2125 3605 2155
rect 3605 2125 3635 2155
rect 3635 2125 3636 2155
rect 3604 2124 3636 2125
rect 3604 2075 3636 2076
rect 3604 2045 3605 2075
rect 3605 2045 3635 2075
rect 3635 2045 3636 2075
rect 3604 2044 3636 2045
rect 3604 1995 3636 1996
rect 3604 1965 3605 1995
rect 3605 1965 3635 1995
rect 3635 1965 3636 1995
rect 3604 1964 3636 1965
rect 3604 1915 3636 1916
rect 3604 1885 3605 1915
rect 3605 1885 3635 1915
rect 3635 1885 3636 1915
rect 3604 1884 3636 1885
rect 3604 1835 3636 1836
rect 3604 1805 3605 1835
rect 3605 1805 3635 1835
rect 3635 1805 3636 1835
rect 3604 1804 3636 1805
rect 3604 1755 3636 1756
rect 3604 1725 3605 1755
rect 3605 1725 3635 1755
rect 3635 1725 3636 1755
rect 3604 1724 3636 1725
rect 3684 2475 3716 2476
rect 3684 2445 3685 2475
rect 3685 2445 3715 2475
rect 3715 2445 3716 2475
rect 3684 2444 3716 2445
rect 3684 2364 3716 2396
rect 3684 2315 3716 2316
rect 3684 2285 3685 2315
rect 3685 2285 3715 2315
rect 3715 2285 3716 2315
rect 3684 2284 3716 2285
rect 3684 2204 3716 2236
rect 3684 2155 3716 2156
rect 3684 2125 3685 2155
rect 3685 2125 3715 2155
rect 3715 2125 3716 2155
rect 3684 2124 3716 2125
rect 3684 2075 3716 2076
rect 3684 2045 3685 2075
rect 3685 2045 3715 2075
rect 3715 2045 3716 2075
rect 3684 2044 3716 2045
rect 3684 1995 3716 1996
rect 3684 1965 3685 1995
rect 3685 1965 3715 1995
rect 3715 1965 3716 1995
rect 3684 1964 3716 1965
rect 3684 1915 3716 1916
rect 3684 1885 3685 1915
rect 3685 1885 3715 1915
rect 3715 1885 3716 1915
rect 3684 1884 3716 1885
rect 3684 1835 3716 1836
rect 3684 1805 3685 1835
rect 3685 1805 3715 1835
rect 3715 1805 3716 1835
rect 3684 1804 3716 1805
rect 3684 1755 3716 1756
rect 3684 1725 3685 1755
rect 3685 1725 3715 1755
rect 3715 1725 3716 1755
rect 3684 1724 3716 1725
rect 3764 2475 3796 2476
rect 3764 2445 3765 2475
rect 3765 2445 3795 2475
rect 3795 2445 3796 2475
rect 3764 2444 3796 2445
rect 3764 2364 3796 2396
rect 3764 2315 3796 2316
rect 3764 2285 3765 2315
rect 3765 2285 3795 2315
rect 3795 2285 3796 2315
rect 3764 2284 3796 2285
rect 3764 2204 3796 2236
rect 3764 2155 3796 2156
rect 3764 2125 3765 2155
rect 3765 2125 3795 2155
rect 3795 2125 3796 2155
rect 3764 2124 3796 2125
rect 3764 2075 3796 2076
rect 3764 2045 3765 2075
rect 3765 2045 3795 2075
rect 3795 2045 3796 2075
rect 3764 2044 3796 2045
rect 3764 1995 3796 1996
rect 3764 1965 3765 1995
rect 3765 1965 3795 1995
rect 3795 1965 3796 1995
rect 3764 1964 3796 1965
rect 3764 1915 3796 1916
rect 3764 1885 3765 1915
rect 3765 1885 3795 1915
rect 3795 1885 3796 1915
rect 3764 1884 3796 1885
rect 3764 1835 3796 1836
rect 3764 1805 3765 1835
rect 3765 1805 3795 1835
rect 3795 1805 3796 1835
rect 3764 1804 3796 1805
rect 3764 1755 3796 1756
rect 3764 1725 3765 1755
rect 3765 1725 3795 1755
rect 3795 1725 3796 1755
rect 3764 1724 3796 1725
rect 3844 2475 3876 2476
rect 3844 2445 3845 2475
rect 3845 2445 3875 2475
rect 3875 2445 3876 2475
rect 3844 2444 3876 2445
rect 3844 2364 3876 2396
rect 3844 2315 3876 2316
rect 3844 2285 3845 2315
rect 3845 2285 3875 2315
rect 3875 2285 3876 2315
rect 3844 2284 3876 2285
rect 3844 2204 3876 2236
rect 3844 2155 3876 2156
rect 3844 2125 3845 2155
rect 3845 2125 3875 2155
rect 3875 2125 3876 2155
rect 3844 2124 3876 2125
rect 3844 2075 3876 2076
rect 3844 2045 3845 2075
rect 3845 2045 3875 2075
rect 3875 2045 3876 2075
rect 3844 2044 3876 2045
rect 3844 1995 3876 1996
rect 3844 1965 3845 1995
rect 3845 1965 3875 1995
rect 3875 1965 3876 1995
rect 3844 1964 3876 1965
rect 3844 1915 3876 1916
rect 3844 1885 3845 1915
rect 3845 1885 3875 1915
rect 3875 1885 3876 1915
rect 3844 1884 3876 1885
rect 3844 1835 3876 1836
rect 3844 1805 3845 1835
rect 3845 1805 3875 1835
rect 3875 1805 3876 1835
rect 3844 1804 3876 1805
rect 3844 1755 3876 1756
rect 3844 1725 3845 1755
rect 3845 1725 3875 1755
rect 3875 1725 3876 1755
rect 3844 1724 3876 1725
rect 3924 2475 3956 2476
rect 3924 2445 3925 2475
rect 3925 2445 3955 2475
rect 3955 2445 3956 2475
rect 3924 2444 3956 2445
rect 3924 2364 3956 2396
rect 3924 2315 3956 2316
rect 3924 2285 3925 2315
rect 3925 2285 3955 2315
rect 3955 2285 3956 2315
rect 3924 2284 3956 2285
rect 3924 2204 3956 2236
rect 3924 2155 3956 2156
rect 3924 2125 3925 2155
rect 3925 2125 3955 2155
rect 3955 2125 3956 2155
rect 3924 2124 3956 2125
rect 3924 2075 3956 2076
rect 3924 2045 3925 2075
rect 3925 2045 3955 2075
rect 3955 2045 3956 2075
rect 3924 2044 3956 2045
rect 3924 1995 3956 1996
rect 3924 1965 3925 1995
rect 3925 1965 3955 1995
rect 3955 1965 3956 1995
rect 3924 1964 3956 1965
rect 3924 1915 3956 1916
rect 3924 1885 3925 1915
rect 3925 1885 3955 1915
rect 3955 1885 3956 1915
rect 3924 1884 3956 1885
rect 3924 1835 3956 1836
rect 3924 1805 3925 1835
rect 3925 1805 3955 1835
rect 3955 1805 3956 1835
rect 3924 1804 3956 1805
rect 3924 1755 3956 1756
rect 3924 1725 3925 1755
rect 3925 1725 3955 1755
rect 3955 1725 3956 1755
rect 3924 1724 3956 1725
rect 4004 2475 4036 2476
rect 4004 2445 4005 2475
rect 4005 2445 4035 2475
rect 4035 2445 4036 2475
rect 4004 2444 4036 2445
rect 4004 2364 4036 2396
rect 4004 2315 4036 2316
rect 4004 2285 4005 2315
rect 4005 2285 4035 2315
rect 4035 2285 4036 2315
rect 4004 2284 4036 2285
rect 4004 2204 4036 2236
rect 4004 2155 4036 2156
rect 4004 2125 4005 2155
rect 4005 2125 4035 2155
rect 4035 2125 4036 2155
rect 4004 2124 4036 2125
rect 4004 2075 4036 2076
rect 4004 2045 4005 2075
rect 4005 2045 4035 2075
rect 4035 2045 4036 2075
rect 4004 2044 4036 2045
rect 4004 1995 4036 1996
rect 4004 1965 4005 1995
rect 4005 1965 4035 1995
rect 4035 1965 4036 1995
rect 4004 1964 4036 1965
rect 4004 1915 4036 1916
rect 4004 1885 4005 1915
rect 4005 1885 4035 1915
rect 4035 1885 4036 1915
rect 4004 1884 4036 1885
rect 4004 1835 4036 1836
rect 4004 1805 4005 1835
rect 4005 1805 4035 1835
rect 4035 1805 4036 1835
rect 4004 1804 4036 1805
rect 4004 1755 4036 1756
rect 4004 1725 4005 1755
rect 4005 1725 4035 1755
rect 4035 1725 4036 1755
rect 4004 1724 4036 1725
rect 4084 2475 4116 2476
rect 4084 2445 4085 2475
rect 4085 2445 4115 2475
rect 4115 2445 4116 2475
rect 4084 2444 4116 2445
rect 4084 2364 4116 2396
rect 4084 2315 4116 2316
rect 4084 2285 4085 2315
rect 4085 2285 4115 2315
rect 4115 2285 4116 2315
rect 4084 2284 4116 2285
rect 4084 2204 4116 2236
rect 4084 2155 4116 2156
rect 4084 2125 4085 2155
rect 4085 2125 4115 2155
rect 4115 2125 4116 2155
rect 4084 2124 4116 2125
rect 4084 2075 4116 2076
rect 4084 2045 4085 2075
rect 4085 2045 4115 2075
rect 4115 2045 4116 2075
rect 4084 2044 4116 2045
rect 4084 1995 4116 1996
rect 4084 1965 4085 1995
rect 4085 1965 4115 1995
rect 4115 1965 4116 1995
rect 4084 1964 4116 1965
rect 4084 1915 4116 1916
rect 4084 1885 4085 1915
rect 4085 1885 4115 1915
rect 4115 1885 4116 1915
rect 4084 1884 4116 1885
rect 4084 1835 4116 1836
rect 4084 1805 4085 1835
rect 4085 1805 4115 1835
rect 4115 1805 4116 1835
rect 4084 1804 4116 1805
rect 4084 1755 4116 1756
rect 4084 1725 4085 1755
rect 4085 1725 4115 1755
rect 4115 1725 4116 1755
rect 4084 1724 4116 1725
rect 4164 2475 4196 2476
rect 4164 2445 4165 2475
rect 4165 2445 4195 2475
rect 4195 2445 4196 2475
rect 4164 2444 4196 2445
rect 4164 2364 4196 2396
rect 4164 2315 4196 2316
rect 4164 2285 4165 2315
rect 4165 2285 4195 2315
rect 4195 2285 4196 2315
rect 4164 2284 4196 2285
rect 4164 2204 4196 2236
rect 4164 2155 4196 2156
rect 4164 2125 4165 2155
rect 4165 2125 4195 2155
rect 4195 2125 4196 2155
rect 4164 2124 4196 2125
rect 4164 2075 4196 2076
rect 4164 2045 4165 2075
rect 4165 2045 4195 2075
rect 4195 2045 4196 2075
rect 4164 2044 4196 2045
rect 4164 1995 4196 1996
rect 4164 1965 4165 1995
rect 4165 1965 4195 1995
rect 4195 1965 4196 1995
rect 4164 1964 4196 1965
rect 4164 1915 4196 1916
rect 4164 1885 4165 1915
rect 4165 1885 4195 1915
rect 4195 1885 4196 1915
rect 4164 1884 4196 1885
rect 4164 1835 4196 1836
rect 4164 1805 4165 1835
rect 4165 1805 4195 1835
rect 4195 1805 4196 1835
rect 4164 1804 4196 1805
rect 4164 1755 4196 1756
rect 4164 1725 4165 1755
rect 4165 1725 4195 1755
rect 4195 1725 4196 1755
rect 4164 1724 4196 1725
rect 4244 2475 4276 2476
rect 4244 2445 4245 2475
rect 4245 2445 4275 2475
rect 4275 2445 4276 2475
rect 4244 2444 4276 2445
rect 4244 2364 4276 2396
rect 4244 2315 4276 2316
rect 4244 2285 4245 2315
rect 4245 2285 4275 2315
rect 4275 2285 4276 2315
rect 4244 2284 4276 2285
rect 4244 2204 4276 2236
rect 4244 2155 4276 2156
rect 4244 2125 4245 2155
rect 4245 2125 4275 2155
rect 4275 2125 4276 2155
rect 4244 2124 4276 2125
rect 4244 2075 4276 2076
rect 4244 2045 4245 2075
rect 4245 2045 4275 2075
rect 4275 2045 4276 2075
rect 4244 2044 4276 2045
rect 4244 1995 4276 1996
rect 4244 1965 4245 1995
rect 4245 1965 4275 1995
rect 4275 1965 4276 1995
rect 4244 1964 4276 1965
rect 4244 1915 4276 1916
rect 4244 1885 4245 1915
rect 4245 1885 4275 1915
rect 4275 1885 4276 1915
rect 4244 1884 4276 1885
rect 4244 1835 4276 1836
rect 4244 1805 4245 1835
rect 4245 1805 4275 1835
rect 4275 1805 4276 1835
rect 4244 1804 4276 1805
rect 4244 1755 4276 1756
rect 4244 1725 4245 1755
rect 4245 1725 4275 1755
rect 4275 1725 4276 1755
rect 4244 1724 4276 1725
rect 4324 2475 4356 2476
rect 4324 2445 4325 2475
rect 4325 2445 4355 2475
rect 4355 2445 4356 2475
rect 4324 2444 4356 2445
rect 4324 2364 4356 2396
rect 4324 2315 4356 2316
rect 4324 2285 4325 2315
rect 4325 2285 4355 2315
rect 4355 2285 4356 2315
rect 4324 2284 4356 2285
rect 4324 2204 4356 2236
rect 4324 2155 4356 2156
rect 4324 2125 4325 2155
rect 4325 2125 4355 2155
rect 4355 2125 4356 2155
rect 4324 2124 4356 2125
rect 4324 2075 4356 2076
rect 4324 2045 4325 2075
rect 4325 2045 4355 2075
rect 4355 2045 4356 2075
rect 4324 2044 4356 2045
rect 4324 1995 4356 1996
rect 4324 1965 4325 1995
rect 4325 1965 4355 1995
rect 4355 1965 4356 1995
rect 4324 1964 4356 1965
rect 4324 1915 4356 1916
rect 4324 1885 4325 1915
rect 4325 1885 4355 1915
rect 4355 1885 4356 1915
rect 4324 1884 4356 1885
rect 4324 1835 4356 1836
rect 4324 1805 4325 1835
rect 4325 1805 4355 1835
rect 4355 1805 4356 1835
rect 4324 1804 4356 1805
rect 4324 1755 4356 1756
rect 4324 1725 4325 1755
rect 4325 1725 4355 1755
rect 4355 1725 4356 1755
rect 4324 1724 4356 1725
rect 4404 2475 4436 2476
rect 4404 2445 4405 2475
rect 4405 2445 4435 2475
rect 4435 2445 4436 2475
rect 4404 2444 4436 2445
rect 4404 2364 4436 2396
rect 4404 2315 4436 2316
rect 4404 2285 4405 2315
rect 4405 2285 4435 2315
rect 4435 2285 4436 2315
rect 4404 2284 4436 2285
rect 4404 2204 4436 2236
rect 4404 2155 4436 2156
rect 4404 2125 4405 2155
rect 4405 2125 4435 2155
rect 4435 2125 4436 2155
rect 4404 2124 4436 2125
rect 4404 2075 4436 2076
rect 4404 2045 4405 2075
rect 4405 2045 4435 2075
rect 4435 2045 4436 2075
rect 4404 2044 4436 2045
rect 4404 1995 4436 1996
rect 4404 1965 4405 1995
rect 4405 1965 4435 1995
rect 4435 1965 4436 1995
rect 4404 1964 4436 1965
rect 4404 1915 4436 1916
rect 4404 1885 4405 1915
rect 4405 1885 4435 1915
rect 4435 1885 4436 1915
rect 4404 1884 4436 1885
rect 4404 1835 4436 1836
rect 4404 1805 4405 1835
rect 4405 1805 4435 1835
rect 4435 1805 4436 1835
rect 4404 1804 4436 1805
rect 4404 1755 4436 1756
rect 4404 1725 4405 1755
rect 4405 1725 4435 1755
rect 4435 1725 4436 1755
rect 4404 1724 4436 1725
rect 4484 2475 4516 2476
rect 4484 2445 4485 2475
rect 4485 2445 4515 2475
rect 4515 2445 4516 2475
rect 4484 2444 4516 2445
rect 4484 2364 4516 2396
rect 4484 2315 4516 2316
rect 4484 2285 4485 2315
rect 4485 2285 4515 2315
rect 4515 2285 4516 2315
rect 4484 2284 4516 2285
rect 4484 2204 4516 2236
rect 4484 2155 4516 2156
rect 4484 2125 4485 2155
rect 4485 2125 4515 2155
rect 4515 2125 4516 2155
rect 4484 2124 4516 2125
rect 4484 2075 4516 2076
rect 4484 2045 4485 2075
rect 4485 2045 4515 2075
rect 4515 2045 4516 2075
rect 4484 2044 4516 2045
rect 4484 1995 4516 1996
rect 4484 1965 4485 1995
rect 4485 1965 4515 1995
rect 4515 1965 4516 1995
rect 4484 1964 4516 1965
rect 4484 1915 4516 1916
rect 4484 1885 4485 1915
rect 4485 1885 4515 1915
rect 4515 1885 4516 1915
rect 4484 1884 4516 1885
rect 4484 1835 4516 1836
rect 4484 1805 4485 1835
rect 4485 1805 4515 1835
rect 4515 1805 4516 1835
rect 4484 1804 4516 1805
rect 4484 1755 4516 1756
rect 4484 1725 4485 1755
rect 4485 1725 4515 1755
rect 4515 1725 4516 1755
rect 4484 1724 4516 1725
rect 4564 2475 4596 2476
rect 4564 2445 4565 2475
rect 4565 2445 4595 2475
rect 4595 2445 4596 2475
rect 4564 2444 4596 2445
rect 4564 2364 4596 2396
rect 4564 2315 4596 2316
rect 4564 2285 4565 2315
rect 4565 2285 4595 2315
rect 4595 2285 4596 2315
rect 4564 2284 4596 2285
rect 4564 2204 4596 2236
rect 4564 2155 4596 2156
rect 4564 2125 4565 2155
rect 4565 2125 4595 2155
rect 4595 2125 4596 2155
rect 4564 2124 4596 2125
rect 4564 2075 4596 2076
rect 4564 2045 4565 2075
rect 4565 2045 4595 2075
rect 4595 2045 4596 2075
rect 4564 2044 4596 2045
rect 4564 1995 4596 1996
rect 4564 1965 4565 1995
rect 4565 1965 4595 1995
rect 4595 1965 4596 1995
rect 4564 1964 4596 1965
rect 4564 1915 4596 1916
rect 4564 1885 4565 1915
rect 4565 1885 4595 1915
rect 4595 1885 4596 1915
rect 4564 1884 4596 1885
rect 4564 1835 4596 1836
rect 4564 1805 4565 1835
rect 4565 1805 4595 1835
rect 4595 1805 4596 1835
rect 4564 1804 4596 1805
rect 4564 1755 4596 1756
rect 4564 1725 4565 1755
rect 4565 1725 4595 1755
rect 4595 1725 4596 1755
rect 4564 1724 4596 1725
rect 4644 2475 4676 2476
rect 4644 2445 4645 2475
rect 4645 2445 4675 2475
rect 4675 2445 4676 2475
rect 4644 2444 4676 2445
rect 4644 2364 4676 2396
rect 4644 2315 4676 2316
rect 4644 2285 4645 2315
rect 4645 2285 4675 2315
rect 4675 2285 4676 2315
rect 4644 2284 4676 2285
rect 4644 2204 4676 2236
rect 4644 2155 4676 2156
rect 4644 2125 4645 2155
rect 4645 2125 4675 2155
rect 4675 2125 4676 2155
rect 4644 2124 4676 2125
rect 4644 2075 4676 2076
rect 4644 2045 4645 2075
rect 4645 2045 4675 2075
rect 4675 2045 4676 2075
rect 4644 2044 4676 2045
rect 4644 1995 4676 1996
rect 4644 1965 4645 1995
rect 4645 1965 4675 1995
rect 4675 1965 4676 1995
rect 4644 1964 4676 1965
rect 4644 1915 4676 1916
rect 4644 1885 4645 1915
rect 4645 1885 4675 1915
rect 4675 1885 4676 1915
rect 4644 1884 4676 1885
rect 4644 1835 4676 1836
rect 4644 1805 4645 1835
rect 4645 1805 4675 1835
rect 4675 1805 4676 1835
rect 4644 1804 4676 1805
rect 4644 1755 4676 1756
rect 4644 1725 4645 1755
rect 4645 1725 4675 1755
rect 4675 1725 4676 1755
rect 4644 1724 4676 1725
rect 4724 2475 4756 2476
rect 4724 2445 4725 2475
rect 4725 2445 4755 2475
rect 4755 2445 4756 2475
rect 4724 2444 4756 2445
rect 4724 2364 4756 2396
rect 4724 2315 4756 2316
rect 4724 2285 4725 2315
rect 4725 2285 4755 2315
rect 4755 2285 4756 2315
rect 4724 2284 4756 2285
rect 4724 2204 4756 2236
rect 4724 2155 4756 2156
rect 4724 2125 4725 2155
rect 4725 2125 4755 2155
rect 4755 2125 4756 2155
rect 4724 2124 4756 2125
rect 4724 2075 4756 2076
rect 4724 2045 4725 2075
rect 4725 2045 4755 2075
rect 4755 2045 4756 2075
rect 4724 2044 4756 2045
rect 4724 1995 4756 1996
rect 4724 1965 4725 1995
rect 4725 1965 4755 1995
rect 4755 1965 4756 1995
rect 4724 1964 4756 1965
rect 4724 1915 4756 1916
rect 4724 1885 4725 1915
rect 4725 1885 4755 1915
rect 4755 1885 4756 1915
rect 4724 1884 4756 1885
rect 4724 1835 4756 1836
rect 4724 1805 4725 1835
rect 4725 1805 4755 1835
rect 4755 1805 4756 1835
rect 4724 1804 4756 1805
rect 4724 1755 4756 1756
rect 4724 1725 4725 1755
rect 4725 1725 4755 1755
rect 4755 1725 4756 1755
rect 4724 1724 4756 1725
rect 4804 2475 4836 2476
rect 4804 2445 4805 2475
rect 4805 2445 4835 2475
rect 4835 2445 4836 2475
rect 4804 2444 4836 2445
rect 4804 2364 4836 2396
rect 4804 2315 4836 2316
rect 4804 2285 4805 2315
rect 4805 2285 4835 2315
rect 4835 2285 4836 2315
rect 4804 2284 4836 2285
rect 4804 2204 4836 2236
rect 4804 2155 4836 2156
rect 4804 2125 4805 2155
rect 4805 2125 4835 2155
rect 4835 2125 4836 2155
rect 4804 2124 4836 2125
rect 4804 2075 4836 2076
rect 4804 2045 4805 2075
rect 4805 2045 4835 2075
rect 4835 2045 4836 2075
rect 4804 2044 4836 2045
rect 4804 1995 4836 1996
rect 4804 1965 4805 1995
rect 4805 1965 4835 1995
rect 4835 1965 4836 1995
rect 4804 1964 4836 1965
rect 4804 1915 4836 1916
rect 4804 1885 4805 1915
rect 4805 1885 4835 1915
rect 4835 1885 4836 1915
rect 4804 1884 4836 1885
rect 4804 1835 4836 1836
rect 4804 1805 4805 1835
rect 4805 1805 4835 1835
rect 4835 1805 4836 1835
rect 4804 1804 4836 1805
rect 4804 1755 4836 1756
rect 4804 1725 4805 1755
rect 4805 1725 4835 1755
rect 4835 1725 4836 1755
rect 4804 1724 4836 1725
rect 4884 2475 4916 2476
rect 4884 2445 4885 2475
rect 4885 2445 4915 2475
rect 4915 2445 4916 2475
rect 4884 2444 4916 2445
rect 4884 2364 4916 2396
rect 4884 2315 4916 2316
rect 4884 2285 4885 2315
rect 4885 2285 4915 2315
rect 4915 2285 4916 2315
rect 4884 2284 4916 2285
rect 4884 2204 4916 2236
rect 4884 2155 4916 2156
rect 4884 2125 4885 2155
rect 4885 2125 4915 2155
rect 4915 2125 4916 2155
rect 4884 2124 4916 2125
rect 4884 2075 4916 2076
rect 4884 2045 4885 2075
rect 4885 2045 4915 2075
rect 4915 2045 4916 2075
rect 4884 2044 4916 2045
rect 4884 1995 4916 1996
rect 4884 1965 4885 1995
rect 4885 1965 4915 1995
rect 4915 1965 4916 1995
rect 4884 1964 4916 1965
rect 4884 1915 4916 1916
rect 4884 1885 4885 1915
rect 4885 1885 4915 1915
rect 4915 1885 4916 1915
rect 4884 1884 4916 1885
rect 4884 1835 4916 1836
rect 4884 1805 4885 1835
rect 4885 1805 4915 1835
rect 4915 1805 4916 1835
rect 4884 1804 4916 1805
rect 4884 1755 4916 1756
rect 4884 1725 4885 1755
rect 4885 1725 4915 1755
rect 4915 1725 4916 1755
rect 4884 1724 4916 1725
rect -876 1675 -844 1676
rect -876 1645 -875 1675
rect -875 1645 -845 1675
rect -845 1645 -844 1675
rect -876 1644 -844 1645
rect -876 1595 -844 1596
rect -876 1565 -875 1595
rect -875 1565 -845 1595
rect -845 1565 -844 1595
rect -876 1564 -844 1565
rect -876 1484 -844 1516
rect -876 1435 -844 1436
rect -876 1405 -875 1435
rect -875 1405 -845 1435
rect -845 1405 -844 1435
rect -876 1404 -844 1405
rect -876 1355 -844 1356
rect -876 1325 -875 1355
rect -875 1325 -845 1355
rect -845 1325 -844 1355
rect -876 1324 -844 1325
rect -876 1275 -844 1276
rect -876 1245 -875 1275
rect -875 1245 -845 1275
rect -845 1245 -844 1275
rect -876 1244 -844 1245
rect -876 1195 -844 1196
rect -876 1165 -875 1195
rect -875 1165 -845 1195
rect -845 1165 -844 1195
rect -876 1164 -844 1165
rect -876 1084 -844 1116
rect -876 1035 -844 1036
rect -876 1005 -875 1035
rect -875 1005 -845 1035
rect -845 1005 -844 1035
rect -876 1004 -844 1005
rect -876 955 -844 956
rect -876 925 -875 955
rect -875 925 -845 955
rect -845 925 -844 955
rect -876 924 -844 925
rect -796 1675 -764 1676
rect -796 1645 -795 1675
rect -795 1645 -765 1675
rect -765 1645 -764 1675
rect -796 1644 -764 1645
rect -796 1595 -764 1596
rect -796 1565 -795 1595
rect -795 1565 -765 1595
rect -765 1565 -764 1595
rect -796 1564 -764 1565
rect -796 1484 -764 1516
rect -796 1435 -764 1436
rect -796 1405 -795 1435
rect -795 1405 -765 1435
rect -765 1405 -764 1435
rect -796 1404 -764 1405
rect -796 1355 -764 1356
rect -796 1325 -795 1355
rect -795 1325 -765 1355
rect -765 1325 -764 1355
rect -796 1324 -764 1325
rect -796 1275 -764 1276
rect -796 1245 -795 1275
rect -795 1245 -765 1275
rect -765 1245 -764 1275
rect -796 1244 -764 1245
rect -796 1195 -764 1196
rect -796 1165 -795 1195
rect -795 1165 -765 1195
rect -765 1165 -764 1195
rect -796 1164 -764 1165
rect -796 1084 -764 1116
rect -796 1035 -764 1036
rect -796 1005 -795 1035
rect -795 1005 -765 1035
rect -765 1005 -764 1035
rect -796 1004 -764 1005
rect -796 955 -764 956
rect -796 925 -795 955
rect -795 925 -765 955
rect -765 925 -764 955
rect -796 924 -764 925
rect -716 1675 -684 1676
rect -716 1645 -715 1675
rect -715 1645 -685 1675
rect -685 1645 -684 1675
rect -716 1644 -684 1645
rect -716 1595 -684 1596
rect -716 1565 -715 1595
rect -715 1565 -685 1595
rect -685 1565 -684 1595
rect -716 1564 -684 1565
rect -716 1484 -684 1516
rect -716 1435 -684 1436
rect -716 1405 -715 1435
rect -715 1405 -685 1435
rect -685 1405 -684 1435
rect -716 1404 -684 1405
rect -716 1355 -684 1356
rect -716 1325 -715 1355
rect -715 1325 -685 1355
rect -685 1325 -684 1355
rect -716 1324 -684 1325
rect -716 1275 -684 1276
rect -716 1245 -715 1275
rect -715 1245 -685 1275
rect -685 1245 -684 1275
rect -716 1244 -684 1245
rect -716 1195 -684 1196
rect -716 1165 -715 1195
rect -715 1165 -685 1195
rect -685 1165 -684 1195
rect -716 1164 -684 1165
rect -716 1084 -684 1116
rect -716 1035 -684 1036
rect -716 1005 -715 1035
rect -715 1005 -685 1035
rect -685 1005 -684 1035
rect -716 1004 -684 1005
rect -716 955 -684 956
rect -716 925 -715 955
rect -715 925 -685 955
rect -685 925 -684 955
rect -716 924 -684 925
rect -636 1675 -604 1676
rect -636 1645 -635 1675
rect -635 1645 -605 1675
rect -605 1645 -604 1675
rect -636 1644 -604 1645
rect -636 1595 -604 1596
rect -636 1565 -635 1595
rect -635 1565 -605 1595
rect -605 1565 -604 1595
rect -636 1564 -604 1565
rect -636 1484 -604 1516
rect -636 1435 -604 1436
rect -636 1405 -635 1435
rect -635 1405 -605 1435
rect -605 1405 -604 1435
rect -636 1404 -604 1405
rect -636 1355 -604 1356
rect -636 1325 -635 1355
rect -635 1325 -605 1355
rect -605 1325 -604 1355
rect -636 1324 -604 1325
rect -636 1275 -604 1276
rect -636 1245 -635 1275
rect -635 1245 -605 1275
rect -605 1245 -604 1275
rect -636 1244 -604 1245
rect -636 1195 -604 1196
rect -636 1165 -635 1195
rect -635 1165 -605 1195
rect -605 1165 -604 1195
rect -636 1164 -604 1165
rect -636 1084 -604 1116
rect -636 1035 -604 1036
rect -636 1005 -635 1035
rect -635 1005 -605 1035
rect -605 1005 -604 1035
rect -636 1004 -604 1005
rect -636 955 -604 956
rect -636 925 -635 955
rect -635 925 -605 955
rect -605 925 -604 955
rect -636 924 -604 925
rect -556 1675 -524 1676
rect -556 1645 -555 1675
rect -555 1645 -525 1675
rect -525 1645 -524 1675
rect -556 1644 -524 1645
rect -556 1595 -524 1596
rect -556 1565 -555 1595
rect -555 1565 -525 1595
rect -525 1565 -524 1595
rect -556 1564 -524 1565
rect -556 1484 -524 1516
rect -556 1435 -524 1436
rect -556 1405 -555 1435
rect -555 1405 -525 1435
rect -525 1405 -524 1435
rect -556 1404 -524 1405
rect -556 1355 -524 1356
rect -556 1325 -555 1355
rect -555 1325 -525 1355
rect -525 1325 -524 1355
rect -556 1324 -524 1325
rect -556 1275 -524 1276
rect -556 1245 -555 1275
rect -555 1245 -525 1275
rect -525 1245 -524 1275
rect -556 1244 -524 1245
rect -556 1195 -524 1196
rect -556 1165 -555 1195
rect -555 1165 -525 1195
rect -525 1165 -524 1195
rect -556 1164 -524 1165
rect -556 1084 -524 1116
rect -556 1035 -524 1036
rect -556 1005 -555 1035
rect -555 1005 -525 1035
rect -525 1005 -524 1035
rect -556 1004 -524 1005
rect -556 955 -524 956
rect -556 925 -555 955
rect -555 925 -525 955
rect -525 925 -524 955
rect -556 924 -524 925
rect -476 1675 -444 1676
rect -476 1645 -475 1675
rect -475 1645 -445 1675
rect -445 1645 -444 1675
rect -476 1644 -444 1645
rect -476 1595 -444 1596
rect -476 1565 -475 1595
rect -475 1565 -445 1595
rect -445 1565 -444 1595
rect -476 1564 -444 1565
rect -476 1484 -444 1516
rect -476 1435 -444 1436
rect -476 1405 -475 1435
rect -475 1405 -445 1435
rect -445 1405 -444 1435
rect -476 1404 -444 1405
rect -476 1355 -444 1356
rect -476 1325 -475 1355
rect -475 1325 -445 1355
rect -445 1325 -444 1355
rect -476 1324 -444 1325
rect -476 1275 -444 1276
rect -476 1245 -475 1275
rect -475 1245 -445 1275
rect -445 1245 -444 1275
rect -476 1244 -444 1245
rect -476 1195 -444 1196
rect -476 1165 -475 1195
rect -475 1165 -445 1195
rect -445 1165 -444 1195
rect -476 1164 -444 1165
rect -476 1084 -444 1116
rect -476 1035 -444 1036
rect -476 1005 -475 1035
rect -475 1005 -445 1035
rect -445 1005 -444 1035
rect -476 1004 -444 1005
rect -476 955 -444 956
rect -476 925 -475 955
rect -475 925 -445 955
rect -445 925 -444 955
rect -476 924 -444 925
rect -396 1675 -364 1676
rect -396 1645 -395 1675
rect -395 1645 -365 1675
rect -365 1645 -364 1675
rect -396 1644 -364 1645
rect -396 1595 -364 1596
rect -396 1565 -395 1595
rect -395 1565 -365 1595
rect -365 1565 -364 1595
rect -396 1564 -364 1565
rect -396 1484 -364 1516
rect -396 1435 -364 1436
rect -396 1405 -395 1435
rect -395 1405 -365 1435
rect -365 1405 -364 1435
rect -396 1404 -364 1405
rect -396 1355 -364 1356
rect -396 1325 -395 1355
rect -395 1325 -365 1355
rect -365 1325 -364 1355
rect -396 1324 -364 1325
rect -396 1275 -364 1276
rect -396 1245 -395 1275
rect -395 1245 -365 1275
rect -365 1245 -364 1275
rect -396 1244 -364 1245
rect -396 1195 -364 1196
rect -396 1165 -395 1195
rect -395 1165 -365 1195
rect -365 1165 -364 1195
rect -396 1164 -364 1165
rect -396 1084 -364 1116
rect -396 1035 -364 1036
rect -396 1005 -395 1035
rect -395 1005 -365 1035
rect -365 1005 -364 1035
rect -396 1004 -364 1005
rect -396 955 -364 956
rect -396 925 -395 955
rect -395 925 -365 955
rect -365 925 -364 955
rect -396 924 -364 925
rect -316 1675 -284 1676
rect -316 1645 -315 1675
rect -315 1645 -285 1675
rect -285 1645 -284 1675
rect -316 1644 -284 1645
rect -316 1595 -284 1596
rect -316 1565 -315 1595
rect -315 1565 -285 1595
rect -285 1565 -284 1595
rect -316 1564 -284 1565
rect -316 1484 -284 1516
rect -316 1435 -284 1436
rect -316 1405 -315 1435
rect -315 1405 -285 1435
rect -285 1405 -284 1435
rect -316 1404 -284 1405
rect -316 1355 -284 1356
rect -316 1325 -315 1355
rect -315 1325 -285 1355
rect -285 1325 -284 1355
rect -316 1324 -284 1325
rect -316 1275 -284 1276
rect -316 1245 -315 1275
rect -315 1245 -285 1275
rect -285 1245 -284 1275
rect -316 1244 -284 1245
rect -316 1195 -284 1196
rect -316 1165 -315 1195
rect -315 1165 -285 1195
rect -285 1165 -284 1195
rect -316 1164 -284 1165
rect -316 1084 -284 1116
rect -316 1035 -284 1036
rect -316 1005 -315 1035
rect -315 1005 -285 1035
rect -285 1005 -284 1035
rect -316 1004 -284 1005
rect -316 955 -284 956
rect -316 925 -315 955
rect -315 925 -285 955
rect -285 925 -284 955
rect -316 924 -284 925
rect -236 1675 -204 1676
rect -236 1645 -235 1675
rect -235 1645 -205 1675
rect -205 1645 -204 1675
rect -236 1644 -204 1645
rect -236 1595 -204 1596
rect -236 1565 -235 1595
rect -235 1565 -205 1595
rect -205 1565 -204 1595
rect -236 1564 -204 1565
rect -236 1484 -204 1516
rect -236 1435 -204 1436
rect -236 1405 -235 1435
rect -235 1405 -205 1435
rect -205 1405 -204 1435
rect -236 1404 -204 1405
rect -236 1355 -204 1356
rect -236 1325 -235 1355
rect -235 1325 -205 1355
rect -205 1325 -204 1355
rect -236 1324 -204 1325
rect -236 1275 -204 1276
rect -236 1245 -235 1275
rect -235 1245 -205 1275
rect -205 1245 -204 1275
rect -236 1244 -204 1245
rect -236 1195 -204 1196
rect -236 1165 -235 1195
rect -235 1165 -205 1195
rect -205 1165 -204 1195
rect -236 1164 -204 1165
rect -236 1084 -204 1116
rect -236 1035 -204 1036
rect -236 1005 -235 1035
rect -235 1005 -205 1035
rect -205 1005 -204 1035
rect -236 1004 -204 1005
rect -236 955 -204 956
rect -236 925 -235 955
rect -235 925 -205 955
rect -205 925 -204 955
rect -236 924 -204 925
rect -156 1675 -124 1676
rect -156 1645 -155 1675
rect -155 1645 -125 1675
rect -125 1645 -124 1675
rect -156 1644 -124 1645
rect -156 1595 -124 1596
rect -156 1565 -155 1595
rect -155 1565 -125 1595
rect -125 1565 -124 1595
rect -156 1564 -124 1565
rect -156 1484 -124 1516
rect -156 1435 -124 1436
rect -156 1405 -155 1435
rect -155 1405 -125 1435
rect -125 1405 -124 1435
rect -156 1404 -124 1405
rect -156 1355 -124 1356
rect -156 1325 -155 1355
rect -155 1325 -125 1355
rect -125 1325 -124 1355
rect -156 1324 -124 1325
rect -156 1275 -124 1276
rect -156 1245 -155 1275
rect -155 1245 -125 1275
rect -125 1245 -124 1275
rect -156 1244 -124 1245
rect -156 1195 -124 1196
rect -156 1165 -155 1195
rect -155 1165 -125 1195
rect -125 1165 -124 1195
rect -156 1164 -124 1165
rect -156 1084 -124 1116
rect -156 1035 -124 1036
rect -156 1005 -155 1035
rect -155 1005 -125 1035
rect -125 1005 -124 1035
rect -156 1004 -124 1005
rect -156 955 -124 956
rect -156 925 -155 955
rect -155 925 -125 955
rect -125 925 -124 955
rect -156 924 -124 925
rect -76 1675 -44 1676
rect -76 1645 -75 1675
rect -75 1645 -45 1675
rect -45 1645 -44 1675
rect -76 1644 -44 1645
rect -76 1595 -44 1596
rect -76 1565 -75 1595
rect -75 1565 -45 1595
rect -45 1565 -44 1595
rect -76 1564 -44 1565
rect -76 1484 -44 1516
rect -76 1435 -44 1436
rect -76 1405 -75 1435
rect -75 1405 -45 1435
rect -45 1405 -44 1435
rect -76 1404 -44 1405
rect -76 1355 -44 1356
rect -76 1325 -75 1355
rect -75 1325 -45 1355
rect -45 1325 -44 1355
rect -76 1324 -44 1325
rect -76 1275 -44 1276
rect -76 1245 -75 1275
rect -75 1245 -45 1275
rect -45 1245 -44 1275
rect -76 1244 -44 1245
rect -76 1195 -44 1196
rect -76 1165 -75 1195
rect -75 1165 -45 1195
rect -45 1165 -44 1195
rect -76 1164 -44 1165
rect -76 1084 -44 1116
rect -76 1035 -44 1036
rect -76 1005 -75 1035
rect -75 1005 -45 1035
rect -45 1005 -44 1035
rect -76 1004 -44 1005
rect -76 955 -44 956
rect -76 925 -75 955
rect -75 925 -45 955
rect -45 925 -44 955
rect -76 924 -44 925
rect 4 1675 36 1676
rect 4 1645 5 1675
rect 5 1645 35 1675
rect 35 1645 36 1675
rect 4 1644 36 1645
rect 4 1595 36 1596
rect 4 1565 5 1595
rect 5 1565 35 1595
rect 35 1565 36 1595
rect 4 1564 36 1565
rect 4 1484 36 1516
rect 4 1435 36 1436
rect 4 1405 5 1435
rect 5 1405 35 1435
rect 35 1405 36 1435
rect 4 1404 36 1405
rect 4 1355 36 1356
rect 4 1325 5 1355
rect 5 1325 35 1355
rect 35 1325 36 1355
rect 4 1324 36 1325
rect 4 1275 36 1276
rect 4 1245 5 1275
rect 5 1245 35 1275
rect 35 1245 36 1275
rect 4 1244 36 1245
rect 4 1195 36 1196
rect 4 1165 5 1195
rect 5 1165 35 1195
rect 35 1165 36 1195
rect 4 1164 36 1165
rect 4 1084 36 1116
rect 4 1035 36 1036
rect 4 1005 5 1035
rect 5 1005 35 1035
rect 35 1005 36 1035
rect 4 1004 36 1005
rect 4 955 36 956
rect 4 925 5 955
rect 5 925 35 955
rect 35 925 36 955
rect 4 924 36 925
rect 84 1675 116 1676
rect 84 1645 85 1675
rect 85 1645 115 1675
rect 115 1645 116 1675
rect 84 1644 116 1645
rect 84 1595 116 1596
rect 84 1565 85 1595
rect 85 1565 115 1595
rect 115 1565 116 1595
rect 84 1564 116 1565
rect 84 1484 116 1516
rect 84 1435 116 1436
rect 84 1405 85 1435
rect 85 1405 115 1435
rect 115 1405 116 1435
rect 84 1404 116 1405
rect 84 1355 116 1356
rect 84 1325 85 1355
rect 85 1325 115 1355
rect 115 1325 116 1355
rect 84 1324 116 1325
rect 84 1275 116 1276
rect 84 1245 85 1275
rect 85 1245 115 1275
rect 115 1245 116 1275
rect 84 1244 116 1245
rect 84 1195 116 1196
rect 84 1165 85 1195
rect 85 1165 115 1195
rect 115 1165 116 1195
rect 84 1164 116 1165
rect 84 1084 116 1116
rect 84 1035 116 1036
rect 84 1005 85 1035
rect 85 1005 115 1035
rect 115 1005 116 1035
rect 84 1004 116 1005
rect 84 955 116 956
rect 84 925 85 955
rect 85 925 115 955
rect 115 925 116 955
rect 84 924 116 925
rect 164 1675 196 1676
rect 164 1645 165 1675
rect 165 1645 195 1675
rect 195 1645 196 1675
rect 164 1644 196 1645
rect 164 1595 196 1596
rect 164 1565 165 1595
rect 165 1565 195 1595
rect 195 1565 196 1595
rect 164 1564 196 1565
rect 164 1484 196 1516
rect 164 1435 196 1436
rect 164 1405 165 1435
rect 165 1405 195 1435
rect 195 1405 196 1435
rect 164 1404 196 1405
rect 164 1355 196 1356
rect 164 1325 165 1355
rect 165 1325 195 1355
rect 195 1325 196 1355
rect 164 1324 196 1325
rect 164 1275 196 1276
rect 164 1245 165 1275
rect 165 1245 195 1275
rect 195 1245 196 1275
rect 164 1244 196 1245
rect 164 1195 196 1196
rect 164 1165 165 1195
rect 165 1165 195 1195
rect 195 1165 196 1195
rect 164 1164 196 1165
rect 164 1084 196 1116
rect 164 1035 196 1036
rect 164 1005 165 1035
rect 165 1005 195 1035
rect 195 1005 196 1035
rect 164 1004 196 1005
rect 164 955 196 956
rect 164 925 165 955
rect 165 925 195 955
rect 195 925 196 955
rect 164 924 196 925
rect 244 1675 276 1676
rect 244 1645 245 1675
rect 245 1645 275 1675
rect 275 1645 276 1675
rect 244 1644 276 1645
rect 244 1595 276 1596
rect 244 1565 245 1595
rect 245 1565 275 1595
rect 275 1565 276 1595
rect 244 1564 276 1565
rect 244 1484 276 1516
rect 244 1435 276 1436
rect 244 1405 245 1435
rect 245 1405 275 1435
rect 275 1405 276 1435
rect 244 1404 276 1405
rect 244 1355 276 1356
rect 244 1325 245 1355
rect 245 1325 275 1355
rect 275 1325 276 1355
rect 244 1324 276 1325
rect 244 1275 276 1276
rect 244 1245 245 1275
rect 245 1245 275 1275
rect 275 1245 276 1275
rect 244 1244 276 1245
rect 244 1195 276 1196
rect 244 1165 245 1195
rect 245 1165 275 1195
rect 275 1165 276 1195
rect 244 1164 276 1165
rect 244 1084 276 1116
rect 244 1035 276 1036
rect 244 1005 245 1035
rect 245 1005 275 1035
rect 275 1005 276 1035
rect 244 1004 276 1005
rect 244 955 276 956
rect 244 925 245 955
rect 245 925 275 955
rect 275 925 276 955
rect 244 924 276 925
rect 324 1675 356 1676
rect 324 1645 325 1675
rect 325 1645 355 1675
rect 355 1645 356 1675
rect 324 1644 356 1645
rect 324 1595 356 1596
rect 324 1565 325 1595
rect 325 1565 355 1595
rect 355 1565 356 1595
rect 324 1564 356 1565
rect 324 1484 356 1516
rect 324 1435 356 1436
rect 324 1405 325 1435
rect 325 1405 355 1435
rect 355 1405 356 1435
rect 324 1404 356 1405
rect 324 1355 356 1356
rect 324 1325 325 1355
rect 325 1325 355 1355
rect 355 1325 356 1355
rect 324 1324 356 1325
rect 324 1275 356 1276
rect 324 1245 325 1275
rect 325 1245 355 1275
rect 355 1245 356 1275
rect 324 1244 356 1245
rect 324 1195 356 1196
rect 324 1165 325 1195
rect 325 1165 355 1195
rect 355 1165 356 1195
rect 324 1164 356 1165
rect 324 1084 356 1116
rect 324 1035 356 1036
rect 324 1005 325 1035
rect 325 1005 355 1035
rect 355 1005 356 1035
rect 324 1004 356 1005
rect 324 955 356 956
rect 324 925 325 955
rect 325 925 355 955
rect 355 925 356 955
rect 324 924 356 925
rect 404 1675 436 1676
rect 404 1645 405 1675
rect 405 1645 435 1675
rect 435 1645 436 1675
rect 404 1644 436 1645
rect 404 1595 436 1596
rect 404 1565 405 1595
rect 405 1565 435 1595
rect 435 1565 436 1595
rect 404 1564 436 1565
rect 404 1484 436 1516
rect 404 1435 436 1436
rect 404 1405 405 1435
rect 405 1405 435 1435
rect 435 1405 436 1435
rect 404 1404 436 1405
rect 404 1355 436 1356
rect 404 1325 405 1355
rect 405 1325 435 1355
rect 435 1325 436 1355
rect 404 1324 436 1325
rect 404 1275 436 1276
rect 404 1245 405 1275
rect 405 1245 435 1275
rect 435 1245 436 1275
rect 404 1244 436 1245
rect 404 1195 436 1196
rect 404 1165 405 1195
rect 405 1165 435 1195
rect 435 1165 436 1195
rect 404 1164 436 1165
rect 404 1084 436 1116
rect 404 1035 436 1036
rect 404 1005 405 1035
rect 405 1005 435 1035
rect 435 1005 436 1035
rect 404 1004 436 1005
rect 404 955 436 956
rect 404 925 405 955
rect 405 925 435 955
rect 435 925 436 955
rect 404 924 436 925
rect 484 1675 516 1676
rect 484 1645 485 1675
rect 485 1645 515 1675
rect 515 1645 516 1675
rect 484 1644 516 1645
rect 484 1595 516 1596
rect 484 1565 485 1595
rect 485 1565 515 1595
rect 515 1565 516 1595
rect 484 1564 516 1565
rect 484 1484 516 1516
rect 484 1435 516 1436
rect 484 1405 485 1435
rect 485 1405 515 1435
rect 515 1405 516 1435
rect 484 1404 516 1405
rect 484 1355 516 1356
rect 484 1325 485 1355
rect 485 1325 515 1355
rect 515 1325 516 1355
rect 484 1324 516 1325
rect 484 1275 516 1276
rect 484 1245 485 1275
rect 485 1245 515 1275
rect 515 1245 516 1275
rect 484 1244 516 1245
rect 484 1195 516 1196
rect 484 1165 485 1195
rect 485 1165 515 1195
rect 515 1165 516 1195
rect 484 1164 516 1165
rect 484 1084 516 1116
rect 484 1035 516 1036
rect 484 1005 485 1035
rect 485 1005 515 1035
rect 515 1005 516 1035
rect 484 1004 516 1005
rect 484 955 516 956
rect 484 925 485 955
rect 485 925 515 955
rect 515 925 516 955
rect 484 924 516 925
rect 564 1675 596 1676
rect 564 1645 565 1675
rect 565 1645 595 1675
rect 595 1645 596 1675
rect 564 1644 596 1645
rect 564 1595 596 1596
rect 564 1565 565 1595
rect 565 1565 595 1595
rect 595 1565 596 1595
rect 564 1564 596 1565
rect 564 1484 596 1516
rect 564 1435 596 1436
rect 564 1405 565 1435
rect 565 1405 595 1435
rect 595 1405 596 1435
rect 564 1404 596 1405
rect 564 1355 596 1356
rect 564 1325 565 1355
rect 565 1325 595 1355
rect 595 1325 596 1355
rect 564 1324 596 1325
rect 564 1275 596 1276
rect 564 1245 565 1275
rect 565 1245 595 1275
rect 595 1245 596 1275
rect 564 1244 596 1245
rect 564 1195 596 1196
rect 564 1165 565 1195
rect 565 1165 595 1195
rect 595 1165 596 1195
rect 564 1164 596 1165
rect 564 1084 596 1116
rect 564 1035 596 1036
rect 564 1005 565 1035
rect 565 1005 595 1035
rect 595 1005 596 1035
rect 564 1004 596 1005
rect 564 955 596 956
rect 564 925 565 955
rect 565 925 595 955
rect 595 925 596 955
rect 564 924 596 925
rect 644 1675 676 1676
rect 644 1645 645 1675
rect 645 1645 675 1675
rect 675 1645 676 1675
rect 644 1644 676 1645
rect 644 1595 676 1596
rect 644 1565 645 1595
rect 645 1565 675 1595
rect 675 1565 676 1595
rect 644 1564 676 1565
rect 644 1484 676 1516
rect 644 1435 676 1436
rect 644 1405 645 1435
rect 645 1405 675 1435
rect 675 1405 676 1435
rect 644 1404 676 1405
rect 644 1355 676 1356
rect 644 1325 645 1355
rect 645 1325 675 1355
rect 675 1325 676 1355
rect 644 1324 676 1325
rect 644 1275 676 1276
rect 644 1245 645 1275
rect 645 1245 675 1275
rect 675 1245 676 1275
rect 644 1244 676 1245
rect 644 1195 676 1196
rect 644 1165 645 1195
rect 645 1165 675 1195
rect 675 1165 676 1195
rect 644 1164 676 1165
rect 644 1084 676 1116
rect 644 1035 676 1036
rect 644 1005 645 1035
rect 645 1005 675 1035
rect 675 1005 676 1035
rect 644 1004 676 1005
rect 644 955 676 956
rect 644 925 645 955
rect 645 925 675 955
rect 675 925 676 955
rect 644 924 676 925
rect 724 1675 756 1676
rect 724 1645 725 1675
rect 725 1645 755 1675
rect 755 1645 756 1675
rect 724 1644 756 1645
rect 724 1595 756 1596
rect 724 1565 725 1595
rect 725 1565 755 1595
rect 755 1565 756 1595
rect 724 1564 756 1565
rect 724 1484 756 1516
rect 724 1435 756 1436
rect 724 1405 725 1435
rect 725 1405 755 1435
rect 755 1405 756 1435
rect 724 1404 756 1405
rect 724 1355 756 1356
rect 724 1325 725 1355
rect 725 1325 755 1355
rect 755 1325 756 1355
rect 724 1324 756 1325
rect 724 1275 756 1276
rect 724 1245 725 1275
rect 725 1245 755 1275
rect 755 1245 756 1275
rect 724 1244 756 1245
rect 724 1195 756 1196
rect 724 1165 725 1195
rect 725 1165 755 1195
rect 755 1165 756 1195
rect 724 1164 756 1165
rect 724 1084 756 1116
rect 724 1035 756 1036
rect 724 1005 725 1035
rect 725 1005 755 1035
rect 755 1005 756 1035
rect 724 1004 756 1005
rect 724 955 756 956
rect 724 925 725 955
rect 725 925 755 955
rect 755 925 756 955
rect 724 924 756 925
rect 804 1675 836 1676
rect 804 1645 805 1675
rect 805 1645 835 1675
rect 835 1645 836 1675
rect 804 1644 836 1645
rect 804 1595 836 1596
rect 804 1565 805 1595
rect 805 1565 835 1595
rect 835 1565 836 1595
rect 804 1564 836 1565
rect 804 1484 836 1516
rect 804 1435 836 1436
rect 804 1405 805 1435
rect 805 1405 835 1435
rect 835 1405 836 1435
rect 804 1404 836 1405
rect 804 1355 836 1356
rect 804 1325 805 1355
rect 805 1325 835 1355
rect 835 1325 836 1355
rect 804 1324 836 1325
rect 804 1275 836 1276
rect 804 1245 805 1275
rect 805 1245 835 1275
rect 835 1245 836 1275
rect 804 1244 836 1245
rect 804 1195 836 1196
rect 804 1165 805 1195
rect 805 1165 835 1195
rect 835 1165 836 1195
rect 804 1164 836 1165
rect 804 1084 836 1116
rect 804 1035 836 1036
rect 804 1005 805 1035
rect 805 1005 835 1035
rect 835 1005 836 1035
rect 804 1004 836 1005
rect 804 955 836 956
rect 804 925 805 955
rect 805 925 835 955
rect 835 925 836 955
rect 804 924 836 925
rect 884 1675 916 1676
rect 884 1645 885 1675
rect 885 1645 915 1675
rect 915 1645 916 1675
rect 884 1644 916 1645
rect 884 1595 916 1596
rect 884 1565 885 1595
rect 885 1565 915 1595
rect 915 1565 916 1595
rect 884 1564 916 1565
rect 884 1484 916 1516
rect 884 1435 916 1436
rect 884 1405 885 1435
rect 885 1405 915 1435
rect 915 1405 916 1435
rect 884 1404 916 1405
rect 884 1355 916 1356
rect 884 1325 885 1355
rect 885 1325 915 1355
rect 915 1325 916 1355
rect 884 1324 916 1325
rect 884 1275 916 1276
rect 884 1245 885 1275
rect 885 1245 915 1275
rect 915 1245 916 1275
rect 884 1244 916 1245
rect 884 1195 916 1196
rect 884 1165 885 1195
rect 885 1165 915 1195
rect 915 1165 916 1195
rect 884 1164 916 1165
rect 884 1084 916 1116
rect 884 1035 916 1036
rect 884 1005 885 1035
rect 885 1005 915 1035
rect 915 1005 916 1035
rect 884 1004 916 1005
rect 884 955 916 956
rect 884 925 885 955
rect 885 925 915 955
rect 915 925 916 955
rect 884 924 916 925
rect 964 1675 996 1676
rect 964 1645 965 1675
rect 965 1645 995 1675
rect 995 1645 996 1675
rect 964 1644 996 1645
rect 964 1595 996 1596
rect 964 1565 965 1595
rect 965 1565 995 1595
rect 995 1565 996 1595
rect 964 1564 996 1565
rect 964 1484 996 1516
rect 964 1435 996 1436
rect 964 1405 965 1435
rect 965 1405 995 1435
rect 995 1405 996 1435
rect 964 1404 996 1405
rect 964 1355 996 1356
rect 964 1325 965 1355
rect 965 1325 995 1355
rect 995 1325 996 1355
rect 964 1324 996 1325
rect 964 1275 996 1276
rect 964 1245 965 1275
rect 965 1245 995 1275
rect 995 1245 996 1275
rect 964 1244 996 1245
rect 964 1195 996 1196
rect 964 1165 965 1195
rect 965 1165 995 1195
rect 995 1165 996 1195
rect 964 1164 996 1165
rect 964 1084 996 1116
rect 964 1035 996 1036
rect 964 1005 965 1035
rect 965 1005 995 1035
rect 995 1005 996 1035
rect 964 1004 996 1005
rect 964 955 996 956
rect 964 925 965 955
rect 965 925 995 955
rect 995 925 996 955
rect 964 924 996 925
rect 1044 1675 1076 1676
rect 1044 1645 1045 1675
rect 1045 1645 1075 1675
rect 1075 1645 1076 1675
rect 1044 1644 1076 1645
rect 1044 1595 1076 1596
rect 1044 1565 1045 1595
rect 1045 1565 1075 1595
rect 1075 1565 1076 1595
rect 1044 1564 1076 1565
rect 1044 1484 1076 1516
rect 1044 1435 1076 1436
rect 1044 1405 1045 1435
rect 1045 1405 1075 1435
rect 1075 1405 1076 1435
rect 1044 1404 1076 1405
rect 1044 1355 1076 1356
rect 1044 1325 1045 1355
rect 1045 1325 1075 1355
rect 1075 1325 1076 1355
rect 1044 1324 1076 1325
rect 1044 1275 1076 1276
rect 1044 1245 1045 1275
rect 1045 1245 1075 1275
rect 1075 1245 1076 1275
rect 1044 1244 1076 1245
rect 1044 1195 1076 1196
rect 1044 1165 1045 1195
rect 1045 1165 1075 1195
rect 1075 1165 1076 1195
rect 1044 1164 1076 1165
rect 1044 1084 1076 1116
rect 1044 1035 1076 1036
rect 1044 1005 1045 1035
rect 1045 1005 1075 1035
rect 1075 1005 1076 1035
rect 1044 1004 1076 1005
rect 1044 955 1076 956
rect 1044 925 1045 955
rect 1045 925 1075 955
rect 1075 925 1076 955
rect 1044 924 1076 925
rect 1124 1675 1156 1676
rect 1124 1645 1125 1675
rect 1125 1645 1155 1675
rect 1155 1645 1156 1675
rect 1124 1644 1156 1645
rect 1124 1595 1156 1596
rect 1124 1565 1125 1595
rect 1125 1565 1155 1595
rect 1155 1565 1156 1595
rect 1124 1564 1156 1565
rect 1124 1484 1156 1516
rect 1124 1435 1156 1436
rect 1124 1405 1125 1435
rect 1125 1405 1155 1435
rect 1155 1405 1156 1435
rect 1124 1404 1156 1405
rect 1124 1355 1156 1356
rect 1124 1325 1125 1355
rect 1125 1325 1155 1355
rect 1155 1325 1156 1355
rect 1124 1324 1156 1325
rect 1124 1275 1156 1276
rect 1124 1245 1125 1275
rect 1125 1245 1155 1275
rect 1155 1245 1156 1275
rect 1124 1244 1156 1245
rect 1124 1195 1156 1196
rect 1124 1165 1125 1195
rect 1125 1165 1155 1195
rect 1155 1165 1156 1195
rect 1124 1164 1156 1165
rect 1124 1084 1156 1116
rect 1124 1035 1156 1036
rect 1124 1005 1125 1035
rect 1125 1005 1155 1035
rect 1155 1005 1156 1035
rect 1124 1004 1156 1005
rect 1124 955 1156 956
rect 1124 925 1125 955
rect 1125 925 1155 955
rect 1155 925 1156 955
rect 1124 924 1156 925
rect 1204 1675 1236 1676
rect 1204 1645 1205 1675
rect 1205 1645 1235 1675
rect 1235 1645 1236 1675
rect 1204 1644 1236 1645
rect 1204 1595 1236 1596
rect 1204 1565 1205 1595
rect 1205 1565 1235 1595
rect 1235 1565 1236 1595
rect 1204 1564 1236 1565
rect 1204 1484 1236 1516
rect 1204 1435 1236 1436
rect 1204 1405 1205 1435
rect 1205 1405 1235 1435
rect 1235 1405 1236 1435
rect 1204 1404 1236 1405
rect 1204 1355 1236 1356
rect 1204 1325 1205 1355
rect 1205 1325 1235 1355
rect 1235 1325 1236 1355
rect 1204 1324 1236 1325
rect 1204 1275 1236 1276
rect 1204 1245 1205 1275
rect 1205 1245 1235 1275
rect 1235 1245 1236 1275
rect 1204 1244 1236 1245
rect 1204 1195 1236 1196
rect 1204 1165 1205 1195
rect 1205 1165 1235 1195
rect 1235 1165 1236 1195
rect 1204 1164 1236 1165
rect 1204 1084 1236 1116
rect 1204 1035 1236 1036
rect 1204 1005 1205 1035
rect 1205 1005 1235 1035
rect 1235 1005 1236 1035
rect 1204 1004 1236 1005
rect 1204 955 1236 956
rect 1204 925 1205 955
rect 1205 925 1235 955
rect 1235 925 1236 955
rect 1204 924 1236 925
rect 1284 1675 1316 1676
rect 1284 1645 1285 1675
rect 1285 1645 1315 1675
rect 1315 1645 1316 1675
rect 1284 1644 1316 1645
rect 1284 1595 1316 1596
rect 1284 1565 1285 1595
rect 1285 1565 1315 1595
rect 1315 1565 1316 1595
rect 1284 1564 1316 1565
rect 1284 1484 1316 1516
rect 1284 1435 1316 1436
rect 1284 1405 1285 1435
rect 1285 1405 1315 1435
rect 1315 1405 1316 1435
rect 1284 1404 1316 1405
rect 1284 1355 1316 1356
rect 1284 1325 1285 1355
rect 1285 1325 1315 1355
rect 1315 1325 1316 1355
rect 1284 1324 1316 1325
rect 1284 1275 1316 1276
rect 1284 1245 1285 1275
rect 1285 1245 1315 1275
rect 1315 1245 1316 1275
rect 1284 1244 1316 1245
rect 1284 1195 1316 1196
rect 1284 1165 1285 1195
rect 1285 1165 1315 1195
rect 1315 1165 1316 1195
rect 1284 1164 1316 1165
rect 1284 1084 1316 1116
rect 1284 1035 1316 1036
rect 1284 1005 1285 1035
rect 1285 1005 1315 1035
rect 1315 1005 1316 1035
rect 1284 1004 1316 1005
rect 1284 955 1316 956
rect 1284 925 1285 955
rect 1285 925 1315 955
rect 1315 925 1316 955
rect 1284 924 1316 925
rect 1364 1675 1396 1676
rect 1364 1645 1365 1675
rect 1365 1645 1395 1675
rect 1395 1645 1396 1675
rect 1364 1644 1396 1645
rect 1364 1595 1396 1596
rect 1364 1565 1365 1595
rect 1365 1565 1395 1595
rect 1395 1565 1396 1595
rect 1364 1564 1396 1565
rect 1364 1484 1396 1516
rect 1364 1435 1396 1436
rect 1364 1405 1365 1435
rect 1365 1405 1395 1435
rect 1395 1405 1396 1435
rect 1364 1404 1396 1405
rect 1364 1355 1396 1356
rect 1364 1325 1365 1355
rect 1365 1325 1395 1355
rect 1395 1325 1396 1355
rect 1364 1324 1396 1325
rect 1364 1275 1396 1276
rect 1364 1245 1365 1275
rect 1365 1245 1395 1275
rect 1395 1245 1396 1275
rect 1364 1244 1396 1245
rect 1364 1195 1396 1196
rect 1364 1165 1365 1195
rect 1365 1165 1395 1195
rect 1395 1165 1396 1195
rect 1364 1164 1396 1165
rect 1364 1084 1396 1116
rect 1364 1035 1396 1036
rect 1364 1005 1365 1035
rect 1365 1005 1395 1035
rect 1395 1005 1396 1035
rect 1364 1004 1396 1005
rect 1364 955 1396 956
rect 1364 925 1365 955
rect 1365 925 1395 955
rect 1395 925 1396 955
rect 1364 924 1396 925
rect 1444 1675 1476 1676
rect 1444 1645 1445 1675
rect 1445 1645 1475 1675
rect 1475 1645 1476 1675
rect 1444 1644 1476 1645
rect 1444 1595 1476 1596
rect 1444 1565 1445 1595
rect 1445 1565 1475 1595
rect 1475 1565 1476 1595
rect 1444 1564 1476 1565
rect 1444 1484 1476 1516
rect 1444 1435 1476 1436
rect 1444 1405 1445 1435
rect 1445 1405 1475 1435
rect 1475 1405 1476 1435
rect 1444 1404 1476 1405
rect 1444 1355 1476 1356
rect 1444 1325 1445 1355
rect 1445 1325 1475 1355
rect 1475 1325 1476 1355
rect 1444 1324 1476 1325
rect 1444 1275 1476 1276
rect 1444 1245 1445 1275
rect 1445 1245 1475 1275
rect 1475 1245 1476 1275
rect 1444 1244 1476 1245
rect 1444 1195 1476 1196
rect 1444 1165 1445 1195
rect 1445 1165 1475 1195
rect 1475 1165 1476 1195
rect 1444 1164 1476 1165
rect 1444 1084 1476 1116
rect 1444 1035 1476 1036
rect 1444 1005 1445 1035
rect 1445 1005 1475 1035
rect 1475 1005 1476 1035
rect 1444 1004 1476 1005
rect 1444 955 1476 956
rect 1444 925 1445 955
rect 1445 925 1475 955
rect 1475 925 1476 955
rect 1444 924 1476 925
rect 1524 1675 1556 1676
rect 1524 1645 1525 1675
rect 1525 1645 1555 1675
rect 1555 1645 1556 1675
rect 1524 1644 1556 1645
rect 1524 1595 1556 1596
rect 1524 1565 1525 1595
rect 1525 1565 1555 1595
rect 1555 1565 1556 1595
rect 1524 1564 1556 1565
rect 1524 1484 1556 1516
rect 1524 1435 1556 1436
rect 1524 1405 1525 1435
rect 1525 1405 1555 1435
rect 1555 1405 1556 1435
rect 1524 1404 1556 1405
rect 1524 1355 1556 1356
rect 1524 1325 1525 1355
rect 1525 1325 1555 1355
rect 1555 1325 1556 1355
rect 1524 1324 1556 1325
rect 1524 1275 1556 1276
rect 1524 1245 1525 1275
rect 1525 1245 1555 1275
rect 1555 1245 1556 1275
rect 1524 1244 1556 1245
rect 1524 1195 1556 1196
rect 1524 1165 1525 1195
rect 1525 1165 1555 1195
rect 1555 1165 1556 1195
rect 1524 1164 1556 1165
rect 1524 1084 1556 1116
rect 1524 1035 1556 1036
rect 1524 1005 1525 1035
rect 1525 1005 1555 1035
rect 1555 1005 1556 1035
rect 1524 1004 1556 1005
rect 1524 955 1556 956
rect 1524 925 1525 955
rect 1525 925 1555 955
rect 1555 925 1556 955
rect 1524 924 1556 925
rect 1604 1675 1636 1676
rect 1604 1645 1605 1675
rect 1605 1645 1635 1675
rect 1635 1645 1636 1675
rect 1604 1644 1636 1645
rect 1604 1595 1636 1596
rect 1604 1565 1605 1595
rect 1605 1565 1635 1595
rect 1635 1565 1636 1595
rect 1604 1564 1636 1565
rect 1604 1484 1636 1516
rect 1604 1435 1636 1436
rect 1604 1405 1605 1435
rect 1605 1405 1635 1435
rect 1635 1405 1636 1435
rect 1604 1404 1636 1405
rect 1604 1355 1636 1356
rect 1604 1325 1605 1355
rect 1605 1325 1635 1355
rect 1635 1325 1636 1355
rect 1604 1324 1636 1325
rect 1604 1275 1636 1276
rect 1604 1245 1605 1275
rect 1605 1245 1635 1275
rect 1635 1245 1636 1275
rect 1604 1244 1636 1245
rect 1604 1195 1636 1196
rect 1604 1165 1605 1195
rect 1605 1165 1635 1195
rect 1635 1165 1636 1195
rect 1604 1164 1636 1165
rect 1604 1084 1636 1116
rect 1604 1035 1636 1036
rect 1604 1005 1605 1035
rect 1605 1005 1635 1035
rect 1635 1005 1636 1035
rect 1604 1004 1636 1005
rect 1604 955 1636 956
rect 1604 925 1605 955
rect 1605 925 1635 955
rect 1635 925 1636 955
rect 1604 924 1636 925
rect 1684 1675 1716 1676
rect 1684 1645 1685 1675
rect 1685 1645 1715 1675
rect 1715 1645 1716 1675
rect 1684 1644 1716 1645
rect 1684 1595 1716 1596
rect 1684 1565 1685 1595
rect 1685 1565 1715 1595
rect 1715 1565 1716 1595
rect 1684 1564 1716 1565
rect 1684 1484 1716 1516
rect 1684 1435 1716 1436
rect 1684 1405 1685 1435
rect 1685 1405 1715 1435
rect 1715 1405 1716 1435
rect 1684 1404 1716 1405
rect 1684 1355 1716 1356
rect 1684 1325 1685 1355
rect 1685 1325 1715 1355
rect 1715 1325 1716 1355
rect 1684 1324 1716 1325
rect 1684 1275 1716 1276
rect 1684 1245 1685 1275
rect 1685 1245 1715 1275
rect 1715 1245 1716 1275
rect 1684 1244 1716 1245
rect 1684 1195 1716 1196
rect 1684 1165 1685 1195
rect 1685 1165 1715 1195
rect 1715 1165 1716 1195
rect 1684 1164 1716 1165
rect 1684 1084 1716 1116
rect 1684 1035 1716 1036
rect 1684 1005 1685 1035
rect 1685 1005 1715 1035
rect 1715 1005 1716 1035
rect 1684 1004 1716 1005
rect 1684 955 1716 956
rect 1684 925 1685 955
rect 1685 925 1715 955
rect 1715 925 1716 955
rect 1684 924 1716 925
rect 1764 1675 1796 1676
rect 1764 1645 1765 1675
rect 1765 1645 1795 1675
rect 1795 1645 1796 1675
rect 1764 1644 1796 1645
rect 1764 1595 1796 1596
rect 1764 1565 1765 1595
rect 1765 1565 1795 1595
rect 1795 1565 1796 1595
rect 1764 1564 1796 1565
rect 1764 1484 1796 1516
rect 1764 1435 1796 1436
rect 1764 1405 1765 1435
rect 1765 1405 1795 1435
rect 1795 1405 1796 1435
rect 1764 1404 1796 1405
rect 1764 1355 1796 1356
rect 1764 1325 1765 1355
rect 1765 1325 1795 1355
rect 1795 1325 1796 1355
rect 1764 1324 1796 1325
rect 1764 1275 1796 1276
rect 1764 1245 1765 1275
rect 1765 1245 1795 1275
rect 1795 1245 1796 1275
rect 1764 1244 1796 1245
rect 1764 1195 1796 1196
rect 1764 1165 1765 1195
rect 1765 1165 1795 1195
rect 1795 1165 1796 1195
rect 1764 1164 1796 1165
rect 1764 1084 1796 1116
rect 1764 1035 1796 1036
rect 1764 1005 1765 1035
rect 1765 1005 1795 1035
rect 1795 1005 1796 1035
rect 1764 1004 1796 1005
rect 1764 955 1796 956
rect 1764 925 1765 955
rect 1765 925 1795 955
rect 1795 925 1796 955
rect 1764 924 1796 925
rect 1844 1675 1876 1676
rect 1844 1645 1845 1675
rect 1845 1645 1875 1675
rect 1875 1645 1876 1675
rect 1844 1644 1876 1645
rect 1844 1595 1876 1596
rect 1844 1565 1845 1595
rect 1845 1565 1875 1595
rect 1875 1565 1876 1595
rect 1844 1564 1876 1565
rect 1844 1484 1876 1516
rect 1844 1435 1876 1436
rect 1844 1405 1845 1435
rect 1845 1405 1875 1435
rect 1875 1405 1876 1435
rect 1844 1404 1876 1405
rect 1844 1355 1876 1356
rect 1844 1325 1845 1355
rect 1845 1325 1875 1355
rect 1875 1325 1876 1355
rect 1844 1324 1876 1325
rect 1844 1275 1876 1276
rect 1844 1245 1845 1275
rect 1845 1245 1875 1275
rect 1875 1245 1876 1275
rect 1844 1244 1876 1245
rect 1844 1195 1876 1196
rect 1844 1165 1845 1195
rect 1845 1165 1875 1195
rect 1875 1165 1876 1195
rect 1844 1164 1876 1165
rect 1844 1084 1876 1116
rect 1844 1035 1876 1036
rect 1844 1005 1845 1035
rect 1845 1005 1875 1035
rect 1875 1005 1876 1035
rect 1844 1004 1876 1005
rect 1844 955 1876 956
rect 1844 925 1845 955
rect 1845 925 1875 955
rect 1875 925 1876 955
rect 1844 924 1876 925
rect 1924 1675 1956 1676
rect 1924 1645 1925 1675
rect 1925 1645 1955 1675
rect 1955 1645 1956 1675
rect 1924 1644 1956 1645
rect 1924 1595 1956 1596
rect 1924 1565 1925 1595
rect 1925 1565 1955 1595
rect 1955 1565 1956 1595
rect 1924 1564 1956 1565
rect 1924 1484 1956 1516
rect 1924 1435 1956 1436
rect 1924 1405 1925 1435
rect 1925 1405 1955 1435
rect 1955 1405 1956 1435
rect 1924 1404 1956 1405
rect 1924 1355 1956 1356
rect 1924 1325 1925 1355
rect 1925 1325 1955 1355
rect 1955 1325 1956 1355
rect 1924 1324 1956 1325
rect 1924 1275 1956 1276
rect 1924 1245 1925 1275
rect 1925 1245 1955 1275
rect 1955 1245 1956 1275
rect 1924 1244 1956 1245
rect 1924 1195 1956 1196
rect 1924 1165 1925 1195
rect 1925 1165 1955 1195
rect 1955 1165 1956 1195
rect 1924 1164 1956 1165
rect 1924 1084 1956 1116
rect 1924 1035 1956 1036
rect 1924 1005 1925 1035
rect 1925 1005 1955 1035
rect 1955 1005 1956 1035
rect 1924 1004 1956 1005
rect 1924 955 1956 956
rect 1924 925 1925 955
rect 1925 925 1955 955
rect 1955 925 1956 955
rect 1924 924 1956 925
rect 2004 1675 2036 1676
rect 2004 1645 2005 1675
rect 2005 1645 2035 1675
rect 2035 1645 2036 1675
rect 2004 1644 2036 1645
rect 2004 1595 2036 1596
rect 2004 1565 2005 1595
rect 2005 1565 2035 1595
rect 2035 1565 2036 1595
rect 2004 1564 2036 1565
rect 2004 1484 2036 1516
rect 2004 1435 2036 1436
rect 2004 1405 2005 1435
rect 2005 1405 2035 1435
rect 2035 1405 2036 1435
rect 2004 1404 2036 1405
rect 2004 1355 2036 1356
rect 2004 1325 2005 1355
rect 2005 1325 2035 1355
rect 2035 1325 2036 1355
rect 2004 1324 2036 1325
rect 2004 1275 2036 1276
rect 2004 1245 2005 1275
rect 2005 1245 2035 1275
rect 2035 1245 2036 1275
rect 2004 1244 2036 1245
rect 2004 1195 2036 1196
rect 2004 1165 2005 1195
rect 2005 1165 2035 1195
rect 2035 1165 2036 1195
rect 2004 1164 2036 1165
rect 2004 1084 2036 1116
rect 2004 1035 2036 1036
rect 2004 1005 2005 1035
rect 2005 1005 2035 1035
rect 2035 1005 2036 1035
rect 2004 1004 2036 1005
rect 2004 955 2036 956
rect 2004 925 2005 955
rect 2005 925 2035 955
rect 2035 925 2036 955
rect 2004 924 2036 925
rect 2084 1675 2116 1676
rect 2084 1645 2085 1675
rect 2085 1645 2115 1675
rect 2115 1645 2116 1675
rect 2084 1644 2116 1645
rect 2084 1595 2116 1596
rect 2084 1565 2085 1595
rect 2085 1565 2115 1595
rect 2115 1565 2116 1595
rect 2084 1564 2116 1565
rect 2084 1484 2116 1516
rect 2084 1435 2116 1436
rect 2084 1405 2085 1435
rect 2085 1405 2115 1435
rect 2115 1405 2116 1435
rect 2084 1404 2116 1405
rect 2084 1355 2116 1356
rect 2084 1325 2085 1355
rect 2085 1325 2115 1355
rect 2115 1325 2116 1355
rect 2084 1324 2116 1325
rect 2084 1275 2116 1276
rect 2084 1245 2085 1275
rect 2085 1245 2115 1275
rect 2115 1245 2116 1275
rect 2084 1244 2116 1245
rect 2084 1195 2116 1196
rect 2084 1165 2085 1195
rect 2085 1165 2115 1195
rect 2115 1165 2116 1195
rect 2084 1164 2116 1165
rect 2084 1084 2116 1116
rect 2084 1035 2116 1036
rect 2084 1005 2085 1035
rect 2085 1005 2115 1035
rect 2115 1005 2116 1035
rect 2084 1004 2116 1005
rect 2084 955 2116 956
rect 2084 925 2085 955
rect 2085 925 2115 955
rect 2115 925 2116 955
rect 2084 924 2116 925
rect 2164 1675 2196 1676
rect 2164 1645 2165 1675
rect 2165 1645 2195 1675
rect 2195 1645 2196 1675
rect 2164 1644 2196 1645
rect 2164 1595 2196 1596
rect 2164 1565 2165 1595
rect 2165 1565 2195 1595
rect 2195 1565 2196 1595
rect 2164 1564 2196 1565
rect 2164 1484 2196 1516
rect 2164 1435 2196 1436
rect 2164 1405 2165 1435
rect 2165 1405 2195 1435
rect 2195 1405 2196 1435
rect 2164 1404 2196 1405
rect 2164 1355 2196 1356
rect 2164 1325 2165 1355
rect 2165 1325 2195 1355
rect 2195 1325 2196 1355
rect 2164 1324 2196 1325
rect 2164 1275 2196 1276
rect 2164 1245 2165 1275
rect 2165 1245 2195 1275
rect 2195 1245 2196 1275
rect 2164 1244 2196 1245
rect 2164 1195 2196 1196
rect 2164 1165 2165 1195
rect 2165 1165 2195 1195
rect 2195 1165 2196 1195
rect 2164 1164 2196 1165
rect 2164 1084 2196 1116
rect 2164 1035 2196 1036
rect 2164 1005 2165 1035
rect 2165 1005 2195 1035
rect 2195 1005 2196 1035
rect 2164 1004 2196 1005
rect 2164 955 2196 956
rect 2164 925 2165 955
rect 2165 925 2195 955
rect 2195 925 2196 955
rect 2164 924 2196 925
rect 2244 1675 2276 1676
rect 2244 1645 2245 1675
rect 2245 1645 2275 1675
rect 2275 1645 2276 1675
rect 2244 1644 2276 1645
rect 2244 1595 2276 1596
rect 2244 1565 2245 1595
rect 2245 1565 2275 1595
rect 2275 1565 2276 1595
rect 2244 1564 2276 1565
rect 2244 1484 2276 1516
rect 2244 1435 2276 1436
rect 2244 1405 2245 1435
rect 2245 1405 2275 1435
rect 2275 1405 2276 1435
rect 2244 1404 2276 1405
rect 2244 1355 2276 1356
rect 2244 1325 2245 1355
rect 2245 1325 2275 1355
rect 2275 1325 2276 1355
rect 2244 1324 2276 1325
rect 2244 1275 2276 1276
rect 2244 1245 2245 1275
rect 2245 1245 2275 1275
rect 2275 1245 2276 1275
rect 2244 1244 2276 1245
rect 2244 1195 2276 1196
rect 2244 1165 2245 1195
rect 2245 1165 2275 1195
rect 2275 1165 2276 1195
rect 2244 1164 2276 1165
rect 2244 1084 2276 1116
rect 2244 1035 2276 1036
rect 2244 1005 2245 1035
rect 2245 1005 2275 1035
rect 2275 1005 2276 1035
rect 2244 1004 2276 1005
rect 2244 955 2276 956
rect 2244 925 2245 955
rect 2245 925 2275 955
rect 2275 925 2276 955
rect 2244 924 2276 925
rect 2324 1675 2356 1676
rect 2324 1645 2325 1675
rect 2325 1645 2355 1675
rect 2355 1645 2356 1675
rect 2324 1644 2356 1645
rect 2324 1595 2356 1596
rect 2324 1565 2325 1595
rect 2325 1565 2355 1595
rect 2355 1565 2356 1595
rect 2324 1564 2356 1565
rect 2324 1484 2356 1516
rect 2324 1435 2356 1436
rect 2324 1405 2325 1435
rect 2325 1405 2355 1435
rect 2355 1405 2356 1435
rect 2324 1404 2356 1405
rect 2324 1355 2356 1356
rect 2324 1325 2325 1355
rect 2325 1325 2355 1355
rect 2355 1325 2356 1355
rect 2324 1324 2356 1325
rect 2324 1275 2356 1276
rect 2324 1245 2325 1275
rect 2325 1245 2355 1275
rect 2355 1245 2356 1275
rect 2324 1244 2356 1245
rect 2324 1195 2356 1196
rect 2324 1165 2325 1195
rect 2325 1165 2355 1195
rect 2355 1165 2356 1195
rect 2324 1164 2356 1165
rect 2324 1084 2356 1116
rect 2324 1035 2356 1036
rect 2324 1005 2325 1035
rect 2325 1005 2355 1035
rect 2355 1005 2356 1035
rect 2324 1004 2356 1005
rect 2324 955 2356 956
rect 2324 925 2325 955
rect 2325 925 2355 955
rect 2355 925 2356 955
rect 2324 924 2356 925
rect 2404 1675 2436 1676
rect 2404 1645 2405 1675
rect 2405 1645 2435 1675
rect 2435 1645 2436 1675
rect 2404 1644 2436 1645
rect 2404 1595 2436 1596
rect 2404 1565 2405 1595
rect 2405 1565 2435 1595
rect 2435 1565 2436 1595
rect 2404 1564 2436 1565
rect 2404 1484 2436 1516
rect 2404 1435 2436 1436
rect 2404 1405 2405 1435
rect 2405 1405 2435 1435
rect 2435 1405 2436 1435
rect 2404 1404 2436 1405
rect 2404 1355 2436 1356
rect 2404 1325 2405 1355
rect 2405 1325 2435 1355
rect 2435 1325 2436 1355
rect 2404 1324 2436 1325
rect 2404 1275 2436 1276
rect 2404 1245 2405 1275
rect 2405 1245 2435 1275
rect 2435 1245 2436 1275
rect 2404 1244 2436 1245
rect 2404 1195 2436 1196
rect 2404 1165 2405 1195
rect 2405 1165 2435 1195
rect 2435 1165 2436 1195
rect 2404 1164 2436 1165
rect 2404 1084 2436 1116
rect 2404 1035 2436 1036
rect 2404 1005 2405 1035
rect 2405 1005 2435 1035
rect 2435 1005 2436 1035
rect 2404 1004 2436 1005
rect 2404 955 2436 956
rect 2404 925 2405 955
rect 2405 925 2435 955
rect 2435 925 2436 955
rect 2404 924 2436 925
rect 2484 1675 2516 1676
rect 2484 1645 2485 1675
rect 2485 1645 2515 1675
rect 2515 1645 2516 1675
rect 2484 1644 2516 1645
rect 2484 1595 2516 1596
rect 2484 1565 2485 1595
rect 2485 1565 2515 1595
rect 2515 1565 2516 1595
rect 2484 1564 2516 1565
rect 2484 1484 2516 1516
rect 2484 1435 2516 1436
rect 2484 1405 2485 1435
rect 2485 1405 2515 1435
rect 2515 1405 2516 1435
rect 2484 1404 2516 1405
rect 2484 1355 2516 1356
rect 2484 1325 2485 1355
rect 2485 1325 2515 1355
rect 2515 1325 2516 1355
rect 2484 1324 2516 1325
rect 2484 1275 2516 1276
rect 2484 1245 2485 1275
rect 2485 1245 2515 1275
rect 2515 1245 2516 1275
rect 2484 1244 2516 1245
rect 2484 1195 2516 1196
rect 2484 1165 2485 1195
rect 2485 1165 2515 1195
rect 2515 1165 2516 1195
rect 2484 1164 2516 1165
rect 2484 1084 2516 1116
rect 2484 1035 2516 1036
rect 2484 1005 2485 1035
rect 2485 1005 2515 1035
rect 2515 1005 2516 1035
rect 2484 1004 2516 1005
rect 2484 955 2516 956
rect 2484 925 2485 955
rect 2485 925 2515 955
rect 2515 925 2516 955
rect 2484 924 2516 925
rect 2564 1675 2596 1676
rect 2564 1645 2565 1675
rect 2565 1645 2595 1675
rect 2595 1645 2596 1675
rect 2564 1644 2596 1645
rect 2564 1595 2596 1596
rect 2564 1565 2565 1595
rect 2565 1565 2595 1595
rect 2595 1565 2596 1595
rect 2564 1564 2596 1565
rect 2564 1484 2596 1516
rect 2564 1435 2596 1436
rect 2564 1405 2565 1435
rect 2565 1405 2595 1435
rect 2595 1405 2596 1435
rect 2564 1404 2596 1405
rect 2564 1355 2596 1356
rect 2564 1325 2565 1355
rect 2565 1325 2595 1355
rect 2595 1325 2596 1355
rect 2564 1324 2596 1325
rect 2564 1275 2596 1276
rect 2564 1245 2565 1275
rect 2565 1245 2595 1275
rect 2595 1245 2596 1275
rect 2564 1244 2596 1245
rect 2564 1195 2596 1196
rect 2564 1165 2565 1195
rect 2565 1165 2595 1195
rect 2595 1165 2596 1195
rect 2564 1164 2596 1165
rect 2564 1084 2596 1116
rect 2564 1035 2596 1036
rect 2564 1005 2565 1035
rect 2565 1005 2595 1035
rect 2595 1005 2596 1035
rect 2564 1004 2596 1005
rect 2564 955 2596 956
rect 2564 925 2565 955
rect 2565 925 2595 955
rect 2595 925 2596 955
rect 2564 924 2596 925
rect 2644 1675 2676 1676
rect 2644 1645 2645 1675
rect 2645 1645 2675 1675
rect 2675 1645 2676 1675
rect 2644 1644 2676 1645
rect 2644 1595 2676 1596
rect 2644 1565 2645 1595
rect 2645 1565 2675 1595
rect 2675 1565 2676 1595
rect 2644 1564 2676 1565
rect 2644 1484 2676 1516
rect 2644 1435 2676 1436
rect 2644 1405 2645 1435
rect 2645 1405 2675 1435
rect 2675 1405 2676 1435
rect 2644 1404 2676 1405
rect 2644 1355 2676 1356
rect 2644 1325 2645 1355
rect 2645 1325 2675 1355
rect 2675 1325 2676 1355
rect 2644 1324 2676 1325
rect 2644 1275 2676 1276
rect 2644 1245 2645 1275
rect 2645 1245 2675 1275
rect 2675 1245 2676 1275
rect 2644 1244 2676 1245
rect 2644 1195 2676 1196
rect 2644 1165 2645 1195
rect 2645 1165 2675 1195
rect 2675 1165 2676 1195
rect 2644 1164 2676 1165
rect 2644 1084 2676 1116
rect 2644 1035 2676 1036
rect 2644 1005 2645 1035
rect 2645 1005 2675 1035
rect 2675 1005 2676 1035
rect 2644 1004 2676 1005
rect 2644 955 2676 956
rect 2644 925 2645 955
rect 2645 925 2675 955
rect 2675 925 2676 955
rect 2644 924 2676 925
rect 2724 1675 2756 1676
rect 2724 1645 2725 1675
rect 2725 1645 2755 1675
rect 2755 1645 2756 1675
rect 2724 1644 2756 1645
rect 2724 1595 2756 1596
rect 2724 1565 2725 1595
rect 2725 1565 2755 1595
rect 2755 1565 2756 1595
rect 2724 1564 2756 1565
rect 2724 1484 2756 1516
rect 2724 1435 2756 1436
rect 2724 1405 2725 1435
rect 2725 1405 2755 1435
rect 2755 1405 2756 1435
rect 2724 1404 2756 1405
rect 2724 1355 2756 1356
rect 2724 1325 2725 1355
rect 2725 1325 2755 1355
rect 2755 1325 2756 1355
rect 2724 1324 2756 1325
rect 2724 1275 2756 1276
rect 2724 1245 2725 1275
rect 2725 1245 2755 1275
rect 2755 1245 2756 1275
rect 2724 1244 2756 1245
rect 2724 1195 2756 1196
rect 2724 1165 2725 1195
rect 2725 1165 2755 1195
rect 2755 1165 2756 1195
rect 2724 1164 2756 1165
rect 2724 1084 2756 1116
rect 2724 1035 2756 1036
rect 2724 1005 2725 1035
rect 2725 1005 2755 1035
rect 2755 1005 2756 1035
rect 2724 1004 2756 1005
rect 2724 955 2756 956
rect 2724 925 2725 955
rect 2725 925 2755 955
rect 2755 925 2756 955
rect 2724 924 2756 925
rect 2804 1675 2836 1676
rect 2804 1645 2805 1675
rect 2805 1645 2835 1675
rect 2835 1645 2836 1675
rect 2804 1644 2836 1645
rect 2804 1595 2836 1596
rect 2804 1565 2805 1595
rect 2805 1565 2835 1595
rect 2835 1565 2836 1595
rect 2804 1564 2836 1565
rect 2804 1484 2836 1516
rect 2804 1435 2836 1436
rect 2804 1405 2805 1435
rect 2805 1405 2835 1435
rect 2835 1405 2836 1435
rect 2804 1404 2836 1405
rect 2804 1355 2836 1356
rect 2804 1325 2805 1355
rect 2805 1325 2835 1355
rect 2835 1325 2836 1355
rect 2804 1324 2836 1325
rect 2804 1275 2836 1276
rect 2804 1245 2805 1275
rect 2805 1245 2835 1275
rect 2835 1245 2836 1275
rect 2804 1244 2836 1245
rect 2804 1195 2836 1196
rect 2804 1165 2805 1195
rect 2805 1165 2835 1195
rect 2835 1165 2836 1195
rect 2804 1164 2836 1165
rect 2804 1084 2836 1116
rect 2804 1035 2836 1036
rect 2804 1005 2805 1035
rect 2805 1005 2835 1035
rect 2835 1005 2836 1035
rect 2804 1004 2836 1005
rect 2804 955 2836 956
rect 2804 925 2805 955
rect 2805 925 2835 955
rect 2835 925 2836 955
rect 2804 924 2836 925
rect 2884 1675 2916 1676
rect 2884 1645 2885 1675
rect 2885 1645 2915 1675
rect 2915 1645 2916 1675
rect 2884 1644 2916 1645
rect 2884 1595 2916 1596
rect 2884 1565 2885 1595
rect 2885 1565 2915 1595
rect 2915 1565 2916 1595
rect 2884 1564 2916 1565
rect 2884 1484 2916 1516
rect 2884 1435 2916 1436
rect 2884 1405 2885 1435
rect 2885 1405 2915 1435
rect 2915 1405 2916 1435
rect 2884 1404 2916 1405
rect 2884 1355 2916 1356
rect 2884 1325 2885 1355
rect 2885 1325 2915 1355
rect 2915 1325 2916 1355
rect 2884 1324 2916 1325
rect 2884 1275 2916 1276
rect 2884 1245 2885 1275
rect 2885 1245 2915 1275
rect 2915 1245 2916 1275
rect 2884 1244 2916 1245
rect 2884 1195 2916 1196
rect 2884 1165 2885 1195
rect 2885 1165 2915 1195
rect 2915 1165 2916 1195
rect 2884 1164 2916 1165
rect 2884 1084 2916 1116
rect 2884 1035 2916 1036
rect 2884 1005 2885 1035
rect 2885 1005 2915 1035
rect 2915 1005 2916 1035
rect 2884 1004 2916 1005
rect 2884 955 2916 956
rect 2884 925 2885 955
rect 2885 925 2915 955
rect 2915 925 2916 955
rect 2884 924 2916 925
rect 2964 1675 2996 1676
rect 2964 1645 2965 1675
rect 2965 1645 2995 1675
rect 2995 1645 2996 1675
rect 2964 1644 2996 1645
rect 2964 1595 2996 1596
rect 2964 1565 2965 1595
rect 2965 1565 2995 1595
rect 2995 1565 2996 1595
rect 2964 1564 2996 1565
rect 2964 1484 2996 1516
rect 2964 1435 2996 1436
rect 2964 1405 2965 1435
rect 2965 1405 2995 1435
rect 2995 1405 2996 1435
rect 2964 1404 2996 1405
rect 2964 1355 2996 1356
rect 2964 1325 2965 1355
rect 2965 1325 2995 1355
rect 2995 1325 2996 1355
rect 2964 1324 2996 1325
rect 2964 1275 2996 1276
rect 2964 1245 2965 1275
rect 2965 1245 2995 1275
rect 2995 1245 2996 1275
rect 2964 1244 2996 1245
rect 2964 1195 2996 1196
rect 2964 1165 2965 1195
rect 2965 1165 2995 1195
rect 2995 1165 2996 1195
rect 2964 1164 2996 1165
rect 2964 1084 2996 1116
rect 2964 1035 2996 1036
rect 2964 1005 2965 1035
rect 2965 1005 2995 1035
rect 2995 1005 2996 1035
rect 2964 1004 2996 1005
rect 2964 955 2996 956
rect 2964 925 2965 955
rect 2965 925 2995 955
rect 2995 925 2996 955
rect 2964 924 2996 925
rect 3044 1675 3076 1676
rect 3044 1645 3045 1675
rect 3045 1645 3075 1675
rect 3075 1645 3076 1675
rect 3044 1644 3076 1645
rect 3044 1595 3076 1596
rect 3044 1565 3045 1595
rect 3045 1565 3075 1595
rect 3075 1565 3076 1595
rect 3044 1564 3076 1565
rect 3044 1484 3076 1516
rect 3044 1435 3076 1436
rect 3044 1405 3045 1435
rect 3045 1405 3075 1435
rect 3075 1405 3076 1435
rect 3044 1404 3076 1405
rect 3044 1355 3076 1356
rect 3044 1325 3045 1355
rect 3045 1325 3075 1355
rect 3075 1325 3076 1355
rect 3044 1324 3076 1325
rect 3044 1275 3076 1276
rect 3044 1245 3045 1275
rect 3045 1245 3075 1275
rect 3075 1245 3076 1275
rect 3044 1244 3076 1245
rect 3044 1195 3076 1196
rect 3044 1165 3045 1195
rect 3045 1165 3075 1195
rect 3075 1165 3076 1195
rect 3044 1164 3076 1165
rect 3044 1084 3076 1116
rect 3044 1035 3076 1036
rect 3044 1005 3045 1035
rect 3045 1005 3075 1035
rect 3075 1005 3076 1035
rect 3044 1004 3076 1005
rect 3044 955 3076 956
rect 3044 925 3045 955
rect 3045 925 3075 955
rect 3075 925 3076 955
rect 3044 924 3076 925
rect 3124 1675 3156 1676
rect 3124 1645 3125 1675
rect 3125 1645 3155 1675
rect 3155 1645 3156 1675
rect 3124 1644 3156 1645
rect 3124 1595 3156 1596
rect 3124 1565 3125 1595
rect 3125 1565 3155 1595
rect 3155 1565 3156 1595
rect 3124 1564 3156 1565
rect 3124 1484 3156 1516
rect 3124 1435 3156 1436
rect 3124 1405 3125 1435
rect 3125 1405 3155 1435
rect 3155 1405 3156 1435
rect 3124 1404 3156 1405
rect 3124 1355 3156 1356
rect 3124 1325 3125 1355
rect 3125 1325 3155 1355
rect 3155 1325 3156 1355
rect 3124 1324 3156 1325
rect 3124 1275 3156 1276
rect 3124 1245 3125 1275
rect 3125 1245 3155 1275
rect 3155 1245 3156 1275
rect 3124 1244 3156 1245
rect 3124 1195 3156 1196
rect 3124 1165 3125 1195
rect 3125 1165 3155 1195
rect 3155 1165 3156 1195
rect 3124 1164 3156 1165
rect 3124 1084 3156 1116
rect 3124 1035 3156 1036
rect 3124 1005 3125 1035
rect 3125 1005 3155 1035
rect 3155 1005 3156 1035
rect 3124 1004 3156 1005
rect 3124 955 3156 956
rect 3124 925 3125 955
rect 3125 925 3155 955
rect 3155 925 3156 955
rect 3124 924 3156 925
rect 3204 1675 3236 1676
rect 3204 1645 3205 1675
rect 3205 1645 3235 1675
rect 3235 1645 3236 1675
rect 3204 1644 3236 1645
rect 3204 1595 3236 1596
rect 3204 1565 3205 1595
rect 3205 1565 3235 1595
rect 3235 1565 3236 1595
rect 3204 1564 3236 1565
rect 3204 1484 3236 1516
rect 3204 1435 3236 1436
rect 3204 1405 3205 1435
rect 3205 1405 3235 1435
rect 3235 1405 3236 1435
rect 3204 1404 3236 1405
rect 3204 1355 3236 1356
rect 3204 1325 3205 1355
rect 3205 1325 3235 1355
rect 3235 1325 3236 1355
rect 3204 1324 3236 1325
rect 3204 1275 3236 1276
rect 3204 1245 3205 1275
rect 3205 1245 3235 1275
rect 3235 1245 3236 1275
rect 3204 1244 3236 1245
rect 3204 1195 3236 1196
rect 3204 1165 3205 1195
rect 3205 1165 3235 1195
rect 3235 1165 3236 1195
rect 3204 1164 3236 1165
rect 3204 1084 3236 1116
rect 3204 1035 3236 1036
rect 3204 1005 3205 1035
rect 3205 1005 3235 1035
rect 3235 1005 3236 1035
rect 3204 1004 3236 1005
rect 3204 955 3236 956
rect 3204 925 3205 955
rect 3205 925 3235 955
rect 3235 925 3236 955
rect 3204 924 3236 925
rect 3284 1675 3316 1676
rect 3284 1645 3285 1675
rect 3285 1645 3315 1675
rect 3315 1645 3316 1675
rect 3284 1644 3316 1645
rect 3284 1595 3316 1596
rect 3284 1565 3285 1595
rect 3285 1565 3315 1595
rect 3315 1565 3316 1595
rect 3284 1564 3316 1565
rect 3284 1484 3316 1516
rect 3284 1435 3316 1436
rect 3284 1405 3285 1435
rect 3285 1405 3315 1435
rect 3315 1405 3316 1435
rect 3284 1404 3316 1405
rect 3284 1355 3316 1356
rect 3284 1325 3285 1355
rect 3285 1325 3315 1355
rect 3315 1325 3316 1355
rect 3284 1324 3316 1325
rect 3284 1275 3316 1276
rect 3284 1245 3285 1275
rect 3285 1245 3315 1275
rect 3315 1245 3316 1275
rect 3284 1244 3316 1245
rect 3284 1195 3316 1196
rect 3284 1165 3285 1195
rect 3285 1165 3315 1195
rect 3315 1165 3316 1195
rect 3284 1164 3316 1165
rect 3284 1084 3316 1116
rect 3284 1035 3316 1036
rect 3284 1005 3285 1035
rect 3285 1005 3315 1035
rect 3315 1005 3316 1035
rect 3284 1004 3316 1005
rect 3284 955 3316 956
rect 3284 925 3285 955
rect 3285 925 3315 955
rect 3315 925 3316 955
rect 3284 924 3316 925
rect 3364 1675 3396 1676
rect 3364 1645 3365 1675
rect 3365 1645 3395 1675
rect 3395 1645 3396 1675
rect 3364 1644 3396 1645
rect 3364 1595 3396 1596
rect 3364 1565 3365 1595
rect 3365 1565 3395 1595
rect 3395 1565 3396 1595
rect 3364 1564 3396 1565
rect 3364 1484 3396 1516
rect 3364 1435 3396 1436
rect 3364 1405 3365 1435
rect 3365 1405 3395 1435
rect 3395 1405 3396 1435
rect 3364 1404 3396 1405
rect 3364 1355 3396 1356
rect 3364 1325 3365 1355
rect 3365 1325 3395 1355
rect 3395 1325 3396 1355
rect 3364 1324 3396 1325
rect 3364 1275 3396 1276
rect 3364 1245 3365 1275
rect 3365 1245 3395 1275
rect 3395 1245 3396 1275
rect 3364 1244 3396 1245
rect 3364 1195 3396 1196
rect 3364 1165 3365 1195
rect 3365 1165 3395 1195
rect 3395 1165 3396 1195
rect 3364 1164 3396 1165
rect 3364 1084 3396 1116
rect 3364 1035 3396 1036
rect 3364 1005 3365 1035
rect 3365 1005 3395 1035
rect 3395 1005 3396 1035
rect 3364 1004 3396 1005
rect 3364 955 3396 956
rect 3364 925 3365 955
rect 3365 925 3395 955
rect 3395 925 3396 955
rect 3364 924 3396 925
rect 3444 1675 3476 1676
rect 3444 1645 3445 1675
rect 3445 1645 3475 1675
rect 3475 1645 3476 1675
rect 3444 1644 3476 1645
rect 3444 1595 3476 1596
rect 3444 1565 3445 1595
rect 3445 1565 3475 1595
rect 3475 1565 3476 1595
rect 3444 1564 3476 1565
rect 3444 1484 3476 1516
rect 3444 1435 3476 1436
rect 3444 1405 3445 1435
rect 3445 1405 3475 1435
rect 3475 1405 3476 1435
rect 3444 1404 3476 1405
rect 3444 1355 3476 1356
rect 3444 1325 3445 1355
rect 3445 1325 3475 1355
rect 3475 1325 3476 1355
rect 3444 1324 3476 1325
rect 3444 1275 3476 1276
rect 3444 1245 3445 1275
rect 3445 1245 3475 1275
rect 3475 1245 3476 1275
rect 3444 1244 3476 1245
rect 3444 1195 3476 1196
rect 3444 1165 3445 1195
rect 3445 1165 3475 1195
rect 3475 1165 3476 1195
rect 3444 1164 3476 1165
rect 3444 1084 3476 1116
rect 3444 1035 3476 1036
rect 3444 1005 3445 1035
rect 3445 1005 3475 1035
rect 3475 1005 3476 1035
rect 3444 1004 3476 1005
rect 3444 955 3476 956
rect 3444 925 3445 955
rect 3445 925 3475 955
rect 3475 925 3476 955
rect 3444 924 3476 925
rect 3524 1675 3556 1676
rect 3524 1645 3525 1675
rect 3525 1645 3555 1675
rect 3555 1645 3556 1675
rect 3524 1644 3556 1645
rect 3524 1595 3556 1596
rect 3524 1565 3525 1595
rect 3525 1565 3555 1595
rect 3555 1565 3556 1595
rect 3524 1564 3556 1565
rect 3524 1484 3556 1516
rect 3524 1435 3556 1436
rect 3524 1405 3525 1435
rect 3525 1405 3555 1435
rect 3555 1405 3556 1435
rect 3524 1404 3556 1405
rect 3524 1355 3556 1356
rect 3524 1325 3525 1355
rect 3525 1325 3555 1355
rect 3555 1325 3556 1355
rect 3524 1324 3556 1325
rect 3524 1275 3556 1276
rect 3524 1245 3525 1275
rect 3525 1245 3555 1275
rect 3555 1245 3556 1275
rect 3524 1244 3556 1245
rect 3524 1195 3556 1196
rect 3524 1165 3525 1195
rect 3525 1165 3555 1195
rect 3555 1165 3556 1195
rect 3524 1164 3556 1165
rect 3524 1084 3556 1116
rect 3524 1035 3556 1036
rect 3524 1005 3525 1035
rect 3525 1005 3555 1035
rect 3555 1005 3556 1035
rect 3524 1004 3556 1005
rect 3524 955 3556 956
rect 3524 925 3525 955
rect 3525 925 3555 955
rect 3555 925 3556 955
rect 3524 924 3556 925
rect 3604 1675 3636 1676
rect 3604 1645 3605 1675
rect 3605 1645 3635 1675
rect 3635 1645 3636 1675
rect 3604 1644 3636 1645
rect 3604 1595 3636 1596
rect 3604 1565 3605 1595
rect 3605 1565 3635 1595
rect 3635 1565 3636 1595
rect 3604 1564 3636 1565
rect 3604 1484 3636 1516
rect 3604 1435 3636 1436
rect 3604 1405 3605 1435
rect 3605 1405 3635 1435
rect 3635 1405 3636 1435
rect 3604 1404 3636 1405
rect 3604 1355 3636 1356
rect 3604 1325 3605 1355
rect 3605 1325 3635 1355
rect 3635 1325 3636 1355
rect 3604 1324 3636 1325
rect 3604 1275 3636 1276
rect 3604 1245 3605 1275
rect 3605 1245 3635 1275
rect 3635 1245 3636 1275
rect 3604 1244 3636 1245
rect 3604 1195 3636 1196
rect 3604 1165 3605 1195
rect 3605 1165 3635 1195
rect 3635 1165 3636 1195
rect 3604 1164 3636 1165
rect 3604 1084 3636 1116
rect 3604 1035 3636 1036
rect 3604 1005 3605 1035
rect 3605 1005 3635 1035
rect 3635 1005 3636 1035
rect 3604 1004 3636 1005
rect 3604 955 3636 956
rect 3604 925 3605 955
rect 3605 925 3635 955
rect 3635 925 3636 955
rect 3604 924 3636 925
rect 3684 1675 3716 1676
rect 3684 1645 3685 1675
rect 3685 1645 3715 1675
rect 3715 1645 3716 1675
rect 3684 1644 3716 1645
rect 3684 1595 3716 1596
rect 3684 1565 3685 1595
rect 3685 1565 3715 1595
rect 3715 1565 3716 1595
rect 3684 1564 3716 1565
rect 3684 1484 3716 1516
rect 3684 1435 3716 1436
rect 3684 1405 3685 1435
rect 3685 1405 3715 1435
rect 3715 1405 3716 1435
rect 3684 1404 3716 1405
rect 3684 1355 3716 1356
rect 3684 1325 3685 1355
rect 3685 1325 3715 1355
rect 3715 1325 3716 1355
rect 3684 1324 3716 1325
rect 3684 1275 3716 1276
rect 3684 1245 3685 1275
rect 3685 1245 3715 1275
rect 3715 1245 3716 1275
rect 3684 1244 3716 1245
rect 3684 1195 3716 1196
rect 3684 1165 3685 1195
rect 3685 1165 3715 1195
rect 3715 1165 3716 1195
rect 3684 1164 3716 1165
rect 3684 1084 3716 1116
rect 3684 1035 3716 1036
rect 3684 1005 3685 1035
rect 3685 1005 3715 1035
rect 3715 1005 3716 1035
rect 3684 1004 3716 1005
rect 3684 955 3716 956
rect 3684 925 3685 955
rect 3685 925 3715 955
rect 3715 925 3716 955
rect 3684 924 3716 925
rect 3764 1675 3796 1676
rect 3764 1645 3765 1675
rect 3765 1645 3795 1675
rect 3795 1645 3796 1675
rect 3764 1644 3796 1645
rect 3764 1595 3796 1596
rect 3764 1565 3765 1595
rect 3765 1565 3795 1595
rect 3795 1565 3796 1595
rect 3764 1564 3796 1565
rect 3764 1484 3796 1516
rect 3764 1435 3796 1436
rect 3764 1405 3765 1435
rect 3765 1405 3795 1435
rect 3795 1405 3796 1435
rect 3764 1404 3796 1405
rect 3764 1355 3796 1356
rect 3764 1325 3765 1355
rect 3765 1325 3795 1355
rect 3795 1325 3796 1355
rect 3764 1324 3796 1325
rect 3764 1275 3796 1276
rect 3764 1245 3765 1275
rect 3765 1245 3795 1275
rect 3795 1245 3796 1275
rect 3764 1244 3796 1245
rect 3764 1195 3796 1196
rect 3764 1165 3765 1195
rect 3765 1165 3795 1195
rect 3795 1165 3796 1195
rect 3764 1164 3796 1165
rect 3764 1084 3796 1116
rect 3764 1035 3796 1036
rect 3764 1005 3765 1035
rect 3765 1005 3795 1035
rect 3795 1005 3796 1035
rect 3764 1004 3796 1005
rect 3764 955 3796 956
rect 3764 925 3765 955
rect 3765 925 3795 955
rect 3795 925 3796 955
rect 3764 924 3796 925
rect 3844 1675 3876 1676
rect 3844 1645 3845 1675
rect 3845 1645 3875 1675
rect 3875 1645 3876 1675
rect 3844 1644 3876 1645
rect 3844 1595 3876 1596
rect 3844 1565 3845 1595
rect 3845 1565 3875 1595
rect 3875 1565 3876 1595
rect 3844 1564 3876 1565
rect 3844 1484 3876 1516
rect 3844 1435 3876 1436
rect 3844 1405 3845 1435
rect 3845 1405 3875 1435
rect 3875 1405 3876 1435
rect 3844 1404 3876 1405
rect 3844 1355 3876 1356
rect 3844 1325 3845 1355
rect 3845 1325 3875 1355
rect 3875 1325 3876 1355
rect 3844 1324 3876 1325
rect 3844 1275 3876 1276
rect 3844 1245 3845 1275
rect 3845 1245 3875 1275
rect 3875 1245 3876 1275
rect 3844 1244 3876 1245
rect 3844 1195 3876 1196
rect 3844 1165 3845 1195
rect 3845 1165 3875 1195
rect 3875 1165 3876 1195
rect 3844 1164 3876 1165
rect 3844 1084 3876 1116
rect 3844 1035 3876 1036
rect 3844 1005 3845 1035
rect 3845 1005 3875 1035
rect 3875 1005 3876 1035
rect 3844 1004 3876 1005
rect 3844 955 3876 956
rect 3844 925 3845 955
rect 3845 925 3875 955
rect 3875 925 3876 955
rect 3844 924 3876 925
rect 3924 1675 3956 1676
rect 3924 1645 3925 1675
rect 3925 1645 3955 1675
rect 3955 1645 3956 1675
rect 3924 1644 3956 1645
rect 3924 1595 3956 1596
rect 3924 1565 3925 1595
rect 3925 1565 3955 1595
rect 3955 1565 3956 1595
rect 3924 1564 3956 1565
rect 3924 1484 3956 1516
rect 3924 1435 3956 1436
rect 3924 1405 3925 1435
rect 3925 1405 3955 1435
rect 3955 1405 3956 1435
rect 3924 1404 3956 1405
rect 3924 1355 3956 1356
rect 3924 1325 3925 1355
rect 3925 1325 3955 1355
rect 3955 1325 3956 1355
rect 3924 1324 3956 1325
rect 3924 1275 3956 1276
rect 3924 1245 3925 1275
rect 3925 1245 3955 1275
rect 3955 1245 3956 1275
rect 3924 1244 3956 1245
rect 3924 1195 3956 1196
rect 3924 1165 3925 1195
rect 3925 1165 3955 1195
rect 3955 1165 3956 1195
rect 3924 1164 3956 1165
rect 3924 1084 3956 1116
rect 3924 1035 3956 1036
rect 3924 1005 3925 1035
rect 3925 1005 3955 1035
rect 3955 1005 3956 1035
rect 3924 1004 3956 1005
rect 3924 955 3956 956
rect 3924 925 3925 955
rect 3925 925 3955 955
rect 3955 925 3956 955
rect 3924 924 3956 925
rect 4004 1675 4036 1676
rect 4004 1645 4005 1675
rect 4005 1645 4035 1675
rect 4035 1645 4036 1675
rect 4004 1644 4036 1645
rect 4004 1595 4036 1596
rect 4004 1565 4005 1595
rect 4005 1565 4035 1595
rect 4035 1565 4036 1595
rect 4004 1564 4036 1565
rect 4004 1484 4036 1516
rect 4004 1435 4036 1436
rect 4004 1405 4005 1435
rect 4005 1405 4035 1435
rect 4035 1405 4036 1435
rect 4004 1404 4036 1405
rect 4004 1355 4036 1356
rect 4004 1325 4005 1355
rect 4005 1325 4035 1355
rect 4035 1325 4036 1355
rect 4004 1324 4036 1325
rect 4004 1275 4036 1276
rect 4004 1245 4005 1275
rect 4005 1245 4035 1275
rect 4035 1245 4036 1275
rect 4004 1244 4036 1245
rect 4004 1195 4036 1196
rect 4004 1165 4005 1195
rect 4005 1165 4035 1195
rect 4035 1165 4036 1195
rect 4004 1164 4036 1165
rect 4004 1084 4036 1116
rect 4004 1035 4036 1036
rect 4004 1005 4005 1035
rect 4005 1005 4035 1035
rect 4035 1005 4036 1035
rect 4004 1004 4036 1005
rect 4004 955 4036 956
rect 4004 925 4005 955
rect 4005 925 4035 955
rect 4035 925 4036 955
rect 4004 924 4036 925
rect 4084 1675 4116 1676
rect 4084 1645 4085 1675
rect 4085 1645 4115 1675
rect 4115 1645 4116 1675
rect 4084 1644 4116 1645
rect 4084 1595 4116 1596
rect 4084 1565 4085 1595
rect 4085 1565 4115 1595
rect 4115 1565 4116 1595
rect 4084 1564 4116 1565
rect 4084 1484 4116 1516
rect 4084 1435 4116 1436
rect 4084 1405 4085 1435
rect 4085 1405 4115 1435
rect 4115 1405 4116 1435
rect 4084 1404 4116 1405
rect 4084 1355 4116 1356
rect 4084 1325 4085 1355
rect 4085 1325 4115 1355
rect 4115 1325 4116 1355
rect 4084 1324 4116 1325
rect 4084 1275 4116 1276
rect 4084 1245 4085 1275
rect 4085 1245 4115 1275
rect 4115 1245 4116 1275
rect 4084 1244 4116 1245
rect 4084 1195 4116 1196
rect 4084 1165 4085 1195
rect 4085 1165 4115 1195
rect 4115 1165 4116 1195
rect 4084 1164 4116 1165
rect 4084 1084 4116 1116
rect 4084 1035 4116 1036
rect 4084 1005 4085 1035
rect 4085 1005 4115 1035
rect 4115 1005 4116 1035
rect 4084 1004 4116 1005
rect 4084 955 4116 956
rect 4084 925 4085 955
rect 4085 925 4115 955
rect 4115 925 4116 955
rect 4084 924 4116 925
rect 4164 1675 4196 1676
rect 4164 1645 4165 1675
rect 4165 1645 4195 1675
rect 4195 1645 4196 1675
rect 4164 1644 4196 1645
rect 4164 1595 4196 1596
rect 4164 1565 4165 1595
rect 4165 1565 4195 1595
rect 4195 1565 4196 1595
rect 4164 1564 4196 1565
rect 4164 1484 4196 1516
rect 4164 1435 4196 1436
rect 4164 1405 4165 1435
rect 4165 1405 4195 1435
rect 4195 1405 4196 1435
rect 4164 1404 4196 1405
rect 4164 1355 4196 1356
rect 4164 1325 4165 1355
rect 4165 1325 4195 1355
rect 4195 1325 4196 1355
rect 4164 1324 4196 1325
rect 4164 1275 4196 1276
rect 4164 1245 4165 1275
rect 4165 1245 4195 1275
rect 4195 1245 4196 1275
rect 4164 1244 4196 1245
rect 4164 1195 4196 1196
rect 4164 1165 4165 1195
rect 4165 1165 4195 1195
rect 4195 1165 4196 1195
rect 4164 1164 4196 1165
rect 4164 1084 4196 1116
rect 4164 1035 4196 1036
rect 4164 1005 4165 1035
rect 4165 1005 4195 1035
rect 4195 1005 4196 1035
rect 4164 1004 4196 1005
rect 4164 955 4196 956
rect 4164 925 4165 955
rect 4165 925 4195 955
rect 4195 925 4196 955
rect 4164 924 4196 925
rect 4244 1675 4276 1676
rect 4244 1645 4245 1675
rect 4245 1645 4275 1675
rect 4275 1645 4276 1675
rect 4244 1644 4276 1645
rect 4244 1595 4276 1596
rect 4244 1565 4245 1595
rect 4245 1565 4275 1595
rect 4275 1565 4276 1595
rect 4244 1564 4276 1565
rect 4244 1484 4276 1516
rect 4244 1435 4276 1436
rect 4244 1405 4245 1435
rect 4245 1405 4275 1435
rect 4275 1405 4276 1435
rect 4244 1404 4276 1405
rect 4244 1355 4276 1356
rect 4244 1325 4245 1355
rect 4245 1325 4275 1355
rect 4275 1325 4276 1355
rect 4244 1324 4276 1325
rect 4244 1275 4276 1276
rect 4244 1245 4245 1275
rect 4245 1245 4275 1275
rect 4275 1245 4276 1275
rect 4244 1244 4276 1245
rect 4244 1195 4276 1196
rect 4244 1165 4245 1195
rect 4245 1165 4275 1195
rect 4275 1165 4276 1195
rect 4244 1164 4276 1165
rect 4244 1084 4276 1116
rect 4244 1035 4276 1036
rect 4244 1005 4245 1035
rect 4245 1005 4275 1035
rect 4275 1005 4276 1035
rect 4244 1004 4276 1005
rect 4244 955 4276 956
rect 4244 925 4245 955
rect 4245 925 4275 955
rect 4275 925 4276 955
rect 4244 924 4276 925
rect 4324 1675 4356 1676
rect 4324 1645 4325 1675
rect 4325 1645 4355 1675
rect 4355 1645 4356 1675
rect 4324 1644 4356 1645
rect 4324 1595 4356 1596
rect 4324 1565 4325 1595
rect 4325 1565 4355 1595
rect 4355 1565 4356 1595
rect 4324 1564 4356 1565
rect 4324 1484 4356 1516
rect 4324 1435 4356 1436
rect 4324 1405 4325 1435
rect 4325 1405 4355 1435
rect 4355 1405 4356 1435
rect 4324 1404 4356 1405
rect 4324 1355 4356 1356
rect 4324 1325 4325 1355
rect 4325 1325 4355 1355
rect 4355 1325 4356 1355
rect 4324 1324 4356 1325
rect 4324 1275 4356 1276
rect 4324 1245 4325 1275
rect 4325 1245 4355 1275
rect 4355 1245 4356 1275
rect 4324 1244 4356 1245
rect 4324 1195 4356 1196
rect 4324 1165 4325 1195
rect 4325 1165 4355 1195
rect 4355 1165 4356 1195
rect 4324 1164 4356 1165
rect 4324 1084 4356 1116
rect 4324 1035 4356 1036
rect 4324 1005 4325 1035
rect 4325 1005 4355 1035
rect 4355 1005 4356 1035
rect 4324 1004 4356 1005
rect 4324 955 4356 956
rect 4324 925 4325 955
rect 4325 925 4355 955
rect 4355 925 4356 955
rect 4324 924 4356 925
rect 4404 1675 4436 1676
rect 4404 1645 4405 1675
rect 4405 1645 4435 1675
rect 4435 1645 4436 1675
rect 4404 1644 4436 1645
rect 4404 1595 4436 1596
rect 4404 1565 4405 1595
rect 4405 1565 4435 1595
rect 4435 1565 4436 1595
rect 4404 1564 4436 1565
rect 4404 1484 4436 1516
rect 4404 1435 4436 1436
rect 4404 1405 4405 1435
rect 4405 1405 4435 1435
rect 4435 1405 4436 1435
rect 4404 1404 4436 1405
rect 4404 1355 4436 1356
rect 4404 1325 4405 1355
rect 4405 1325 4435 1355
rect 4435 1325 4436 1355
rect 4404 1324 4436 1325
rect 4404 1275 4436 1276
rect 4404 1245 4405 1275
rect 4405 1245 4435 1275
rect 4435 1245 4436 1275
rect 4404 1244 4436 1245
rect 4404 1195 4436 1196
rect 4404 1165 4405 1195
rect 4405 1165 4435 1195
rect 4435 1165 4436 1195
rect 4404 1164 4436 1165
rect 4404 1084 4436 1116
rect 4404 1035 4436 1036
rect 4404 1005 4405 1035
rect 4405 1005 4435 1035
rect 4435 1005 4436 1035
rect 4404 1004 4436 1005
rect 4404 955 4436 956
rect 4404 925 4405 955
rect 4405 925 4435 955
rect 4435 925 4436 955
rect 4404 924 4436 925
rect 4484 1675 4516 1676
rect 4484 1645 4485 1675
rect 4485 1645 4515 1675
rect 4515 1645 4516 1675
rect 4484 1644 4516 1645
rect 4484 1595 4516 1596
rect 4484 1565 4485 1595
rect 4485 1565 4515 1595
rect 4515 1565 4516 1595
rect 4484 1564 4516 1565
rect 4484 1484 4516 1516
rect 4484 1435 4516 1436
rect 4484 1405 4485 1435
rect 4485 1405 4515 1435
rect 4515 1405 4516 1435
rect 4484 1404 4516 1405
rect 4484 1355 4516 1356
rect 4484 1325 4485 1355
rect 4485 1325 4515 1355
rect 4515 1325 4516 1355
rect 4484 1324 4516 1325
rect 4484 1275 4516 1276
rect 4484 1245 4485 1275
rect 4485 1245 4515 1275
rect 4515 1245 4516 1275
rect 4484 1244 4516 1245
rect 4484 1195 4516 1196
rect 4484 1165 4485 1195
rect 4485 1165 4515 1195
rect 4515 1165 4516 1195
rect 4484 1164 4516 1165
rect 4484 1084 4516 1116
rect 4484 1035 4516 1036
rect 4484 1005 4485 1035
rect 4485 1005 4515 1035
rect 4515 1005 4516 1035
rect 4484 1004 4516 1005
rect 4484 955 4516 956
rect 4484 925 4485 955
rect 4485 925 4515 955
rect 4515 925 4516 955
rect 4484 924 4516 925
rect 4564 1675 4596 1676
rect 4564 1645 4565 1675
rect 4565 1645 4595 1675
rect 4595 1645 4596 1675
rect 4564 1644 4596 1645
rect 4564 1595 4596 1596
rect 4564 1565 4565 1595
rect 4565 1565 4595 1595
rect 4595 1565 4596 1595
rect 4564 1564 4596 1565
rect 4564 1484 4596 1516
rect 4564 1435 4596 1436
rect 4564 1405 4565 1435
rect 4565 1405 4595 1435
rect 4595 1405 4596 1435
rect 4564 1404 4596 1405
rect 4564 1355 4596 1356
rect 4564 1325 4565 1355
rect 4565 1325 4595 1355
rect 4595 1325 4596 1355
rect 4564 1324 4596 1325
rect 4564 1275 4596 1276
rect 4564 1245 4565 1275
rect 4565 1245 4595 1275
rect 4595 1245 4596 1275
rect 4564 1244 4596 1245
rect 4564 1195 4596 1196
rect 4564 1165 4565 1195
rect 4565 1165 4595 1195
rect 4595 1165 4596 1195
rect 4564 1164 4596 1165
rect 4564 1084 4596 1116
rect 4564 1035 4596 1036
rect 4564 1005 4565 1035
rect 4565 1005 4595 1035
rect 4595 1005 4596 1035
rect 4564 1004 4596 1005
rect 4564 955 4596 956
rect 4564 925 4565 955
rect 4565 925 4595 955
rect 4595 925 4596 955
rect 4564 924 4596 925
rect 4644 1675 4676 1676
rect 4644 1645 4645 1675
rect 4645 1645 4675 1675
rect 4675 1645 4676 1675
rect 4644 1644 4676 1645
rect 4644 1595 4676 1596
rect 4644 1565 4645 1595
rect 4645 1565 4675 1595
rect 4675 1565 4676 1595
rect 4644 1564 4676 1565
rect 4644 1484 4676 1516
rect 4644 1435 4676 1436
rect 4644 1405 4645 1435
rect 4645 1405 4675 1435
rect 4675 1405 4676 1435
rect 4644 1404 4676 1405
rect 4644 1355 4676 1356
rect 4644 1325 4645 1355
rect 4645 1325 4675 1355
rect 4675 1325 4676 1355
rect 4644 1324 4676 1325
rect 4644 1275 4676 1276
rect 4644 1245 4645 1275
rect 4645 1245 4675 1275
rect 4675 1245 4676 1275
rect 4644 1244 4676 1245
rect 4644 1195 4676 1196
rect 4644 1165 4645 1195
rect 4645 1165 4675 1195
rect 4675 1165 4676 1195
rect 4644 1164 4676 1165
rect 4644 1084 4676 1116
rect 4644 1035 4676 1036
rect 4644 1005 4645 1035
rect 4645 1005 4675 1035
rect 4675 1005 4676 1035
rect 4644 1004 4676 1005
rect 4644 955 4676 956
rect 4644 925 4645 955
rect 4645 925 4675 955
rect 4675 925 4676 955
rect 4644 924 4676 925
rect 4724 1675 4756 1676
rect 4724 1645 4725 1675
rect 4725 1645 4755 1675
rect 4755 1645 4756 1675
rect 4724 1644 4756 1645
rect 4724 1595 4756 1596
rect 4724 1565 4725 1595
rect 4725 1565 4755 1595
rect 4755 1565 4756 1595
rect 4724 1564 4756 1565
rect 4724 1484 4756 1516
rect 4724 1435 4756 1436
rect 4724 1405 4725 1435
rect 4725 1405 4755 1435
rect 4755 1405 4756 1435
rect 4724 1404 4756 1405
rect 4724 1355 4756 1356
rect 4724 1325 4725 1355
rect 4725 1325 4755 1355
rect 4755 1325 4756 1355
rect 4724 1324 4756 1325
rect 4724 1275 4756 1276
rect 4724 1245 4725 1275
rect 4725 1245 4755 1275
rect 4755 1245 4756 1275
rect 4724 1244 4756 1245
rect 4724 1195 4756 1196
rect 4724 1165 4725 1195
rect 4725 1165 4755 1195
rect 4755 1165 4756 1195
rect 4724 1164 4756 1165
rect 4724 1084 4756 1116
rect 4724 1035 4756 1036
rect 4724 1005 4725 1035
rect 4725 1005 4755 1035
rect 4755 1005 4756 1035
rect 4724 1004 4756 1005
rect 4724 955 4756 956
rect 4724 925 4725 955
rect 4725 925 4755 955
rect 4755 925 4756 955
rect 4724 924 4756 925
rect 4804 1675 4836 1676
rect 4804 1645 4805 1675
rect 4805 1645 4835 1675
rect 4835 1645 4836 1675
rect 4804 1644 4836 1645
rect 4804 1595 4836 1596
rect 4804 1565 4805 1595
rect 4805 1565 4835 1595
rect 4835 1565 4836 1595
rect 4804 1564 4836 1565
rect 4804 1484 4836 1516
rect 4804 1435 4836 1436
rect 4804 1405 4805 1435
rect 4805 1405 4835 1435
rect 4835 1405 4836 1435
rect 4804 1404 4836 1405
rect 4804 1355 4836 1356
rect 4804 1325 4805 1355
rect 4805 1325 4835 1355
rect 4835 1325 4836 1355
rect 4804 1324 4836 1325
rect 4804 1275 4836 1276
rect 4804 1245 4805 1275
rect 4805 1245 4835 1275
rect 4835 1245 4836 1275
rect 4804 1244 4836 1245
rect 4804 1195 4836 1196
rect 4804 1165 4805 1195
rect 4805 1165 4835 1195
rect 4835 1165 4836 1195
rect 4804 1164 4836 1165
rect 4804 1084 4836 1116
rect 4804 1035 4836 1036
rect 4804 1005 4805 1035
rect 4805 1005 4835 1035
rect 4835 1005 4836 1035
rect 4804 1004 4836 1005
rect 4804 955 4836 956
rect 4804 925 4805 955
rect 4805 925 4835 955
rect 4835 925 4836 955
rect 4804 924 4836 925
rect 4884 1675 4916 1676
rect 4884 1645 4885 1675
rect 4885 1645 4915 1675
rect 4915 1645 4916 1675
rect 4884 1644 4916 1645
rect 4884 1595 4916 1596
rect 4884 1565 4885 1595
rect 4885 1565 4915 1595
rect 4915 1565 4916 1595
rect 4884 1564 4916 1565
rect 4884 1515 4916 1516
rect 4884 1485 4885 1515
rect 4885 1485 4915 1515
rect 4915 1485 4916 1515
rect 4884 1484 4916 1485
rect 4884 1435 4916 1436
rect 4884 1405 4885 1435
rect 4885 1405 4915 1435
rect 4915 1405 4916 1435
rect 4884 1404 4916 1405
rect 4884 1355 4916 1356
rect 4884 1325 4885 1355
rect 4885 1325 4915 1355
rect 4915 1325 4916 1355
rect 4884 1324 4916 1325
rect 4884 1275 4916 1276
rect 4884 1245 4885 1275
rect 4885 1245 4915 1275
rect 4915 1245 4916 1275
rect 4884 1244 4916 1245
rect 4884 1195 4916 1196
rect 4884 1165 4885 1195
rect 4885 1165 4915 1195
rect 4915 1165 4916 1195
rect 4884 1164 4916 1165
rect 4884 1115 4916 1116
rect 4884 1085 4885 1115
rect 4885 1085 4915 1115
rect 4915 1085 4916 1115
rect 4884 1084 4916 1085
rect 4884 1035 4916 1036
rect 4884 1005 4885 1035
rect 4885 1005 4915 1035
rect 4915 1005 4916 1035
rect 4884 1004 4916 1005
rect 4884 955 4916 956
rect 4884 925 4885 955
rect 4885 925 4915 955
rect 4915 925 4916 955
rect 4884 924 4916 925
rect -876 875 -844 876
rect -876 845 -875 875
rect -875 845 -845 875
rect -845 845 -844 875
rect -876 844 -844 845
rect -876 795 -844 796
rect -876 765 -875 795
rect -875 765 -845 795
rect -845 765 -844 795
rect -876 764 -844 765
rect -876 715 -844 716
rect -876 685 -875 715
rect -875 685 -845 715
rect -845 685 -844 715
rect -876 684 -844 685
rect -876 635 -844 636
rect -876 605 -875 635
rect -875 605 -845 635
rect -845 605 -844 635
rect -876 604 -844 605
rect -876 555 -844 556
rect -876 525 -875 555
rect -875 525 -845 555
rect -845 525 -844 555
rect -876 524 -844 525
rect -876 475 -844 476
rect -876 445 -875 475
rect -875 445 -845 475
rect -845 445 -844 475
rect -876 444 -844 445
rect -876 395 -844 396
rect -876 365 -875 395
rect -875 365 -845 395
rect -845 365 -844 395
rect -876 364 -844 365
rect -876 315 -844 316
rect -876 285 -875 315
rect -875 285 -845 315
rect -845 285 -844 315
rect -876 284 -844 285
rect -876 235 -844 236
rect -876 205 -875 235
rect -875 205 -845 235
rect -845 205 -844 235
rect -876 204 -844 205
rect -876 155 -844 156
rect -876 125 -875 155
rect -875 125 -845 155
rect -845 125 -844 155
rect -876 124 -844 125
rect -876 75 -844 76
rect -876 45 -875 75
rect -875 45 -845 75
rect -845 45 -844 75
rect -876 44 -844 45
rect -876 -5 -844 -4
rect -876 -35 -875 -5
rect -875 -35 -845 -5
rect -845 -35 -844 -5
rect -876 -36 -844 -35
rect -876 -85 -844 -84
rect -876 -115 -875 -85
rect -875 -115 -845 -85
rect -845 -115 -844 -85
rect -876 -116 -844 -115
rect -796 875 -764 876
rect -796 845 -795 875
rect -795 845 -765 875
rect -765 845 -764 875
rect -796 844 -764 845
rect -796 764 -764 796
rect -796 715 -764 716
rect -796 685 -795 715
rect -795 685 -765 715
rect -765 685 -764 715
rect -796 684 -764 685
rect -796 604 -764 636
rect -796 555 -764 556
rect -796 525 -795 555
rect -795 525 -765 555
rect -765 525 -764 555
rect -796 524 -764 525
rect -796 444 -764 476
rect -796 395 -764 396
rect -796 365 -795 395
rect -795 365 -765 395
rect -765 365 -764 395
rect -796 364 -764 365
rect -796 284 -764 316
rect -796 235 -764 236
rect -796 205 -795 235
rect -795 205 -765 235
rect -765 205 -764 235
rect -796 204 -764 205
rect -796 155 -764 156
rect -796 125 -795 155
rect -795 125 -765 155
rect -765 125 -764 155
rect -796 124 -764 125
rect -796 75 -764 76
rect -796 45 -795 75
rect -795 45 -765 75
rect -765 45 -764 75
rect -796 44 -764 45
rect -796 -5 -764 -4
rect -796 -35 -795 -5
rect -795 -35 -765 -5
rect -765 -35 -764 -5
rect -796 -36 -764 -35
rect -796 -85 -764 -84
rect -796 -115 -795 -85
rect -795 -115 -765 -85
rect -765 -115 -764 -85
rect -796 -116 -764 -115
rect -716 875 -684 876
rect -716 845 -715 875
rect -715 845 -685 875
rect -685 845 -684 875
rect -716 844 -684 845
rect -716 764 -684 796
rect -716 715 -684 716
rect -716 685 -715 715
rect -715 685 -685 715
rect -685 685 -684 715
rect -716 684 -684 685
rect -716 604 -684 636
rect -716 555 -684 556
rect -716 525 -715 555
rect -715 525 -685 555
rect -685 525 -684 555
rect -716 524 -684 525
rect -716 444 -684 476
rect -716 395 -684 396
rect -716 365 -715 395
rect -715 365 -685 395
rect -685 365 -684 395
rect -716 364 -684 365
rect -716 284 -684 316
rect -716 235 -684 236
rect -716 205 -715 235
rect -715 205 -685 235
rect -685 205 -684 235
rect -716 204 -684 205
rect -716 155 -684 156
rect -716 125 -715 155
rect -715 125 -685 155
rect -685 125 -684 155
rect -716 124 -684 125
rect -716 75 -684 76
rect -716 45 -715 75
rect -715 45 -685 75
rect -685 45 -684 75
rect -716 44 -684 45
rect -716 -5 -684 -4
rect -716 -35 -715 -5
rect -715 -35 -685 -5
rect -685 -35 -684 -5
rect -716 -36 -684 -35
rect -716 -85 -684 -84
rect -716 -115 -715 -85
rect -715 -115 -685 -85
rect -685 -115 -684 -85
rect -716 -116 -684 -115
rect -636 875 -604 876
rect -636 845 -635 875
rect -635 845 -605 875
rect -605 845 -604 875
rect -636 844 -604 845
rect -636 764 -604 796
rect -636 715 -604 716
rect -636 685 -635 715
rect -635 685 -605 715
rect -605 685 -604 715
rect -636 684 -604 685
rect -636 604 -604 636
rect -636 555 -604 556
rect -636 525 -635 555
rect -635 525 -605 555
rect -605 525 -604 555
rect -636 524 -604 525
rect -636 444 -604 476
rect -636 395 -604 396
rect -636 365 -635 395
rect -635 365 -605 395
rect -605 365 -604 395
rect -636 364 -604 365
rect -636 284 -604 316
rect -636 235 -604 236
rect -636 205 -635 235
rect -635 205 -605 235
rect -605 205 -604 235
rect -636 204 -604 205
rect -636 155 -604 156
rect -636 125 -635 155
rect -635 125 -605 155
rect -605 125 -604 155
rect -636 124 -604 125
rect -636 75 -604 76
rect -636 45 -635 75
rect -635 45 -605 75
rect -605 45 -604 75
rect -636 44 -604 45
rect -636 -5 -604 -4
rect -636 -35 -635 -5
rect -635 -35 -605 -5
rect -605 -35 -604 -5
rect -636 -36 -604 -35
rect -636 -85 -604 -84
rect -636 -115 -635 -85
rect -635 -115 -605 -85
rect -605 -115 -604 -85
rect -636 -116 -604 -115
rect -556 875 -524 876
rect -556 845 -555 875
rect -555 845 -525 875
rect -525 845 -524 875
rect -556 844 -524 845
rect -556 764 -524 796
rect -556 715 -524 716
rect -556 685 -555 715
rect -555 685 -525 715
rect -525 685 -524 715
rect -556 684 -524 685
rect -556 604 -524 636
rect -556 555 -524 556
rect -556 525 -555 555
rect -555 525 -525 555
rect -525 525 -524 555
rect -556 524 -524 525
rect -556 444 -524 476
rect -556 395 -524 396
rect -556 365 -555 395
rect -555 365 -525 395
rect -525 365 -524 395
rect -556 364 -524 365
rect -556 284 -524 316
rect -556 235 -524 236
rect -556 205 -555 235
rect -555 205 -525 235
rect -525 205 -524 235
rect -556 204 -524 205
rect -556 155 -524 156
rect -556 125 -555 155
rect -555 125 -525 155
rect -525 125 -524 155
rect -556 124 -524 125
rect -556 75 -524 76
rect -556 45 -555 75
rect -555 45 -525 75
rect -525 45 -524 75
rect -556 44 -524 45
rect -556 -5 -524 -4
rect -556 -35 -555 -5
rect -555 -35 -525 -5
rect -525 -35 -524 -5
rect -556 -36 -524 -35
rect -556 -85 -524 -84
rect -556 -115 -555 -85
rect -555 -115 -525 -85
rect -525 -115 -524 -85
rect -556 -116 -524 -115
rect -476 875 -444 876
rect -476 845 -475 875
rect -475 845 -445 875
rect -445 845 -444 875
rect -476 844 -444 845
rect -476 764 -444 796
rect -476 715 -444 716
rect -476 685 -475 715
rect -475 685 -445 715
rect -445 685 -444 715
rect -476 684 -444 685
rect -476 604 -444 636
rect -476 555 -444 556
rect -476 525 -475 555
rect -475 525 -445 555
rect -445 525 -444 555
rect -476 524 -444 525
rect -476 444 -444 476
rect -476 395 -444 396
rect -476 365 -475 395
rect -475 365 -445 395
rect -445 365 -444 395
rect -476 364 -444 365
rect -476 284 -444 316
rect -476 235 -444 236
rect -476 205 -475 235
rect -475 205 -445 235
rect -445 205 -444 235
rect -476 204 -444 205
rect -476 155 -444 156
rect -476 125 -475 155
rect -475 125 -445 155
rect -445 125 -444 155
rect -476 124 -444 125
rect -476 75 -444 76
rect -476 45 -475 75
rect -475 45 -445 75
rect -445 45 -444 75
rect -476 44 -444 45
rect -476 -5 -444 -4
rect -476 -35 -475 -5
rect -475 -35 -445 -5
rect -445 -35 -444 -5
rect -476 -36 -444 -35
rect -476 -85 -444 -84
rect -476 -115 -475 -85
rect -475 -115 -445 -85
rect -445 -115 -444 -85
rect -476 -116 -444 -115
rect -396 875 -364 876
rect -396 845 -395 875
rect -395 845 -365 875
rect -365 845 -364 875
rect -396 844 -364 845
rect -396 764 -364 796
rect -396 715 -364 716
rect -396 685 -395 715
rect -395 685 -365 715
rect -365 685 -364 715
rect -396 684 -364 685
rect -396 604 -364 636
rect -396 555 -364 556
rect -396 525 -395 555
rect -395 525 -365 555
rect -365 525 -364 555
rect -396 524 -364 525
rect -396 444 -364 476
rect -396 395 -364 396
rect -396 365 -395 395
rect -395 365 -365 395
rect -365 365 -364 395
rect -396 364 -364 365
rect -396 284 -364 316
rect -396 235 -364 236
rect -396 205 -395 235
rect -395 205 -365 235
rect -365 205 -364 235
rect -396 204 -364 205
rect -396 155 -364 156
rect -396 125 -395 155
rect -395 125 -365 155
rect -365 125 -364 155
rect -396 124 -364 125
rect -396 75 -364 76
rect -396 45 -395 75
rect -395 45 -365 75
rect -365 45 -364 75
rect -396 44 -364 45
rect -396 -5 -364 -4
rect -396 -35 -395 -5
rect -395 -35 -365 -5
rect -365 -35 -364 -5
rect -396 -36 -364 -35
rect -396 -85 -364 -84
rect -396 -115 -395 -85
rect -395 -115 -365 -85
rect -365 -115 -364 -85
rect -396 -116 -364 -115
rect -316 875 -284 876
rect -316 845 -315 875
rect -315 845 -285 875
rect -285 845 -284 875
rect -316 844 -284 845
rect -316 764 -284 796
rect -316 715 -284 716
rect -316 685 -315 715
rect -315 685 -285 715
rect -285 685 -284 715
rect -316 684 -284 685
rect -316 604 -284 636
rect -316 555 -284 556
rect -316 525 -315 555
rect -315 525 -285 555
rect -285 525 -284 555
rect -316 524 -284 525
rect -316 444 -284 476
rect -316 395 -284 396
rect -316 365 -315 395
rect -315 365 -285 395
rect -285 365 -284 395
rect -316 364 -284 365
rect -316 284 -284 316
rect -316 235 -284 236
rect -316 205 -315 235
rect -315 205 -285 235
rect -285 205 -284 235
rect -316 204 -284 205
rect -316 155 -284 156
rect -316 125 -315 155
rect -315 125 -285 155
rect -285 125 -284 155
rect -316 124 -284 125
rect -316 75 -284 76
rect -316 45 -315 75
rect -315 45 -285 75
rect -285 45 -284 75
rect -316 44 -284 45
rect -316 -5 -284 -4
rect -316 -35 -315 -5
rect -315 -35 -285 -5
rect -285 -35 -284 -5
rect -316 -36 -284 -35
rect -316 -85 -284 -84
rect -316 -115 -315 -85
rect -315 -115 -285 -85
rect -285 -115 -284 -85
rect -316 -116 -284 -115
rect -236 875 -204 876
rect -236 845 -235 875
rect -235 845 -205 875
rect -205 845 -204 875
rect -236 844 -204 845
rect -236 764 -204 796
rect -236 715 -204 716
rect -236 685 -235 715
rect -235 685 -205 715
rect -205 685 -204 715
rect -236 684 -204 685
rect -236 604 -204 636
rect -236 555 -204 556
rect -236 525 -235 555
rect -235 525 -205 555
rect -205 525 -204 555
rect -236 524 -204 525
rect -236 444 -204 476
rect -236 395 -204 396
rect -236 365 -235 395
rect -235 365 -205 395
rect -205 365 -204 395
rect -236 364 -204 365
rect -236 284 -204 316
rect -236 235 -204 236
rect -236 205 -235 235
rect -235 205 -205 235
rect -205 205 -204 235
rect -236 204 -204 205
rect -236 155 -204 156
rect -236 125 -235 155
rect -235 125 -205 155
rect -205 125 -204 155
rect -236 124 -204 125
rect -236 75 -204 76
rect -236 45 -235 75
rect -235 45 -205 75
rect -205 45 -204 75
rect -236 44 -204 45
rect -236 -5 -204 -4
rect -236 -35 -235 -5
rect -235 -35 -205 -5
rect -205 -35 -204 -5
rect -236 -36 -204 -35
rect -236 -85 -204 -84
rect -236 -115 -235 -85
rect -235 -115 -205 -85
rect -205 -115 -204 -85
rect -236 -116 -204 -115
rect -156 875 -124 876
rect -156 845 -155 875
rect -155 845 -125 875
rect -125 845 -124 875
rect -156 844 -124 845
rect -156 764 -124 796
rect -156 715 -124 716
rect -156 685 -155 715
rect -155 685 -125 715
rect -125 685 -124 715
rect -156 684 -124 685
rect -156 604 -124 636
rect -156 555 -124 556
rect -156 525 -155 555
rect -155 525 -125 555
rect -125 525 -124 555
rect -156 524 -124 525
rect -156 444 -124 476
rect -156 395 -124 396
rect -156 365 -155 395
rect -155 365 -125 395
rect -125 365 -124 395
rect -156 364 -124 365
rect -156 284 -124 316
rect -156 235 -124 236
rect -156 205 -155 235
rect -155 205 -125 235
rect -125 205 -124 235
rect -156 204 -124 205
rect -156 155 -124 156
rect -156 125 -155 155
rect -155 125 -125 155
rect -125 125 -124 155
rect -156 124 -124 125
rect -156 75 -124 76
rect -156 45 -155 75
rect -155 45 -125 75
rect -125 45 -124 75
rect -156 44 -124 45
rect -156 -5 -124 -4
rect -156 -35 -155 -5
rect -155 -35 -125 -5
rect -125 -35 -124 -5
rect -156 -36 -124 -35
rect -156 -85 -124 -84
rect -156 -115 -155 -85
rect -155 -115 -125 -85
rect -125 -115 -124 -85
rect -156 -116 -124 -115
rect -76 875 -44 876
rect -76 845 -75 875
rect -75 845 -45 875
rect -45 845 -44 875
rect -76 844 -44 845
rect -76 764 -44 796
rect -76 715 -44 716
rect -76 685 -75 715
rect -75 685 -45 715
rect -45 685 -44 715
rect -76 684 -44 685
rect -76 604 -44 636
rect -76 555 -44 556
rect -76 525 -75 555
rect -75 525 -45 555
rect -45 525 -44 555
rect -76 524 -44 525
rect -76 444 -44 476
rect -76 395 -44 396
rect -76 365 -75 395
rect -75 365 -45 395
rect -45 365 -44 395
rect -76 364 -44 365
rect -76 284 -44 316
rect -76 235 -44 236
rect -76 205 -75 235
rect -75 205 -45 235
rect -45 205 -44 235
rect -76 204 -44 205
rect -76 155 -44 156
rect -76 125 -75 155
rect -75 125 -45 155
rect -45 125 -44 155
rect -76 124 -44 125
rect -76 75 -44 76
rect -76 45 -75 75
rect -75 45 -45 75
rect -45 45 -44 75
rect -76 44 -44 45
rect -76 -5 -44 -4
rect -76 -35 -75 -5
rect -75 -35 -45 -5
rect -45 -35 -44 -5
rect -76 -36 -44 -35
rect -76 -85 -44 -84
rect -76 -115 -75 -85
rect -75 -115 -45 -85
rect -45 -115 -44 -85
rect -76 -116 -44 -115
rect 4 875 36 876
rect 4 845 5 875
rect 5 845 35 875
rect 35 845 36 875
rect 4 844 36 845
rect 4 764 36 796
rect 4 715 36 716
rect 4 685 5 715
rect 5 685 35 715
rect 35 685 36 715
rect 4 684 36 685
rect 4 604 36 636
rect 4 555 36 556
rect 4 525 5 555
rect 5 525 35 555
rect 35 525 36 555
rect 4 524 36 525
rect 4 444 36 476
rect 4 395 36 396
rect 4 365 5 395
rect 5 365 35 395
rect 35 365 36 395
rect 4 364 36 365
rect 4 284 36 316
rect 4 235 36 236
rect 4 205 5 235
rect 5 205 35 235
rect 35 205 36 235
rect 4 204 36 205
rect 4 155 36 156
rect 4 125 5 155
rect 5 125 35 155
rect 35 125 36 155
rect 4 124 36 125
rect 4 75 36 76
rect 4 45 5 75
rect 5 45 35 75
rect 35 45 36 75
rect 4 44 36 45
rect 4 -5 36 -4
rect 4 -35 5 -5
rect 5 -35 35 -5
rect 35 -35 36 -5
rect 4 -36 36 -35
rect 4 -85 36 -84
rect 4 -115 5 -85
rect 5 -115 35 -85
rect 35 -115 36 -85
rect 4 -116 36 -115
rect 84 875 116 876
rect 84 845 85 875
rect 85 845 115 875
rect 115 845 116 875
rect 84 844 116 845
rect 84 764 116 796
rect 84 715 116 716
rect 84 685 85 715
rect 85 685 115 715
rect 115 685 116 715
rect 84 684 116 685
rect 84 604 116 636
rect 84 555 116 556
rect 84 525 85 555
rect 85 525 115 555
rect 115 525 116 555
rect 84 524 116 525
rect 84 444 116 476
rect 84 395 116 396
rect 84 365 85 395
rect 85 365 115 395
rect 115 365 116 395
rect 84 364 116 365
rect 84 284 116 316
rect 84 235 116 236
rect 84 205 85 235
rect 85 205 115 235
rect 115 205 116 235
rect 84 204 116 205
rect 84 155 116 156
rect 84 125 85 155
rect 85 125 115 155
rect 115 125 116 155
rect 84 124 116 125
rect 84 75 116 76
rect 84 45 85 75
rect 85 45 115 75
rect 115 45 116 75
rect 84 44 116 45
rect 84 -5 116 -4
rect 84 -35 85 -5
rect 85 -35 115 -5
rect 115 -35 116 -5
rect 84 -36 116 -35
rect 84 -85 116 -84
rect 84 -115 85 -85
rect 85 -115 115 -85
rect 115 -115 116 -85
rect 84 -116 116 -115
rect 164 875 196 876
rect 164 845 165 875
rect 165 845 195 875
rect 195 845 196 875
rect 164 844 196 845
rect 164 764 196 796
rect 164 715 196 716
rect 164 685 165 715
rect 165 685 195 715
rect 195 685 196 715
rect 164 684 196 685
rect 164 604 196 636
rect 164 555 196 556
rect 164 525 165 555
rect 165 525 195 555
rect 195 525 196 555
rect 164 524 196 525
rect 164 444 196 476
rect 164 395 196 396
rect 164 365 165 395
rect 165 365 195 395
rect 195 365 196 395
rect 164 364 196 365
rect 164 284 196 316
rect 164 235 196 236
rect 164 205 165 235
rect 165 205 195 235
rect 195 205 196 235
rect 164 204 196 205
rect 164 155 196 156
rect 164 125 165 155
rect 165 125 195 155
rect 195 125 196 155
rect 164 124 196 125
rect 164 75 196 76
rect 164 45 165 75
rect 165 45 195 75
rect 195 45 196 75
rect 164 44 196 45
rect 164 -5 196 -4
rect 164 -35 165 -5
rect 165 -35 195 -5
rect 195 -35 196 -5
rect 164 -36 196 -35
rect 164 -85 196 -84
rect 164 -115 165 -85
rect 165 -115 195 -85
rect 195 -115 196 -85
rect 164 -116 196 -115
rect 244 875 276 876
rect 244 845 245 875
rect 245 845 275 875
rect 275 845 276 875
rect 244 844 276 845
rect 244 764 276 796
rect 244 715 276 716
rect 244 685 245 715
rect 245 685 275 715
rect 275 685 276 715
rect 244 684 276 685
rect 244 604 276 636
rect 244 555 276 556
rect 244 525 245 555
rect 245 525 275 555
rect 275 525 276 555
rect 244 524 276 525
rect 244 444 276 476
rect 244 395 276 396
rect 244 365 245 395
rect 245 365 275 395
rect 275 365 276 395
rect 244 364 276 365
rect 244 284 276 316
rect 244 235 276 236
rect 244 205 245 235
rect 245 205 275 235
rect 275 205 276 235
rect 244 204 276 205
rect 244 155 276 156
rect 244 125 245 155
rect 245 125 275 155
rect 275 125 276 155
rect 244 124 276 125
rect 244 75 276 76
rect 244 45 245 75
rect 245 45 275 75
rect 275 45 276 75
rect 244 44 276 45
rect 244 -5 276 -4
rect 244 -35 245 -5
rect 245 -35 275 -5
rect 275 -35 276 -5
rect 244 -36 276 -35
rect 244 -85 276 -84
rect 244 -115 245 -85
rect 245 -115 275 -85
rect 275 -115 276 -85
rect 244 -116 276 -115
rect 324 875 356 876
rect 324 845 325 875
rect 325 845 355 875
rect 355 845 356 875
rect 324 844 356 845
rect 324 764 356 796
rect 324 715 356 716
rect 324 685 325 715
rect 325 685 355 715
rect 355 685 356 715
rect 324 684 356 685
rect 324 604 356 636
rect 324 555 356 556
rect 324 525 325 555
rect 325 525 355 555
rect 355 525 356 555
rect 324 524 356 525
rect 324 444 356 476
rect 324 395 356 396
rect 324 365 325 395
rect 325 365 355 395
rect 355 365 356 395
rect 324 364 356 365
rect 324 284 356 316
rect 324 235 356 236
rect 324 205 325 235
rect 325 205 355 235
rect 355 205 356 235
rect 324 204 356 205
rect 324 155 356 156
rect 324 125 325 155
rect 325 125 355 155
rect 355 125 356 155
rect 324 124 356 125
rect 324 75 356 76
rect 324 45 325 75
rect 325 45 355 75
rect 355 45 356 75
rect 324 44 356 45
rect 324 -5 356 -4
rect 324 -35 325 -5
rect 325 -35 355 -5
rect 355 -35 356 -5
rect 324 -36 356 -35
rect 324 -85 356 -84
rect 324 -115 325 -85
rect 325 -115 355 -85
rect 355 -115 356 -85
rect 324 -116 356 -115
rect 404 875 436 876
rect 404 845 405 875
rect 405 845 435 875
rect 435 845 436 875
rect 404 844 436 845
rect 404 764 436 796
rect 404 715 436 716
rect 404 685 405 715
rect 405 685 435 715
rect 435 685 436 715
rect 404 684 436 685
rect 404 604 436 636
rect 404 555 436 556
rect 404 525 405 555
rect 405 525 435 555
rect 435 525 436 555
rect 404 524 436 525
rect 404 444 436 476
rect 404 395 436 396
rect 404 365 405 395
rect 405 365 435 395
rect 435 365 436 395
rect 404 364 436 365
rect 404 284 436 316
rect 404 235 436 236
rect 404 205 405 235
rect 405 205 435 235
rect 435 205 436 235
rect 404 204 436 205
rect 404 155 436 156
rect 404 125 405 155
rect 405 125 435 155
rect 435 125 436 155
rect 404 124 436 125
rect 404 75 436 76
rect 404 45 405 75
rect 405 45 435 75
rect 435 45 436 75
rect 404 44 436 45
rect 404 -5 436 -4
rect 404 -35 405 -5
rect 405 -35 435 -5
rect 435 -35 436 -5
rect 404 -36 436 -35
rect 404 -85 436 -84
rect 404 -115 405 -85
rect 405 -115 435 -85
rect 435 -115 436 -85
rect 404 -116 436 -115
rect 484 875 516 876
rect 484 845 485 875
rect 485 845 515 875
rect 515 845 516 875
rect 484 844 516 845
rect 484 764 516 796
rect 484 715 516 716
rect 484 685 485 715
rect 485 685 515 715
rect 515 685 516 715
rect 484 684 516 685
rect 484 604 516 636
rect 484 555 516 556
rect 484 525 485 555
rect 485 525 515 555
rect 515 525 516 555
rect 484 524 516 525
rect 484 444 516 476
rect 484 395 516 396
rect 484 365 485 395
rect 485 365 515 395
rect 515 365 516 395
rect 484 364 516 365
rect 484 284 516 316
rect 484 235 516 236
rect 484 205 485 235
rect 485 205 515 235
rect 515 205 516 235
rect 484 204 516 205
rect 484 155 516 156
rect 484 125 485 155
rect 485 125 515 155
rect 515 125 516 155
rect 484 124 516 125
rect 484 75 516 76
rect 484 45 485 75
rect 485 45 515 75
rect 515 45 516 75
rect 484 44 516 45
rect 484 -5 516 -4
rect 484 -35 485 -5
rect 485 -35 515 -5
rect 515 -35 516 -5
rect 484 -36 516 -35
rect 484 -85 516 -84
rect 484 -115 485 -85
rect 485 -115 515 -85
rect 515 -115 516 -85
rect 484 -116 516 -115
rect 564 875 596 876
rect 564 845 565 875
rect 565 845 595 875
rect 595 845 596 875
rect 564 844 596 845
rect 564 764 596 796
rect 564 715 596 716
rect 564 685 565 715
rect 565 685 595 715
rect 595 685 596 715
rect 564 684 596 685
rect 564 604 596 636
rect 564 555 596 556
rect 564 525 565 555
rect 565 525 595 555
rect 595 525 596 555
rect 564 524 596 525
rect 564 444 596 476
rect 564 395 596 396
rect 564 365 565 395
rect 565 365 595 395
rect 595 365 596 395
rect 564 364 596 365
rect 564 284 596 316
rect 564 235 596 236
rect 564 205 565 235
rect 565 205 595 235
rect 595 205 596 235
rect 564 204 596 205
rect 564 155 596 156
rect 564 125 565 155
rect 565 125 595 155
rect 595 125 596 155
rect 564 124 596 125
rect 564 75 596 76
rect 564 45 565 75
rect 565 45 595 75
rect 595 45 596 75
rect 564 44 596 45
rect 564 -5 596 -4
rect 564 -35 565 -5
rect 565 -35 595 -5
rect 595 -35 596 -5
rect 564 -36 596 -35
rect 564 -85 596 -84
rect 564 -115 565 -85
rect 565 -115 595 -85
rect 595 -115 596 -85
rect 564 -116 596 -115
rect 644 875 676 876
rect 644 845 645 875
rect 645 845 675 875
rect 675 845 676 875
rect 644 844 676 845
rect 644 764 676 796
rect 644 715 676 716
rect 644 685 645 715
rect 645 685 675 715
rect 675 685 676 715
rect 644 684 676 685
rect 644 604 676 636
rect 644 555 676 556
rect 644 525 645 555
rect 645 525 675 555
rect 675 525 676 555
rect 644 524 676 525
rect 644 444 676 476
rect 644 395 676 396
rect 644 365 645 395
rect 645 365 675 395
rect 675 365 676 395
rect 644 364 676 365
rect 644 284 676 316
rect 644 235 676 236
rect 644 205 645 235
rect 645 205 675 235
rect 675 205 676 235
rect 644 204 676 205
rect 644 155 676 156
rect 644 125 645 155
rect 645 125 675 155
rect 675 125 676 155
rect 644 124 676 125
rect 644 75 676 76
rect 644 45 645 75
rect 645 45 675 75
rect 675 45 676 75
rect 644 44 676 45
rect 644 -5 676 -4
rect 644 -35 645 -5
rect 645 -35 675 -5
rect 675 -35 676 -5
rect 644 -36 676 -35
rect 644 -85 676 -84
rect 644 -115 645 -85
rect 645 -115 675 -85
rect 675 -115 676 -85
rect 644 -116 676 -115
rect 724 875 756 876
rect 724 845 725 875
rect 725 845 755 875
rect 755 845 756 875
rect 724 844 756 845
rect 724 764 756 796
rect 724 715 756 716
rect 724 685 725 715
rect 725 685 755 715
rect 755 685 756 715
rect 724 684 756 685
rect 724 604 756 636
rect 724 555 756 556
rect 724 525 725 555
rect 725 525 755 555
rect 755 525 756 555
rect 724 524 756 525
rect 724 444 756 476
rect 724 395 756 396
rect 724 365 725 395
rect 725 365 755 395
rect 755 365 756 395
rect 724 364 756 365
rect 724 284 756 316
rect 724 235 756 236
rect 724 205 725 235
rect 725 205 755 235
rect 755 205 756 235
rect 724 204 756 205
rect 724 155 756 156
rect 724 125 725 155
rect 725 125 755 155
rect 755 125 756 155
rect 724 124 756 125
rect 724 75 756 76
rect 724 45 725 75
rect 725 45 755 75
rect 755 45 756 75
rect 724 44 756 45
rect 724 -5 756 -4
rect 724 -35 725 -5
rect 725 -35 755 -5
rect 755 -35 756 -5
rect 724 -36 756 -35
rect 724 -85 756 -84
rect 724 -115 725 -85
rect 725 -115 755 -85
rect 755 -115 756 -85
rect 724 -116 756 -115
rect 804 875 836 876
rect 804 845 805 875
rect 805 845 835 875
rect 835 845 836 875
rect 804 844 836 845
rect 804 764 836 796
rect 804 715 836 716
rect 804 685 805 715
rect 805 685 835 715
rect 835 685 836 715
rect 804 684 836 685
rect 804 604 836 636
rect 804 555 836 556
rect 804 525 805 555
rect 805 525 835 555
rect 835 525 836 555
rect 804 524 836 525
rect 804 444 836 476
rect 804 395 836 396
rect 804 365 805 395
rect 805 365 835 395
rect 835 365 836 395
rect 804 364 836 365
rect 804 284 836 316
rect 804 235 836 236
rect 804 205 805 235
rect 805 205 835 235
rect 835 205 836 235
rect 804 204 836 205
rect 804 155 836 156
rect 804 125 805 155
rect 805 125 835 155
rect 835 125 836 155
rect 804 124 836 125
rect 804 75 836 76
rect 804 45 805 75
rect 805 45 835 75
rect 835 45 836 75
rect 804 44 836 45
rect 804 -5 836 -4
rect 804 -35 805 -5
rect 805 -35 835 -5
rect 835 -35 836 -5
rect 804 -36 836 -35
rect 804 -85 836 -84
rect 804 -115 805 -85
rect 805 -115 835 -85
rect 835 -115 836 -85
rect 804 -116 836 -115
rect 884 875 916 876
rect 884 845 885 875
rect 885 845 915 875
rect 915 845 916 875
rect 884 844 916 845
rect 884 764 916 796
rect 884 715 916 716
rect 884 685 885 715
rect 885 685 915 715
rect 915 685 916 715
rect 884 684 916 685
rect 884 604 916 636
rect 884 555 916 556
rect 884 525 885 555
rect 885 525 915 555
rect 915 525 916 555
rect 884 524 916 525
rect 884 444 916 476
rect 884 395 916 396
rect 884 365 885 395
rect 885 365 915 395
rect 915 365 916 395
rect 884 364 916 365
rect 884 284 916 316
rect 884 235 916 236
rect 884 205 885 235
rect 885 205 915 235
rect 915 205 916 235
rect 884 204 916 205
rect 884 155 916 156
rect 884 125 885 155
rect 885 125 915 155
rect 915 125 916 155
rect 884 124 916 125
rect 884 75 916 76
rect 884 45 885 75
rect 885 45 915 75
rect 915 45 916 75
rect 884 44 916 45
rect 884 -5 916 -4
rect 884 -35 885 -5
rect 885 -35 915 -5
rect 915 -35 916 -5
rect 884 -36 916 -35
rect 884 -85 916 -84
rect 884 -115 885 -85
rect 885 -115 915 -85
rect 915 -115 916 -85
rect 884 -116 916 -115
rect 964 875 996 876
rect 964 845 965 875
rect 965 845 995 875
rect 995 845 996 875
rect 964 844 996 845
rect 964 764 996 796
rect 964 715 996 716
rect 964 685 965 715
rect 965 685 995 715
rect 995 685 996 715
rect 964 684 996 685
rect 964 604 996 636
rect 964 555 996 556
rect 964 525 965 555
rect 965 525 995 555
rect 995 525 996 555
rect 964 524 996 525
rect 964 444 996 476
rect 964 395 996 396
rect 964 365 965 395
rect 965 365 995 395
rect 995 365 996 395
rect 964 364 996 365
rect 964 284 996 316
rect 964 235 996 236
rect 964 205 965 235
rect 965 205 995 235
rect 995 205 996 235
rect 964 204 996 205
rect 964 155 996 156
rect 964 125 965 155
rect 965 125 995 155
rect 995 125 996 155
rect 964 124 996 125
rect 964 75 996 76
rect 964 45 965 75
rect 965 45 995 75
rect 995 45 996 75
rect 964 44 996 45
rect 964 -5 996 -4
rect 964 -35 965 -5
rect 965 -35 995 -5
rect 995 -35 996 -5
rect 964 -36 996 -35
rect 964 -85 996 -84
rect 964 -115 965 -85
rect 965 -115 995 -85
rect 995 -115 996 -85
rect 964 -116 996 -115
rect 1044 875 1076 876
rect 1044 845 1045 875
rect 1045 845 1075 875
rect 1075 845 1076 875
rect 1044 844 1076 845
rect 1044 764 1076 796
rect 1044 715 1076 716
rect 1044 685 1045 715
rect 1045 685 1075 715
rect 1075 685 1076 715
rect 1044 684 1076 685
rect 1044 604 1076 636
rect 1044 555 1076 556
rect 1044 525 1045 555
rect 1045 525 1075 555
rect 1075 525 1076 555
rect 1044 524 1076 525
rect 1044 444 1076 476
rect 1044 395 1076 396
rect 1044 365 1045 395
rect 1045 365 1075 395
rect 1075 365 1076 395
rect 1044 364 1076 365
rect 1044 284 1076 316
rect 1044 235 1076 236
rect 1044 205 1045 235
rect 1045 205 1075 235
rect 1075 205 1076 235
rect 1044 204 1076 205
rect 1044 155 1076 156
rect 1044 125 1045 155
rect 1045 125 1075 155
rect 1075 125 1076 155
rect 1044 124 1076 125
rect 1044 75 1076 76
rect 1044 45 1045 75
rect 1045 45 1075 75
rect 1075 45 1076 75
rect 1044 44 1076 45
rect 1044 -5 1076 -4
rect 1044 -35 1045 -5
rect 1045 -35 1075 -5
rect 1075 -35 1076 -5
rect 1044 -36 1076 -35
rect 1044 -85 1076 -84
rect 1044 -115 1045 -85
rect 1045 -115 1075 -85
rect 1075 -115 1076 -85
rect 1044 -116 1076 -115
rect 1124 875 1156 876
rect 1124 845 1125 875
rect 1125 845 1155 875
rect 1155 845 1156 875
rect 1124 844 1156 845
rect 1124 764 1156 796
rect 1124 715 1156 716
rect 1124 685 1125 715
rect 1125 685 1155 715
rect 1155 685 1156 715
rect 1124 684 1156 685
rect 1124 604 1156 636
rect 1124 555 1156 556
rect 1124 525 1125 555
rect 1125 525 1155 555
rect 1155 525 1156 555
rect 1124 524 1156 525
rect 1124 444 1156 476
rect 1124 395 1156 396
rect 1124 365 1125 395
rect 1125 365 1155 395
rect 1155 365 1156 395
rect 1124 364 1156 365
rect 1124 284 1156 316
rect 1124 235 1156 236
rect 1124 205 1125 235
rect 1125 205 1155 235
rect 1155 205 1156 235
rect 1124 204 1156 205
rect 1124 155 1156 156
rect 1124 125 1125 155
rect 1125 125 1155 155
rect 1155 125 1156 155
rect 1124 124 1156 125
rect 1124 75 1156 76
rect 1124 45 1125 75
rect 1125 45 1155 75
rect 1155 45 1156 75
rect 1124 44 1156 45
rect 1124 -5 1156 -4
rect 1124 -35 1125 -5
rect 1125 -35 1155 -5
rect 1155 -35 1156 -5
rect 1124 -36 1156 -35
rect 1124 -85 1156 -84
rect 1124 -115 1125 -85
rect 1125 -115 1155 -85
rect 1155 -115 1156 -85
rect 1124 -116 1156 -115
rect 1204 875 1236 876
rect 1204 845 1205 875
rect 1205 845 1235 875
rect 1235 845 1236 875
rect 1204 844 1236 845
rect 1204 764 1236 796
rect 1204 715 1236 716
rect 1204 685 1205 715
rect 1205 685 1235 715
rect 1235 685 1236 715
rect 1204 684 1236 685
rect 1204 604 1236 636
rect 1204 555 1236 556
rect 1204 525 1205 555
rect 1205 525 1235 555
rect 1235 525 1236 555
rect 1204 524 1236 525
rect 1204 444 1236 476
rect 1204 395 1236 396
rect 1204 365 1205 395
rect 1205 365 1235 395
rect 1235 365 1236 395
rect 1204 364 1236 365
rect 1204 284 1236 316
rect 1204 235 1236 236
rect 1204 205 1205 235
rect 1205 205 1235 235
rect 1235 205 1236 235
rect 1204 204 1236 205
rect 1204 155 1236 156
rect 1204 125 1205 155
rect 1205 125 1235 155
rect 1235 125 1236 155
rect 1204 124 1236 125
rect 1204 75 1236 76
rect 1204 45 1205 75
rect 1205 45 1235 75
rect 1235 45 1236 75
rect 1204 44 1236 45
rect 1204 -5 1236 -4
rect 1204 -35 1205 -5
rect 1205 -35 1235 -5
rect 1235 -35 1236 -5
rect 1204 -36 1236 -35
rect 1204 -85 1236 -84
rect 1204 -115 1205 -85
rect 1205 -115 1235 -85
rect 1235 -115 1236 -85
rect 1204 -116 1236 -115
rect 1284 875 1316 876
rect 1284 845 1285 875
rect 1285 845 1315 875
rect 1315 845 1316 875
rect 1284 844 1316 845
rect 1284 764 1316 796
rect 1284 715 1316 716
rect 1284 685 1285 715
rect 1285 685 1315 715
rect 1315 685 1316 715
rect 1284 684 1316 685
rect 1284 604 1316 636
rect 1284 555 1316 556
rect 1284 525 1285 555
rect 1285 525 1315 555
rect 1315 525 1316 555
rect 1284 524 1316 525
rect 1284 444 1316 476
rect 1284 395 1316 396
rect 1284 365 1285 395
rect 1285 365 1315 395
rect 1315 365 1316 395
rect 1284 364 1316 365
rect 1284 284 1316 316
rect 1284 235 1316 236
rect 1284 205 1285 235
rect 1285 205 1315 235
rect 1315 205 1316 235
rect 1284 204 1316 205
rect 1284 155 1316 156
rect 1284 125 1285 155
rect 1285 125 1315 155
rect 1315 125 1316 155
rect 1284 124 1316 125
rect 1284 75 1316 76
rect 1284 45 1285 75
rect 1285 45 1315 75
rect 1315 45 1316 75
rect 1284 44 1316 45
rect 1284 -5 1316 -4
rect 1284 -35 1285 -5
rect 1285 -35 1315 -5
rect 1315 -35 1316 -5
rect 1284 -36 1316 -35
rect 1284 -85 1316 -84
rect 1284 -115 1285 -85
rect 1285 -115 1315 -85
rect 1315 -115 1316 -85
rect 1284 -116 1316 -115
rect 1364 875 1396 876
rect 1364 845 1365 875
rect 1365 845 1395 875
rect 1395 845 1396 875
rect 1364 844 1396 845
rect 1364 764 1396 796
rect 1364 715 1396 716
rect 1364 685 1365 715
rect 1365 685 1395 715
rect 1395 685 1396 715
rect 1364 684 1396 685
rect 1364 604 1396 636
rect 1364 555 1396 556
rect 1364 525 1365 555
rect 1365 525 1395 555
rect 1395 525 1396 555
rect 1364 524 1396 525
rect 1364 444 1396 476
rect 1364 395 1396 396
rect 1364 365 1365 395
rect 1365 365 1395 395
rect 1395 365 1396 395
rect 1364 364 1396 365
rect 1364 284 1396 316
rect 1364 235 1396 236
rect 1364 205 1365 235
rect 1365 205 1395 235
rect 1395 205 1396 235
rect 1364 204 1396 205
rect 1364 155 1396 156
rect 1364 125 1365 155
rect 1365 125 1395 155
rect 1395 125 1396 155
rect 1364 124 1396 125
rect 1364 75 1396 76
rect 1364 45 1365 75
rect 1365 45 1395 75
rect 1395 45 1396 75
rect 1364 44 1396 45
rect 1364 -5 1396 -4
rect 1364 -35 1365 -5
rect 1365 -35 1395 -5
rect 1395 -35 1396 -5
rect 1364 -36 1396 -35
rect 1364 -85 1396 -84
rect 1364 -115 1365 -85
rect 1365 -115 1395 -85
rect 1395 -115 1396 -85
rect 1364 -116 1396 -115
rect 1444 875 1476 876
rect 1444 845 1445 875
rect 1445 845 1475 875
rect 1475 845 1476 875
rect 1444 844 1476 845
rect 1444 764 1476 796
rect 1444 715 1476 716
rect 1444 685 1445 715
rect 1445 685 1475 715
rect 1475 685 1476 715
rect 1444 684 1476 685
rect 1444 604 1476 636
rect 1444 555 1476 556
rect 1444 525 1445 555
rect 1445 525 1475 555
rect 1475 525 1476 555
rect 1444 524 1476 525
rect 1444 444 1476 476
rect 1444 395 1476 396
rect 1444 365 1445 395
rect 1445 365 1475 395
rect 1475 365 1476 395
rect 1444 364 1476 365
rect 1444 284 1476 316
rect 1444 235 1476 236
rect 1444 205 1445 235
rect 1445 205 1475 235
rect 1475 205 1476 235
rect 1444 204 1476 205
rect 1444 155 1476 156
rect 1444 125 1445 155
rect 1445 125 1475 155
rect 1475 125 1476 155
rect 1444 124 1476 125
rect 1444 75 1476 76
rect 1444 45 1445 75
rect 1445 45 1475 75
rect 1475 45 1476 75
rect 1444 44 1476 45
rect 1444 -5 1476 -4
rect 1444 -35 1445 -5
rect 1445 -35 1475 -5
rect 1475 -35 1476 -5
rect 1444 -36 1476 -35
rect 1444 -85 1476 -84
rect 1444 -115 1445 -85
rect 1445 -115 1475 -85
rect 1475 -115 1476 -85
rect 1444 -116 1476 -115
rect 1524 875 1556 876
rect 1524 845 1525 875
rect 1525 845 1555 875
rect 1555 845 1556 875
rect 1524 844 1556 845
rect 1524 764 1556 796
rect 1524 715 1556 716
rect 1524 685 1525 715
rect 1525 685 1555 715
rect 1555 685 1556 715
rect 1524 684 1556 685
rect 1524 604 1556 636
rect 1524 555 1556 556
rect 1524 525 1525 555
rect 1525 525 1555 555
rect 1555 525 1556 555
rect 1524 524 1556 525
rect 1524 444 1556 476
rect 1524 395 1556 396
rect 1524 365 1525 395
rect 1525 365 1555 395
rect 1555 365 1556 395
rect 1524 364 1556 365
rect 1524 284 1556 316
rect 1524 235 1556 236
rect 1524 205 1525 235
rect 1525 205 1555 235
rect 1555 205 1556 235
rect 1524 204 1556 205
rect 1524 155 1556 156
rect 1524 125 1525 155
rect 1525 125 1555 155
rect 1555 125 1556 155
rect 1524 124 1556 125
rect 1524 75 1556 76
rect 1524 45 1525 75
rect 1525 45 1555 75
rect 1555 45 1556 75
rect 1524 44 1556 45
rect 1524 -5 1556 -4
rect 1524 -35 1525 -5
rect 1525 -35 1555 -5
rect 1555 -35 1556 -5
rect 1524 -36 1556 -35
rect 1524 -85 1556 -84
rect 1524 -115 1525 -85
rect 1525 -115 1555 -85
rect 1555 -115 1556 -85
rect 1524 -116 1556 -115
rect 1604 875 1636 876
rect 1604 845 1605 875
rect 1605 845 1635 875
rect 1635 845 1636 875
rect 1604 844 1636 845
rect 1604 764 1636 796
rect 1604 715 1636 716
rect 1604 685 1605 715
rect 1605 685 1635 715
rect 1635 685 1636 715
rect 1604 684 1636 685
rect 1604 604 1636 636
rect 1604 555 1636 556
rect 1604 525 1605 555
rect 1605 525 1635 555
rect 1635 525 1636 555
rect 1604 524 1636 525
rect 1604 444 1636 476
rect 1604 395 1636 396
rect 1604 365 1605 395
rect 1605 365 1635 395
rect 1635 365 1636 395
rect 1604 364 1636 365
rect 1604 284 1636 316
rect 1604 235 1636 236
rect 1604 205 1605 235
rect 1605 205 1635 235
rect 1635 205 1636 235
rect 1604 204 1636 205
rect 1604 155 1636 156
rect 1604 125 1605 155
rect 1605 125 1635 155
rect 1635 125 1636 155
rect 1604 124 1636 125
rect 1604 75 1636 76
rect 1604 45 1605 75
rect 1605 45 1635 75
rect 1635 45 1636 75
rect 1604 44 1636 45
rect 1604 -5 1636 -4
rect 1604 -35 1605 -5
rect 1605 -35 1635 -5
rect 1635 -35 1636 -5
rect 1604 -36 1636 -35
rect 1604 -85 1636 -84
rect 1604 -115 1605 -85
rect 1605 -115 1635 -85
rect 1635 -115 1636 -85
rect 1604 -116 1636 -115
rect 1684 875 1716 876
rect 1684 845 1685 875
rect 1685 845 1715 875
rect 1715 845 1716 875
rect 1684 844 1716 845
rect 1684 764 1716 796
rect 1684 715 1716 716
rect 1684 685 1685 715
rect 1685 685 1715 715
rect 1715 685 1716 715
rect 1684 684 1716 685
rect 1684 604 1716 636
rect 1684 555 1716 556
rect 1684 525 1685 555
rect 1685 525 1715 555
rect 1715 525 1716 555
rect 1684 524 1716 525
rect 1684 444 1716 476
rect 1684 395 1716 396
rect 1684 365 1685 395
rect 1685 365 1715 395
rect 1715 365 1716 395
rect 1684 364 1716 365
rect 1684 284 1716 316
rect 1684 235 1716 236
rect 1684 205 1685 235
rect 1685 205 1715 235
rect 1715 205 1716 235
rect 1684 204 1716 205
rect 1684 155 1716 156
rect 1684 125 1685 155
rect 1685 125 1715 155
rect 1715 125 1716 155
rect 1684 124 1716 125
rect 1684 75 1716 76
rect 1684 45 1685 75
rect 1685 45 1715 75
rect 1715 45 1716 75
rect 1684 44 1716 45
rect 1684 -5 1716 -4
rect 1684 -35 1685 -5
rect 1685 -35 1715 -5
rect 1715 -35 1716 -5
rect 1684 -36 1716 -35
rect 1684 -85 1716 -84
rect 1684 -115 1685 -85
rect 1685 -115 1715 -85
rect 1715 -115 1716 -85
rect 1684 -116 1716 -115
rect 1764 875 1796 876
rect 1764 845 1765 875
rect 1765 845 1795 875
rect 1795 845 1796 875
rect 1764 844 1796 845
rect 1764 764 1796 796
rect 1764 715 1796 716
rect 1764 685 1765 715
rect 1765 685 1795 715
rect 1795 685 1796 715
rect 1764 684 1796 685
rect 1764 604 1796 636
rect 1764 555 1796 556
rect 1764 525 1765 555
rect 1765 525 1795 555
rect 1795 525 1796 555
rect 1764 524 1796 525
rect 1764 444 1796 476
rect 1764 395 1796 396
rect 1764 365 1765 395
rect 1765 365 1795 395
rect 1795 365 1796 395
rect 1764 364 1796 365
rect 1764 284 1796 316
rect 1764 235 1796 236
rect 1764 205 1765 235
rect 1765 205 1795 235
rect 1795 205 1796 235
rect 1764 204 1796 205
rect 1764 155 1796 156
rect 1764 125 1765 155
rect 1765 125 1795 155
rect 1795 125 1796 155
rect 1764 124 1796 125
rect 1764 75 1796 76
rect 1764 45 1765 75
rect 1765 45 1795 75
rect 1795 45 1796 75
rect 1764 44 1796 45
rect 1764 -5 1796 -4
rect 1764 -35 1765 -5
rect 1765 -35 1795 -5
rect 1795 -35 1796 -5
rect 1764 -36 1796 -35
rect 1764 -85 1796 -84
rect 1764 -115 1765 -85
rect 1765 -115 1795 -85
rect 1795 -115 1796 -85
rect 1764 -116 1796 -115
rect 1844 875 1876 876
rect 1844 845 1845 875
rect 1845 845 1875 875
rect 1875 845 1876 875
rect 1844 844 1876 845
rect 1844 764 1876 796
rect 1844 715 1876 716
rect 1844 685 1845 715
rect 1845 685 1875 715
rect 1875 685 1876 715
rect 1844 684 1876 685
rect 1844 604 1876 636
rect 1844 555 1876 556
rect 1844 525 1845 555
rect 1845 525 1875 555
rect 1875 525 1876 555
rect 1844 524 1876 525
rect 1844 444 1876 476
rect 1844 395 1876 396
rect 1844 365 1845 395
rect 1845 365 1875 395
rect 1875 365 1876 395
rect 1844 364 1876 365
rect 1844 284 1876 316
rect 1844 235 1876 236
rect 1844 205 1845 235
rect 1845 205 1875 235
rect 1875 205 1876 235
rect 1844 204 1876 205
rect 1844 155 1876 156
rect 1844 125 1845 155
rect 1845 125 1875 155
rect 1875 125 1876 155
rect 1844 124 1876 125
rect 1844 75 1876 76
rect 1844 45 1845 75
rect 1845 45 1875 75
rect 1875 45 1876 75
rect 1844 44 1876 45
rect 1844 -5 1876 -4
rect 1844 -35 1845 -5
rect 1845 -35 1875 -5
rect 1875 -35 1876 -5
rect 1844 -36 1876 -35
rect 1844 -85 1876 -84
rect 1844 -115 1845 -85
rect 1845 -115 1875 -85
rect 1875 -115 1876 -85
rect 1844 -116 1876 -115
rect 1924 875 1956 876
rect 1924 845 1925 875
rect 1925 845 1955 875
rect 1955 845 1956 875
rect 1924 844 1956 845
rect 1924 764 1956 796
rect 1924 715 1956 716
rect 1924 685 1925 715
rect 1925 685 1955 715
rect 1955 685 1956 715
rect 1924 684 1956 685
rect 1924 604 1956 636
rect 1924 555 1956 556
rect 1924 525 1925 555
rect 1925 525 1955 555
rect 1955 525 1956 555
rect 1924 524 1956 525
rect 1924 444 1956 476
rect 1924 395 1956 396
rect 1924 365 1925 395
rect 1925 365 1955 395
rect 1955 365 1956 395
rect 1924 364 1956 365
rect 1924 284 1956 316
rect 1924 235 1956 236
rect 1924 205 1925 235
rect 1925 205 1955 235
rect 1955 205 1956 235
rect 1924 204 1956 205
rect 1924 155 1956 156
rect 1924 125 1925 155
rect 1925 125 1955 155
rect 1955 125 1956 155
rect 1924 124 1956 125
rect 1924 75 1956 76
rect 1924 45 1925 75
rect 1925 45 1955 75
rect 1955 45 1956 75
rect 1924 44 1956 45
rect 1924 -5 1956 -4
rect 1924 -35 1925 -5
rect 1925 -35 1955 -5
rect 1955 -35 1956 -5
rect 1924 -36 1956 -35
rect 1924 -85 1956 -84
rect 1924 -115 1925 -85
rect 1925 -115 1955 -85
rect 1955 -115 1956 -85
rect 1924 -116 1956 -115
rect 2004 875 2036 876
rect 2004 845 2005 875
rect 2005 845 2035 875
rect 2035 845 2036 875
rect 2004 844 2036 845
rect 2004 764 2036 796
rect 2004 715 2036 716
rect 2004 685 2005 715
rect 2005 685 2035 715
rect 2035 685 2036 715
rect 2004 684 2036 685
rect 2004 604 2036 636
rect 2004 555 2036 556
rect 2004 525 2005 555
rect 2005 525 2035 555
rect 2035 525 2036 555
rect 2004 524 2036 525
rect 2004 444 2036 476
rect 2004 395 2036 396
rect 2004 365 2005 395
rect 2005 365 2035 395
rect 2035 365 2036 395
rect 2004 364 2036 365
rect 2004 284 2036 316
rect 2004 235 2036 236
rect 2004 205 2005 235
rect 2005 205 2035 235
rect 2035 205 2036 235
rect 2004 204 2036 205
rect 2004 155 2036 156
rect 2004 125 2005 155
rect 2005 125 2035 155
rect 2035 125 2036 155
rect 2004 124 2036 125
rect 2004 75 2036 76
rect 2004 45 2005 75
rect 2005 45 2035 75
rect 2035 45 2036 75
rect 2004 44 2036 45
rect 2004 -5 2036 -4
rect 2004 -35 2005 -5
rect 2005 -35 2035 -5
rect 2035 -35 2036 -5
rect 2004 -36 2036 -35
rect 2004 -85 2036 -84
rect 2004 -115 2005 -85
rect 2005 -115 2035 -85
rect 2035 -115 2036 -85
rect 2004 -116 2036 -115
rect 2084 875 2116 876
rect 2084 845 2085 875
rect 2085 845 2115 875
rect 2115 845 2116 875
rect 2084 844 2116 845
rect 2084 764 2116 796
rect 2084 715 2116 716
rect 2084 685 2085 715
rect 2085 685 2115 715
rect 2115 685 2116 715
rect 2084 684 2116 685
rect 2084 604 2116 636
rect 2084 555 2116 556
rect 2084 525 2085 555
rect 2085 525 2115 555
rect 2115 525 2116 555
rect 2084 524 2116 525
rect 2084 444 2116 476
rect 2084 395 2116 396
rect 2084 365 2085 395
rect 2085 365 2115 395
rect 2115 365 2116 395
rect 2084 364 2116 365
rect 2084 284 2116 316
rect 2084 235 2116 236
rect 2084 205 2085 235
rect 2085 205 2115 235
rect 2115 205 2116 235
rect 2084 204 2116 205
rect 2084 155 2116 156
rect 2084 125 2085 155
rect 2085 125 2115 155
rect 2115 125 2116 155
rect 2084 124 2116 125
rect 2084 75 2116 76
rect 2084 45 2085 75
rect 2085 45 2115 75
rect 2115 45 2116 75
rect 2084 44 2116 45
rect 2084 -5 2116 -4
rect 2084 -35 2085 -5
rect 2085 -35 2115 -5
rect 2115 -35 2116 -5
rect 2084 -36 2116 -35
rect 2084 -85 2116 -84
rect 2084 -115 2085 -85
rect 2085 -115 2115 -85
rect 2115 -115 2116 -85
rect 2084 -116 2116 -115
rect 2164 875 2196 876
rect 2164 845 2165 875
rect 2165 845 2195 875
rect 2195 845 2196 875
rect 2164 844 2196 845
rect 2164 764 2196 796
rect 2164 715 2196 716
rect 2164 685 2165 715
rect 2165 685 2195 715
rect 2195 685 2196 715
rect 2164 684 2196 685
rect 2164 604 2196 636
rect 2164 555 2196 556
rect 2164 525 2165 555
rect 2165 525 2195 555
rect 2195 525 2196 555
rect 2164 524 2196 525
rect 2164 444 2196 476
rect 2164 395 2196 396
rect 2164 365 2165 395
rect 2165 365 2195 395
rect 2195 365 2196 395
rect 2164 364 2196 365
rect 2164 284 2196 316
rect 2164 235 2196 236
rect 2164 205 2165 235
rect 2165 205 2195 235
rect 2195 205 2196 235
rect 2164 204 2196 205
rect 2164 155 2196 156
rect 2164 125 2165 155
rect 2165 125 2195 155
rect 2195 125 2196 155
rect 2164 124 2196 125
rect 2164 75 2196 76
rect 2164 45 2165 75
rect 2165 45 2195 75
rect 2195 45 2196 75
rect 2164 44 2196 45
rect 2164 -5 2196 -4
rect 2164 -35 2165 -5
rect 2165 -35 2195 -5
rect 2195 -35 2196 -5
rect 2164 -36 2196 -35
rect 2164 -85 2196 -84
rect 2164 -115 2165 -85
rect 2165 -115 2195 -85
rect 2195 -115 2196 -85
rect 2164 -116 2196 -115
rect 2244 875 2276 876
rect 2244 845 2245 875
rect 2245 845 2275 875
rect 2275 845 2276 875
rect 2244 844 2276 845
rect 2244 764 2276 796
rect 2244 715 2276 716
rect 2244 685 2245 715
rect 2245 685 2275 715
rect 2275 685 2276 715
rect 2244 684 2276 685
rect 2244 604 2276 636
rect 2244 555 2276 556
rect 2244 525 2245 555
rect 2245 525 2275 555
rect 2275 525 2276 555
rect 2244 524 2276 525
rect 2244 444 2276 476
rect 2244 395 2276 396
rect 2244 365 2245 395
rect 2245 365 2275 395
rect 2275 365 2276 395
rect 2244 364 2276 365
rect 2244 284 2276 316
rect 2244 235 2276 236
rect 2244 205 2245 235
rect 2245 205 2275 235
rect 2275 205 2276 235
rect 2244 204 2276 205
rect 2244 155 2276 156
rect 2244 125 2245 155
rect 2245 125 2275 155
rect 2275 125 2276 155
rect 2244 124 2276 125
rect 2244 75 2276 76
rect 2244 45 2245 75
rect 2245 45 2275 75
rect 2275 45 2276 75
rect 2244 44 2276 45
rect 2244 -5 2276 -4
rect 2244 -35 2245 -5
rect 2245 -35 2275 -5
rect 2275 -35 2276 -5
rect 2244 -36 2276 -35
rect 2244 -85 2276 -84
rect 2244 -115 2245 -85
rect 2245 -115 2275 -85
rect 2275 -115 2276 -85
rect 2244 -116 2276 -115
rect 2324 875 2356 876
rect 2324 845 2325 875
rect 2325 845 2355 875
rect 2355 845 2356 875
rect 2324 844 2356 845
rect 2324 764 2356 796
rect 2324 715 2356 716
rect 2324 685 2325 715
rect 2325 685 2355 715
rect 2355 685 2356 715
rect 2324 684 2356 685
rect 2324 604 2356 636
rect 2324 555 2356 556
rect 2324 525 2325 555
rect 2325 525 2355 555
rect 2355 525 2356 555
rect 2324 524 2356 525
rect 2324 444 2356 476
rect 2324 395 2356 396
rect 2324 365 2325 395
rect 2325 365 2355 395
rect 2355 365 2356 395
rect 2324 364 2356 365
rect 2324 284 2356 316
rect 2324 235 2356 236
rect 2324 205 2325 235
rect 2325 205 2355 235
rect 2355 205 2356 235
rect 2324 204 2356 205
rect 2324 155 2356 156
rect 2324 125 2325 155
rect 2325 125 2355 155
rect 2355 125 2356 155
rect 2324 124 2356 125
rect 2324 75 2356 76
rect 2324 45 2325 75
rect 2325 45 2355 75
rect 2355 45 2356 75
rect 2324 44 2356 45
rect 2324 -5 2356 -4
rect 2324 -35 2325 -5
rect 2325 -35 2355 -5
rect 2355 -35 2356 -5
rect 2324 -36 2356 -35
rect 2324 -85 2356 -84
rect 2324 -115 2325 -85
rect 2325 -115 2355 -85
rect 2355 -115 2356 -85
rect 2324 -116 2356 -115
rect 2404 875 2436 876
rect 2404 845 2405 875
rect 2405 845 2435 875
rect 2435 845 2436 875
rect 2404 844 2436 845
rect 2404 764 2436 796
rect 2404 715 2436 716
rect 2404 685 2405 715
rect 2405 685 2435 715
rect 2435 685 2436 715
rect 2404 684 2436 685
rect 2404 604 2436 636
rect 2404 555 2436 556
rect 2404 525 2405 555
rect 2405 525 2435 555
rect 2435 525 2436 555
rect 2404 524 2436 525
rect 2404 444 2436 476
rect 2404 395 2436 396
rect 2404 365 2405 395
rect 2405 365 2435 395
rect 2435 365 2436 395
rect 2404 364 2436 365
rect 2404 284 2436 316
rect 2404 235 2436 236
rect 2404 205 2405 235
rect 2405 205 2435 235
rect 2435 205 2436 235
rect 2404 204 2436 205
rect 2404 155 2436 156
rect 2404 125 2405 155
rect 2405 125 2435 155
rect 2435 125 2436 155
rect 2404 124 2436 125
rect 2404 75 2436 76
rect 2404 45 2405 75
rect 2405 45 2435 75
rect 2435 45 2436 75
rect 2404 44 2436 45
rect 2404 -5 2436 -4
rect 2404 -35 2405 -5
rect 2405 -35 2435 -5
rect 2435 -35 2436 -5
rect 2404 -36 2436 -35
rect 2404 -85 2436 -84
rect 2404 -115 2405 -85
rect 2405 -115 2435 -85
rect 2435 -115 2436 -85
rect 2404 -116 2436 -115
rect 2484 875 2516 876
rect 2484 845 2485 875
rect 2485 845 2515 875
rect 2515 845 2516 875
rect 2484 844 2516 845
rect 2484 764 2516 796
rect 2484 715 2516 716
rect 2484 685 2485 715
rect 2485 685 2515 715
rect 2515 685 2516 715
rect 2484 684 2516 685
rect 2484 604 2516 636
rect 2484 555 2516 556
rect 2484 525 2485 555
rect 2485 525 2515 555
rect 2515 525 2516 555
rect 2484 524 2516 525
rect 2484 444 2516 476
rect 2484 395 2516 396
rect 2484 365 2485 395
rect 2485 365 2515 395
rect 2515 365 2516 395
rect 2484 364 2516 365
rect 2484 284 2516 316
rect 2484 235 2516 236
rect 2484 205 2485 235
rect 2485 205 2515 235
rect 2515 205 2516 235
rect 2484 204 2516 205
rect 2484 155 2516 156
rect 2484 125 2485 155
rect 2485 125 2515 155
rect 2515 125 2516 155
rect 2484 124 2516 125
rect 2484 75 2516 76
rect 2484 45 2485 75
rect 2485 45 2515 75
rect 2515 45 2516 75
rect 2484 44 2516 45
rect 2484 -5 2516 -4
rect 2484 -35 2485 -5
rect 2485 -35 2515 -5
rect 2515 -35 2516 -5
rect 2484 -36 2516 -35
rect 2484 -85 2516 -84
rect 2484 -115 2485 -85
rect 2485 -115 2515 -85
rect 2515 -115 2516 -85
rect 2484 -116 2516 -115
rect 2564 875 2596 876
rect 2564 845 2565 875
rect 2565 845 2595 875
rect 2595 845 2596 875
rect 2564 844 2596 845
rect 2564 764 2596 796
rect 2564 715 2596 716
rect 2564 685 2565 715
rect 2565 685 2595 715
rect 2595 685 2596 715
rect 2564 684 2596 685
rect 2564 604 2596 636
rect 2564 555 2596 556
rect 2564 525 2565 555
rect 2565 525 2595 555
rect 2595 525 2596 555
rect 2564 524 2596 525
rect 2564 444 2596 476
rect 2564 395 2596 396
rect 2564 365 2565 395
rect 2565 365 2595 395
rect 2595 365 2596 395
rect 2564 364 2596 365
rect 2564 284 2596 316
rect 2564 235 2596 236
rect 2564 205 2565 235
rect 2565 205 2595 235
rect 2595 205 2596 235
rect 2564 204 2596 205
rect 2564 155 2596 156
rect 2564 125 2565 155
rect 2565 125 2595 155
rect 2595 125 2596 155
rect 2564 124 2596 125
rect 2564 75 2596 76
rect 2564 45 2565 75
rect 2565 45 2595 75
rect 2595 45 2596 75
rect 2564 44 2596 45
rect 2564 -5 2596 -4
rect 2564 -35 2565 -5
rect 2565 -35 2595 -5
rect 2595 -35 2596 -5
rect 2564 -36 2596 -35
rect 2564 -85 2596 -84
rect 2564 -115 2565 -85
rect 2565 -115 2595 -85
rect 2595 -115 2596 -85
rect 2564 -116 2596 -115
rect 2644 875 2676 876
rect 2644 845 2645 875
rect 2645 845 2675 875
rect 2675 845 2676 875
rect 2644 844 2676 845
rect 2644 764 2676 796
rect 2644 715 2676 716
rect 2644 685 2645 715
rect 2645 685 2675 715
rect 2675 685 2676 715
rect 2644 684 2676 685
rect 2644 604 2676 636
rect 2644 555 2676 556
rect 2644 525 2645 555
rect 2645 525 2675 555
rect 2675 525 2676 555
rect 2644 524 2676 525
rect 2644 444 2676 476
rect 2644 395 2676 396
rect 2644 365 2645 395
rect 2645 365 2675 395
rect 2675 365 2676 395
rect 2644 364 2676 365
rect 2644 284 2676 316
rect 2644 235 2676 236
rect 2644 205 2645 235
rect 2645 205 2675 235
rect 2675 205 2676 235
rect 2644 204 2676 205
rect 2644 155 2676 156
rect 2644 125 2645 155
rect 2645 125 2675 155
rect 2675 125 2676 155
rect 2644 124 2676 125
rect 2644 75 2676 76
rect 2644 45 2645 75
rect 2645 45 2675 75
rect 2675 45 2676 75
rect 2644 44 2676 45
rect 2644 -5 2676 -4
rect 2644 -35 2645 -5
rect 2645 -35 2675 -5
rect 2675 -35 2676 -5
rect 2644 -36 2676 -35
rect 2644 -85 2676 -84
rect 2644 -115 2645 -85
rect 2645 -115 2675 -85
rect 2675 -115 2676 -85
rect 2644 -116 2676 -115
rect 2724 875 2756 876
rect 2724 845 2725 875
rect 2725 845 2755 875
rect 2755 845 2756 875
rect 2724 844 2756 845
rect 2724 764 2756 796
rect 2724 715 2756 716
rect 2724 685 2725 715
rect 2725 685 2755 715
rect 2755 685 2756 715
rect 2724 684 2756 685
rect 2724 604 2756 636
rect 2724 555 2756 556
rect 2724 525 2725 555
rect 2725 525 2755 555
rect 2755 525 2756 555
rect 2724 524 2756 525
rect 2724 444 2756 476
rect 2724 395 2756 396
rect 2724 365 2725 395
rect 2725 365 2755 395
rect 2755 365 2756 395
rect 2724 364 2756 365
rect 2724 284 2756 316
rect 2724 235 2756 236
rect 2724 205 2725 235
rect 2725 205 2755 235
rect 2755 205 2756 235
rect 2724 204 2756 205
rect 2724 155 2756 156
rect 2724 125 2725 155
rect 2725 125 2755 155
rect 2755 125 2756 155
rect 2724 124 2756 125
rect 2724 75 2756 76
rect 2724 45 2725 75
rect 2725 45 2755 75
rect 2755 45 2756 75
rect 2724 44 2756 45
rect 2724 -5 2756 -4
rect 2724 -35 2725 -5
rect 2725 -35 2755 -5
rect 2755 -35 2756 -5
rect 2724 -36 2756 -35
rect 2724 -85 2756 -84
rect 2724 -115 2725 -85
rect 2725 -115 2755 -85
rect 2755 -115 2756 -85
rect 2724 -116 2756 -115
rect 2804 875 2836 876
rect 2804 845 2805 875
rect 2805 845 2835 875
rect 2835 845 2836 875
rect 2804 844 2836 845
rect 2804 764 2836 796
rect 2804 715 2836 716
rect 2804 685 2805 715
rect 2805 685 2835 715
rect 2835 685 2836 715
rect 2804 684 2836 685
rect 2804 604 2836 636
rect 2804 555 2836 556
rect 2804 525 2805 555
rect 2805 525 2835 555
rect 2835 525 2836 555
rect 2804 524 2836 525
rect 2804 444 2836 476
rect 2804 395 2836 396
rect 2804 365 2805 395
rect 2805 365 2835 395
rect 2835 365 2836 395
rect 2804 364 2836 365
rect 2804 284 2836 316
rect 2804 235 2836 236
rect 2804 205 2805 235
rect 2805 205 2835 235
rect 2835 205 2836 235
rect 2804 204 2836 205
rect 2804 155 2836 156
rect 2804 125 2805 155
rect 2805 125 2835 155
rect 2835 125 2836 155
rect 2804 124 2836 125
rect 2804 75 2836 76
rect 2804 45 2805 75
rect 2805 45 2835 75
rect 2835 45 2836 75
rect 2804 44 2836 45
rect 2804 -5 2836 -4
rect 2804 -35 2805 -5
rect 2805 -35 2835 -5
rect 2835 -35 2836 -5
rect 2804 -36 2836 -35
rect 2804 -85 2836 -84
rect 2804 -115 2805 -85
rect 2805 -115 2835 -85
rect 2835 -115 2836 -85
rect 2804 -116 2836 -115
rect 2884 875 2916 876
rect 2884 845 2885 875
rect 2885 845 2915 875
rect 2915 845 2916 875
rect 2884 844 2916 845
rect 2884 764 2916 796
rect 2884 715 2916 716
rect 2884 685 2885 715
rect 2885 685 2915 715
rect 2915 685 2916 715
rect 2884 684 2916 685
rect 2884 604 2916 636
rect 2884 555 2916 556
rect 2884 525 2885 555
rect 2885 525 2915 555
rect 2915 525 2916 555
rect 2884 524 2916 525
rect 2884 444 2916 476
rect 2884 395 2916 396
rect 2884 365 2885 395
rect 2885 365 2915 395
rect 2915 365 2916 395
rect 2884 364 2916 365
rect 2884 284 2916 316
rect 2884 235 2916 236
rect 2884 205 2885 235
rect 2885 205 2915 235
rect 2915 205 2916 235
rect 2884 204 2916 205
rect 2884 155 2916 156
rect 2884 125 2885 155
rect 2885 125 2915 155
rect 2915 125 2916 155
rect 2884 124 2916 125
rect 2884 75 2916 76
rect 2884 45 2885 75
rect 2885 45 2915 75
rect 2915 45 2916 75
rect 2884 44 2916 45
rect 2884 -5 2916 -4
rect 2884 -35 2885 -5
rect 2885 -35 2915 -5
rect 2915 -35 2916 -5
rect 2884 -36 2916 -35
rect 2884 -85 2916 -84
rect 2884 -115 2885 -85
rect 2885 -115 2915 -85
rect 2915 -115 2916 -85
rect 2884 -116 2916 -115
rect 2964 875 2996 876
rect 2964 845 2965 875
rect 2965 845 2995 875
rect 2995 845 2996 875
rect 2964 844 2996 845
rect 2964 764 2996 796
rect 2964 715 2996 716
rect 2964 685 2965 715
rect 2965 685 2995 715
rect 2995 685 2996 715
rect 2964 684 2996 685
rect 2964 604 2996 636
rect 2964 555 2996 556
rect 2964 525 2965 555
rect 2965 525 2995 555
rect 2995 525 2996 555
rect 2964 524 2996 525
rect 2964 444 2996 476
rect 2964 395 2996 396
rect 2964 365 2965 395
rect 2965 365 2995 395
rect 2995 365 2996 395
rect 2964 364 2996 365
rect 2964 284 2996 316
rect 2964 235 2996 236
rect 2964 205 2965 235
rect 2965 205 2995 235
rect 2995 205 2996 235
rect 2964 204 2996 205
rect 2964 155 2996 156
rect 2964 125 2965 155
rect 2965 125 2995 155
rect 2995 125 2996 155
rect 2964 124 2996 125
rect 2964 75 2996 76
rect 2964 45 2965 75
rect 2965 45 2995 75
rect 2995 45 2996 75
rect 2964 44 2996 45
rect 2964 -5 2996 -4
rect 2964 -35 2965 -5
rect 2965 -35 2995 -5
rect 2995 -35 2996 -5
rect 2964 -36 2996 -35
rect 2964 -85 2996 -84
rect 2964 -115 2965 -85
rect 2965 -115 2995 -85
rect 2995 -115 2996 -85
rect 2964 -116 2996 -115
rect 3044 875 3076 876
rect 3044 845 3045 875
rect 3045 845 3075 875
rect 3075 845 3076 875
rect 3044 844 3076 845
rect 3044 764 3076 796
rect 3044 715 3076 716
rect 3044 685 3045 715
rect 3045 685 3075 715
rect 3075 685 3076 715
rect 3044 684 3076 685
rect 3044 604 3076 636
rect 3044 555 3076 556
rect 3044 525 3045 555
rect 3045 525 3075 555
rect 3075 525 3076 555
rect 3044 524 3076 525
rect 3044 444 3076 476
rect 3044 395 3076 396
rect 3044 365 3045 395
rect 3045 365 3075 395
rect 3075 365 3076 395
rect 3044 364 3076 365
rect 3044 284 3076 316
rect 3044 235 3076 236
rect 3044 205 3045 235
rect 3045 205 3075 235
rect 3075 205 3076 235
rect 3044 204 3076 205
rect 3044 155 3076 156
rect 3044 125 3045 155
rect 3045 125 3075 155
rect 3075 125 3076 155
rect 3044 124 3076 125
rect 3044 75 3076 76
rect 3044 45 3045 75
rect 3045 45 3075 75
rect 3075 45 3076 75
rect 3044 44 3076 45
rect 3044 -5 3076 -4
rect 3044 -35 3045 -5
rect 3045 -35 3075 -5
rect 3075 -35 3076 -5
rect 3044 -36 3076 -35
rect 3044 -85 3076 -84
rect 3044 -115 3045 -85
rect 3045 -115 3075 -85
rect 3075 -115 3076 -85
rect 3044 -116 3076 -115
rect 3124 875 3156 876
rect 3124 845 3125 875
rect 3125 845 3155 875
rect 3155 845 3156 875
rect 3124 844 3156 845
rect 3124 764 3156 796
rect 3124 715 3156 716
rect 3124 685 3125 715
rect 3125 685 3155 715
rect 3155 685 3156 715
rect 3124 684 3156 685
rect 3124 604 3156 636
rect 3124 555 3156 556
rect 3124 525 3125 555
rect 3125 525 3155 555
rect 3155 525 3156 555
rect 3124 524 3156 525
rect 3124 444 3156 476
rect 3124 395 3156 396
rect 3124 365 3125 395
rect 3125 365 3155 395
rect 3155 365 3156 395
rect 3124 364 3156 365
rect 3124 284 3156 316
rect 3124 235 3156 236
rect 3124 205 3125 235
rect 3125 205 3155 235
rect 3155 205 3156 235
rect 3124 204 3156 205
rect 3124 155 3156 156
rect 3124 125 3125 155
rect 3125 125 3155 155
rect 3155 125 3156 155
rect 3124 124 3156 125
rect 3124 75 3156 76
rect 3124 45 3125 75
rect 3125 45 3155 75
rect 3155 45 3156 75
rect 3124 44 3156 45
rect 3124 -5 3156 -4
rect 3124 -35 3125 -5
rect 3125 -35 3155 -5
rect 3155 -35 3156 -5
rect 3124 -36 3156 -35
rect 3124 -85 3156 -84
rect 3124 -115 3125 -85
rect 3125 -115 3155 -85
rect 3155 -115 3156 -85
rect 3124 -116 3156 -115
rect 3204 875 3236 876
rect 3204 845 3205 875
rect 3205 845 3235 875
rect 3235 845 3236 875
rect 3204 844 3236 845
rect 3204 764 3236 796
rect 3204 715 3236 716
rect 3204 685 3205 715
rect 3205 685 3235 715
rect 3235 685 3236 715
rect 3204 684 3236 685
rect 3204 604 3236 636
rect 3204 555 3236 556
rect 3204 525 3205 555
rect 3205 525 3235 555
rect 3235 525 3236 555
rect 3204 524 3236 525
rect 3204 444 3236 476
rect 3204 395 3236 396
rect 3204 365 3205 395
rect 3205 365 3235 395
rect 3235 365 3236 395
rect 3204 364 3236 365
rect 3204 284 3236 316
rect 3204 235 3236 236
rect 3204 205 3205 235
rect 3205 205 3235 235
rect 3235 205 3236 235
rect 3204 204 3236 205
rect 3204 155 3236 156
rect 3204 125 3205 155
rect 3205 125 3235 155
rect 3235 125 3236 155
rect 3204 124 3236 125
rect 3204 75 3236 76
rect 3204 45 3205 75
rect 3205 45 3235 75
rect 3235 45 3236 75
rect 3204 44 3236 45
rect 3204 -5 3236 -4
rect 3204 -35 3205 -5
rect 3205 -35 3235 -5
rect 3235 -35 3236 -5
rect 3204 -36 3236 -35
rect 3204 -85 3236 -84
rect 3204 -115 3205 -85
rect 3205 -115 3235 -85
rect 3235 -115 3236 -85
rect 3204 -116 3236 -115
rect 3284 875 3316 876
rect 3284 845 3285 875
rect 3285 845 3315 875
rect 3315 845 3316 875
rect 3284 844 3316 845
rect 3284 764 3316 796
rect 3284 715 3316 716
rect 3284 685 3285 715
rect 3285 685 3315 715
rect 3315 685 3316 715
rect 3284 684 3316 685
rect 3284 604 3316 636
rect 3284 555 3316 556
rect 3284 525 3285 555
rect 3285 525 3315 555
rect 3315 525 3316 555
rect 3284 524 3316 525
rect 3284 444 3316 476
rect 3284 395 3316 396
rect 3284 365 3285 395
rect 3285 365 3315 395
rect 3315 365 3316 395
rect 3284 364 3316 365
rect 3284 284 3316 316
rect 3284 235 3316 236
rect 3284 205 3285 235
rect 3285 205 3315 235
rect 3315 205 3316 235
rect 3284 204 3316 205
rect 3284 155 3316 156
rect 3284 125 3285 155
rect 3285 125 3315 155
rect 3315 125 3316 155
rect 3284 124 3316 125
rect 3284 75 3316 76
rect 3284 45 3285 75
rect 3285 45 3315 75
rect 3315 45 3316 75
rect 3284 44 3316 45
rect 3284 -5 3316 -4
rect 3284 -35 3285 -5
rect 3285 -35 3315 -5
rect 3315 -35 3316 -5
rect 3284 -36 3316 -35
rect 3284 -85 3316 -84
rect 3284 -115 3285 -85
rect 3285 -115 3315 -85
rect 3315 -115 3316 -85
rect 3284 -116 3316 -115
rect 3364 875 3396 876
rect 3364 845 3365 875
rect 3365 845 3395 875
rect 3395 845 3396 875
rect 3364 844 3396 845
rect 3364 764 3396 796
rect 3364 715 3396 716
rect 3364 685 3365 715
rect 3365 685 3395 715
rect 3395 685 3396 715
rect 3364 684 3396 685
rect 3364 604 3396 636
rect 3364 555 3396 556
rect 3364 525 3365 555
rect 3365 525 3395 555
rect 3395 525 3396 555
rect 3364 524 3396 525
rect 3364 444 3396 476
rect 3364 395 3396 396
rect 3364 365 3365 395
rect 3365 365 3395 395
rect 3395 365 3396 395
rect 3364 364 3396 365
rect 3364 284 3396 316
rect 3364 235 3396 236
rect 3364 205 3365 235
rect 3365 205 3395 235
rect 3395 205 3396 235
rect 3364 204 3396 205
rect 3364 155 3396 156
rect 3364 125 3365 155
rect 3365 125 3395 155
rect 3395 125 3396 155
rect 3364 124 3396 125
rect 3364 75 3396 76
rect 3364 45 3365 75
rect 3365 45 3395 75
rect 3395 45 3396 75
rect 3364 44 3396 45
rect 3364 -5 3396 -4
rect 3364 -35 3365 -5
rect 3365 -35 3395 -5
rect 3395 -35 3396 -5
rect 3364 -36 3396 -35
rect 3364 -85 3396 -84
rect 3364 -115 3365 -85
rect 3365 -115 3395 -85
rect 3395 -115 3396 -85
rect 3364 -116 3396 -115
rect 3444 875 3476 876
rect 3444 845 3445 875
rect 3445 845 3475 875
rect 3475 845 3476 875
rect 3444 844 3476 845
rect 3444 764 3476 796
rect 3444 715 3476 716
rect 3444 685 3445 715
rect 3445 685 3475 715
rect 3475 685 3476 715
rect 3444 684 3476 685
rect 3444 604 3476 636
rect 3444 555 3476 556
rect 3444 525 3445 555
rect 3445 525 3475 555
rect 3475 525 3476 555
rect 3444 524 3476 525
rect 3444 444 3476 476
rect 3444 395 3476 396
rect 3444 365 3445 395
rect 3445 365 3475 395
rect 3475 365 3476 395
rect 3444 364 3476 365
rect 3444 284 3476 316
rect 3444 235 3476 236
rect 3444 205 3445 235
rect 3445 205 3475 235
rect 3475 205 3476 235
rect 3444 204 3476 205
rect 3444 155 3476 156
rect 3444 125 3445 155
rect 3445 125 3475 155
rect 3475 125 3476 155
rect 3444 124 3476 125
rect 3444 75 3476 76
rect 3444 45 3445 75
rect 3445 45 3475 75
rect 3475 45 3476 75
rect 3444 44 3476 45
rect 3444 -5 3476 -4
rect 3444 -35 3445 -5
rect 3445 -35 3475 -5
rect 3475 -35 3476 -5
rect 3444 -36 3476 -35
rect 3444 -85 3476 -84
rect 3444 -115 3445 -85
rect 3445 -115 3475 -85
rect 3475 -115 3476 -85
rect 3444 -116 3476 -115
rect 3524 875 3556 876
rect 3524 845 3525 875
rect 3525 845 3555 875
rect 3555 845 3556 875
rect 3524 844 3556 845
rect 3524 764 3556 796
rect 3524 715 3556 716
rect 3524 685 3525 715
rect 3525 685 3555 715
rect 3555 685 3556 715
rect 3524 684 3556 685
rect 3524 604 3556 636
rect 3524 555 3556 556
rect 3524 525 3525 555
rect 3525 525 3555 555
rect 3555 525 3556 555
rect 3524 524 3556 525
rect 3524 444 3556 476
rect 3524 395 3556 396
rect 3524 365 3525 395
rect 3525 365 3555 395
rect 3555 365 3556 395
rect 3524 364 3556 365
rect 3524 284 3556 316
rect 3524 235 3556 236
rect 3524 205 3525 235
rect 3525 205 3555 235
rect 3555 205 3556 235
rect 3524 204 3556 205
rect 3524 155 3556 156
rect 3524 125 3525 155
rect 3525 125 3555 155
rect 3555 125 3556 155
rect 3524 124 3556 125
rect 3524 75 3556 76
rect 3524 45 3525 75
rect 3525 45 3555 75
rect 3555 45 3556 75
rect 3524 44 3556 45
rect 3524 -5 3556 -4
rect 3524 -35 3525 -5
rect 3525 -35 3555 -5
rect 3555 -35 3556 -5
rect 3524 -36 3556 -35
rect 3524 -85 3556 -84
rect 3524 -115 3525 -85
rect 3525 -115 3555 -85
rect 3555 -115 3556 -85
rect 3524 -116 3556 -115
rect 3604 875 3636 876
rect 3604 845 3605 875
rect 3605 845 3635 875
rect 3635 845 3636 875
rect 3604 844 3636 845
rect 3604 764 3636 796
rect 3604 715 3636 716
rect 3604 685 3605 715
rect 3605 685 3635 715
rect 3635 685 3636 715
rect 3604 684 3636 685
rect 3604 604 3636 636
rect 3604 555 3636 556
rect 3604 525 3605 555
rect 3605 525 3635 555
rect 3635 525 3636 555
rect 3604 524 3636 525
rect 3604 444 3636 476
rect 3604 395 3636 396
rect 3604 365 3605 395
rect 3605 365 3635 395
rect 3635 365 3636 395
rect 3604 364 3636 365
rect 3604 284 3636 316
rect 3604 235 3636 236
rect 3604 205 3605 235
rect 3605 205 3635 235
rect 3635 205 3636 235
rect 3604 204 3636 205
rect 3604 155 3636 156
rect 3604 125 3605 155
rect 3605 125 3635 155
rect 3635 125 3636 155
rect 3604 124 3636 125
rect 3604 75 3636 76
rect 3604 45 3605 75
rect 3605 45 3635 75
rect 3635 45 3636 75
rect 3604 44 3636 45
rect 3604 -5 3636 -4
rect 3604 -35 3605 -5
rect 3605 -35 3635 -5
rect 3635 -35 3636 -5
rect 3604 -36 3636 -35
rect 3604 -85 3636 -84
rect 3604 -115 3605 -85
rect 3605 -115 3635 -85
rect 3635 -115 3636 -85
rect 3604 -116 3636 -115
rect 3684 875 3716 876
rect 3684 845 3685 875
rect 3685 845 3715 875
rect 3715 845 3716 875
rect 3684 844 3716 845
rect 3684 764 3716 796
rect 3684 715 3716 716
rect 3684 685 3685 715
rect 3685 685 3715 715
rect 3715 685 3716 715
rect 3684 684 3716 685
rect 3684 604 3716 636
rect 3684 555 3716 556
rect 3684 525 3685 555
rect 3685 525 3715 555
rect 3715 525 3716 555
rect 3684 524 3716 525
rect 3684 444 3716 476
rect 3684 395 3716 396
rect 3684 365 3685 395
rect 3685 365 3715 395
rect 3715 365 3716 395
rect 3684 364 3716 365
rect 3684 284 3716 316
rect 3684 235 3716 236
rect 3684 205 3685 235
rect 3685 205 3715 235
rect 3715 205 3716 235
rect 3684 204 3716 205
rect 3684 155 3716 156
rect 3684 125 3685 155
rect 3685 125 3715 155
rect 3715 125 3716 155
rect 3684 124 3716 125
rect 3684 75 3716 76
rect 3684 45 3685 75
rect 3685 45 3715 75
rect 3715 45 3716 75
rect 3684 44 3716 45
rect 3684 -5 3716 -4
rect 3684 -35 3685 -5
rect 3685 -35 3715 -5
rect 3715 -35 3716 -5
rect 3684 -36 3716 -35
rect 3684 -85 3716 -84
rect 3684 -115 3685 -85
rect 3685 -115 3715 -85
rect 3715 -115 3716 -85
rect 3684 -116 3716 -115
rect 3764 875 3796 876
rect 3764 845 3765 875
rect 3765 845 3795 875
rect 3795 845 3796 875
rect 3764 844 3796 845
rect 3764 764 3796 796
rect 3764 715 3796 716
rect 3764 685 3765 715
rect 3765 685 3795 715
rect 3795 685 3796 715
rect 3764 684 3796 685
rect 3764 604 3796 636
rect 3764 555 3796 556
rect 3764 525 3765 555
rect 3765 525 3795 555
rect 3795 525 3796 555
rect 3764 524 3796 525
rect 3764 444 3796 476
rect 3764 395 3796 396
rect 3764 365 3765 395
rect 3765 365 3795 395
rect 3795 365 3796 395
rect 3764 364 3796 365
rect 3764 284 3796 316
rect 3764 235 3796 236
rect 3764 205 3765 235
rect 3765 205 3795 235
rect 3795 205 3796 235
rect 3764 204 3796 205
rect 3764 155 3796 156
rect 3764 125 3765 155
rect 3765 125 3795 155
rect 3795 125 3796 155
rect 3764 124 3796 125
rect 3764 75 3796 76
rect 3764 45 3765 75
rect 3765 45 3795 75
rect 3795 45 3796 75
rect 3764 44 3796 45
rect 3764 -5 3796 -4
rect 3764 -35 3765 -5
rect 3765 -35 3795 -5
rect 3795 -35 3796 -5
rect 3764 -36 3796 -35
rect 3764 -85 3796 -84
rect 3764 -115 3765 -85
rect 3765 -115 3795 -85
rect 3795 -115 3796 -85
rect 3764 -116 3796 -115
rect 3844 875 3876 876
rect 3844 845 3845 875
rect 3845 845 3875 875
rect 3875 845 3876 875
rect 3844 844 3876 845
rect 3844 764 3876 796
rect 3844 715 3876 716
rect 3844 685 3845 715
rect 3845 685 3875 715
rect 3875 685 3876 715
rect 3844 684 3876 685
rect 3844 604 3876 636
rect 3844 555 3876 556
rect 3844 525 3845 555
rect 3845 525 3875 555
rect 3875 525 3876 555
rect 3844 524 3876 525
rect 3844 444 3876 476
rect 3844 395 3876 396
rect 3844 365 3845 395
rect 3845 365 3875 395
rect 3875 365 3876 395
rect 3844 364 3876 365
rect 3844 284 3876 316
rect 3844 235 3876 236
rect 3844 205 3845 235
rect 3845 205 3875 235
rect 3875 205 3876 235
rect 3844 204 3876 205
rect 3844 155 3876 156
rect 3844 125 3845 155
rect 3845 125 3875 155
rect 3875 125 3876 155
rect 3844 124 3876 125
rect 3844 75 3876 76
rect 3844 45 3845 75
rect 3845 45 3875 75
rect 3875 45 3876 75
rect 3844 44 3876 45
rect 3844 -5 3876 -4
rect 3844 -35 3845 -5
rect 3845 -35 3875 -5
rect 3875 -35 3876 -5
rect 3844 -36 3876 -35
rect 3844 -85 3876 -84
rect 3844 -115 3845 -85
rect 3845 -115 3875 -85
rect 3875 -115 3876 -85
rect 3844 -116 3876 -115
rect 3924 875 3956 876
rect 3924 845 3925 875
rect 3925 845 3955 875
rect 3955 845 3956 875
rect 3924 844 3956 845
rect 3924 764 3956 796
rect 3924 715 3956 716
rect 3924 685 3925 715
rect 3925 685 3955 715
rect 3955 685 3956 715
rect 3924 684 3956 685
rect 3924 604 3956 636
rect 3924 555 3956 556
rect 3924 525 3925 555
rect 3925 525 3955 555
rect 3955 525 3956 555
rect 3924 524 3956 525
rect 3924 444 3956 476
rect 3924 395 3956 396
rect 3924 365 3925 395
rect 3925 365 3955 395
rect 3955 365 3956 395
rect 3924 364 3956 365
rect 3924 284 3956 316
rect 3924 235 3956 236
rect 3924 205 3925 235
rect 3925 205 3955 235
rect 3955 205 3956 235
rect 3924 204 3956 205
rect 3924 155 3956 156
rect 3924 125 3925 155
rect 3925 125 3955 155
rect 3955 125 3956 155
rect 3924 124 3956 125
rect 3924 75 3956 76
rect 3924 45 3925 75
rect 3925 45 3955 75
rect 3955 45 3956 75
rect 3924 44 3956 45
rect 3924 -5 3956 -4
rect 3924 -35 3925 -5
rect 3925 -35 3955 -5
rect 3955 -35 3956 -5
rect 3924 -36 3956 -35
rect 3924 -85 3956 -84
rect 3924 -115 3925 -85
rect 3925 -115 3955 -85
rect 3955 -115 3956 -85
rect 3924 -116 3956 -115
rect 4004 875 4036 876
rect 4004 845 4005 875
rect 4005 845 4035 875
rect 4035 845 4036 875
rect 4004 844 4036 845
rect 4004 764 4036 796
rect 4004 715 4036 716
rect 4004 685 4005 715
rect 4005 685 4035 715
rect 4035 685 4036 715
rect 4004 684 4036 685
rect 4004 604 4036 636
rect 4004 555 4036 556
rect 4004 525 4005 555
rect 4005 525 4035 555
rect 4035 525 4036 555
rect 4004 524 4036 525
rect 4004 444 4036 476
rect 4004 395 4036 396
rect 4004 365 4005 395
rect 4005 365 4035 395
rect 4035 365 4036 395
rect 4004 364 4036 365
rect 4004 284 4036 316
rect 4004 235 4036 236
rect 4004 205 4005 235
rect 4005 205 4035 235
rect 4035 205 4036 235
rect 4004 204 4036 205
rect 4004 155 4036 156
rect 4004 125 4005 155
rect 4005 125 4035 155
rect 4035 125 4036 155
rect 4004 124 4036 125
rect 4004 75 4036 76
rect 4004 45 4005 75
rect 4005 45 4035 75
rect 4035 45 4036 75
rect 4004 44 4036 45
rect 4004 -5 4036 -4
rect 4004 -35 4005 -5
rect 4005 -35 4035 -5
rect 4035 -35 4036 -5
rect 4004 -36 4036 -35
rect 4004 -85 4036 -84
rect 4004 -115 4005 -85
rect 4005 -115 4035 -85
rect 4035 -115 4036 -85
rect 4004 -116 4036 -115
rect 4084 875 4116 876
rect 4084 845 4085 875
rect 4085 845 4115 875
rect 4115 845 4116 875
rect 4084 844 4116 845
rect 4084 764 4116 796
rect 4084 715 4116 716
rect 4084 685 4085 715
rect 4085 685 4115 715
rect 4115 685 4116 715
rect 4084 684 4116 685
rect 4084 604 4116 636
rect 4084 555 4116 556
rect 4084 525 4085 555
rect 4085 525 4115 555
rect 4115 525 4116 555
rect 4084 524 4116 525
rect 4084 444 4116 476
rect 4084 395 4116 396
rect 4084 365 4085 395
rect 4085 365 4115 395
rect 4115 365 4116 395
rect 4084 364 4116 365
rect 4084 284 4116 316
rect 4084 235 4116 236
rect 4084 205 4085 235
rect 4085 205 4115 235
rect 4115 205 4116 235
rect 4084 204 4116 205
rect 4084 155 4116 156
rect 4084 125 4085 155
rect 4085 125 4115 155
rect 4115 125 4116 155
rect 4084 124 4116 125
rect 4084 75 4116 76
rect 4084 45 4085 75
rect 4085 45 4115 75
rect 4115 45 4116 75
rect 4084 44 4116 45
rect 4084 -5 4116 -4
rect 4084 -35 4085 -5
rect 4085 -35 4115 -5
rect 4115 -35 4116 -5
rect 4084 -36 4116 -35
rect 4084 -85 4116 -84
rect 4084 -115 4085 -85
rect 4085 -115 4115 -85
rect 4115 -115 4116 -85
rect 4084 -116 4116 -115
rect 4164 875 4196 876
rect 4164 845 4165 875
rect 4165 845 4195 875
rect 4195 845 4196 875
rect 4164 844 4196 845
rect 4164 764 4196 796
rect 4164 715 4196 716
rect 4164 685 4165 715
rect 4165 685 4195 715
rect 4195 685 4196 715
rect 4164 684 4196 685
rect 4164 604 4196 636
rect 4164 555 4196 556
rect 4164 525 4165 555
rect 4165 525 4195 555
rect 4195 525 4196 555
rect 4164 524 4196 525
rect 4164 444 4196 476
rect 4164 395 4196 396
rect 4164 365 4165 395
rect 4165 365 4195 395
rect 4195 365 4196 395
rect 4164 364 4196 365
rect 4164 284 4196 316
rect 4164 235 4196 236
rect 4164 205 4165 235
rect 4165 205 4195 235
rect 4195 205 4196 235
rect 4164 204 4196 205
rect 4164 155 4196 156
rect 4164 125 4165 155
rect 4165 125 4195 155
rect 4195 125 4196 155
rect 4164 124 4196 125
rect 4164 75 4196 76
rect 4164 45 4165 75
rect 4165 45 4195 75
rect 4195 45 4196 75
rect 4164 44 4196 45
rect 4164 -5 4196 -4
rect 4164 -35 4165 -5
rect 4165 -35 4195 -5
rect 4195 -35 4196 -5
rect 4164 -36 4196 -35
rect 4164 -85 4196 -84
rect 4164 -115 4165 -85
rect 4165 -115 4195 -85
rect 4195 -115 4196 -85
rect 4164 -116 4196 -115
rect 4244 875 4276 876
rect 4244 845 4245 875
rect 4245 845 4275 875
rect 4275 845 4276 875
rect 4244 844 4276 845
rect 4244 764 4276 796
rect 4244 715 4276 716
rect 4244 685 4245 715
rect 4245 685 4275 715
rect 4275 685 4276 715
rect 4244 684 4276 685
rect 4244 604 4276 636
rect 4244 555 4276 556
rect 4244 525 4245 555
rect 4245 525 4275 555
rect 4275 525 4276 555
rect 4244 524 4276 525
rect 4244 444 4276 476
rect 4244 395 4276 396
rect 4244 365 4245 395
rect 4245 365 4275 395
rect 4275 365 4276 395
rect 4244 364 4276 365
rect 4244 284 4276 316
rect 4244 235 4276 236
rect 4244 205 4245 235
rect 4245 205 4275 235
rect 4275 205 4276 235
rect 4244 204 4276 205
rect 4244 155 4276 156
rect 4244 125 4245 155
rect 4245 125 4275 155
rect 4275 125 4276 155
rect 4244 124 4276 125
rect 4244 75 4276 76
rect 4244 45 4245 75
rect 4245 45 4275 75
rect 4275 45 4276 75
rect 4244 44 4276 45
rect 4244 -5 4276 -4
rect 4244 -35 4245 -5
rect 4245 -35 4275 -5
rect 4275 -35 4276 -5
rect 4244 -36 4276 -35
rect 4244 -85 4276 -84
rect 4244 -115 4245 -85
rect 4245 -115 4275 -85
rect 4275 -115 4276 -85
rect 4244 -116 4276 -115
rect 4324 875 4356 876
rect 4324 845 4325 875
rect 4325 845 4355 875
rect 4355 845 4356 875
rect 4324 844 4356 845
rect 4324 764 4356 796
rect 4324 715 4356 716
rect 4324 685 4325 715
rect 4325 685 4355 715
rect 4355 685 4356 715
rect 4324 684 4356 685
rect 4324 604 4356 636
rect 4324 555 4356 556
rect 4324 525 4325 555
rect 4325 525 4355 555
rect 4355 525 4356 555
rect 4324 524 4356 525
rect 4324 444 4356 476
rect 4324 395 4356 396
rect 4324 365 4325 395
rect 4325 365 4355 395
rect 4355 365 4356 395
rect 4324 364 4356 365
rect 4324 284 4356 316
rect 4324 235 4356 236
rect 4324 205 4325 235
rect 4325 205 4355 235
rect 4355 205 4356 235
rect 4324 204 4356 205
rect 4324 155 4356 156
rect 4324 125 4325 155
rect 4325 125 4355 155
rect 4355 125 4356 155
rect 4324 124 4356 125
rect 4324 75 4356 76
rect 4324 45 4325 75
rect 4325 45 4355 75
rect 4355 45 4356 75
rect 4324 44 4356 45
rect 4324 -5 4356 -4
rect 4324 -35 4325 -5
rect 4325 -35 4355 -5
rect 4355 -35 4356 -5
rect 4324 -36 4356 -35
rect 4324 -85 4356 -84
rect 4324 -115 4325 -85
rect 4325 -115 4355 -85
rect 4355 -115 4356 -85
rect 4324 -116 4356 -115
rect 4404 875 4436 876
rect 4404 845 4405 875
rect 4405 845 4435 875
rect 4435 845 4436 875
rect 4404 844 4436 845
rect 4404 764 4436 796
rect 4404 715 4436 716
rect 4404 685 4405 715
rect 4405 685 4435 715
rect 4435 685 4436 715
rect 4404 684 4436 685
rect 4404 604 4436 636
rect 4404 555 4436 556
rect 4404 525 4405 555
rect 4405 525 4435 555
rect 4435 525 4436 555
rect 4404 524 4436 525
rect 4404 444 4436 476
rect 4404 395 4436 396
rect 4404 365 4405 395
rect 4405 365 4435 395
rect 4435 365 4436 395
rect 4404 364 4436 365
rect 4404 284 4436 316
rect 4404 235 4436 236
rect 4404 205 4405 235
rect 4405 205 4435 235
rect 4435 205 4436 235
rect 4404 204 4436 205
rect 4404 155 4436 156
rect 4404 125 4405 155
rect 4405 125 4435 155
rect 4435 125 4436 155
rect 4404 124 4436 125
rect 4404 75 4436 76
rect 4404 45 4405 75
rect 4405 45 4435 75
rect 4435 45 4436 75
rect 4404 44 4436 45
rect 4404 -5 4436 -4
rect 4404 -35 4405 -5
rect 4405 -35 4435 -5
rect 4435 -35 4436 -5
rect 4404 -36 4436 -35
rect 4404 -85 4436 -84
rect 4404 -115 4405 -85
rect 4405 -115 4435 -85
rect 4435 -115 4436 -85
rect 4404 -116 4436 -115
rect 4484 875 4516 876
rect 4484 845 4485 875
rect 4485 845 4515 875
rect 4515 845 4516 875
rect 4484 844 4516 845
rect 4484 764 4516 796
rect 4484 715 4516 716
rect 4484 685 4485 715
rect 4485 685 4515 715
rect 4515 685 4516 715
rect 4484 684 4516 685
rect 4484 604 4516 636
rect 4484 555 4516 556
rect 4484 525 4485 555
rect 4485 525 4515 555
rect 4515 525 4516 555
rect 4484 524 4516 525
rect 4484 444 4516 476
rect 4484 395 4516 396
rect 4484 365 4485 395
rect 4485 365 4515 395
rect 4515 365 4516 395
rect 4484 364 4516 365
rect 4484 284 4516 316
rect 4484 235 4516 236
rect 4484 205 4485 235
rect 4485 205 4515 235
rect 4515 205 4516 235
rect 4484 204 4516 205
rect 4484 155 4516 156
rect 4484 125 4485 155
rect 4485 125 4515 155
rect 4515 125 4516 155
rect 4484 124 4516 125
rect 4484 75 4516 76
rect 4484 45 4485 75
rect 4485 45 4515 75
rect 4515 45 4516 75
rect 4484 44 4516 45
rect 4484 -5 4516 -4
rect 4484 -35 4485 -5
rect 4485 -35 4515 -5
rect 4515 -35 4516 -5
rect 4484 -36 4516 -35
rect 4484 -85 4516 -84
rect 4484 -115 4485 -85
rect 4485 -115 4515 -85
rect 4515 -115 4516 -85
rect 4484 -116 4516 -115
rect 4564 875 4596 876
rect 4564 845 4565 875
rect 4565 845 4595 875
rect 4595 845 4596 875
rect 4564 844 4596 845
rect 4564 764 4596 796
rect 4564 715 4596 716
rect 4564 685 4565 715
rect 4565 685 4595 715
rect 4595 685 4596 715
rect 4564 684 4596 685
rect 4564 604 4596 636
rect 4564 555 4596 556
rect 4564 525 4565 555
rect 4565 525 4595 555
rect 4595 525 4596 555
rect 4564 524 4596 525
rect 4564 444 4596 476
rect 4564 395 4596 396
rect 4564 365 4565 395
rect 4565 365 4595 395
rect 4595 365 4596 395
rect 4564 364 4596 365
rect 4564 284 4596 316
rect 4564 235 4596 236
rect 4564 205 4565 235
rect 4565 205 4595 235
rect 4595 205 4596 235
rect 4564 204 4596 205
rect 4564 155 4596 156
rect 4564 125 4565 155
rect 4565 125 4595 155
rect 4595 125 4596 155
rect 4564 124 4596 125
rect 4564 75 4596 76
rect 4564 45 4565 75
rect 4565 45 4595 75
rect 4595 45 4596 75
rect 4564 44 4596 45
rect 4564 -5 4596 -4
rect 4564 -35 4565 -5
rect 4565 -35 4595 -5
rect 4595 -35 4596 -5
rect 4564 -36 4596 -35
rect 4564 -85 4596 -84
rect 4564 -115 4565 -85
rect 4565 -115 4595 -85
rect 4595 -115 4596 -85
rect 4564 -116 4596 -115
rect 4644 875 4676 876
rect 4644 845 4645 875
rect 4645 845 4675 875
rect 4675 845 4676 875
rect 4644 844 4676 845
rect 4644 764 4676 796
rect 4644 715 4676 716
rect 4644 685 4645 715
rect 4645 685 4675 715
rect 4675 685 4676 715
rect 4644 684 4676 685
rect 4644 604 4676 636
rect 4644 555 4676 556
rect 4644 525 4645 555
rect 4645 525 4675 555
rect 4675 525 4676 555
rect 4644 524 4676 525
rect 4644 444 4676 476
rect 4644 395 4676 396
rect 4644 365 4645 395
rect 4645 365 4675 395
rect 4675 365 4676 395
rect 4644 364 4676 365
rect 4644 284 4676 316
rect 4644 235 4676 236
rect 4644 205 4645 235
rect 4645 205 4675 235
rect 4675 205 4676 235
rect 4644 204 4676 205
rect 4644 155 4676 156
rect 4644 125 4645 155
rect 4645 125 4675 155
rect 4675 125 4676 155
rect 4644 124 4676 125
rect 4644 75 4676 76
rect 4644 45 4645 75
rect 4645 45 4675 75
rect 4675 45 4676 75
rect 4644 44 4676 45
rect 4644 -5 4676 -4
rect 4644 -35 4645 -5
rect 4645 -35 4675 -5
rect 4675 -35 4676 -5
rect 4644 -36 4676 -35
rect 4644 -85 4676 -84
rect 4644 -115 4645 -85
rect 4645 -115 4675 -85
rect 4675 -115 4676 -85
rect 4644 -116 4676 -115
rect 4724 875 4756 876
rect 4724 845 4725 875
rect 4725 845 4755 875
rect 4755 845 4756 875
rect 4724 844 4756 845
rect 4724 764 4756 796
rect 4724 715 4756 716
rect 4724 685 4725 715
rect 4725 685 4755 715
rect 4755 685 4756 715
rect 4724 684 4756 685
rect 4724 604 4756 636
rect 4724 555 4756 556
rect 4724 525 4725 555
rect 4725 525 4755 555
rect 4755 525 4756 555
rect 4724 524 4756 525
rect 4724 444 4756 476
rect 4724 395 4756 396
rect 4724 365 4725 395
rect 4725 365 4755 395
rect 4755 365 4756 395
rect 4724 364 4756 365
rect 4724 284 4756 316
rect 4724 235 4756 236
rect 4724 205 4725 235
rect 4725 205 4755 235
rect 4755 205 4756 235
rect 4724 204 4756 205
rect 4724 155 4756 156
rect 4724 125 4725 155
rect 4725 125 4755 155
rect 4755 125 4756 155
rect 4724 124 4756 125
rect 4724 75 4756 76
rect 4724 45 4725 75
rect 4725 45 4755 75
rect 4755 45 4756 75
rect 4724 44 4756 45
rect 4724 -5 4756 -4
rect 4724 -35 4725 -5
rect 4725 -35 4755 -5
rect 4755 -35 4756 -5
rect 4724 -36 4756 -35
rect 4724 -85 4756 -84
rect 4724 -115 4725 -85
rect 4725 -115 4755 -85
rect 4755 -115 4756 -85
rect 4724 -116 4756 -115
rect 4804 875 4836 876
rect 4804 845 4805 875
rect 4805 845 4835 875
rect 4835 845 4836 875
rect 4804 844 4836 845
rect 4804 764 4836 796
rect 4804 715 4836 716
rect 4804 685 4805 715
rect 4805 685 4835 715
rect 4835 685 4836 715
rect 4804 684 4836 685
rect 4804 604 4836 636
rect 4804 555 4836 556
rect 4804 525 4805 555
rect 4805 525 4835 555
rect 4835 525 4836 555
rect 4804 524 4836 525
rect 4804 444 4836 476
rect 4804 395 4836 396
rect 4804 365 4805 395
rect 4805 365 4835 395
rect 4835 365 4836 395
rect 4804 364 4836 365
rect 4804 284 4836 316
rect 4804 235 4836 236
rect 4804 205 4805 235
rect 4805 205 4835 235
rect 4835 205 4836 235
rect 4804 204 4836 205
rect 4804 155 4836 156
rect 4804 125 4805 155
rect 4805 125 4835 155
rect 4835 125 4836 155
rect 4804 124 4836 125
rect 4804 75 4836 76
rect 4804 45 4805 75
rect 4805 45 4835 75
rect 4835 45 4836 75
rect 4804 44 4836 45
rect 4804 -5 4836 -4
rect 4804 -35 4805 -5
rect 4805 -35 4835 -5
rect 4835 -35 4836 -5
rect 4804 -36 4836 -35
rect 4804 -85 4836 -84
rect 4804 -115 4805 -85
rect 4805 -115 4835 -85
rect 4835 -115 4836 -85
rect 4804 -116 4836 -115
rect 4884 875 4916 876
rect 4884 845 4885 875
rect 4885 845 4915 875
rect 4915 845 4916 875
rect 4884 844 4916 845
rect 4884 764 4916 796
rect 4884 715 4916 716
rect 4884 685 4885 715
rect 4885 685 4915 715
rect 4915 685 4916 715
rect 4884 684 4916 685
rect 4884 604 4916 636
rect 4884 555 4916 556
rect 4884 525 4885 555
rect 4885 525 4915 555
rect 4915 525 4916 555
rect 4884 524 4916 525
rect 4884 444 4916 476
rect 4884 395 4916 396
rect 4884 365 4885 395
rect 4885 365 4915 395
rect 4915 365 4916 395
rect 4884 364 4916 365
rect 4884 284 4916 316
rect 4884 235 4916 236
rect 4884 205 4885 235
rect 4885 205 4915 235
rect 4915 205 4916 235
rect 4884 204 4916 205
rect 4884 155 4916 156
rect 4884 125 4885 155
rect 4885 125 4915 155
rect 4915 125 4916 155
rect 4884 124 4916 125
rect 4884 75 4916 76
rect 4884 45 4885 75
rect 4885 45 4915 75
rect 4915 45 4916 75
rect 4884 44 4916 45
rect 4884 -5 4916 -4
rect 4884 -35 4885 -5
rect 4885 -35 4915 -5
rect 4915 -35 4916 -5
rect 4884 -36 4916 -35
rect 4884 -85 4916 -84
rect 4884 -115 4885 -85
rect 4885 -115 4915 -85
rect 4915 -115 4916 -85
rect 4884 -116 4916 -115
rect 5044 5595 5076 5596
rect 5044 5565 5045 5595
rect 5045 5565 5075 5595
rect 5075 5565 5076 5595
rect 5044 5564 5076 5565
rect 5044 5515 5076 5516
rect 5044 5485 5045 5515
rect 5045 5485 5075 5515
rect 5075 5485 5076 5515
rect 5044 5484 5076 5485
rect 5044 5435 5076 5436
rect 5044 5405 5045 5435
rect 5045 5405 5075 5435
rect 5075 5405 5076 5435
rect 5044 5404 5076 5405
rect 5044 5355 5076 5356
rect 5044 5325 5045 5355
rect 5045 5325 5075 5355
rect 5075 5325 5076 5355
rect 5044 5324 5076 5325
rect 5044 5275 5076 5276
rect 5044 5245 5045 5275
rect 5045 5245 5075 5275
rect 5075 5245 5076 5275
rect 5044 5244 5076 5245
rect 5044 5195 5076 5196
rect 5044 5165 5045 5195
rect 5045 5165 5075 5195
rect 5075 5165 5076 5195
rect 5044 5164 5076 5165
rect 5044 5115 5076 5116
rect 5044 5085 5045 5115
rect 5045 5085 5075 5115
rect 5075 5085 5076 5115
rect 5044 5084 5076 5085
rect 5044 5035 5076 5036
rect 5044 5005 5045 5035
rect 5045 5005 5075 5035
rect 5075 5005 5076 5035
rect 5044 5004 5076 5005
rect 5044 4955 5076 4956
rect 5044 4925 5045 4955
rect 5045 4925 5075 4955
rect 5075 4925 5076 4955
rect 5044 4924 5076 4925
rect 5044 4875 5076 4876
rect 5044 4845 5045 4875
rect 5045 4845 5075 4875
rect 5075 4845 5076 4875
rect 5044 4844 5076 4845
rect 5044 4795 5076 4796
rect 5044 4765 5045 4795
rect 5045 4765 5075 4795
rect 5075 4765 5076 4795
rect 5044 4764 5076 4765
rect 5044 4715 5076 4716
rect 5044 4685 5045 4715
rect 5045 4685 5075 4715
rect 5075 4685 5076 4715
rect 5044 4684 5076 4685
rect 5044 4635 5076 4636
rect 5044 4605 5045 4635
rect 5045 4605 5075 4635
rect 5075 4605 5076 4635
rect 5044 4604 5076 4605
rect 5044 4555 5076 4556
rect 5044 4525 5045 4555
rect 5045 4525 5075 4555
rect 5075 4525 5076 4555
rect 5044 4524 5076 4525
rect 5044 4475 5076 4476
rect 5044 4445 5045 4475
rect 5045 4445 5075 4475
rect 5075 4445 5076 4475
rect 5044 4444 5076 4445
rect 5044 4395 5076 4396
rect 5044 4365 5045 4395
rect 5045 4365 5075 4395
rect 5075 4365 5076 4395
rect 5044 4364 5076 4365
rect 5044 4284 5076 4316
rect 5044 4235 5076 4236
rect 5044 4205 5045 4235
rect 5045 4205 5075 4235
rect 5075 4205 5076 4235
rect 5044 4204 5076 4205
rect 5044 4155 5076 4156
rect 5044 4125 5045 4155
rect 5045 4125 5075 4155
rect 5075 4125 5076 4155
rect 5044 4124 5076 4125
rect 5044 4075 5076 4076
rect 5044 4045 5045 4075
rect 5045 4045 5075 4075
rect 5075 4045 5076 4075
rect 5044 4044 5076 4045
rect 5044 3995 5076 3996
rect 5044 3965 5045 3995
rect 5045 3965 5075 3995
rect 5075 3965 5076 3995
rect 5044 3964 5076 3965
rect 5044 3915 5076 3916
rect 5044 3885 5045 3915
rect 5045 3885 5075 3915
rect 5075 3885 5076 3915
rect 5044 3884 5076 3885
rect 5044 3835 5076 3836
rect 5044 3805 5045 3835
rect 5045 3805 5075 3835
rect 5075 3805 5076 3835
rect 5044 3804 5076 3805
rect 5044 3755 5076 3756
rect 5044 3725 5045 3755
rect 5045 3725 5075 3755
rect 5075 3725 5076 3755
rect 5044 3724 5076 3725
rect 5044 3675 5076 3676
rect 5044 3645 5045 3675
rect 5045 3645 5075 3675
rect 5075 3645 5076 3675
rect 5044 3644 5076 3645
rect 5044 3595 5076 3596
rect 5044 3565 5045 3595
rect 5045 3565 5075 3595
rect 5075 3565 5076 3595
rect 5044 3564 5076 3565
rect 5044 3515 5076 3516
rect 5044 3485 5045 3515
rect 5045 3485 5075 3515
rect 5075 3485 5076 3515
rect 5044 3484 5076 3485
rect 5044 3435 5076 3436
rect 5044 3405 5045 3435
rect 5045 3405 5075 3435
rect 5075 3405 5076 3435
rect 5044 3404 5076 3405
rect 5044 3355 5076 3356
rect 5044 3325 5045 3355
rect 5045 3325 5075 3355
rect 5075 3325 5076 3355
rect 5044 3324 5076 3325
rect 5044 3275 5076 3276
rect 5044 3245 5045 3275
rect 5045 3245 5075 3275
rect 5075 3245 5076 3275
rect 5044 3244 5076 3245
rect 5044 3195 5076 3196
rect 5044 3165 5045 3195
rect 5045 3165 5075 3195
rect 5075 3165 5076 3195
rect 5044 3164 5076 3165
rect 5044 3115 5076 3116
rect 5044 3085 5045 3115
rect 5045 3085 5075 3115
rect 5075 3085 5076 3115
rect 5044 3084 5076 3085
rect 5044 3035 5076 3036
rect 5044 3005 5045 3035
rect 5045 3005 5075 3035
rect 5075 3005 5076 3035
rect 5044 3004 5076 3005
rect 5044 2955 5076 2956
rect 5044 2925 5045 2955
rect 5045 2925 5075 2955
rect 5075 2925 5076 2955
rect 5044 2924 5076 2925
rect 5044 2875 5076 2876
rect 5044 2845 5045 2875
rect 5045 2845 5075 2875
rect 5075 2845 5076 2875
rect 5044 2844 5076 2845
rect 5044 2795 5076 2796
rect 5044 2765 5045 2795
rect 5045 2765 5075 2795
rect 5075 2765 5076 2795
rect 5044 2764 5076 2765
rect 5044 2715 5076 2716
rect 5044 2685 5045 2715
rect 5045 2685 5075 2715
rect 5075 2685 5076 2715
rect 5044 2684 5076 2685
rect 5044 2635 5076 2636
rect 5044 2605 5045 2635
rect 5045 2605 5075 2635
rect 5075 2605 5076 2635
rect 5044 2604 5076 2605
rect 5044 2555 5076 2556
rect 5044 2525 5045 2555
rect 5045 2525 5075 2555
rect 5075 2525 5076 2555
rect 5044 2524 5076 2525
rect 5044 2475 5076 2476
rect 5044 2445 5045 2475
rect 5045 2445 5075 2475
rect 5075 2445 5076 2475
rect 5044 2444 5076 2445
rect 5044 2364 5076 2396
rect 5044 2315 5076 2316
rect 5044 2285 5045 2315
rect 5045 2285 5075 2315
rect 5075 2285 5076 2315
rect 5044 2284 5076 2285
rect 5044 2235 5076 2236
rect 5044 2205 5045 2235
rect 5045 2205 5075 2235
rect 5075 2205 5076 2235
rect 5044 2204 5076 2205
rect 5044 2155 5076 2156
rect 5044 2125 5045 2155
rect 5045 2125 5075 2155
rect 5075 2125 5076 2155
rect 5044 2124 5076 2125
rect 5044 2075 5076 2076
rect 5044 2045 5045 2075
rect 5045 2045 5075 2075
rect 5075 2045 5076 2075
rect 5044 2044 5076 2045
rect 5044 1995 5076 1996
rect 5044 1965 5045 1995
rect 5045 1965 5075 1995
rect 5075 1965 5076 1995
rect 5044 1964 5076 1965
rect 5044 1915 5076 1916
rect 5044 1885 5045 1915
rect 5045 1885 5075 1915
rect 5075 1885 5076 1915
rect 5044 1884 5076 1885
rect 5044 1835 5076 1836
rect 5044 1805 5045 1835
rect 5045 1805 5075 1835
rect 5075 1805 5076 1835
rect 5044 1804 5076 1805
rect 5044 1755 5076 1756
rect 5044 1725 5045 1755
rect 5045 1725 5075 1755
rect 5075 1725 5076 1755
rect 5044 1724 5076 1725
rect 5044 1675 5076 1676
rect 5044 1645 5045 1675
rect 5045 1645 5075 1675
rect 5075 1645 5076 1675
rect 5044 1644 5076 1645
rect 5044 1595 5076 1596
rect 5044 1565 5045 1595
rect 5045 1565 5075 1595
rect 5075 1565 5076 1595
rect 5044 1564 5076 1565
rect 5044 1515 5076 1516
rect 5044 1485 5045 1515
rect 5045 1485 5075 1515
rect 5075 1485 5076 1515
rect 5044 1484 5076 1485
rect 5044 1435 5076 1436
rect 5044 1405 5045 1435
rect 5045 1405 5075 1435
rect 5075 1405 5076 1435
rect 5044 1404 5076 1405
rect 5044 1355 5076 1356
rect 5044 1325 5045 1355
rect 5045 1325 5075 1355
rect 5075 1325 5076 1355
rect 5044 1324 5076 1325
rect 5044 1275 5076 1276
rect 5044 1245 5045 1275
rect 5045 1245 5075 1275
rect 5075 1245 5076 1275
rect 5044 1244 5076 1245
rect 5044 1195 5076 1196
rect 5044 1165 5045 1195
rect 5045 1165 5075 1195
rect 5075 1165 5076 1195
rect 5044 1164 5076 1165
rect 5044 1115 5076 1116
rect 5044 1085 5045 1115
rect 5045 1085 5075 1115
rect 5075 1085 5076 1115
rect 5044 1084 5076 1085
rect 5044 1035 5076 1036
rect 5044 1005 5045 1035
rect 5045 1005 5075 1035
rect 5075 1005 5076 1035
rect 5044 1004 5076 1005
rect 5044 955 5076 956
rect 5044 925 5045 955
rect 5045 925 5075 955
rect 5075 925 5076 955
rect 5044 924 5076 925
rect 5044 875 5076 876
rect 5044 845 5045 875
rect 5045 845 5075 875
rect 5075 845 5076 875
rect 5044 844 5076 845
rect 5044 764 5076 796
rect 5044 715 5076 716
rect 5044 685 5045 715
rect 5045 685 5075 715
rect 5075 685 5076 715
rect 5044 684 5076 685
rect 5044 604 5076 636
rect 5044 555 5076 556
rect 5044 525 5045 555
rect 5045 525 5075 555
rect 5075 525 5076 555
rect 5044 524 5076 525
rect 5044 444 5076 476
rect 5044 395 5076 396
rect 5044 365 5045 395
rect 5045 365 5075 395
rect 5075 365 5076 395
rect 5044 364 5076 365
rect 5044 315 5076 316
rect 5044 285 5045 315
rect 5045 285 5075 315
rect 5075 285 5076 315
rect 5044 284 5076 285
rect 5044 235 5076 236
rect 5044 205 5045 235
rect 5045 205 5075 235
rect 5075 205 5076 235
rect 5044 204 5076 205
rect 5044 155 5076 156
rect 5044 125 5045 155
rect 5045 125 5075 155
rect 5075 125 5076 155
rect 5044 124 5076 125
rect 5044 75 5076 76
rect 5044 45 5045 75
rect 5045 45 5075 75
rect 5075 45 5076 75
rect 5044 44 5076 45
rect 5044 -5 5076 -4
rect 5044 -35 5045 -5
rect 5045 -35 5075 -5
rect 5075 -35 5076 -5
rect 5044 -36 5076 -35
rect 5044 -85 5076 -84
rect 5044 -115 5045 -85
rect 5045 -115 5075 -85
rect 5075 -115 5076 -85
rect 5044 -116 5076 -115
rect 5204 5595 5236 5596
rect 5204 5565 5205 5595
rect 5205 5565 5235 5595
rect 5235 5565 5236 5595
rect 5204 5564 5236 5565
rect 5204 5515 5236 5516
rect 5204 5485 5205 5515
rect 5205 5485 5235 5515
rect 5235 5485 5236 5515
rect 5204 5484 5236 5485
rect 5204 5435 5236 5436
rect 5204 5405 5205 5435
rect 5205 5405 5235 5435
rect 5235 5405 5236 5435
rect 5204 5404 5236 5405
rect 5204 5355 5236 5356
rect 5204 5325 5205 5355
rect 5205 5325 5235 5355
rect 5235 5325 5236 5355
rect 5204 5324 5236 5325
rect 5204 5275 5236 5276
rect 5204 5245 5205 5275
rect 5205 5245 5235 5275
rect 5235 5245 5236 5275
rect 5204 5244 5236 5245
rect 5204 5195 5236 5196
rect 5204 5165 5205 5195
rect 5205 5165 5235 5195
rect 5235 5165 5236 5195
rect 5204 5164 5236 5165
rect 5204 5115 5236 5116
rect 5204 5085 5205 5115
rect 5205 5085 5235 5115
rect 5235 5085 5236 5115
rect 5204 5084 5236 5085
rect 5204 5035 5236 5036
rect 5204 5005 5205 5035
rect 5205 5005 5235 5035
rect 5235 5005 5236 5035
rect 5204 5004 5236 5005
rect 5204 4955 5236 4956
rect 5204 4925 5205 4955
rect 5205 4925 5235 4955
rect 5235 4925 5236 4955
rect 5204 4924 5236 4925
rect 5204 4875 5236 4876
rect 5204 4845 5205 4875
rect 5205 4845 5235 4875
rect 5235 4845 5236 4875
rect 5204 4844 5236 4845
rect 5204 4795 5236 4796
rect 5204 4765 5205 4795
rect 5205 4765 5235 4795
rect 5235 4765 5236 4795
rect 5204 4764 5236 4765
rect 5204 4715 5236 4716
rect 5204 4685 5205 4715
rect 5205 4685 5235 4715
rect 5235 4685 5236 4715
rect 5204 4684 5236 4685
rect 5204 4635 5236 4636
rect 5204 4605 5205 4635
rect 5205 4605 5235 4635
rect 5235 4605 5236 4635
rect 5204 4604 5236 4605
rect 5204 4555 5236 4556
rect 5204 4525 5205 4555
rect 5205 4525 5235 4555
rect 5235 4525 5236 4555
rect 5204 4524 5236 4525
rect 5204 4475 5236 4476
rect 5204 4445 5205 4475
rect 5205 4445 5235 4475
rect 5235 4445 5236 4475
rect 5204 4444 5236 4445
rect 5204 4395 5236 4396
rect 5204 4365 5205 4395
rect 5205 4365 5235 4395
rect 5235 4365 5236 4395
rect 5204 4364 5236 4365
rect 5204 4284 5236 4316
rect 5204 4235 5236 4236
rect 5204 4205 5205 4235
rect 5205 4205 5235 4235
rect 5235 4205 5236 4235
rect 5204 4204 5236 4205
rect 5204 4155 5236 4156
rect 5204 4125 5205 4155
rect 5205 4125 5235 4155
rect 5235 4125 5236 4155
rect 5204 4124 5236 4125
rect 5204 4075 5236 4076
rect 5204 4045 5205 4075
rect 5205 4045 5235 4075
rect 5235 4045 5236 4075
rect 5204 4044 5236 4045
rect 5204 3995 5236 3996
rect 5204 3965 5205 3995
rect 5205 3965 5235 3995
rect 5235 3965 5236 3995
rect 5204 3964 5236 3965
rect 5204 3915 5236 3916
rect 5204 3885 5205 3915
rect 5205 3885 5235 3915
rect 5235 3885 5236 3915
rect 5204 3884 5236 3885
rect 5204 3835 5236 3836
rect 5204 3805 5205 3835
rect 5205 3805 5235 3835
rect 5235 3805 5236 3835
rect 5204 3804 5236 3805
rect 5204 3755 5236 3756
rect 5204 3725 5205 3755
rect 5205 3725 5235 3755
rect 5235 3725 5236 3755
rect 5204 3724 5236 3725
rect 5204 3675 5236 3676
rect 5204 3645 5205 3675
rect 5205 3645 5235 3675
rect 5235 3645 5236 3675
rect 5204 3644 5236 3645
rect 5204 3595 5236 3596
rect 5204 3565 5205 3595
rect 5205 3565 5235 3595
rect 5235 3565 5236 3595
rect 5204 3564 5236 3565
rect 5204 3515 5236 3516
rect 5204 3485 5205 3515
rect 5205 3485 5235 3515
rect 5235 3485 5236 3515
rect 5204 3484 5236 3485
rect 5204 3435 5236 3436
rect 5204 3405 5205 3435
rect 5205 3405 5235 3435
rect 5235 3405 5236 3435
rect 5204 3404 5236 3405
rect 5204 3355 5236 3356
rect 5204 3325 5205 3355
rect 5205 3325 5235 3355
rect 5235 3325 5236 3355
rect 5204 3324 5236 3325
rect 5204 3275 5236 3276
rect 5204 3245 5205 3275
rect 5205 3245 5235 3275
rect 5235 3245 5236 3275
rect 5204 3244 5236 3245
rect 5204 3195 5236 3196
rect 5204 3165 5205 3195
rect 5205 3165 5235 3195
rect 5235 3165 5236 3195
rect 5204 3164 5236 3165
rect 5204 3115 5236 3116
rect 5204 3085 5205 3115
rect 5205 3085 5235 3115
rect 5235 3085 5236 3115
rect 5204 3084 5236 3085
rect 5204 3035 5236 3036
rect 5204 3005 5205 3035
rect 5205 3005 5235 3035
rect 5235 3005 5236 3035
rect 5204 3004 5236 3005
rect 5204 2955 5236 2956
rect 5204 2925 5205 2955
rect 5205 2925 5235 2955
rect 5235 2925 5236 2955
rect 5204 2924 5236 2925
rect 5204 2875 5236 2876
rect 5204 2845 5205 2875
rect 5205 2845 5235 2875
rect 5235 2845 5236 2875
rect 5204 2844 5236 2845
rect 5204 2795 5236 2796
rect 5204 2765 5205 2795
rect 5205 2765 5235 2795
rect 5235 2765 5236 2795
rect 5204 2764 5236 2765
rect 5204 2715 5236 2716
rect 5204 2685 5205 2715
rect 5205 2685 5235 2715
rect 5235 2685 5236 2715
rect 5204 2684 5236 2685
rect 5204 2635 5236 2636
rect 5204 2605 5205 2635
rect 5205 2605 5235 2635
rect 5235 2605 5236 2635
rect 5204 2604 5236 2605
rect 5204 2555 5236 2556
rect 5204 2525 5205 2555
rect 5205 2525 5235 2555
rect 5235 2525 5236 2555
rect 5204 2524 5236 2525
rect 5204 2475 5236 2476
rect 5204 2445 5205 2475
rect 5205 2445 5235 2475
rect 5235 2445 5236 2475
rect 5204 2444 5236 2445
rect 5204 2364 5236 2396
rect 5204 2315 5236 2316
rect 5204 2285 5205 2315
rect 5205 2285 5235 2315
rect 5235 2285 5236 2315
rect 5204 2284 5236 2285
rect 5204 2235 5236 2236
rect 5204 2205 5205 2235
rect 5205 2205 5235 2235
rect 5235 2205 5236 2235
rect 5204 2204 5236 2205
rect 5204 2155 5236 2156
rect 5204 2125 5205 2155
rect 5205 2125 5235 2155
rect 5235 2125 5236 2155
rect 5204 2124 5236 2125
rect 5204 2075 5236 2076
rect 5204 2045 5205 2075
rect 5205 2045 5235 2075
rect 5235 2045 5236 2075
rect 5204 2044 5236 2045
rect 5204 1995 5236 1996
rect 5204 1965 5205 1995
rect 5205 1965 5235 1995
rect 5235 1965 5236 1995
rect 5204 1964 5236 1965
rect 5204 1915 5236 1916
rect 5204 1885 5205 1915
rect 5205 1885 5235 1915
rect 5235 1885 5236 1915
rect 5204 1884 5236 1885
rect 5204 1835 5236 1836
rect 5204 1805 5205 1835
rect 5205 1805 5235 1835
rect 5235 1805 5236 1835
rect 5204 1804 5236 1805
rect 5204 1755 5236 1756
rect 5204 1725 5205 1755
rect 5205 1725 5235 1755
rect 5235 1725 5236 1755
rect 5204 1724 5236 1725
rect 5204 1675 5236 1676
rect 5204 1645 5205 1675
rect 5205 1645 5235 1675
rect 5235 1645 5236 1675
rect 5204 1644 5236 1645
rect 5204 1595 5236 1596
rect 5204 1565 5205 1595
rect 5205 1565 5235 1595
rect 5235 1565 5236 1595
rect 5204 1564 5236 1565
rect 5204 1515 5236 1516
rect 5204 1485 5205 1515
rect 5205 1485 5235 1515
rect 5235 1485 5236 1515
rect 5204 1484 5236 1485
rect 5204 1435 5236 1436
rect 5204 1405 5205 1435
rect 5205 1405 5235 1435
rect 5235 1405 5236 1435
rect 5204 1404 5236 1405
rect 5204 1355 5236 1356
rect 5204 1325 5205 1355
rect 5205 1325 5235 1355
rect 5235 1325 5236 1355
rect 5204 1324 5236 1325
rect 5204 1275 5236 1276
rect 5204 1245 5205 1275
rect 5205 1245 5235 1275
rect 5235 1245 5236 1275
rect 5204 1244 5236 1245
rect 5204 1195 5236 1196
rect 5204 1165 5205 1195
rect 5205 1165 5235 1195
rect 5235 1165 5236 1195
rect 5204 1164 5236 1165
rect 5204 1115 5236 1116
rect 5204 1085 5205 1115
rect 5205 1085 5235 1115
rect 5235 1085 5236 1115
rect 5204 1084 5236 1085
rect 5204 1035 5236 1036
rect 5204 1005 5205 1035
rect 5205 1005 5235 1035
rect 5235 1005 5236 1035
rect 5204 1004 5236 1005
rect 5204 955 5236 956
rect 5204 925 5205 955
rect 5205 925 5235 955
rect 5235 925 5236 955
rect 5204 924 5236 925
rect 5204 875 5236 876
rect 5204 845 5205 875
rect 5205 845 5235 875
rect 5235 845 5236 875
rect 5204 844 5236 845
rect 5204 764 5236 796
rect 5204 715 5236 716
rect 5204 685 5205 715
rect 5205 685 5235 715
rect 5235 685 5236 715
rect 5204 684 5236 685
rect 5204 604 5236 636
rect 5204 555 5236 556
rect 5204 525 5205 555
rect 5205 525 5235 555
rect 5235 525 5236 555
rect 5204 524 5236 525
rect 5204 475 5236 476
rect 5204 445 5205 475
rect 5205 445 5235 475
rect 5235 445 5236 475
rect 5204 444 5236 445
rect 5204 395 5236 396
rect 5204 365 5205 395
rect 5205 365 5235 395
rect 5235 365 5236 395
rect 5204 364 5236 365
rect 5204 315 5236 316
rect 5204 285 5205 315
rect 5205 285 5235 315
rect 5235 285 5236 315
rect 5204 284 5236 285
rect 5204 235 5236 236
rect 5204 205 5205 235
rect 5205 205 5235 235
rect 5235 205 5236 235
rect 5204 204 5236 205
rect 5204 155 5236 156
rect 5204 125 5205 155
rect 5205 125 5235 155
rect 5235 125 5236 155
rect 5204 124 5236 125
rect 5204 75 5236 76
rect 5204 45 5205 75
rect 5205 45 5235 75
rect 5235 45 5236 75
rect 5204 44 5236 45
rect 5204 -5 5236 -4
rect 5204 -35 5205 -5
rect 5205 -35 5235 -5
rect 5235 -35 5236 -5
rect 5204 -36 5236 -35
rect 5204 -85 5236 -84
rect 5204 -115 5205 -85
rect 5205 -115 5235 -85
rect 5235 -115 5236 -85
rect 5204 -116 5236 -115
rect 5364 5595 5396 5596
rect 5364 5565 5365 5595
rect 5365 5565 5395 5595
rect 5395 5565 5396 5595
rect 5364 5564 5396 5565
rect 5364 5515 5396 5516
rect 5364 5485 5365 5515
rect 5365 5485 5395 5515
rect 5395 5485 5396 5515
rect 5364 5484 5396 5485
rect 5364 5435 5396 5436
rect 5364 5405 5365 5435
rect 5365 5405 5395 5435
rect 5395 5405 5396 5435
rect 5364 5404 5396 5405
rect 5364 5355 5396 5356
rect 5364 5325 5365 5355
rect 5365 5325 5395 5355
rect 5395 5325 5396 5355
rect 5364 5324 5396 5325
rect 5364 5275 5396 5276
rect 5364 5245 5365 5275
rect 5365 5245 5395 5275
rect 5395 5245 5396 5275
rect 5364 5244 5396 5245
rect 5364 5195 5396 5196
rect 5364 5165 5365 5195
rect 5365 5165 5395 5195
rect 5395 5165 5396 5195
rect 5364 5164 5396 5165
rect 5364 5115 5396 5116
rect 5364 5085 5365 5115
rect 5365 5085 5395 5115
rect 5395 5085 5396 5115
rect 5364 5084 5396 5085
rect 5364 5035 5396 5036
rect 5364 5005 5365 5035
rect 5365 5005 5395 5035
rect 5395 5005 5396 5035
rect 5364 5004 5396 5005
rect 5364 4955 5396 4956
rect 5364 4925 5365 4955
rect 5365 4925 5395 4955
rect 5395 4925 5396 4955
rect 5364 4924 5396 4925
rect 5364 4875 5396 4876
rect 5364 4845 5365 4875
rect 5365 4845 5395 4875
rect 5395 4845 5396 4875
rect 5364 4844 5396 4845
rect 5364 4795 5396 4796
rect 5364 4765 5365 4795
rect 5365 4765 5395 4795
rect 5395 4765 5396 4795
rect 5364 4764 5396 4765
rect 5364 4715 5396 4716
rect 5364 4685 5365 4715
rect 5365 4685 5395 4715
rect 5395 4685 5396 4715
rect 5364 4684 5396 4685
rect 5364 4635 5396 4636
rect 5364 4605 5365 4635
rect 5365 4605 5395 4635
rect 5395 4605 5396 4635
rect 5364 4604 5396 4605
rect 5364 4555 5396 4556
rect 5364 4525 5365 4555
rect 5365 4525 5395 4555
rect 5395 4525 5396 4555
rect 5364 4524 5396 4525
rect 5364 4475 5396 4476
rect 5364 4445 5365 4475
rect 5365 4445 5395 4475
rect 5395 4445 5396 4475
rect 5364 4444 5396 4445
rect 5364 4395 5396 4396
rect 5364 4365 5365 4395
rect 5365 4365 5395 4395
rect 5395 4365 5396 4395
rect 5364 4364 5396 4365
rect 5364 4284 5396 4316
rect 5364 4235 5396 4236
rect 5364 4205 5365 4235
rect 5365 4205 5395 4235
rect 5395 4205 5396 4235
rect 5364 4204 5396 4205
rect 5364 4155 5396 4156
rect 5364 4125 5365 4155
rect 5365 4125 5395 4155
rect 5395 4125 5396 4155
rect 5364 4124 5396 4125
rect 5364 4075 5396 4076
rect 5364 4045 5365 4075
rect 5365 4045 5395 4075
rect 5395 4045 5396 4075
rect 5364 4044 5396 4045
rect 5364 3995 5396 3996
rect 5364 3965 5365 3995
rect 5365 3965 5395 3995
rect 5395 3965 5396 3995
rect 5364 3964 5396 3965
rect 5364 3915 5396 3916
rect 5364 3885 5365 3915
rect 5365 3885 5395 3915
rect 5395 3885 5396 3915
rect 5364 3884 5396 3885
rect 5364 3835 5396 3836
rect 5364 3805 5365 3835
rect 5365 3805 5395 3835
rect 5395 3805 5396 3835
rect 5364 3804 5396 3805
rect 5364 3755 5396 3756
rect 5364 3725 5365 3755
rect 5365 3725 5395 3755
rect 5395 3725 5396 3755
rect 5364 3724 5396 3725
rect 5364 3675 5396 3676
rect 5364 3645 5365 3675
rect 5365 3645 5395 3675
rect 5395 3645 5396 3675
rect 5364 3644 5396 3645
rect 5364 3595 5396 3596
rect 5364 3565 5365 3595
rect 5365 3565 5395 3595
rect 5395 3565 5396 3595
rect 5364 3564 5396 3565
rect 5364 3515 5396 3516
rect 5364 3485 5365 3515
rect 5365 3485 5395 3515
rect 5395 3485 5396 3515
rect 5364 3484 5396 3485
rect 5364 3435 5396 3436
rect 5364 3405 5365 3435
rect 5365 3405 5395 3435
rect 5395 3405 5396 3435
rect 5364 3404 5396 3405
rect 5364 3355 5396 3356
rect 5364 3325 5365 3355
rect 5365 3325 5395 3355
rect 5395 3325 5396 3355
rect 5364 3324 5396 3325
rect 5364 3275 5396 3276
rect 5364 3245 5365 3275
rect 5365 3245 5395 3275
rect 5395 3245 5396 3275
rect 5364 3244 5396 3245
rect 5364 3195 5396 3196
rect 5364 3165 5365 3195
rect 5365 3165 5395 3195
rect 5395 3165 5396 3195
rect 5364 3164 5396 3165
rect 5364 3115 5396 3116
rect 5364 3085 5365 3115
rect 5365 3085 5395 3115
rect 5395 3085 5396 3115
rect 5364 3084 5396 3085
rect 5364 3035 5396 3036
rect 5364 3005 5365 3035
rect 5365 3005 5395 3035
rect 5395 3005 5396 3035
rect 5364 3004 5396 3005
rect 5364 2955 5396 2956
rect 5364 2925 5365 2955
rect 5365 2925 5395 2955
rect 5395 2925 5396 2955
rect 5364 2924 5396 2925
rect 5364 2875 5396 2876
rect 5364 2845 5365 2875
rect 5365 2845 5395 2875
rect 5395 2845 5396 2875
rect 5364 2844 5396 2845
rect 5364 2795 5396 2796
rect 5364 2765 5365 2795
rect 5365 2765 5395 2795
rect 5395 2765 5396 2795
rect 5364 2764 5396 2765
rect 5364 2715 5396 2716
rect 5364 2685 5365 2715
rect 5365 2685 5395 2715
rect 5395 2685 5396 2715
rect 5364 2684 5396 2685
rect 5364 2635 5396 2636
rect 5364 2605 5365 2635
rect 5365 2605 5395 2635
rect 5395 2605 5396 2635
rect 5364 2604 5396 2605
rect 5364 2555 5396 2556
rect 5364 2525 5365 2555
rect 5365 2525 5395 2555
rect 5395 2525 5396 2555
rect 5364 2524 5396 2525
rect 5364 2475 5396 2476
rect 5364 2445 5365 2475
rect 5365 2445 5395 2475
rect 5395 2445 5396 2475
rect 5364 2444 5396 2445
rect 5364 2364 5396 2396
rect 5364 2315 5396 2316
rect 5364 2285 5365 2315
rect 5365 2285 5395 2315
rect 5395 2285 5396 2315
rect 5364 2284 5396 2285
rect 5364 2235 5396 2236
rect 5364 2205 5365 2235
rect 5365 2205 5395 2235
rect 5395 2205 5396 2235
rect 5364 2204 5396 2205
rect 5364 2155 5396 2156
rect 5364 2125 5365 2155
rect 5365 2125 5395 2155
rect 5395 2125 5396 2155
rect 5364 2124 5396 2125
rect 5364 2075 5396 2076
rect 5364 2045 5365 2075
rect 5365 2045 5395 2075
rect 5395 2045 5396 2075
rect 5364 2044 5396 2045
rect 5364 1995 5396 1996
rect 5364 1965 5365 1995
rect 5365 1965 5395 1995
rect 5395 1965 5396 1995
rect 5364 1964 5396 1965
rect 5364 1915 5396 1916
rect 5364 1885 5365 1915
rect 5365 1885 5395 1915
rect 5395 1885 5396 1915
rect 5364 1884 5396 1885
rect 5364 1835 5396 1836
rect 5364 1805 5365 1835
rect 5365 1805 5395 1835
rect 5395 1805 5396 1835
rect 5364 1804 5396 1805
rect 5364 1755 5396 1756
rect 5364 1725 5365 1755
rect 5365 1725 5395 1755
rect 5395 1725 5396 1755
rect 5364 1724 5396 1725
rect 5364 1675 5396 1676
rect 5364 1645 5365 1675
rect 5365 1645 5395 1675
rect 5395 1645 5396 1675
rect 5364 1644 5396 1645
rect 5364 1595 5396 1596
rect 5364 1565 5365 1595
rect 5365 1565 5395 1595
rect 5395 1565 5396 1595
rect 5364 1564 5396 1565
rect 5364 1515 5396 1516
rect 5364 1485 5365 1515
rect 5365 1485 5395 1515
rect 5395 1485 5396 1515
rect 5364 1484 5396 1485
rect 5364 1435 5396 1436
rect 5364 1405 5365 1435
rect 5365 1405 5395 1435
rect 5395 1405 5396 1435
rect 5364 1404 5396 1405
rect 5364 1355 5396 1356
rect 5364 1325 5365 1355
rect 5365 1325 5395 1355
rect 5395 1325 5396 1355
rect 5364 1324 5396 1325
rect 5364 1275 5396 1276
rect 5364 1245 5365 1275
rect 5365 1245 5395 1275
rect 5395 1245 5396 1275
rect 5364 1244 5396 1245
rect 5364 1195 5396 1196
rect 5364 1165 5365 1195
rect 5365 1165 5395 1195
rect 5395 1165 5396 1195
rect 5364 1164 5396 1165
rect 5364 1115 5396 1116
rect 5364 1085 5365 1115
rect 5365 1085 5395 1115
rect 5395 1085 5396 1115
rect 5364 1084 5396 1085
rect 5364 1035 5396 1036
rect 5364 1005 5365 1035
rect 5365 1005 5395 1035
rect 5395 1005 5396 1035
rect 5364 1004 5396 1005
rect 5364 955 5396 956
rect 5364 925 5365 955
rect 5365 925 5395 955
rect 5395 925 5396 955
rect 5364 924 5396 925
rect 5364 875 5396 876
rect 5364 845 5365 875
rect 5365 845 5395 875
rect 5395 845 5396 875
rect 5364 844 5396 845
rect 5364 764 5396 796
rect 5364 715 5396 716
rect 5364 685 5365 715
rect 5365 685 5395 715
rect 5395 685 5396 715
rect 5364 684 5396 685
rect 5364 635 5396 636
rect 5364 605 5365 635
rect 5365 605 5395 635
rect 5395 605 5396 635
rect 5364 604 5396 605
rect 5364 555 5396 556
rect 5364 525 5365 555
rect 5365 525 5395 555
rect 5395 525 5396 555
rect 5364 524 5396 525
rect 5364 475 5396 476
rect 5364 445 5365 475
rect 5365 445 5395 475
rect 5395 445 5396 475
rect 5364 444 5396 445
rect 5364 395 5396 396
rect 5364 365 5365 395
rect 5365 365 5395 395
rect 5395 365 5396 395
rect 5364 364 5396 365
rect 5364 315 5396 316
rect 5364 285 5365 315
rect 5365 285 5395 315
rect 5395 285 5396 315
rect 5364 284 5396 285
rect 5364 235 5396 236
rect 5364 205 5365 235
rect 5365 205 5395 235
rect 5395 205 5396 235
rect 5364 204 5396 205
rect 5364 155 5396 156
rect 5364 125 5365 155
rect 5365 125 5395 155
rect 5395 125 5396 155
rect 5364 124 5396 125
rect 5364 75 5396 76
rect 5364 45 5365 75
rect 5365 45 5395 75
rect 5395 45 5396 75
rect 5364 44 5396 45
rect 5364 -5 5396 -4
rect 5364 -35 5365 -5
rect 5365 -35 5395 -5
rect 5395 -35 5396 -5
rect 5364 -36 5396 -35
rect 5364 -85 5396 -84
rect 5364 -115 5365 -85
rect 5365 -115 5395 -85
rect 5395 -115 5396 -85
rect 5364 -116 5396 -115
rect 5524 5595 5556 5596
rect 5524 5565 5525 5595
rect 5525 5565 5555 5595
rect 5555 5565 5556 5595
rect 5524 5564 5556 5565
rect 5524 5515 5556 5516
rect 5524 5485 5525 5515
rect 5525 5485 5555 5515
rect 5555 5485 5556 5515
rect 5524 5484 5556 5485
rect 5524 5435 5556 5436
rect 5524 5405 5525 5435
rect 5525 5405 5555 5435
rect 5555 5405 5556 5435
rect 5524 5404 5556 5405
rect 5524 5355 5556 5356
rect 5524 5325 5525 5355
rect 5525 5325 5555 5355
rect 5555 5325 5556 5355
rect 5524 5324 5556 5325
rect 5524 5275 5556 5276
rect 5524 5245 5525 5275
rect 5525 5245 5555 5275
rect 5555 5245 5556 5275
rect 5524 5244 5556 5245
rect 5524 5195 5556 5196
rect 5524 5165 5525 5195
rect 5525 5165 5555 5195
rect 5555 5165 5556 5195
rect 5524 5164 5556 5165
rect 5524 5115 5556 5116
rect 5524 5085 5525 5115
rect 5525 5085 5555 5115
rect 5555 5085 5556 5115
rect 5524 5084 5556 5085
rect 5524 5035 5556 5036
rect 5524 5005 5525 5035
rect 5525 5005 5555 5035
rect 5555 5005 5556 5035
rect 5524 5004 5556 5005
rect 5524 4955 5556 4956
rect 5524 4925 5525 4955
rect 5525 4925 5555 4955
rect 5555 4925 5556 4955
rect 5524 4924 5556 4925
rect 5524 4875 5556 4876
rect 5524 4845 5525 4875
rect 5525 4845 5555 4875
rect 5555 4845 5556 4875
rect 5524 4844 5556 4845
rect 5524 4795 5556 4796
rect 5524 4765 5525 4795
rect 5525 4765 5555 4795
rect 5555 4765 5556 4795
rect 5524 4764 5556 4765
rect 5524 4715 5556 4716
rect 5524 4685 5525 4715
rect 5525 4685 5555 4715
rect 5555 4685 5556 4715
rect 5524 4684 5556 4685
rect 5524 4635 5556 4636
rect 5524 4605 5525 4635
rect 5525 4605 5555 4635
rect 5555 4605 5556 4635
rect 5524 4604 5556 4605
rect 5524 4555 5556 4556
rect 5524 4525 5525 4555
rect 5525 4525 5555 4555
rect 5555 4525 5556 4555
rect 5524 4524 5556 4525
rect 5524 4475 5556 4476
rect 5524 4445 5525 4475
rect 5525 4445 5555 4475
rect 5555 4445 5556 4475
rect 5524 4444 5556 4445
rect 5524 4395 5556 4396
rect 5524 4365 5525 4395
rect 5525 4365 5555 4395
rect 5555 4365 5556 4395
rect 5524 4364 5556 4365
rect 5524 4284 5556 4316
rect 5524 4235 5556 4236
rect 5524 4205 5525 4235
rect 5525 4205 5555 4235
rect 5555 4205 5556 4235
rect 5524 4204 5556 4205
rect 5524 4155 5556 4156
rect 5524 4125 5525 4155
rect 5525 4125 5555 4155
rect 5555 4125 5556 4155
rect 5524 4124 5556 4125
rect 5524 4075 5556 4076
rect 5524 4045 5525 4075
rect 5525 4045 5555 4075
rect 5555 4045 5556 4075
rect 5524 4044 5556 4045
rect 5524 3995 5556 3996
rect 5524 3965 5525 3995
rect 5525 3965 5555 3995
rect 5555 3965 5556 3995
rect 5524 3964 5556 3965
rect 5524 3915 5556 3916
rect 5524 3885 5525 3915
rect 5525 3885 5555 3915
rect 5555 3885 5556 3915
rect 5524 3884 5556 3885
rect 5524 3835 5556 3836
rect 5524 3805 5525 3835
rect 5525 3805 5555 3835
rect 5555 3805 5556 3835
rect 5524 3804 5556 3805
rect 5524 3755 5556 3756
rect 5524 3725 5525 3755
rect 5525 3725 5555 3755
rect 5555 3725 5556 3755
rect 5524 3724 5556 3725
rect 5524 3675 5556 3676
rect 5524 3645 5525 3675
rect 5525 3645 5555 3675
rect 5555 3645 5556 3675
rect 5524 3644 5556 3645
rect 5524 3595 5556 3596
rect 5524 3565 5525 3595
rect 5525 3565 5555 3595
rect 5555 3565 5556 3595
rect 5524 3564 5556 3565
rect 5524 3515 5556 3516
rect 5524 3485 5525 3515
rect 5525 3485 5555 3515
rect 5555 3485 5556 3515
rect 5524 3484 5556 3485
rect 5524 3435 5556 3436
rect 5524 3405 5525 3435
rect 5525 3405 5555 3435
rect 5555 3405 5556 3435
rect 5524 3404 5556 3405
rect 5524 3355 5556 3356
rect 5524 3325 5525 3355
rect 5525 3325 5555 3355
rect 5555 3325 5556 3355
rect 5524 3324 5556 3325
rect 5524 3275 5556 3276
rect 5524 3245 5525 3275
rect 5525 3245 5555 3275
rect 5555 3245 5556 3275
rect 5524 3244 5556 3245
rect 5524 3195 5556 3196
rect 5524 3165 5525 3195
rect 5525 3165 5555 3195
rect 5555 3165 5556 3195
rect 5524 3164 5556 3165
rect 5524 3115 5556 3116
rect 5524 3085 5525 3115
rect 5525 3085 5555 3115
rect 5555 3085 5556 3115
rect 5524 3084 5556 3085
rect 5524 3035 5556 3036
rect 5524 3005 5525 3035
rect 5525 3005 5555 3035
rect 5555 3005 5556 3035
rect 5524 3004 5556 3005
rect 5524 2955 5556 2956
rect 5524 2925 5525 2955
rect 5525 2925 5555 2955
rect 5555 2925 5556 2955
rect 5524 2924 5556 2925
rect 5524 2875 5556 2876
rect 5524 2845 5525 2875
rect 5525 2845 5555 2875
rect 5555 2845 5556 2875
rect 5524 2844 5556 2845
rect 5524 2795 5556 2796
rect 5524 2765 5525 2795
rect 5525 2765 5555 2795
rect 5555 2765 5556 2795
rect 5524 2764 5556 2765
rect 5524 2715 5556 2716
rect 5524 2685 5525 2715
rect 5525 2685 5555 2715
rect 5555 2685 5556 2715
rect 5524 2684 5556 2685
rect 5524 2635 5556 2636
rect 5524 2605 5525 2635
rect 5525 2605 5555 2635
rect 5555 2605 5556 2635
rect 5524 2604 5556 2605
rect 5524 2555 5556 2556
rect 5524 2525 5525 2555
rect 5525 2525 5555 2555
rect 5555 2525 5556 2555
rect 5524 2524 5556 2525
rect 5524 2475 5556 2476
rect 5524 2445 5525 2475
rect 5525 2445 5555 2475
rect 5555 2445 5556 2475
rect 5524 2444 5556 2445
rect 5524 2364 5556 2396
rect 5524 2315 5556 2316
rect 5524 2285 5525 2315
rect 5525 2285 5555 2315
rect 5555 2285 5556 2315
rect 5524 2284 5556 2285
rect 5524 2235 5556 2236
rect 5524 2205 5525 2235
rect 5525 2205 5555 2235
rect 5555 2205 5556 2235
rect 5524 2204 5556 2205
rect 5524 2155 5556 2156
rect 5524 2125 5525 2155
rect 5525 2125 5555 2155
rect 5555 2125 5556 2155
rect 5524 2124 5556 2125
rect 5524 2075 5556 2076
rect 5524 2045 5525 2075
rect 5525 2045 5555 2075
rect 5555 2045 5556 2075
rect 5524 2044 5556 2045
rect 5524 1995 5556 1996
rect 5524 1965 5525 1995
rect 5525 1965 5555 1995
rect 5555 1965 5556 1995
rect 5524 1964 5556 1965
rect 5524 1915 5556 1916
rect 5524 1885 5525 1915
rect 5525 1885 5555 1915
rect 5555 1885 5556 1915
rect 5524 1884 5556 1885
rect 5524 1835 5556 1836
rect 5524 1805 5525 1835
rect 5525 1805 5555 1835
rect 5555 1805 5556 1835
rect 5524 1804 5556 1805
rect 5524 1755 5556 1756
rect 5524 1725 5525 1755
rect 5525 1725 5555 1755
rect 5555 1725 5556 1755
rect 5524 1724 5556 1725
rect 5524 1675 5556 1676
rect 5524 1645 5525 1675
rect 5525 1645 5555 1675
rect 5555 1645 5556 1675
rect 5524 1644 5556 1645
rect 5524 1595 5556 1596
rect 5524 1565 5525 1595
rect 5525 1565 5555 1595
rect 5555 1565 5556 1595
rect 5524 1564 5556 1565
rect 5524 1515 5556 1516
rect 5524 1485 5525 1515
rect 5525 1485 5555 1515
rect 5555 1485 5556 1515
rect 5524 1484 5556 1485
rect 5524 1435 5556 1436
rect 5524 1405 5525 1435
rect 5525 1405 5555 1435
rect 5555 1405 5556 1435
rect 5524 1404 5556 1405
rect 5524 1355 5556 1356
rect 5524 1325 5525 1355
rect 5525 1325 5555 1355
rect 5555 1325 5556 1355
rect 5524 1324 5556 1325
rect 5524 1275 5556 1276
rect 5524 1245 5525 1275
rect 5525 1245 5555 1275
rect 5555 1245 5556 1275
rect 5524 1244 5556 1245
rect 5524 1195 5556 1196
rect 5524 1165 5525 1195
rect 5525 1165 5555 1195
rect 5555 1165 5556 1195
rect 5524 1164 5556 1165
rect 5524 1115 5556 1116
rect 5524 1085 5525 1115
rect 5525 1085 5555 1115
rect 5555 1085 5556 1115
rect 5524 1084 5556 1085
rect 5524 1035 5556 1036
rect 5524 1005 5525 1035
rect 5525 1005 5555 1035
rect 5555 1005 5556 1035
rect 5524 1004 5556 1005
rect 5524 955 5556 956
rect 5524 925 5525 955
rect 5525 925 5555 955
rect 5555 925 5556 955
rect 5524 924 5556 925
rect 5524 875 5556 876
rect 5524 845 5525 875
rect 5525 845 5555 875
rect 5555 845 5556 875
rect 5524 844 5556 845
rect 5524 795 5556 796
rect 5524 765 5525 795
rect 5525 765 5555 795
rect 5555 765 5556 795
rect 5524 764 5556 765
rect 5524 715 5556 716
rect 5524 685 5525 715
rect 5525 685 5555 715
rect 5555 685 5556 715
rect 5524 684 5556 685
rect 5524 635 5556 636
rect 5524 605 5525 635
rect 5525 605 5555 635
rect 5555 605 5556 635
rect 5524 604 5556 605
rect 5524 555 5556 556
rect 5524 525 5525 555
rect 5525 525 5555 555
rect 5555 525 5556 555
rect 5524 524 5556 525
rect 5524 475 5556 476
rect 5524 445 5525 475
rect 5525 445 5555 475
rect 5555 445 5556 475
rect 5524 444 5556 445
rect 5524 395 5556 396
rect 5524 365 5525 395
rect 5525 365 5555 395
rect 5555 365 5556 395
rect 5524 364 5556 365
rect 5524 315 5556 316
rect 5524 285 5525 315
rect 5525 285 5555 315
rect 5555 285 5556 315
rect 5524 284 5556 285
rect 5524 235 5556 236
rect 5524 205 5525 235
rect 5525 205 5555 235
rect 5555 205 5556 235
rect 5524 204 5556 205
rect 5524 155 5556 156
rect 5524 125 5525 155
rect 5525 125 5555 155
rect 5555 125 5556 155
rect 5524 124 5556 125
rect 5524 75 5556 76
rect 5524 45 5525 75
rect 5525 45 5555 75
rect 5555 45 5556 75
rect 5524 44 5556 45
rect 5524 -5 5556 -4
rect 5524 -35 5525 -5
rect 5525 -35 5555 -5
rect 5555 -35 5556 -5
rect 5524 -36 5556 -35
rect 5524 -85 5556 -84
rect 5524 -115 5525 -85
rect 5525 -115 5555 -85
rect 5555 -115 5556 -85
rect 5524 -116 5556 -115
rect 5684 5595 5716 5596
rect 5684 5565 5685 5595
rect 5685 5565 5715 5595
rect 5715 5565 5716 5595
rect 5684 5564 5716 5565
rect 5684 5515 5716 5516
rect 5684 5485 5685 5515
rect 5685 5485 5715 5515
rect 5715 5485 5716 5515
rect 5684 5484 5716 5485
rect 5684 5435 5716 5436
rect 5684 5405 5685 5435
rect 5685 5405 5715 5435
rect 5715 5405 5716 5435
rect 5684 5404 5716 5405
rect 5684 5355 5716 5356
rect 5684 5325 5685 5355
rect 5685 5325 5715 5355
rect 5715 5325 5716 5355
rect 5684 5324 5716 5325
rect 5684 5275 5716 5276
rect 5684 5245 5685 5275
rect 5685 5245 5715 5275
rect 5715 5245 5716 5275
rect 5684 5244 5716 5245
rect 5684 5195 5716 5196
rect 5684 5165 5685 5195
rect 5685 5165 5715 5195
rect 5715 5165 5716 5195
rect 5684 5164 5716 5165
rect 5684 5115 5716 5116
rect 5684 5085 5685 5115
rect 5685 5085 5715 5115
rect 5715 5085 5716 5115
rect 5684 5084 5716 5085
rect 5684 5035 5716 5036
rect 5684 5005 5685 5035
rect 5685 5005 5715 5035
rect 5715 5005 5716 5035
rect 5684 5004 5716 5005
rect 5684 4955 5716 4956
rect 5684 4925 5685 4955
rect 5685 4925 5715 4955
rect 5715 4925 5716 4955
rect 5684 4924 5716 4925
rect 5684 4875 5716 4876
rect 5684 4845 5685 4875
rect 5685 4845 5715 4875
rect 5715 4845 5716 4875
rect 5684 4844 5716 4845
rect 5684 4795 5716 4796
rect 5684 4765 5685 4795
rect 5685 4765 5715 4795
rect 5715 4765 5716 4795
rect 5684 4764 5716 4765
rect 5684 4715 5716 4716
rect 5684 4685 5685 4715
rect 5685 4685 5715 4715
rect 5715 4685 5716 4715
rect 5684 4684 5716 4685
rect 5684 4635 5716 4636
rect 5684 4605 5685 4635
rect 5685 4605 5715 4635
rect 5715 4605 5716 4635
rect 5684 4604 5716 4605
rect 5684 4555 5716 4556
rect 5684 4525 5685 4555
rect 5685 4525 5715 4555
rect 5715 4525 5716 4555
rect 5684 4524 5716 4525
rect 5684 4475 5716 4476
rect 5684 4445 5685 4475
rect 5685 4445 5715 4475
rect 5715 4445 5716 4475
rect 5684 4444 5716 4445
rect 5684 4395 5716 4396
rect 5684 4365 5685 4395
rect 5685 4365 5715 4395
rect 5715 4365 5716 4395
rect 5684 4364 5716 4365
rect 5684 4284 5716 4316
rect 5684 4235 5716 4236
rect 5684 4205 5685 4235
rect 5685 4205 5715 4235
rect 5715 4205 5716 4235
rect 5684 4204 5716 4205
rect 5684 4155 5716 4156
rect 5684 4125 5685 4155
rect 5685 4125 5715 4155
rect 5715 4125 5716 4155
rect 5684 4124 5716 4125
rect 5684 4075 5716 4076
rect 5684 4045 5685 4075
rect 5685 4045 5715 4075
rect 5715 4045 5716 4075
rect 5684 4044 5716 4045
rect 5684 3995 5716 3996
rect 5684 3965 5685 3995
rect 5685 3965 5715 3995
rect 5715 3965 5716 3995
rect 5684 3964 5716 3965
rect 5684 3915 5716 3916
rect 5684 3885 5685 3915
rect 5685 3885 5715 3915
rect 5715 3885 5716 3915
rect 5684 3884 5716 3885
rect 5684 3835 5716 3836
rect 5684 3805 5685 3835
rect 5685 3805 5715 3835
rect 5715 3805 5716 3835
rect 5684 3804 5716 3805
rect 5684 3755 5716 3756
rect 5684 3725 5685 3755
rect 5685 3725 5715 3755
rect 5715 3725 5716 3755
rect 5684 3724 5716 3725
rect 5684 3675 5716 3676
rect 5684 3645 5685 3675
rect 5685 3645 5715 3675
rect 5715 3645 5716 3675
rect 5684 3644 5716 3645
rect 5684 3595 5716 3596
rect 5684 3565 5685 3595
rect 5685 3565 5715 3595
rect 5715 3565 5716 3595
rect 5684 3564 5716 3565
rect 5684 3515 5716 3516
rect 5684 3485 5685 3515
rect 5685 3485 5715 3515
rect 5715 3485 5716 3515
rect 5684 3484 5716 3485
rect 5684 3435 5716 3436
rect 5684 3405 5685 3435
rect 5685 3405 5715 3435
rect 5715 3405 5716 3435
rect 5684 3404 5716 3405
rect 5684 3355 5716 3356
rect 5684 3325 5685 3355
rect 5685 3325 5715 3355
rect 5715 3325 5716 3355
rect 5684 3324 5716 3325
rect 5684 3275 5716 3276
rect 5684 3245 5685 3275
rect 5685 3245 5715 3275
rect 5715 3245 5716 3275
rect 5684 3244 5716 3245
rect 5684 3195 5716 3196
rect 5684 3165 5685 3195
rect 5685 3165 5715 3195
rect 5715 3165 5716 3195
rect 5684 3164 5716 3165
rect 5684 3115 5716 3116
rect 5684 3085 5685 3115
rect 5685 3085 5715 3115
rect 5715 3085 5716 3115
rect 5684 3084 5716 3085
rect 5684 3035 5716 3036
rect 5684 3005 5685 3035
rect 5685 3005 5715 3035
rect 5715 3005 5716 3035
rect 5684 3004 5716 3005
rect 5684 2955 5716 2956
rect 5684 2925 5685 2955
rect 5685 2925 5715 2955
rect 5715 2925 5716 2955
rect 5684 2924 5716 2925
rect 5684 2875 5716 2876
rect 5684 2845 5685 2875
rect 5685 2845 5715 2875
rect 5715 2845 5716 2875
rect 5684 2844 5716 2845
rect 5684 2795 5716 2796
rect 5684 2765 5685 2795
rect 5685 2765 5715 2795
rect 5715 2765 5716 2795
rect 5684 2764 5716 2765
rect 5684 2715 5716 2716
rect 5684 2685 5685 2715
rect 5685 2685 5715 2715
rect 5715 2685 5716 2715
rect 5684 2684 5716 2685
rect 5684 2635 5716 2636
rect 5684 2605 5685 2635
rect 5685 2605 5715 2635
rect 5715 2605 5716 2635
rect 5684 2604 5716 2605
rect 5684 2555 5716 2556
rect 5684 2525 5685 2555
rect 5685 2525 5715 2555
rect 5715 2525 5716 2555
rect 5684 2524 5716 2525
rect 5684 2475 5716 2476
rect 5684 2445 5685 2475
rect 5685 2445 5715 2475
rect 5715 2445 5716 2475
rect 5684 2444 5716 2445
rect 5684 2364 5716 2396
rect 5684 2315 5716 2316
rect 5684 2285 5685 2315
rect 5685 2285 5715 2315
rect 5715 2285 5716 2315
rect 5684 2284 5716 2285
rect 5684 2235 5716 2236
rect 5684 2205 5685 2235
rect 5685 2205 5715 2235
rect 5715 2205 5716 2235
rect 5684 2204 5716 2205
rect 5684 2155 5716 2156
rect 5684 2125 5685 2155
rect 5685 2125 5715 2155
rect 5715 2125 5716 2155
rect 5684 2124 5716 2125
rect 5684 2075 5716 2076
rect 5684 2045 5685 2075
rect 5685 2045 5715 2075
rect 5715 2045 5716 2075
rect 5684 2044 5716 2045
rect 5684 1995 5716 1996
rect 5684 1965 5685 1995
rect 5685 1965 5715 1995
rect 5715 1965 5716 1995
rect 5684 1964 5716 1965
rect 5684 1915 5716 1916
rect 5684 1885 5685 1915
rect 5685 1885 5715 1915
rect 5715 1885 5716 1915
rect 5684 1884 5716 1885
rect 5684 1835 5716 1836
rect 5684 1805 5685 1835
rect 5685 1805 5715 1835
rect 5715 1805 5716 1835
rect 5684 1804 5716 1805
rect 5684 1755 5716 1756
rect 5684 1725 5685 1755
rect 5685 1725 5715 1755
rect 5715 1725 5716 1755
rect 5684 1724 5716 1725
rect 5684 1675 5716 1676
rect 5684 1645 5685 1675
rect 5685 1645 5715 1675
rect 5715 1645 5716 1675
rect 5684 1644 5716 1645
rect 5684 1595 5716 1596
rect 5684 1565 5685 1595
rect 5685 1565 5715 1595
rect 5715 1565 5716 1595
rect 5684 1564 5716 1565
rect 5684 1515 5716 1516
rect 5684 1485 5685 1515
rect 5685 1485 5715 1515
rect 5715 1485 5716 1515
rect 5684 1484 5716 1485
rect 5684 1435 5716 1436
rect 5684 1405 5685 1435
rect 5685 1405 5715 1435
rect 5715 1405 5716 1435
rect 5684 1404 5716 1405
rect 5684 1355 5716 1356
rect 5684 1325 5685 1355
rect 5685 1325 5715 1355
rect 5715 1325 5716 1355
rect 5684 1324 5716 1325
rect 5684 1275 5716 1276
rect 5684 1245 5685 1275
rect 5685 1245 5715 1275
rect 5715 1245 5716 1275
rect 5684 1244 5716 1245
rect 5684 1195 5716 1196
rect 5684 1165 5685 1195
rect 5685 1165 5715 1195
rect 5715 1165 5716 1195
rect 5684 1164 5716 1165
rect 5684 1115 5716 1116
rect 5684 1085 5685 1115
rect 5685 1085 5715 1115
rect 5715 1085 5716 1115
rect 5684 1084 5716 1085
rect 5684 1035 5716 1036
rect 5684 1005 5685 1035
rect 5685 1005 5715 1035
rect 5715 1005 5716 1035
rect 5684 1004 5716 1005
rect 5684 955 5716 956
rect 5684 925 5685 955
rect 5685 925 5715 955
rect 5715 925 5716 955
rect 5684 924 5716 925
rect 5684 875 5716 876
rect 5684 845 5685 875
rect 5685 845 5715 875
rect 5715 845 5716 875
rect 5684 844 5716 845
rect 5684 795 5716 796
rect 5684 765 5685 795
rect 5685 765 5715 795
rect 5715 765 5716 795
rect 5684 764 5716 765
rect 5684 715 5716 716
rect 5684 685 5685 715
rect 5685 685 5715 715
rect 5715 685 5716 715
rect 5684 684 5716 685
rect 5684 635 5716 636
rect 5684 605 5685 635
rect 5685 605 5715 635
rect 5715 605 5716 635
rect 5684 604 5716 605
rect 5684 555 5716 556
rect 5684 525 5685 555
rect 5685 525 5715 555
rect 5715 525 5716 555
rect 5684 524 5716 525
rect 5684 475 5716 476
rect 5684 445 5685 475
rect 5685 445 5715 475
rect 5715 445 5716 475
rect 5684 444 5716 445
rect 5684 395 5716 396
rect 5684 365 5685 395
rect 5685 365 5715 395
rect 5715 365 5716 395
rect 5684 364 5716 365
rect 5684 315 5716 316
rect 5684 285 5685 315
rect 5685 285 5715 315
rect 5715 285 5716 315
rect 5684 284 5716 285
rect 5684 235 5716 236
rect 5684 205 5685 235
rect 5685 205 5715 235
rect 5715 205 5716 235
rect 5684 204 5716 205
rect 5684 155 5716 156
rect 5684 125 5685 155
rect 5685 125 5715 155
rect 5715 125 5716 155
rect 5684 124 5716 125
rect 5684 75 5716 76
rect 5684 45 5685 75
rect 5685 45 5715 75
rect 5715 45 5716 75
rect 5684 44 5716 45
rect 5684 -5 5716 -4
rect 5684 -35 5685 -5
rect 5685 -35 5715 -5
rect 5715 -35 5716 -5
rect 5684 -36 5716 -35
rect 5684 -85 5716 -84
rect 5684 -115 5685 -85
rect 5685 -115 5715 -85
rect 5715 -115 5716 -85
rect 5684 -116 5716 -115
<< metal4 >>
rect -1520 5596 -840 5600
rect -1520 5564 -1516 5596
rect -1484 5564 -1356 5596
rect -1324 5564 -1196 5596
rect -1164 5564 -1036 5596
rect -1004 5564 -876 5596
rect -844 5564 -840 5596
rect -1520 5560 -840 5564
rect -800 5596 5720 5600
rect -800 5564 4884 5596
rect 4916 5564 5044 5596
rect 5076 5564 5204 5596
rect 5236 5564 5364 5596
rect 5396 5564 5524 5596
rect 5556 5564 5684 5596
rect 5716 5564 5720 5596
rect -800 5560 5720 5564
rect -1520 5516 -840 5520
rect -1520 5484 -1516 5516
rect -1484 5484 -1356 5516
rect -1324 5484 -1196 5516
rect -1164 5484 -1036 5516
rect -1004 5484 -876 5516
rect -844 5484 -840 5516
rect -1520 5480 -840 5484
rect -800 5516 4840 5520
rect -800 5484 -796 5516
rect -764 5484 -716 5516
rect -684 5484 -636 5516
rect -604 5484 -556 5516
rect -524 5484 -476 5516
rect -444 5484 -396 5516
rect -364 5484 -316 5516
rect -284 5484 -236 5516
rect -204 5484 -156 5516
rect -124 5484 -76 5516
rect -44 5484 4 5516
rect 36 5484 84 5516
rect 116 5484 164 5516
rect 196 5484 244 5516
rect 276 5484 324 5516
rect 356 5484 404 5516
rect 436 5484 484 5516
rect 516 5484 564 5516
rect 596 5484 644 5516
rect 676 5484 724 5516
rect 756 5484 804 5516
rect 836 5484 884 5516
rect 916 5484 964 5516
rect 996 5484 1044 5516
rect 1076 5484 1124 5516
rect 1156 5484 1204 5516
rect 1236 5484 1284 5516
rect 1316 5484 1364 5516
rect 1396 5484 1444 5516
rect 1476 5484 1524 5516
rect 1556 5484 1604 5516
rect 1636 5484 1684 5516
rect 1716 5484 1764 5516
rect 1796 5484 1844 5516
rect 1876 5484 1924 5516
rect 1956 5484 2004 5516
rect 2036 5484 2084 5516
rect 2116 5484 2164 5516
rect 2196 5484 2244 5516
rect 2276 5484 2324 5516
rect 2356 5484 2404 5516
rect 2436 5484 2484 5516
rect 2516 5484 2564 5516
rect 2596 5484 2644 5516
rect 2676 5484 2724 5516
rect 2756 5484 2804 5516
rect 2836 5484 2884 5516
rect 2916 5484 2964 5516
rect 2996 5484 3044 5516
rect 3076 5484 3124 5516
rect 3156 5484 3204 5516
rect 3236 5484 3284 5516
rect 3316 5484 3364 5516
rect 3396 5484 3444 5516
rect 3476 5484 3524 5516
rect 3556 5484 3604 5516
rect 3636 5484 3684 5516
rect 3716 5484 3764 5516
rect 3796 5484 3844 5516
rect 3876 5484 3924 5516
rect 3956 5484 4004 5516
rect 4036 5484 4084 5516
rect 4116 5484 4164 5516
rect 4196 5484 4244 5516
rect 4276 5484 4324 5516
rect 4356 5484 4404 5516
rect 4436 5484 4484 5516
rect 4516 5484 4564 5516
rect 4596 5484 4644 5516
rect 4676 5484 4724 5516
rect 4756 5484 4804 5516
rect 4836 5484 4840 5516
rect -800 5480 4840 5484
rect 4880 5516 5720 5520
rect 4880 5484 4884 5516
rect 4916 5484 5044 5516
rect 5076 5484 5204 5516
rect 5236 5484 5364 5516
rect 5396 5484 5524 5516
rect 5556 5484 5684 5516
rect 5716 5484 5720 5516
rect 4880 5480 5720 5484
rect -1520 5436 -840 5440
rect -1520 5404 -1516 5436
rect -1484 5404 -1356 5436
rect -1324 5404 -1196 5436
rect -1164 5404 -1036 5436
rect -1004 5404 -876 5436
rect -844 5404 -840 5436
rect -1520 5400 -840 5404
rect -800 5436 4840 5440
rect -800 5404 -796 5436
rect -764 5404 -716 5436
rect -684 5404 -636 5436
rect -604 5404 -556 5436
rect -524 5404 -476 5436
rect -444 5404 -396 5436
rect -364 5404 -316 5436
rect -284 5404 -236 5436
rect -204 5404 -156 5436
rect -124 5404 -76 5436
rect -44 5404 4 5436
rect 36 5404 84 5436
rect 116 5404 164 5436
rect 196 5404 244 5436
rect 276 5404 324 5436
rect 356 5404 404 5436
rect 436 5404 484 5436
rect 516 5404 564 5436
rect 596 5404 644 5436
rect 676 5404 724 5436
rect 756 5404 804 5436
rect 836 5404 884 5436
rect 916 5404 964 5436
rect 996 5404 1044 5436
rect 1076 5404 1124 5436
rect 1156 5404 1204 5436
rect 1236 5404 1284 5436
rect 1316 5404 1364 5436
rect 1396 5404 1444 5436
rect 1476 5404 1524 5436
rect 1556 5404 1604 5436
rect 1636 5404 1684 5436
rect 1716 5404 1764 5436
rect 1796 5404 1844 5436
rect 1876 5404 1924 5436
rect 1956 5404 2004 5436
rect 2036 5404 2084 5436
rect 2116 5404 2164 5436
rect 2196 5404 2244 5436
rect 2276 5404 2324 5436
rect 2356 5404 2404 5436
rect 2436 5404 2484 5436
rect 2516 5404 2564 5436
rect 2596 5404 2644 5436
rect 2676 5404 2724 5436
rect 2756 5404 2804 5436
rect 2836 5404 2884 5436
rect 2916 5404 2964 5436
rect 2996 5404 3044 5436
rect 3076 5404 3124 5436
rect 3156 5404 3204 5436
rect 3236 5404 3284 5436
rect 3316 5404 3364 5436
rect 3396 5404 3444 5436
rect 3476 5404 3524 5436
rect 3556 5404 3604 5436
rect 3636 5404 3684 5436
rect 3716 5404 3764 5436
rect 3796 5404 3844 5436
rect 3876 5404 3924 5436
rect 3956 5404 4004 5436
rect 4036 5404 4084 5436
rect 4116 5404 4164 5436
rect 4196 5404 4244 5436
rect 4276 5404 4324 5436
rect 4356 5404 4404 5436
rect 4436 5404 4484 5436
rect 4516 5404 4564 5436
rect 4596 5404 4644 5436
rect 4676 5404 4724 5436
rect 4756 5404 4804 5436
rect 4836 5404 4840 5436
rect -800 5400 4840 5404
rect 4880 5436 5720 5440
rect 4880 5404 4884 5436
rect 4916 5404 5044 5436
rect 5076 5404 5204 5436
rect 5236 5404 5364 5436
rect 5396 5404 5524 5436
rect 5556 5404 5684 5436
rect 5716 5404 5720 5436
rect 4880 5400 5720 5404
rect -1520 5356 -840 5360
rect -1520 5324 -1516 5356
rect -1484 5324 -1356 5356
rect -1324 5324 -1196 5356
rect -1164 5324 -1036 5356
rect -1004 5324 -876 5356
rect -844 5324 -840 5356
rect -1520 5320 -840 5324
rect -800 5356 4840 5360
rect -800 5324 -796 5356
rect -764 5324 -716 5356
rect -684 5324 -636 5356
rect -604 5324 -556 5356
rect -524 5324 -476 5356
rect -444 5324 -396 5356
rect -364 5324 -316 5356
rect -284 5324 -236 5356
rect -204 5324 -156 5356
rect -124 5324 -76 5356
rect -44 5324 4 5356
rect 36 5324 84 5356
rect 116 5324 164 5356
rect 196 5324 244 5356
rect 276 5324 324 5356
rect 356 5324 404 5356
rect 436 5324 484 5356
rect 516 5324 564 5356
rect 596 5324 644 5356
rect 676 5324 724 5356
rect 756 5324 804 5356
rect 836 5324 884 5356
rect 916 5324 964 5356
rect 996 5324 1044 5356
rect 1076 5324 1124 5356
rect 1156 5324 1204 5356
rect 1236 5324 1284 5356
rect 1316 5324 1364 5356
rect 1396 5324 1444 5356
rect 1476 5324 1524 5356
rect 1556 5324 1604 5356
rect 1636 5324 1684 5356
rect 1716 5324 1764 5356
rect 1796 5324 1844 5356
rect 1876 5324 1924 5356
rect 1956 5324 2004 5356
rect 2036 5324 2084 5356
rect 2116 5324 2164 5356
rect 2196 5324 2244 5356
rect 2276 5324 2324 5356
rect 2356 5324 2404 5356
rect 2436 5324 2484 5356
rect 2516 5324 2564 5356
rect 2596 5324 2644 5356
rect 2676 5324 2724 5356
rect 2756 5324 2804 5356
rect 2836 5324 2884 5356
rect 2916 5324 2964 5356
rect 2996 5324 3044 5356
rect 3076 5324 3124 5356
rect 3156 5324 3204 5356
rect 3236 5324 3284 5356
rect 3316 5324 3364 5356
rect 3396 5324 3444 5356
rect 3476 5324 3524 5356
rect 3556 5324 3604 5356
rect 3636 5324 3684 5356
rect 3716 5324 3764 5356
rect 3796 5324 3844 5356
rect 3876 5324 3924 5356
rect 3956 5324 4004 5356
rect 4036 5324 4084 5356
rect 4116 5324 4164 5356
rect 4196 5324 4244 5356
rect 4276 5324 4324 5356
rect 4356 5324 4404 5356
rect 4436 5324 4484 5356
rect 4516 5324 4564 5356
rect 4596 5324 4644 5356
rect 4676 5324 4724 5356
rect 4756 5324 4804 5356
rect 4836 5324 4840 5356
rect -800 5320 4840 5324
rect 4880 5356 5720 5360
rect 4880 5324 4884 5356
rect 4916 5324 5044 5356
rect 5076 5324 5204 5356
rect 5236 5324 5364 5356
rect 5396 5324 5524 5356
rect 5556 5324 5684 5356
rect 5716 5324 5720 5356
rect 4880 5320 5720 5324
rect -1520 5276 -840 5280
rect -1520 5244 -1516 5276
rect -1484 5244 -1356 5276
rect -1324 5244 -1196 5276
rect -1164 5244 -1036 5276
rect -1004 5244 -876 5276
rect -844 5244 -840 5276
rect -1520 5240 -840 5244
rect -800 5276 4840 5280
rect -800 5244 -796 5276
rect -764 5244 -716 5276
rect -684 5244 -636 5276
rect -604 5244 -556 5276
rect -524 5244 -476 5276
rect -444 5244 -396 5276
rect -364 5244 -316 5276
rect -284 5244 -236 5276
rect -204 5244 -156 5276
rect -124 5244 -76 5276
rect -44 5244 4 5276
rect 36 5244 84 5276
rect 116 5244 164 5276
rect 196 5244 244 5276
rect 276 5244 324 5276
rect 356 5244 404 5276
rect 436 5244 484 5276
rect 516 5244 564 5276
rect 596 5244 644 5276
rect 676 5244 724 5276
rect 756 5244 804 5276
rect 836 5244 884 5276
rect 916 5244 964 5276
rect 996 5244 1044 5276
rect 1076 5244 1124 5276
rect 1156 5244 1204 5276
rect 1236 5244 1284 5276
rect 1316 5244 1364 5276
rect 1396 5244 1444 5276
rect 1476 5244 1524 5276
rect 1556 5244 1604 5276
rect 1636 5244 1684 5276
rect 1716 5244 1764 5276
rect 1796 5244 1844 5276
rect 1876 5244 1924 5276
rect 1956 5244 2004 5276
rect 2036 5244 2084 5276
rect 2116 5244 2164 5276
rect 2196 5244 2244 5276
rect 2276 5244 2324 5276
rect 2356 5244 2404 5276
rect 2436 5244 2484 5276
rect 2516 5244 2564 5276
rect 2596 5244 2644 5276
rect 2676 5244 2724 5276
rect 2756 5244 2804 5276
rect 2836 5244 2884 5276
rect 2916 5244 2964 5276
rect 2996 5244 3044 5276
rect 3076 5244 3124 5276
rect 3156 5244 3204 5276
rect 3236 5244 3284 5276
rect 3316 5244 3364 5276
rect 3396 5244 3444 5276
rect 3476 5244 3524 5276
rect 3556 5244 3604 5276
rect 3636 5244 3684 5276
rect 3716 5244 3764 5276
rect 3796 5244 3844 5276
rect 3876 5244 3924 5276
rect 3956 5244 4004 5276
rect 4036 5244 4084 5276
rect 4116 5244 4164 5276
rect 4196 5244 4244 5276
rect 4276 5244 4324 5276
rect 4356 5244 4404 5276
rect 4436 5244 4484 5276
rect 4516 5244 4564 5276
rect 4596 5244 4644 5276
rect 4676 5244 4724 5276
rect 4756 5244 4804 5276
rect 4836 5244 4840 5276
rect -800 5240 4840 5244
rect 4880 5276 5720 5280
rect 4880 5244 4884 5276
rect 4916 5244 5044 5276
rect 5076 5244 5204 5276
rect 5236 5244 5364 5276
rect 5396 5244 5524 5276
rect 5556 5244 5684 5276
rect 5716 5244 5720 5276
rect 4880 5240 5720 5244
rect -1520 5196 -840 5200
rect -1520 5164 -1516 5196
rect -1484 5164 -1356 5196
rect -1324 5164 -1196 5196
rect -1164 5164 -1036 5196
rect -1004 5164 -876 5196
rect -844 5164 -840 5196
rect -1520 5160 -840 5164
rect -800 5196 4840 5200
rect -800 5164 -796 5196
rect -764 5164 -716 5196
rect -684 5164 -636 5196
rect -604 5164 -556 5196
rect -524 5164 -476 5196
rect -444 5164 -396 5196
rect -364 5164 -316 5196
rect -284 5164 -236 5196
rect -204 5164 -156 5196
rect -124 5164 -76 5196
rect -44 5164 4 5196
rect 36 5164 84 5196
rect 116 5164 164 5196
rect 196 5164 244 5196
rect 276 5164 324 5196
rect 356 5164 404 5196
rect 436 5164 484 5196
rect 516 5164 564 5196
rect 596 5164 644 5196
rect 676 5164 724 5196
rect 756 5164 804 5196
rect 836 5164 884 5196
rect 916 5164 964 5196
rect 996 5164 1044 5196
rect 1076 5164 1124 5196
rect 1156 5164 1204 5196
rect 1236 5164 1284 5196
rect 1316 5164 1364 5196
rect 1396 5164 1444 5196
rect 1476 5164 1524 5196
rect 1556 5164 1604 5196
rect 1636 5164 1684 5196
rect 1716 5164 1764 5196
rect 1796 5164 1844 5196
rect 1876 5164 1924 5196
rect 1956 5164 2004 5196
rect 2036 5164 2084 5196
rect 2116 5164 2164 5196
rect 2196 5164 2244 5196
rect 2276 5164 2324 5196
rect 2356 5164 2404 5196
rect 2436 5164 2484 5196
rect 2516 5164 2564 5196
rect 2596 5164 2644 5196
rect 2676 5164 2724 5196
rect 2756 5164 2804 5196
rect 2836 5164 2884 5196
rect 2916 5164 2964 5196
rect 2996 5164 3044 5196
rect 3076 5164 3124 5196
rect 3156 5164 3204 5196
rect 3236 5164 3284 5196
rect 3316 5164 3364 5196
rect 3396 5164 3444 5196
rect 3476 5164 3524 5196
rect 3556 5164 3604 5196
rect 3636 5164 3684 5196
rect 3716 5164 3764 5196
rect 3796 5164 3844 5196
rect 3876 5164 3924 5196
rect 3956 5164 4004 5196
rect 4036 5164 4084 5196
rect 4116 5164 4164 5196
rect 4196 5164 4244 5196
rect 4276 5164 4324 5196
rect 4356 5164 4404 5196
rect 4436 5164 4484 5196
rect 4516 5164 4564 5196
rect 4596 5164 4644 5196
rect 4676 5164 4724 5196
rect 4756 5164 4804 5196
rect 4836 5164 4840 5196
rect -800 5160 4840 5164
rect 4880 5196 5720 5200
rect 4880 5164 4884 5196
rect 4916 5164 5044 5196
rect 5076 5164 5204 5196
rect 5236 5164 5364 5196
rect 5396 5164 5524 5196
rect 5556 5164 5684 5196
rect 5716 5164 5720 5196
rect 4880 5160 5720 5164
rect -1520 5116 -840 5120
rect -1520 5084 -1516 5116
rect -1484 5084 -1356 5116
rect -1324 5084 -1196 5116
rect -1164 5084 -1036 5116
rect -1004 5084 -876 5116
rect -844 5084 -840 5116
rect -1520 5080 -840 5084
rect -800 5116 4840 5120
rect -800 5084 -796 5116
rect -764 5084 -716 5116
rect -684 5084 -636 5116
rect -604 5084 -556 5116
rect -524 5084 -476 5116
rect -444 5084 -396 5116
rect -364 5084 -316 5116
rect -284 5084 -236 5116
rect -204 5084 -156 5116
rect -124 5084 -76 5116
rect -44 5084 4 5116
rect 36 5084 84 5116
rect 116 5084 164 5116
rect 196 5084 244 5116
rect 276 5084 324 5116
rect 356 5084 404 5116
rect 436 5084 484 5116
rect 516 5084 564 5116
rect 596 5084 644 5116
rect 676 5084 724 5116
rect 756 5084 804 5116
rect 836 5084 884 5116
rect 916 5084 964 5116
rect 996 5084 1044 5116
rect 1076 5084 1124 5116
rect 1156 5084 1204 5116
rect 1236 5084 1284 5116
rect 1316 5084 1364 5116
rect 1396 5084 1444 5116
rect 1476 5084 1524 5116
rect 1556 5084 1604 5116
rect 1636 5084 1684 5116
rect 1716 5084 1764 5116
rect 1796 5084 1844 5116
rect 1876 5084 1924 5116
rect 1956 5084 2004 5116
rect 2036 5084 2084 5116
rect 2116 5084 2164 5116
rect 2196 5084 2244 5116
rect 2276 5084 2324 5116
rect 2356 5084 2404 5116
rect 2436 5084 2484 5116
rect 2516 5084 2564 5116
rect 2596 5084 2644 5116
rect 2676 5084 2724 5116
rect 2756 5084 2804 5116
rect 2836 5084 2884 5116
rect 2916 5084 2964 5116
rect 2996 5084 3044 5116
rect 3076 5084 3124 5116
rect 3156 5084 3204 5116
rect 3236 5084 3284 5116
rect 3316 5084 3364 5116
rect 3396 5084 3444 5116
rect 3476 5084 3524 5116
rect 3556 5084 3604 5116
rect 3636 5084 3684 5116
rect 3716 5084 3764 5116
rect 3796 5084 3844 5116
rect 3876 5084 3924 5116
rect 3956 5084 4004 5116
rect 4036 5084 4084 5116
rect 4116 5084 4164 5116
rect 4196 5084 4244 5116
rect 4276 5084 4324 5116
rect 4356 5084 4404 5116
rect 4436 5084 4484 5116
rect 4516 5084 4564 5116
rect 4596 5084 4644 5116
rect 4676 5084 4724 5116
rect 4756 5084 4804 5116
rect 4836 5084 4840 5116
rect -800 5080 4840 5084
rect 4880 5116 5720 5120
rect 4880 5084 4884 5116
rect 4916 5084 5044 5116
rect 5076 5084 5204 5116
rect 5236 5084 5364 5116
rect 5396 5084 5524 5116
rect 5556 5084 5684 5116
rect 5716 5084 5720 5116
rect 4880 5080 5720 5084
rect -1520 5036 -840 5040
rect -1520 5004 -1516 5036
rect -1484 5004 -1356 5036
rect -1324 5004 -1196 5036
rect -1164 5004 -1036 5036
rect -1004 5004 -876 5036
rect -844 5004 -840 5036
rect -1520 5000 -840 5004
rect -800 5036 4840 5040
rect -800 5004 -796 5036
rect -764 5004 -716 5036
rect -684 5004 -636 5036
rect -604 5004 -556 5036
rect -524 5004 -476 5036
rect -444 5004 -396 5036
rect -364 5004 -316 5036
rect -284 5004 -236 5036
rect -204 5004 -156 5036
rect -124 5004 -76 5036
rect -44 5004 4 5036
rect 36 5004 84 5036
rect 116 5004 164 5036
rect 196 5004 244 5036
rect 276 5004 324 5036
rect 356 5004 404 5036
rect 436 5004 484 5036
rect 516 5004 564 5036
rect 596 5004 644 5036
rect 676 5004 724 5036
rect 756 5004 804 5036
rect 836 5004 884 5036
rect 916 5004 964 5036
rect 996 5004 1044 5036
rect 1076 5004 1124 5036
rect 1156 5004 1204 5036
rect 1236 5004 1284 5036
rect 1316 5004 1364 5036
rect 1396 5004 1444 5036
rect 1476 5004 1524 5036
rect 1556 5004 1604 5036
rect 1636 5004 1684 5036
rect 1716 5004 1764 5036
rect 1796 5004 1844 5036
rect 1876 5004 1924 5036
rect 1956 5004 2004 5036
rect 2036 5004 2084 5036
rect 2116 5004 2164 5036
rect 2196 5004 2244 5036
rect 2276 5004 2324 5036
rect 2356 5004 2404 5036
rect 2436 5004 2484 5036
rect 2516 5004 2564 5036
rect 2596 5004 2644 5036
rect 2676 5004 2724 5036
rect 2756 5004 2804 5036
rect 2836 5004 2884 5036
rect 2916 5004 2964 5036
rect 2996 5004 3044 5036
rect 3076 5004 3124 5036
rect 3156 5004 3204 5036
rect 3236 5004 3284 5036
rect 3316 5004 3364 5036
rect 3396 5004 3444 5036
rect 3476 5004 3524 5036
rect 3556 5004 3604 5036
rect 3636 5004 3684 5036
rect 3716 5004 3764 5036
rect 3796 5004 3844 5036
rect 3876 5004 3924 5036
rect 3956 5004 4004 5036
rect 4036 5004 4084 5036
rect 4116 5004 4164 5036
rect 4196 5004 4244 5036
rect 4276 5004 4324 5036
rect 4356 5004 4404 5036
rect 4436 5004 4484 5036
rect 4516 5004 4564 5036
rect 4596 5004 4644 5036
rect 4676 5004 4724 5036
rect 4756 5004 4804 5036
rect 4836 5004 4840 5036
rect -800 5000 4840 5004
rect 4880 5036 5720 5040
rect 4880 5004 4884 5036
rect 4916 5004 5044 5036
rect 5076 5004 5204 5036
rect 5236 5004 5364 5036
rect 5396 5004 5524 5036
rect 5556 5004 5684 5036
rect 5716 5004 5720 5036
rect 4880 5000 5720 5004
rect -1520 4956 -840 4960
rect -1520 4924 -1516 4956
rect -1484 4924 -1356 4956
rect -1324 4924 -1196 4956
rect -1164 4924 -1036 4956
rect -1004 4924 -876 4956
rect -844 4924 -840 4956
rect -1520 4920 -840 4924
rect -800 4956 4840 4960
rect -800 4924 -796 4956
rect -764 4924 -716 4956
rect -684 4924 -636 4956
rect -604 4924 -556 4956
rect -524 4924 -476 4956
rect -444 4924 -396 4956
rect -364 4924 -316 4956
rect -284 4924 -236 4956
rect -204 4924 -156 4956
rect -124 4924 -76 4956
rect -44 4924 4 4956
rect 36 4924 84 4956
rect 116 4924 164 4956
rect 196 4924 244 4956
rect 276 4924 324 4956
rect 356 4924 404 4956
rect 436 4924 484 4956
rect 516 4924 564 4956
rect 596 4924 644 4956
rect 676 4924 724 4956
rect 756 4924 804 4956
rect 836 4924 884 4956
rect 916 4924 964 4956
rect 996 4924 1044 4956
rect 1076 4924 1124 4956
rect 1156 4924 1204 4956
rect 1236 4924 1284 4956
rect 1316 4924 1364 4956
rect 1396 4924 1444 4956
rect 1476 4924 1524 4956
rect 1556 4924 1604 4956
rect 1636 4924 1684 4956
rect 1716 4924 1764 4956
rect 1796 4924 1844 4956
rect 1876 4924 1924 4956
rect 1956 4924 2004 4956
rect 2036 4924 2084 4956
rect 2116 4924 2164 4956
rect 2196 4924 2244 4956
rect 2276 4924 2324 4956
rect 2356 4924 2404 4956
rect 2436 4924 2484 4956
rect 2516 4924 2564 4956
rect 2596 4924 2644 4956
rect 2676 4924 2724 4956
rect 2756 4924 2804 4956
rect 2836 4924 2884 4956
rect 2916 4924 2964 4956
rect 2996 4924 3044 4956
rect 3076 4924 3124 4956
rect 3156 4924 3204 4956
rect 3236 4924 3284 4956
rect 3316 4924 3364 4956
rect 3396 4924 3444 4956
rect 3476 4924 3524 4956
rect 3556 4924 3604 4956
rect 3636 4924 3684 4956
rect 3716 4924 3764 4956
rect 3796 4924 3844 4956
rect 3876 4924 3924 4956
rect 3956 4924 4004 4956
rect 4036 4924 4084 4956
rect 4116 4924 4164 4956
rect 4196 4924 4244 4956
rect 4276 4924 4324 4956
rect 4356 4924 4404 4956
rect 4436 4924 4484 4956
rect 4516 4924 4564 4956
rect 4596 4924 4644 4956
rect 4676 4924 4724 4956
rect 4756 4924 4804 4956
rect 4836 4924 4840 4956
rect -800 4920 4840 4924
rect 4880 4956 5720 4960
rect 4880 4924 4884 4956
rect 4916 4924 5044 4956
rect 5076 4924 5204 4956
rect 5236 4924 5364 4956
rect 5396 4924 5524 4956
rect 5556 4924 5684 4956
rect 5716 4924 5720 4956
rect 4880 4920 5720 4924
rect -1520 4876 -840 4880
rect -1520 4844 -1516 4876
rect -1484 4844 -1356 4876
rect -1324 4844 -1196 4876
rect -1164 4844 -1036 4876
rect -1004 4844 -876 4876
rect -844 4844 -840 4876
rect -1520 4840 -840 4844
rect -800 4876 4840 4880
rect -800 4844 -796 4876
rect -764 4844 -716 4876
rect -684 4844 -636 4876
rect -604 4844 -556 4876
rect -524 4844 -476 4876
rect -444 4844 -396 4876
rect -364 4844 -316 4876
rect -284 4844 -236 4876
rect -204 4844 -156 4876
rect -124 4844 -76 4876
rect -44 4844 4 4876
rect 36 4844 84 4876
rect 116 4844 164 4876
rect 196 4844 244 4876
rect 276 4844 324 4876
rect 356 4844 404 4876
rect 436 4844 484 4876
rect 516 4844 564 4876
rect 596 4844 644 4876
rect 676 4844 724 4876
rect 756 4844 804 4876
rect 836 4844 884 4876
rect 916 4844 964 4876
rect 996 4844 1044 4876
rect 1076 4844 1124 4876
rect 1156 4844 1204 4876
rect 1236 4844 1284 4876
rect 1316 4844 1364 4876
rect 1396 4844 1444 4876
rect 1476 4844 1524 4876
rect 1556 4844 1604 4876
rect 1636 4844 1684 4876
rect 1716 4844 1764 4876
rect 1796 4844 1844 4876
rect 1876 4844 1924 4876
rect 1956 4844 2004 4876
rect 2036 4844 2084 4876
rect 2116 4844 2164 4876
rect 2196 4844 2244 4876
rect 2276 4844 2324 4876
rect 2356 4844 2404 4876
rect 2436 4844 2484 4876
rect 2516 4844 2564 4876
rect 2596 4844 2644 4876
rect 2676 4844 2724 4876
rect 2756 4844 2804 4876
rect 2836 4844 2884 4876
rect 2916 4844 2964 4876
rect 2996 4844 3044 4876
rect 3076 4844 3124 4876
rect 3156 4844 3204 4876
rect 3236 4844 3284 4876
rect 3316 4844 3364 4876
rect 3396 4844 3444 4876
rect 3476 4844 3524 4876
rect 3556 4844 3604 4876
rect 3636 4844 3684 4876
rect 3716 4844 3764 4876
rect 3796 4844 3844 4876
rect 3876 4844 3924 4876
rect 3956 4844 4004 4876
rect 4036 4844 4084 4876
rect 4116 4844 4164 4876
rect 4196 4844 4244 4876
rect 4276 4844 4324 4876
rect 4356 4844 4404 4876
rect 4436 4844 4484 4876
rect 4516 4844 4564 4876
rect 4596 4844 4644 4876
rect 4676 4844 4724 4876
rect 4756 4844 4804 4876
rect 4836 4844 4840 4876
rect -800 4840 4840 4844
rect 4880 4876 5720 4880
rect 4880 4844 4884 4876
rect 4916 4844 5044 4876
rect 5076 4844 5204 4876
rect 5236 4844 5364 4876
rect 5396 4844 5524 4876
rect 5556 4844 5684 4876
rect 5716 4844 5720 4876
rect 4880 4840 5720 4844
rect -1520 4796 -840 4800
rect -1520 4764 -1516 4796
rect -1484 4764 -1356 4796
rect -1324 4764 -1196 4796
rect -1164 4764 -1036 4796
rect -1004 4764 -876 4796
rect -844 4764 -840 4796
rect -1520 4760 -840 4764
rect -800 4796 4840 4800
rect -800 4764 -796 4796
rect -764 4764 -716 4796
rect -684 4764 -636 4796
rect -604 4764 -556 4796
rect -524 4764 -476 4796
rect -444 4764 -396 4796
rect -364 4764 -316 4796
rect -284 4764 -236 4796
rect -204 4764 -156 4796
rect -124 4764 -76 4796
rect -44 4764 4 4796
rect 36 4764 84 4796
rect 116 4764 164 4796
rect 196 4764 244 4796
rect 276 4764 324 4796
rect 356 4764 404 4796
rect 436 4764 484 4796
rect 516 4764 564 4796
rect 596 4764 644 4796
rect 676 4764 724 4796
rect 756 4764 804 4796
rect 836 4764 884 4796
rect 916 4764 964 4796
rect 996 4764 1044 4796
rect 1076 4764 1124 4796
rect 1156 4764 1204 4796
rect 1236 4764 1284 4796
rect 1316 4764 1364 4796
rect 1396 4764 1444 4796
rect 1476 4764 1524 4796
rect 1556 4764 1604 4796
rect 1636 4764 1684 4796
rect 1716 4764 1764 4796
rect 1796 4764 1844 4796
rect 1876 4764 1924 4796
rect 1956 4764 2004 4796
rect 2036 4764 2084 4796
rect 2116 4764 2164 4796
rect 2196 4764 2244 4796
rect 2276 4764 2324 4796
rect 2356 4764 2404 4796
rect 2436 4764 2484 4796
rect 2516 4764 2564 4796
rect 2596 4764 2644 4796
rect 2676 4764 2724 4796
rect 2756 4764 2804 4796
rect 2836 4764 2884 4796
rect 2916 4764 2964 4796
rect 2996 4764 3044 4796
rect 3076 4764 3124 4796
rect 3156 4764 3204 4796
rect 3236 4764 3284 4796
rect 3316 4764 3364 4796
rect 3396 4764 3444 4796
rect 3476 4764 3524 4796
rect 3556 4764 3604 4796
rect 3636 4764 3684 4796
rect 3716 4764 3764 4796
rect 3796 4764 3844 4796
rect 3876 4764 3924 4796
rect 3956 4764 4004 4796
rect 4036 4764 4084 4796
rect 4116 4764 4164 4796
rect 4196 4764 4244 4796
rect 4276 4764 4324 4796
rect 4356 4764 4404 4796
rect 4436 4764 4484 4796
rect 4516 4764 4564 4796
rect 4596 4764 4644 4796
rect 4676 4764 4724 4796
rect 4756 4764 4804 4796
rect 4836 4764 4840 4796
rect -800 4760 4840 4764
rect 4880 4796 5720 4800
rect 4880 4764 4884 4796
rect 4916 4764 5044 4796
rect 5076 4764 5204 4796
rect 5236 4764 5364 4796
rect 5396 4764 5524 4796
rect 5556 4764 5684 4796
rect 5716 4764 5720 4796
rect 4880 4760 5720 4764
rect -1520 4716 -840 4720
rect -1520 4684 -1516 4716
rect -1484 4684 -1356 4716
rect -1324 4684 -1196 4716
rect -1164 4684 -1036 4716
rect -1004 4684 -876 4716
rect -844 4684 -840 4716
rect -1520 4680 -840 4684
rect -800 4716 4840 4720
rect -800 4684 -796 4716
rect -764 4684 -716 4716
rect -684 4684 -636 4716
rect -604 4684 -556 4716
rect -524 4684 -476 4716
rect -444 4684 -396 4716
rect -364 4684 -316 4716
rect -284 4684 -236 4716
rect -204 4684 -156 4716
rect -124 4684 -76 4716
rect -44 4684 4 4716
rect 36 4684 84 4716
rect 116 4684 164 4716
rect 196 4684 244 4716
rect 276 4684 324 4716
rect 356 4684 404 4716
rect 436 4684 484 4716
rect 516 4684 564 4716
rect 596 4684 644 4716
rect 676 4684 724 4716
rect 756 4684 804 4716
rect 836 4684 884 4716
rect 916 4684 964 4716
rect 996 4684 1044 4716
rect 1076 4684 1124 4716
rect 1156 4684 1204 4716
rect 1236 4684 1284 4716
rect 1316 4684 1364 4716
rect 1396 4684 1444 4716
rect 1476 4684 1524 4716
rect 1556 4684 1604 4716
rect 1636 4684 1684 4716
rect 1716 4684 1764 4716
rect 1796 4684 1844 4716
rect 1876 4684 1924 4716
rect 1956 4684 2004 4716
rect 2036 4684 2084 4716
rect 2116 4684 2164 4716
rect 2196 4684 2244 4716
rect 2276 4684 2324 4716
rect 2356 4684 2404 4716
rect 2436 4684 2484 4716
rect 2516 4684 2564 4716
rect 2596 4684 2644 4716
rect 2676 4684 2724 4716
rect 2756 4684 2804 4716
rect 2836 4684 2884 4716
rect 2916 4684 2964 4716
rect 2996 4684 3044 4716
rect 3076 4684 3124 4716
rect 3156 4684 3204 4716
rect 3236 4684 3284 4716
rect 3316 4684 3364 4716
rect 3396 4684 3444 4716
rect 3476 4684 3524 4716
rect 3556 4684 3604 4716
rect 3636 4684 3684 4716
rect 3716 4684 3764 4716
rect 3796 4684 3844 4716
rect 3876 4684 3924 4716
rect 3956 4684 4004 4716
rect 4036 4684 4084 4716
rect 4116 4684 4164 4716
rect 4196 4684 4244 4716
rect 4276 4684 4324 4716
rect 4356 4684 4404 4716
rect 4436 4684 4484 4716
rect 4516 4684 4564 4716
rect 4596 4684 4644 4716
rect 4676 4684 4724 4716
rect 4756 4684 4804 4716
rect 4836 4684 4840 4716
rect -800 4680 4840 4684
rect 4880 4716 5720 4720
rect 4880 4684 4884 4716
rect 4916 4684 5044 4716
rect 5076 4684 5204 4716
rect 5236 4684 5364 4716
rect 5396 4684 5524 4716
rect 5556 4684 5684 4716
rect 5716 4684 5720 4716
rect 4880 4680 5720 4684
rect -1520 4636 -840 4640
rect -1520 4604 -1516 4636
rect -1484 4604 -1356 4636
rect -1324 4604 -1196 4636
rect -1164 4604 -1036 4636
rect -1004 4604 -876 4636
rect -844 4604 -840 4636
rect -1520 4600 -840 4604
rect -800 4636 4840 4640
rect -800 4604 -796 4636
rect -764 4604 -716 4636
rect -684 4604 -636 4636
rect -604 4604 -556 4636
rect -524 4604 -476 4636
rect -444 4604 -396 4636
rect -364 4604 -316 4636
rect -284 4604 -236 4636
rect -204 4604 -156 4636
rect -124 4604 -76 4636
rect -44 4604 4 4636
rect 36 4604 84 4636
rect 116 4604 164 4636
rect 196 4604 244 4636
rect 276 4604 324 4636
rect 356 4604 404 4636
rect 436 4604 484 4636
rect 516 4604 564 4636
rect 596 4604 644 4636
rect 676 4604 724 4636
rect 756 4604 804 4636
rect 836 4604 884 4636
rect 916 4604 964 4636
rect 996 4604 1044 4636
rect 1076 4604 1124 4636
rect 1156 4604 1204 4636
rect 1236 4604 1284 4636
rect 1316 4604 1364 4636
rect 1396 4604 1444 4636
rect 1476 4604 1524 4636
rect 1556 4604 1604 4636
rect 1636 4604 1684 4636
rect 1716 4604 1764 4636
rect 1796 4604 1844 4636
rect 1876 4604 1924 4636
rect 1956 4604 2004 4636
rect 2036 4604 2084 4636
rect 2116 4604 2164 4636
rect 2196 4604 2244 4636
rect 2276 4604 2324 4636
rect 2356 4604 2404 4636
rect 2436 4604 2484 4636
rect 2516 4604 2564 4636
rect 2596 4604 2644 4636
rect 2676 4604 2724 4636
rect 2756 4604 2804 4636
rect 2836 4604 2884 4636
rect 2916 4604 2964 4636
rect 2996 4604 3044 4636
rect 3076 4604 3124 4636
rect 3156 4604 3204 4636
rect 3236 4604 3284 4636
rect 3316 4604 3364 4636
rect 3396 4604 3444 4636
rect 3476 4604 3524 4636
rect 3556 4604 3604 4636
rect 3636 4604 3684 4636
rect 3716 4604 3764 4636
rect 3796 4604 3844 4636
rect 3876 4604 3924 4636
rect 3956 4604 4004 4636
rect 4036 4604 4084 4636
rect 4116 4604 4164 4636
rect 4196 4604 4244 4636
rect 4276 4604 4324 4636
rect 4356 4604 4404 4636
rect 4436 4604 4484 4636
rect 4516 4604 4564 4636
rect 4596 4604 4644 4636
rect 4676 4604 4724 4636
rect 4756 4604 4804 4636
rect 4836 4604 4840 4636
rect -800 4600 4840 4604
rect 4880 4636 5720 4640
rect 4880 4604 4884 4636
rect 4916 4604 5044 4636
rect 5076 4604 5204 4636
rect 5236 4604 5364 4636
rect 5396 4604 5524 4636
rect 5556 4604 5684 4636
rect 5716 4604 5720 4636
rect 4880 4600 5720 4604
rect -1520 4556 -840 4560
rect -1520 4524 -1516 4556
rect -1484 4524 -1356 4556
rect -1324 4524 -1196 4556
rect -1164 4524 -1036 4556
rect -1004 4524 -876 4556
rect -844 4524 -840 4556
rect -1520 4520 -840 4524
rect -800 4556 4840 4560
rect -800 4524 -796 4556
rect -764 4524 -716 4556
rect -684 4524 -636 4556
rect -604 4524 -556 4556
rect -524 4524 -476 4556
rect -444 4524 -396 4556
rect -364 4524 -316 4556
rect -284 4524 -236 4556
rect -204 4524 -156 4556
rect -124 4524 -76 4556
rect -44 4524 4 4556
rect 36 4524 84 4556
rect 116 4524 164 4556
rect 196 4524 244 4556
rect 276 4524 324 4556
rect 356 4524 404 4556
rect 436 4524 484 4556
rect 516 4524 564 4556
rect 596 4524 644 4556
rect 676 4524 724 4556
rect 756 4524 804 4556
rect 836 4524 884 4556
rect 916 4524 964 4556
rect 996 4524 1044 4556
rect 1076 4524 1124 4556
rect 1156 4524 1204 4556
rect 1236 4524 1284 4556
rect 1316 4524 1364 4556
rect 1396 4524 1444 4556
rect 1476 4524 1524 4556
rect 1556 4524 1604 4556
rect 1636 4524 1684 4556
rect 1716 4524 1764 4556
rect 1796 4524 1844 4556
rect 1876 4524 1924 4556
rect 1956 4524 2004 4556
rect 2036 4524 2084 4556
rect 2116 4524 2164 4556
rect 2196 4524 2244 4556
rect 2276 4524 2324 4556
rect 2356 4524 2404 4556
rect 2436 4524 2484 4556
rect 2516 4524 2564 4556
rect 2596 4524 2644 4556
rect 2676 4524 2724 4556
rect 2756 4524 2804 4556
rect 2836 4524 2884 4556
rect 2916 4524 2964 4556
rect 2996 4524 3044 4556
rect 3076 4524 3124 4556
rect 3156 4524 3204 4556
rect 3236 4524 3284 4556
rect 3316 4524 3364 4556
rect 3396 4524 3444 4556
rect 3476 4524 3524 4556
rect 3556 4524 3604 4556
rect 3636 4524 3684 4556
rect 3716 4524 3764 4556
rect 3796 4524 3844 4556
rect 3876 4524 3924 4556
rect 3956 4524 4004 4556
rect 4036 4524 4084 4556
rect 4116 4524 4164 4556
rect 4196 4524 4244 4556
rect 4276 4524 4324 4556
rect 4356 4524 4404 4556
rect 4436 4524 4484 4556
rect 4516 4524 4564 4556
rect 4596 4524 4644 4556
rect 4676 4524 4724 4556
rect 4756 4524 4804 4556
rect 4836 4524 4840 4556
rect -800 4520 4840 4524
rect 4880 4556 5720 4560
rect 4880 4524 4884 4556
rect 4916 4524 5044 4556
rect 5076 4524 5204 4556
rect 5236 4524 5364 4556
rect 5396 4524 5524 4556
rect 5556 4524 5684 4556
rect 5716 4524 5720 4556
rect 4880 4520 5720 4524
rect -1520 4476 -840 4480
rect -1520 4444 -1516 4476
rect -1484 4444 -1356 4476
rect -1324 4444 -1196 4476
rect -1164 4444 -1036 4476
rect -1004 4444 -876 4476
rect -844 4444 -840 4476
rect -1520 4440 -840 4444
rect -800 4476 4840 4480
rect -800 4444 -796 4476
rect -764 4444 -716 4476
rect -684 4444 -636 4476
rect -604 4444 -556 4476
rect -524 4444 -476 4476
rect -444 4444 -396 4476
rect -364 4444 -316 4476
rect -284 4444 -236 4476
rect -204 4444 -156 4476
rect -124 4444 -76 4476
rect -44 4444 4 4476
rect 36 4444 84 4476
rect 116 4444 164 4476
rect 196 4444 244 4476
rect 276 4444 324 4476
rect 356 4444 404 4476
rect 436 4444 484 4476
rect 516 4444 564 4476
rect 596 4444 644 4476
rect 676 4444 724 4476
rect 756 4444 804 4476
rect 836 4444 884 4476
rect 916 4444 964 4476
rect 996 4444 1044 4476
rect 1076 4444 1124 4476
rect 1156 4444 1204 4476
rect 1236 4444 1284 4476
rect 1316 4444 1364 4476
rect 1396 4444 1444 4476
rect 1476 4444 1524 4476
rect 1556 4444 1604 4476
rect 1636 4444 1684 4476
rect 1716 4444 1764 4476
rect 1796 4444 1844 4476
rect 1876 4444 1924 4476
rect 1956 4444 2004 4476
rect 2036 4444 2084 4476
rect 2116 4444 2164 4476
rect 2196 4444 2244 4476
rect 2276 4444 2324 4476
rect 2356 4444 2404 4476
rect 2436 4444 2484 4476
rect 2516 4444 2564 4476
rect 2596 4444 2644 4476
rect 2676 4444 2724 4476
rect 2756 4444 2804 4476
rect 2836 4444 2884 4476
rect 2916 4444 2964 4476
rect 2996 4444 3044 4476
rect 3076 4444 3124 4476
rect 3156 4444 3204 4476
rect 3236 4444 3284 4476
rect 3316 4444 3364 4476
rect 3396 4444 3444 4476
rect 3476 4444 3524 4476
rect 3556 4444 3604 4476
rect 3636 4444 3684 4476
rect 3716 4444 3764 4476
rect 3796 4444 3844 4476
rect 3876 4444 3924 4476
rect 3956 4444 4004 4476
rect 4036 4444 4084 4476
rect 4116 4444 4164 4476
rect 4196 4444 4244 4476
rect 4276 4444 4324 4476
rect 4356 4444 4404 4476
rect 4436 4444 4484 4476
rect 4516 4444 4564 4476
rect 4596 4444 4644 4476
rect 4676 4444 4724 4476
rect 4756 4444 4804 4476
rect 4836 4444 4840 4476
rect -800 4440 4840 4444
rect 4880 4476 5720 4480
rect 4880 4444 4884 4476
rect 4916 4444 5044 4476
rect 5076 4444 5204 4476
rect 5236 4444 5364 4476
rect 5396 4444 5524 4476
rect 5556 4444 5684 4476
rect 5716 4444 5720 4476
rect 4880 4440 5720 4444
rect -1520 4396 -840 4400
rect -1520 4364 -1516 4396
rect -1484 4364 -1356 4396
rect -1324 4364 -1196 4396
rect -1164 4364 -1036 4396
rect -1004 4364 -876 4396
rect -844 4364 -840 4396
rect -1520 4360 -840 4364
rect -800 4396 4840 4400
rect -800 4364 -796 4396
rect -764 4364 -716 4396
rect -684 4364 -636 4396
rect -604 4364 -556 4396
rect -524 4364 -476 4396
rect -444 4364 -396 4396
rect -364 4364 -316 4396
rect -284 4364 -236 4396
rect -204 4364 -156 4396
rect -124 4364 -76 4396
rect -44 4364 4 4396
rect 36 4364 84 4396
rect 116 4364 164 4396
rect 196 4364 244 4396
rect 276 4364 324 4396
rect 356 4364 404 4396
rect 436 4364 484 4396
rect 516 4364 564 4396
rect 596 4364 644 4396
rect 676 4364 724 4396
rect 756 4364 804 4396
rect 836 4364 884 4396
rect 916 4364 964 4396
rect 996 4364 1044 4396
rect 1076 4364 1124 4396
rect 1156 4364 1204 4396
rect 1236 4364 1284 4396
rect 1316 4364 1364 4396
rect 1396 4364 1444 4396
rect 1476 4364 1524 4396
rect 1556 4364 1604 4396
rect 1636 4364 1684 4396
rect 1716 4364 1764 4396
rect 1796 4364 1844 4396
rect 1876 4364 1924 4396
rect 1956 4364 2004 4396
rect 2036 4364 2084 4396
rect 2116 4364 2164 4396
rect 2196 4364 2244 4396
rect 2276 4364 2324 4396
rect 2356 4364 2404 4396
rect 2436 4364 2484 4396
rect 2516 4364 2564 4396
rect 2596 4364 2644 4396
rect 2676 4364 2724 4396
rect 2756 4364 2804 4396
rect 2836 4364 2884 4396
rect 2916 4364 2964 4396
rect 2996 4364 3044 4396
rect 3076 4364 3124 4396
rect 3156 4364 3204 4396
rect 3236 4364 3284 4396
rect 3316 4364 3364 4396
rect 3396 4364 3444 4396
rect 3476 4364 3524 4396
rect 3556 4364 3604 4396
rect 3636 4364 3684 4396
rect 3716 4364 3764 4396
rect 3796 4364 3844 4396
rect 3876 4364 3924 4396
rect 3956 4364 4004 4396
rect 4036 4364 4084 4396
rect 4116 4364 4164 4396
rect 4196 4364 4244 4396
rect 4276 4364 4324 4396
rect 4356 4364 4404 4396
rect 4436 4364 4484 4396
rect 4516 4364 4564 4396
rect 4596 4364 4644 4396
rect 4676 4364 4724 4396
rect 4756 4364 4804 4396
rect 4836 4364 4840 4396
rect -800 4360 4840 4364
rect 4880 4396 5720 4400
rect 4880 4364 4884 4396
rect 4916 4364 5044 4396
rect 5076 4364 5204 4396
rect 5236 4364 5364 4396
rect 5396 4364 5524 4396
rect 5556 4364 5684 4396
rect 5716 4364 5720 4396
rect 4880 4360 5720 4364
rect -1520 4316 -840 4320
rect -1520 4284 -1516 4316
rect -1484 4284 -1356 4316
rect -1324 4284 -1196 4316
rect -1164 4284 -1036 4316
rect -1004 4284 -876 4316
rect -844 4284 -840 4316
rect -1520 4280 -840 4284
rect -800 4316 4840 4320
rect -800 4284 -796 4316
rect -764 4284 -716 4316
rect -684 4284 -636 4316
rect -604 4284 -556 4316
rect -524 4284 -476 4316
rect -444 4284 -396 4316
rect -364 4284 -316 4316
rect -284 4284 -236 4316
rect -204 4284 -156 4316
rect -124 4284 -76 4316
rect -44 4284 4 4316
rect 36 4284 84 4316
rect 116 4284 164 4316
rect 196 4284 244 4316
rect 276 4284 324 4316
rect 356 4284 404 4316
rect 436 4284 484 4316
rect 516 4284 564 4316
rect 596 4284 644 4316
rect 676 4284 724 4316
rect 756 4284 804 4316
rect 836 4284 884 4316
rect 916 4284 964 4316
rect 996 4284 1044 4316
rect 1076 4284 1124 4316
rect 1156 4284 1204 4316
rect 1236 4284 1284 4316
rect 1316 4284 1364 4316
rect 1396 4284 1444 4316
rect 1476 4284 1524 4316
rect 1556 4284 1604 4316
rect 1636 4284 1684 4316
rect 1716 4284 1764 4316
rect 1796 4284 1844 4316
rect 1876 4284 1924 4316
rect 1956 4284 2004 4316
rect 2036 4284 2084 4316
rect 2116 4284 2164 4316
rect 2196 4284 2244 4316
rect 2276 4284 2324 4316
rect 2356 4284 2404 4316
rect 2436 4284 2484 4316
rect 2516 4284 2564 4316
rect 2596 4284 2644 4316
rect 2676 4284 2724 4316
rect 2756 4284 2804 4316
rect 2836 4284 2884 4316
rect 2916 4284 2964 4316
rect 2996 4284 3044 4316
rect 3076 4284 3124 4316
rect 3156 4284 3204 4316
rect 3236 4284 3284 4316
rect 3316 4284 3364 4316
rect 3396 4284 3444 4316
rect 3476 4284 3524 4316
rect 3556 4284 3604 4316
rect 3636 4284 3684 4316
rect 3716 4284 3764 4316
rect 3796 4284 3844 4316
rect 3876 4284 3924 4316
rect 3956 4284 4004 4316
rect 4036 4284 4084 4316
rect 4116 4284 4164 4316
rect 4196 4284 4244 4316
rect 4276 4284 4324 4316
rect 4356 4284 4404 4316
rect 4436 4284 4484 4316
rect 4516 4284 4564 4316
rect 4596 4284 4644 4316
rect 4676 4284 4724 4316
rect 4756 4284 4804 4316
rect 4836 4284 4840 4316
rect -800 4280 4840 4284
rect 4880 4316 5720 4320
rect 4880 4284 4884 4316
rect 4916 4284 5044 4316
rect 5076 4284 5204 4316
rect 5236 4284 5364 4316
rect 5396 4284 5524 4316
rect 5556 4284 5684 4316
rect 5716 4284 5720 4316
rect 4880 4280 5720 4284
rect -1520 4236 -840 4240
rect -1520 4204 -1516 4236
rect -1484 4204 -1356 4236
rect -1324 4204 -1196 4236
rect -1164 4204 -1036 4236
rect -1004 4204 -876 4236
rect -844 4204 -840 4236
rect -1520 4200 -840 4204
rect -800 4236 4840 4240
rect -800 4204 -796 4236
rect -764 4204 -716 4236
rect -684 4204 -636 4236
rect -604 4204 -556 4236
rect -524 4204 -476 4236
rect -444 4204 -396 4236
rect -364 4204 -316 4236
rect -284 4204 -236 4236
rect -204 4204 -156 4236
rect -124 4204 -76 4236
rect -44 4204 4 4236
rect 36 4204 84 4236
rect 116 4204 164 4236
rect 196 4204 244 4236
rect 276 4204 324 4236
rect 356 4204 404 4236
rect 436 4204 484 4236
rect 516 4204 564 4236
rect 596 4204 644 4236
rect 676 4204 724 4236
rect 756 4204 804 4236
rect 836 4204 884 4236
rect 916 4204 964 4236
rect 996 4204 1044 4236
rect 1076 4204 1124 4236
rect 1156 4204 1204 4236
rect 1236 4204 1284 4236
rect 1316 4204 1364 4236
rect 1396 4204 1444 4236
rect 1476 4204 1524 4236
rect 1556 4204 1604 4236
rect 1636 4204 1684 4236
rect 1716 4204 1764 4236
rect 1796 4204 1844 4236
rect 1876 4204 1924 4236
rect 1956 4204 2004 4236
rect 2036 4204 2084 4236
rect 2116 4204 2164 4236
rect 2196 4204 2244 4236
rect 2276 4204 2324 4236
rect 2356 4204 2404 4236
rect 2436 4204 2484 4236
rect 2516 4204 2564 4236
rect 2596 4204 2644 4236
rect 2676 4204 2724 4236
rect 2756 4204 2804 4236
rect 2836 4204 2884 4236
rect 2916 4204 2964 4236
rect 2996 4204 3044 4236
rect 3076 4204 3124 4236
rect 3156 4204 3204 4236
rect 3236 4204 3284 4236
rect 3316 4204 3364 4236
rect 3396 4204 3444 4236
rect 3476 4204 3524 4236
rect 3556 4204 3604 4236
rect 3636 4204 3684 4236
rect 3716 4204 3764 4236
rect 3796 4204 3844 4236
rect 3876 4204 3924 4236
rect 3956 4204 4004 4236
rect 4036 4204 4084 4236
rect 4116 4204 4164 4236
rect 4196 4204 4244 4236
rect 4276 4204 4324 4236
rect 4356 4204 4404 4236
rect 4436 4204 4484 4236
rect 4516 4204 4564 4236
rect 4596 4204 4644 4236
rect 4676 4204 4724 4236
rect 4756 4204 4804 4236
rect 4836 4204 4840 4236
rect -800 4200 4840 4204
rect 4880 4236 5720 4240
rect 4880 4204 4884 4236
rect 4916 4204 5044 4236
rect 5076 4204 5204 4236
rect 5236 4204 5364 4236
rect 5396 4204 5524 4236
rect 5556 4204 5684 4236
rect 5716 4204 5720 4236
rect 4880 4200 5720 4204
rect -1520 4156 -840 4160
rect -1520 4124 -1516 4156
rect -1484 4124 -1356 4156
rect -1324 4124 -1196 4156
rect -1164 4124 -1036 4156
rect -1004 4124 -876 4156
rect -844 4124 -840 4156
rect -1520 4120 -840 4124
rect -800 4156 4840 4160
rect -800 4124 -796 4156
rect -764 4124 -716 4156
rect -684 4124 -636 4156
rect -604 4124 -556 4156
rect -524 4124 -476 4156
rect -444 4124 -396 4156
rect -364 4124 -316 4156
rect -284 4124 -236 4156
rect -204 4124 -156 4156
rect -124 4124 -76 4156
rect -44 4124 4 4156
rect 36 4124 84 4156
rect 116 4124 164 4156
rect 196 4124 244 4156
rect 276 4124 324 4156
rect 356 4124 404 4156
rect 436 4124 484 4156
rect 516 4124 564 4156
rect 596 4124 644 4156
rect 676 4124 724 4156
rect 756 4124 804 4156
rect 836 4124 884 4156
rect 916 4124 964 4156
rect 996 4124 1044 4156
rect 1076 4124 1124 4156
rect 1156 4124 1204 4156
rect 1236 4124 1284 4156
rect 1316 4124 1364 4156
rect 1396 4124 1444 4156
rect 1476 4124 1524 4156
rect 1556 4124 1604 4156
rect 1636 4124 1684 4156
rect 1716 4124 1764 4156
rect 1796 4124 1844 4156
rect 1876 4124 1924 4156
rect 1956 4124 2004 4156
rect 2036 4124 2084 4156
rect 2116 4124 2164 4156
rect 2196 4124 2244 4156
rect 2276 4124 2324 4156
rect 2356 4124 2404 4156
rect 2436 4124 2484 4156
rect 2516 4124 2564 4156
rect 2596 4124 2644 4156
rect 2676 4124 2724 4156
rect 2756 4124 2804 4156
rect 2836 4124 2884 4156
rect 2916 4124 2964 4156
rect 2996 4124 3044 4156
rect 3076 4124 3124 4156
rect 3156 4124 3204 4156
rect 3236 4124 3284 4156
rect 3316 4124 3364 4156
rect 3396 4124 3444 4156
rect 3476 4124 3524 4156
rect 3556 4124 3604 4156
rect 3636 4124 3684 4156
rect 3716 4124 3764 4156
rect 3796 4124 3844 4156
rect 3876 4124 3924 4156
rect 3956 4124 4004 4156
rect 4036 4124 4084 4156
rect 4116 4124 4164 4156
rect 4196 4124 4244 4156
rect 4276 4124 4324 4156
rect 4356 4124 4404 4156
rect 4436 4124 4484 4156
rect 4516 4124 4564 4156
rect 4596 4124 4644 4156
rect 4676 4124 4724 4156
rect 4756 4124 4804 4156
rect 4836 4124 4840 4156
rect -800 4120 4840 4124
rect 4880 4156 5720 4160
rect 4880 4124 4884 4156
rect 4916 4124 5044 4156
rect 5076 4124 5204 4156
rect 5236 4124 5364 4156
rect 5396 4124 5524 4156
rect 5556 4124 5684 4156
rect 5716 4124 5720 4156
rect 4880 4120 5720 4124
rect -1520 4076 -840 4080
rect -1520 4044 -1516 4076
rect -1484 4044 -1356 4076
rect -1324 4044 -1196 4076
rect -1164 4044 -1036 4076
rect -1004 4044 -876 4076
rect -844 4044 -840 4076
rect -1520 4040 -840 4044
rect -800 4076 4840 4080
rect -800 4044 -796 4076
rect -764 4044 -716 4076
rect -684 4044 -636 4076
rect -604 4044 -556 4076
rect -524 4044 -476 4076
rect -444 4044 -396 4076
rect -364 4044 -316 4076
rect -284 4044 -236 4076
rect -204 4044 -156 4076
rect -124 4044 -76 4076
rect -44 4044 4 4076
rect 36 4044 84 4076
rect 116 4044 164 4076
rect 196 4044 244 4076
rect 276 4044 324 4076
rect 356 4044 404 4076
rect 436 4044 484 4076
rect 516 4044 564 4076
rect 596 4044 644 4076
rect 676 4044 724 4076
rect 756 4044 804 4076
rect 836 4044 884 4076
rect 916 4044 964 4076
rect 996 4044 1044 4076
rect 1076 4044 1124 4076
rect 1156 4044 1204 4076
rect 1236 4044 1284 4076
rect 1316 4044 1364 4076
rect 1396 4044 1444 4076
rect 1476 4044 1524 4076
rect 1556 4044 1604 4076
rect 1636 4044 1684 4076
rect 1716 4044 1764 4076
rect 1796 4044 1844 4076
rect 1876 4044 1924 4076
rect 1956 4044 2004 4076
rect 2036 4044 2084 4076
rect 2116 4044 2164 4076
rect 2196 4044 2244 4076
rect 2276 4044 2324 4076
rect 2356 4044 2404 4076
rect 2436 4044 2484 4076
rect 2516 4044 2564 4076
rect 2596 4044 2644 4076
rect 2676 4044 2724 4076
rect 2756 4044 2804 4076
rect 2836 4044 2884 4076
rect 2916 4044 2964 4076
rect 2996 4044 3044 4076
rect 3076 4044 3124 4076
rect 3156 4044 3204 4076
rect 3236 4044 3284 4076
rect 3316 4044 3364 4076
rect 3396 4044 3444 4076
rect 3476 4044 3524 4076
rect 3556 4044 3604 4076
rect 3636 4044 3684 4076
rect 3716 4044 3764 4076
rect 3796 4044 3844 4076
rect 3876 4044 3924 4076
rect 3956 4044 4004 4076
rect 4036 4044 4084 4076
rect 4116 4044 4164 4076
rect 4196 4044 4244 4076
rect 4276 4044 4324 4076
rect 4356 4044 4404 4076
rect 4436 4044 4484 4076
rect 4516 4044 4564 4076
rect 4596 4044 4644 4076
rect 4676 4044 4724 4076
rect 4756 4044 4804 4076
rect 4836 4044 4840 4076
rect -800 4040 4840 4044
rect 4880 4076 5720 4080
rect 4880 4044 4884 4076
rect 4916 4044 5044 4076
rect 5076 4044 5204 4076
rect 5236 4044 5364 4076
rect 5396 4044 5524 4076
rect 5556 4044 5684 4076
rect 5716 4044 5720 4076
rect 4880 4040 5720 4044
rect -1520 3996 -840 4000
rect -1520 3964 -1516 3996
rect -1484 3964 -1356 3996
rect -1324 3964 -1196 3996
rect -1164 3964 -1036 3996
rect -1004 3964 -876 3996
rect -844 3964 -840 3996
rect -1520 3960 -840 3964
rect -800 3996 4840 4000
rect -800 3964 -796 3996
rect -764 3964 -716 3996
rect -684 3964 -636 3996
rect -604 3964 -556 3996
rect -524 3964 -476 3996
rect -444 3964 -396 3996
rect -364 3964 -316 3996
rect -284 3964 -236 3996
rect -204 3964 -156 3996
rect -124 3964 -76 3996
rect -44 3964 4 3996
rect 36 3964 84 3996
rect 116 3964 164 3996
rect 196 3964 244 3996
rect 276 3964 324 3996
rect 356 3964 404 3996
rect 436 3964 484 3996
rect 516 3964 564 3996
rect 596 3964 644 3996
rect 676 3964 724 3996
rect 756 3964 804 3996
rect 836 3964 884 3996
rect 916 3964 964 3996
rect 996 3964 1044 3996
rect 1076 3964 1124 3996
rect 1156 3964 1204 3996
rect 1236 3964 1284 3996
rect 1316 3964 1364 3996
rect 1396 3964 1444 3996
rect 1476 3964 1524 3996
rect 1556 3964 1604 3996
rect 1636 3964 1684 3996
rect 1716 3964 1764 3996
rect 1796 3964 1844 3996
rect 1876 3964 1924 3996
rect 1956 3964 2004 3996
rect 2036 3964 2084 3996
rect 2116 3964 2164 3996
rect 2196 3964 2244 3996
rect 2276 3964 2324 3996
rect 2356 3964 2404 3996
rect 2436 3964 2484 3996
rect 2516 3964 2564 3996
rect 2596 3964 2644 3996
rect 2676 3964 2724 3996
rect 2756 3964 2804 3996
rect 2836 3964 2884 3996
rect 2916 3964 2964 3996
rect 2996 3964 3044 3996
rect 3076 3964 3124 3996
rect 3156 3964 3204 3996
rect 3236 3964 3284 3996
rect 3316 3964 3364 3996
rect 3396 3964 3444 3996
rect 3476 3964 3524 3996
rect 3556 3964 3604 3996
rect 3636 3964 3684 3996
rect 3716 3964 3764 3996
rect 3796 3964 3844 3996
rect 3876 3964 3924 3996
rect 3956 3964 4004 3996
rect 4036 3964 4084 3996
rect 4116 3964 4164 3996
rect 4196 3964 4244 3996
rect 4276 3964 4324 3996
rect 4356 3964 4404 3996
rect 4436 3964 4484 3996
rect 4516 3964 4564 3996
rect 4596 3964 4644 3996
rect 4676 3964 4724 3996
rect 4756 3964 4804 3996
rect 4836 3964 4840 3996
rect -800 3960 4840 3964
rect 4880 3996 5720 4000
rect 4880 3964 4884 3996
rect 4916 3964 5044 3996
rect 5076 3964 5204 3996
rect 5236 3964 5364 3996
rect 5396 3964 5524 3996
rect 5556 3964 5684 3996
rect 5716 3964 5720 3996
rect 4880 3960 5720 3964
rect -1520 3916 -840 3920
rect -1520 3884 -1516 3916
rect -1484 3884 -1356 3916
rect -1324 3884 -1196 3916
rect -1164 3884 -1036 3916
rect -1004 3884 -876 3916
rect -844 3884 -840 3916
rect -1520 3880 -840 3884
rect -800 3916 4840 3920
rect -800 3884 -796 3916
rect -764 3884 -716 3916
rect -684 3884 -636 3916
rect -604 3884 -556 3916
rect -524 3884 -476 3916
rect -444 3884 -396 3916
rect -364 3884 -316 3916
rect -284 3884 -236 3916
rect -204 3884 -156 3916
rect -124 3884 -76 3916
rect -44 3884 4 3916
rect 36 3884 84 3916
rect 116 3884 164 3916
rect 196 3884 244 3916
rect 276 3884 324 3916
rect 356 3884 404 3916
rect 436 3884 484 3916
rect 516 3884 564 3916
rect 596 3884 644 3916
rect 676 3884 724 3916
rect 756 3884 804 3916
rect 836 3884 884 3916
rect 916 3884 964 3916
rect 996 3884 1044 3916
rect 1076 3884 1124 3916
rect 1156 3884 1204 3916
rect 1236 3884 1284 3916
rect 1316 3884 1364 3916
rect 1396 3884 1444 3916
rect 1476 3884 1524 3916
rect 1556 3884 1604 3916
rect 1636 3884 1684 3916
rect 1716 3884 1764 3916
rect 1796 3884 1844 3916
rect 1876 3884 1924 3916
rect 1956 3884 2004 3916
rect 2036 3884 2084 3916
rect 2116 3884 2164 3916
rect 2196 3884 2244 3916
rect 2276 3884 2324 3916
rect 2356 3884 2404 3916
rect 2436 3884 2484 3916
rect 2516 3884 2564 3916
rect 2596 3884 2644 3916
rect 2676 3884 2724 3916
rect 2756 3884 2804 3916
rect 2836 3884 2884 3916
rect 2916 3884 2964 3916
rect 2996 3884 3044 3916
rect 3076 3884 3124 3916
rect 3156 3884 3204 3916
rect 3236 3884 3284 3916
rect 3316 3884 3364 3916
rect 3396 3884 3444 3916
rect 3476 3884 3524 3916
rect 3556 3884 3604 3916
rect 3636 3884 3684 3916
rect 3716 3884 3764 3916
rect 3796 3884 3844 3916
rect 3876 3884 3924 3916
rect 3956 3884 4004 3916
rect 4036 3884 4084 3916
rect 4116 3884 4164 3916
rect 4196 3884 4244 3916
rect 4276 3884 4324 3916
rect 4356 3884 4404 3916
rect 4436 3884 4484 3916
rect 4516 3884 4564 3916
rect 4596 3884 4644 3916
rect 4676 3884 4724 3916
rect 4756 3884 4804 3916
rect 4836 3884 4840 3916
rect -800 3880 4840 3884
rect 4880 3916 5720 3920
rect 4880 3884 4884 3916
rect 4916 3884 5044 3916
rect 5076 3884 5204 3916
rect 5236 3884 5364 3916
rect 5396 3884 5524 3916
rect 5556 3884 5684 3916
rect 5716 3884 5720 3916
rect 4880 3880 5720 3884
rect -1520 3836 -840 3840
rect -1520 3804 -1516 3836
rect -1484 3804 -1356 3836
rect -1324 3804 -1196 3836
rect -1164 3804 -1036 3836
rect -1004 3804 -876 3836
rect -844 3804 -840 3836
rect -1520 3800 -840 3804
rect -800 3836 4840 3840
rect -800 3804 -796 3836
rect -764 3804 -716 3836
rect -684 3804 -636 3836
rect -604 3804 -556 3836
rect -524 3804 -476 3836
rect -444 3804 -396 3836
rect -364 3804 -316 3836
rect -284 3804 -236 3836
rect -204 3804 -156 3836
rect -124 3804 -76 3836
rect -44 3804 4 3836
rect 36 3804 84 3836
rect 116 3804 164 3836
rect 196 3804 244 3836
rect 276 3804 324 3836
rect 356 3804 404 3836
rect 436 3804 484 3836
rect 516 3804 564 3836
rect 596 3804 644 3836
rect 676 3804 724 3836
rect 756 3804 804 3836
rect 836 3804 884 3836
rect 916 3804 964 3836
rect 996 3804 1044 3836
rect 1076 3804 1124 3836
rect 1156 3804 1204 3836
rect 1236 3804 1284 3836
rect 1316 3804 1364 3836
rect 1396 3804 1444 3836
rect 1476 3804 1524 3836
rect 1556 3804 1604 3836
rect 1636 3804 1684 3836
rect 1716 3804 1764 3836
rect 1796 3804 1844 3836
rect 1876 3804 1924 3836
rect 1956 3804 2004 3836
rect 2036 3804 2084 3836
rect 2116 3804 2164 3836
rect 2196 3804 2244 3836
rect 2276 3804 2324 3836
rect 2356 3804 2404 3836
rect 2436 3804 2484 3836
rect 2516 3804 2564 3836
rect 2596 3804 2644 3836
rect 2676 3804 2724 3836
rect 2756 3804 2804 3836
rect 2836 3804 2884 3836
rect 2916 3804 2964 3836
rect 2996 3804 3044 3836
rect 3076 3804 3124 3836
rect 3156 3804 3204 3836
rect 3236 3804 3284 3836
rect 3316 3804 3364 3836
rect 3396 3804 3444 3836
rect 3476 3804 3524 3836
rect 3556 3804 3604 3836
rect 3636 3804 3684 3836
rect 3716 3804 3764 3836
rect 3796 3804 3844 3836
rect 3876 3804 3924 3836
rect 3956 3804 4004 3836
rect 4036 3804 4084 3836
rect 4116 3804 4164 3836
rect 4196 3804 4244 3836
rect 4276 3804 4324 3836
rect 4356 3804 4404 3836
rect 4436 3804 4484 3836
rect 4516 3804 4564 3836
rect 4596 3804 4644 3836
rect 4676 3804 4724 3836
rect 4756 3804 4804 3836
rect 4836 3804 4840 3836
rect -800 3800 4840 3804
rect 4880 3836 5720 3840
rect 4880 3804 4884 3836
rect 4916 3804 5044 3836
rect 5076 3804 5204 3836
rect 5236 3804 5364 3836
rect 5396 3804 5524 3836
rect 5556 3804 5684 3836
rect 5716 3804 5720 3836
rect 4880 3800 5720 3804
rect -1520 3756 -840 3760
rect -1520 3724 -1516 3756
rect -1484 3724 -1356 3756
rect -1324 3724 -1196 3756
rect -1164 3724 -1036 3756
rect -1004 3724 -876 3756
rect -844 3724 -840 3756
rect -1520 3720 -840 3724
rect -800 3756 4840 3760
rect -800 3724 -796 3756
rect -764 3724 -716 3756
rect -684 3724 -636 3756
rect -604 3724 -556 3756
rect -524 3724 -476 3756
rect -444 3724 -396 3756
rect -364 3724 -316 3756
rect -284 3724 -236 3756
rect -204 3724 -156 3756
rect -124 3724 -76 3756
rect -44 3724 4 3756
rect 36 3724 84 3756
rect 116 3724 164 3756
rect 196 3724 244 3756
rect 276 3724 324 3756
rect 356 3724 404 3756
rect 436 3724 484 3756
rect 516 3724 564 3756
rect 596 3724 644 3756
rect 676 3724 724 3756
rect 756 3724 804 3756
rect 836 3724 884 3756
rect 916 3724 964 3756
rect 996 3724 1044 3756
rect 1076 3724 1124 3756
rect 1156 3724 1204 3756
rect 1236 3724 1284 3756
rect 1316 3724 1364 3756
rect 1396 3724 1444 3756
rect 1476 3724 1524 3756
rect 1556 3724 1604 3756
rect 1636 3724 1684 3756
rect 1716 3724 1764 3756
rect 1796 3724 1844 3756
rect 1876 3724 1924 3756
rect 1956 3724 2004 3756
rect 2036 3724 2084 3756
rect 2116 3724 2164 3756
rect 2196 3724 2244 3756
rect 2276 3724 2324 3756
rect 2356 3724 2404 3756
rect 2436 3724 2484 3756
rect 2516 3724 2564 3756
rect 2596 3724 2644 3756
rect 2676 3724 2724 3756
rect 2756 3724 2804 3756
rect 2836 3724 2884 3756
rect 2916 3724 2964 3756
rect 2996 3724 3044 3756
rect 3076 3724 3124 3756
rect 3156 3724 3204 3756
rect 3236 3724 3284 3756
rect 3316 3724 3364 3756
rect 3396 3724 3444 3756
rect 3476 3724 3524 3756
rect 3556 3724 3604 3756
rect 3636 3724 3684 3756
rect 3716 3724 3764 3756
rect 3796 3724 3844 3756
rect 3876 3724 3924 3756
rect 3956 3724 4004 3756
rect 4036 3724 4084 3756
rect 4116 3724 4164 3756
rect 4196 3724 4244 3756
rect 4276 3724 4324 3756
rect 4356 3724 4404 3756
rect 4436 3724 4484 3756
rect 4516 3724 4564 3756
rect 4596 3724 4644 3756
rect 4676 3724 4724 3756
rect 4756 3724 4804 3756
rect 4836 3724 4840 3756
rect -800 3720 4840 3724
rect 4880 3756 5720 3760
rect 4880 3724 4884 3756
rect 4916 3724 5044 3756
rect 5076 3724 5204 3756
rect 5236 3724 5364 3756
rect 5396 3724 5524 3756
rect 5556 3724 5684 3756
rect 5716 3724 5720 3756
rect 4880 3720 5720 3724
rect -1520 3676 -840 3680
rect -1520 3644 -1516 3676
rect -1484 3644 -1356 3676
rect -1324 3644 -1196 3676
rect -1164 3644 -1036 3676
rect -1004 3644 -876 3676
rect -844 3644 -840 3676
rect -1520 3640 -840 3644
rect -800 3676 4840 3680
rect -800 3644 -796 3676
rect -764 3644 -716 3676
rect -684 3644 -636 3676
rect -604 3644 -556 3676
rect -524 3644 -476 3676
rect -444 3644 -396 3676
rect -364 3644 -316 3676
rect -284 3644 -236 3676
rect -204 3644 -156 3676
rect -124 3644 -76 3676
rect -44 3644 4 3676
rect 36 3644 84 3676
rect 116 3644 164 3676
rect 196 3644 244 3676
rect 276 3644 324 3676
rect 356 3644 404 3676
rect 436 3644 484 3676
rect 516 3644 564 3676
rect 596 3644 644 3676
rect 676 3644 724 3676
rect 756 3644 804 3676
rect 836 3644 884 3676
rect 916 3644 964 3676
rect 996 3644 1044 3676
rect 1076 3644 1124 3676
rect 1156 3644 1204 3676
rect 1236 3644 1284 3676
rect 1316 3644 1364 3676
rect 1396 3644 1444 3676
rect 1476 3644 1524 3676
rect 1556 3644 1604 3676
rect 1636 3644 1684 3676
rect 1716 3644 1764 3676
rect 1796 3644 1844 3676
rect 1876 3644 1924 3676
rect 1956 3644 2004 3676
rect 2036 3644 2084 3676
rect 2116 3644 2164 3676
rect 2196 3644 2244 3676
rect 2276 3644 2324 3676
rect 2356 3644 2404 3676
rect 2436 3644 2484 3676
rect 2516 3644 2564 3676
rect 2596 3644 2644 3676
rect 2676 3644 2724 3676
rect 2756 3644 2804 3676
rect 2836 3644 2884 3676
rect 2916 3644 2964 3676
rect 2996 3644 3044 3676
rect 3076 3644 3124 3676
rect 3156 3644 3204 3676
rect 3236 3644 3284 3676
rect 3316 3644 3364 3676
rect 3396 3644 3444 3676
rect 3476 3644 3524 3676
rect 3556 3644 3604 3676
rect 3636 3644 3684 3676
rect 3716 3644 3764 3676
rect 3796 3644 3844 3676
rect 3876 3644 3924 3676
rect 3956 3644 4004 3676
rect 4036 3644 4084 3676
rect 4116 3644 4164 3676
rect 4196 3644 4244 3676
rect 4276 3644 4324 3676
rect 4356 3644 4404 3676
rect 4436 3644 4484 3676
rect 4516 3644 4564 3676
rect 4596 3644 4644 3676
rect 4676 3644 4724 3676
rect 4756 3644 4804 3676
rect 4836 3644 4840 3676
rect -800 3640 4840 3644
rect 4880 3676 5720 3680
rect 4880 3644 4884 3676
rect 4916 3644 5044 3676
rect 5076 3644 5204 3676
rect 5236 3644 5364 3676
rect 5396 3644 5524 3676
rect 5556 3644 5684 3676
rect 5716 3644 5720 3676
rect 4880 3640 5720 3644
rect -1520 3596 -840 3600
rect -1520 3564 -1516 3596
rect -1484 3564 -1356 3596
rect -1324 3564 -1196 3596
rect -1164 3564 -1036 3596
rect -1004 3564 -876 3596
rect -844 3564 -840 3596
rect -1520 3560 -840 3564
rect -800 3596 4840 3600
rect -800 3564 -796 3596
rect -764 3564 -716 3596
rect -684 3564 -636 3596
rect -604 3564 -556 3596
rect -524 3564 -476 3596
rect -444 3564 -396 3596
rect -364 3564 -316 3596
rect -284 3564 -236 3596
rect -204 3564 -156 3596
rect -124 3564 -76 3596
rect -44 3564 4 3596
rect 36 3564 84 3596
rect 116 3564 164 3596
rect 196 3564 244 3596
rect 276 3564 324 3596
rect 356 3564 404 3596
rect 436 3564 484 3596
rect 516 3564 564 3596
rect 596 3564 644 3596
rect 676 3564 724 3596
rect 756 3564 804 3596
rect 836 3564 884 3596
rect 916 3564 964 3596
rect 996 3564 1044 3596
rect 1076 3564 1124 3596
rect 1156 3564 1204 3596
rect 1236 3564 1284 3596
rect 1316 3564 1364 3596
rect 1396 3564 1444 3596
rect 1476 3564 1524 3596
rect 1556 3564 1604 3596
rect 1636 3564 1684 3596
rect 1716 3564 1764 3596
rect 1796 3564 1844 3596
rect 1876 3564 1924 3596
rect 1956 3564 2004 3596
rect 2036 3564 2084 3596
rect 2116 3564 2164 3596
rect 2196 3564 2244 3596
rect 2276 3564 2324 3596
rect 2356 3564 2404 3596
rect 2436 3564 2484 3596
rect 2516 3564 2564 3596
rect 2596 3564 2644 3596
rect 2676 3564 2724 3596
rect 2756 3564 2804 3596
rect 2836 3564 2884 3596
rect 2916 3564 2964 3596
rect 2996 3564 3044 3596
rect 3076 3564 3124 3596
rect 3156 3564 3204 3596
rect 3236 3564 3284 3596
rect 3316 3564 3364 3596
rect 3396 3564 3444 3596
rect 3476 3564 3524 3596
rect 3556 3564 3604 3596
rect 3636 3564 3684 3596
rect 3716 3564 3764 3596
rect 3796 3564 3844 3596
rect 3876 3564 3924 3596
rect 3956 3564 4004 3596
rect 4036 3564 4084 3596
rect 4116 3564 4164 3596
rect 4196 3564 4244 3596
rect 4276 3564 4324 3596
rect 4356 3564 4404 3596
rect 4436 3564 4484 3596
rect 4516 3564 4564 3596
rect 4596 3564 4644 3596
rect 4676 3564 4724 3596
rect 4756 3564 4804 3596
rect 4836 3564 4840 3596
rect -800 3560 4840 3564
rect 4880 3596 5720 3600
rect 4880 3564 4884 3596
rect 4916 3564 5044 3596
rect 5076 3564 5204 3596
rect 5236 3564 5364 3596
rect 5396 3564 5524 3596
rect 5556 3564 5684 3596
rect 5716 3564 5720 3596
rect 4880 3560 5720 3564
rect -1520 3516 -840 3520
rect -1520 3484 -1516 3516
rect -1484 3484 -1356 3516
rect -1324 3484 -1196 3516
rect -1164 3484 -1036 3516
rect -1004 3484 -876 3516
rect -844 3484 -840 3516
rect -1520 3480 -840 3484
rect -800 3516 4840 3520
rect -800 3484 -796 3516
rect -764 3484 -716 3516
rect -684 3484 -636 3516
rect -604 3484 -556 3516
rect -524 3484 -476 3516
rect -444 3484 -396 3516
rect -364 3484 -316 3516
rect -284 3484 -236 3516
rect -204 3484 -156 3516
rect -124 3484 -76 3516
rect -44 3484 4 3516
rect 36 3484 84 3516
rect 116 3484 164 3516
rect 196 3484 244 3516
rect 276 3484 324 3516
rect 356 3484 404 3516
rect 436 3484 484 3516
rect 516 3484 564 3516
rect 596 3484 644 3516
rect 676 3484 724 3516
rect 756 3484 804 3516
rect 836 3484 884 3516
rect 916 3484 964 3516
rect 996 3484 1044 3516
rect 1076 3484 1124 3516
rect 1156 3484 1204 3516
rect 1236 3484 1284 3516
rect 1316 3484 1364 3516
rect 1396 3484 1444 3516
rect 1476 3484 1524 3516
rect 1556 3484 1604 3516
rect 1636 3484 1684 3516
rect 1716 3484 1764 3516
rect 1796 3484 1844 3516
rect 1876 3484 1924 3516
rect 1956 3484 2004 3516
rect 2036 3484 2084 3516
rect 2116 3484 2164 3516
rect 2196 3484 2244 3516
rect 2276 3484 2324 3516
rect 2356 3484 2404 3516
rect 2436 3484 2484 3516
rect 2516 3484 2564 3516
rect 2596 3484 2644 3516
rect 2676 3484 2724 3516
rect 2756 3484 2804 3516
rect 2836 3484 2884 3516
rect 2916 3484 2964 3516
rect 2996 3484 3044 3516
rect 3076 3484 3124 3516
rect 3156 3484 3204 3516
rect 3236 3484 3284 3516
rect 3316 3484 3364 3516
rect 3396 3484 3444 3516
rect 3476 3484 3524 3516
rect 3556 3484 3604 3516
rect 3636 3484 3684 3516
rect 3716 3484 3764 3516
rect 3796 3484 3844 3516
rect 3876 3484 3924 3516
rect 3956 3484 4004 3516
rect 4036 3484 4084 3516
rect 4116 3484 4164 3516
rect 4196 3484 4244 3516
rect 4276 3484 4324 3516
rect 4356 3484 4404 3516
rect 4436 3484 4484 3516
rect 4516 3484 4564 3516
rect 4596 3484 4644 3516
rect 4676 3484 4724 3516
rect 4756 3484 4804 3516
rect 4836 3484 4840 3516
rect -800 3480 4840 3484
rect 4880 3516 5720 3520
rect 4880 3484 4884 3516
rect 4916 3484 5044 3516
rect 5076 3484 5204 3516
rect 5236 3484 5364 3516
rect 5396 3484 5524 3516
rect 5556 3484 5684 3516
rect 5716 3484 5720 3516
rect 4880 3480 5720 3484
rect -1520 3436 -840 3440
rect -1520 3404 -1516 3436
rect -1484 3404 -1356 3436
rect -1324 3404 -1196 3436
rect -1164 3404 -1036 3436
rect -1004 3404 -876 3436
rect -844 3404 -840 3436
rect -1520 3400 -840 3404
rect -800 3436 4840 3440
rect -800 3404 -796 3436
rect -764 3404 -716 3436
rect -684 3404 -636 3436
rect -604 3404 -556 3436
rect -524 3404 -476 3436
rect -444 3404 -396 3436
rect -364 3404 -316 3436
rect -284 3404 -236 3436
rect -204 3404 -156 3436
rect -124 3404 -76 3436
rect -44 3404 4 3436
rect 36 3404 84 3436
rect 116 3404 164 3436
rect 196 3404 244 3436
rect 276 3404 324 3436
rect 356 3404 404 3436
rect 436 3404 484 3436
rect 516 3404 564 3436
rect 596 3404 644 3436
rect 676 3404 724 3436
rect 756 3404 804 3436
rect 836 3404 884 3436
rect 916 3404 964 3436
rect 996 3404 1044 3436
rect 1076 3404 1124 3436
rect 1156 3404 1204 3436
rect 1236 3404 1284 3436
rect 1316 3404 1364 3436
rect 1396 3404 1444 3436
rect 1476 3404 1524 3436
rect 1556 3404 1604 3436
rect 1636 3404 1684 3436
rect 1716 3404 1764 3436
rect 1796 3404 1844 3436
rect 1876 3404 1924 3436
rect 1956 3404 2004 3436
rect 2036 3404 2084 3436
rect 2116 3404 2164 3436
rect 2196 3404 2244 3436
rect 2276 3404 2324 3436
rect 2356 3404 2404 3436
rect 2436 3404 2484 3436
rect 2516 3404 2564 3436
rect 2596 3404 2644 3436
rect 2676 3404 2724 3436
rect 2756 3404 2804 3436
rect 2836 3404 2884 3436
rect 2916 3404 2964 3436
rect 2996 3404 3044 3436
rect 3076 3404 3124 3436
rect 3156 3404 3204 3436
rect 3236 3404 3284 3436
rect 3316 3404 3364 3436
rect 3396 3404 3444 3436
rect 3476 3404 3524 3436
rect 3556 3404 3604 3436
rect 3636 3404 3684 3436
rect 3716 3404 3764 3436
rect 3796 3404 3844 3436
rect 3876 3404 3924 3436
rect 3956 3404 4004 3436
rect 4036 3404 4084 3436
rect 4116 3404 4164 3436
rect 4196 3404 4244 3436
rect 4276 3404 4324 3436
rect 4356 3404 4404 3436
rect 4436 3404 4484 3436
rect 4516 3404 4564 3436
rect 4596 3404 4644 3436
rect 4676 3404 4724 3436
rect 4756 3404 4804 3436
rect 4836 3404 4840 3436
rect -800 3400 4840 3404
rect 4880 3436 5720 3440
rect 4880 3404 4884 3436
rect 4916 3404 5044 3436
rect 5076 3404 5204 3436
rect 5236 3404 5364 3436
rect 5396 3404 5524 3436
rect 5556 3404 5684 3436
rect 5716 3404 5720 3436
rect 4880 3400 5720 3404
rect -1520 3356 -840 3360
rect -1520 3324 -1516 3356
rect -1484 3324 -1356 3356
rect -1324 3324 -1196 3356
rect -1164 3324 -1036 3356
rect -1004 3324 -876 3356
rect -844 3324 -840 3356
rect -1520 3320 -840 3324
rect -800 3356 4840 3360
rect -800 3324 -796 3356
rect -764 3324 -716 3356
rect -684 3324 -636 3356
rect -604 3324 -556 3356
rect -524 3324 -476 3356
rect -444 3324 -396 3356
rect -364 3324 -316 3356
rect -284 3324 -236 3356
rect -204 3324 -156 3356
rect -124 3324 -76 3356
rect -44 3324 4 3356
rect 36 3324 84 3356
rect 116 3324 164 3356
rect 196 3324 244 3356
rect 276 3324 324 3356
rect 356 3324 404 3356
rect 436 3324 484 3356
rect 516 3324 564 3356
rect 596 3324 644 3356
rect 676 3324 724 3356
rect 756 3324 804 3356
rect 836 3324 884 3356
rect 916 3324 964 3356
rect 996 3324 1044 3356
rect 1076 3324 1124 3356
rect 1156 3324 1204 3356
rect 1236 3324 1284 3356
rect 1316 3324 1364 3356
rect 1396 3324 1444 3356
rect 1476 3324 1524 3356
rect 1556 3324 1604 3356
rect 1636 3324 1684 3356
rect 1716 3324 1764 3356
rect 1796 3324 1844 3356
rect 1876 3324 1924 3356
rect 1956 3324 2004 3356
rect 2036 3324 2084 3356
rect 2116 3324 2164 3356
rect 2196 3324 2244 3356
rect 2276 3324 2324 3356
rect 2356 3324 2404 3356
rect 2436 3324 2484 3356
rect 2516 3324 2564 3356
rect 2596 3324 2644 3356
rect 2676 3324 2724 3356
rect 2756 3324 2804 3356
rect 2836 3324 2884 3356
rect 2916 3324 2964 3356
rect 2996 3324 3044 3356
rect 3076 3324 3124 3356
rect 3156 3324 3204 3356
rect 3236 3324 3284 3356
rect 3316 3324 3364 3356
rect 3396 3324 3444 3356
rect 3476 3324 3524 3356
rect 3556 3324 3604 3356
rect 3636 3324 3684 3356
rect 3716 3324 3764 3356
rect 3796 3324 3844 3356
rect 3876 3324 3924 3356
rect 3956 3324 4004 3356
rect 4036 3324 4084 3356
rect 4116 3324 4164 3356
rect 4196 3324 4244 3356
rect 4276 3324 4324 3356
rect 4356 3324 4404 3356
rect 4436 3324 4484 3356
rect 4516 3324 4564 3356
rect 4596 3324 4644 3356
rect 4676 3324 4724 3356
rect 4756 3324 4804 3356
rect 4836 3324 4840 3356
rect -800 3320 4840 3324
rect 4880 3356 5720 3360
rect 4880 3324 4884 3356
rect 4916 3324 5044 3356
rect 5076 3324 5204 3356
rect 5236 3324 5364 3356
rect 5396 3324 5524 3356
rect 5556 3324 5684 3356
rect 5716 3324 5720 3356
rect 4880 3320 5720 3324
rect -1520 3276 -840 3280
rect -1520 3244 -1516 3276
rect -1484 3244 -1356 3276
rect -1324 3244 -1196 3276
rect -1164 3244 -1036 3276
rect -1004 3244 -876 3276
rect -844 3244 -840 3276
rect -1520 3240 -840 3244
rect -800 3276 4840 3280
rect -800 3244 -796 3276
rect -764 3244 -716 3276
rect -684 3244 -636 3276
rect -604 3244 -556 3276
rect -524 3244 -476 3276
rect -444 3244 -396 3276
rect -364 3244 -316 3276
rect -284 3244 -236 3276
rect -204 3244 -156 3276
rect -124 3244 -76 3276
rect -44 3244 4 3276
rect 36 3244 84 3276
rect 116 3244 164 3276
rect 196 3244 244 3276
rect 276 3244 324 3276
rect 356 3244 404 3276
rect 436 3244 484 3276
rect 516 3244 564 3276
rect 596 3244 644 3276
rect 676 3244 724 3276
rect 756 3244 804 3276
rect 836 3244 884 3276
rect 916 3244 964 3276
rect 996 3244 1044 3276
rect 1076 3244 1124 3276
rect 1156 3244 1204 3276
rect 1236 3244 1284 3276
rect 1316 3244 1364 3276
rect 1396 3244 1444 3276
rect 1476 3244 1524 3276
rect 1556 3244 1604 3276
rect 1636 3244 1684 3276
rect 1716 3244 1764 3276
rect 1796 3244 1844 3276
rect 1876 3244 1924 3276
rect 1956 3244 2004 3276
rect 2036 3244 2084 3276
rect 2116 3244 2164 3276
rect 2196 3244 2244 3276
rect 2276 3244 2324 3276
rect 2356 3244 2404 3276
rect 2436 3244 2484 3276
rect 2516 3244 2564 3276
rect 2596 3244 2644 3276
rect 2676 3244 2724 3276
rect 2756 3244 2804 3276
rect 2836 3244 2884 3276
rect 2916 3244 2964 3276
rect 2996 3244 3044 3276
rect 3076 3244 3124 3276
rect 3156 3244 3204 3276
rect 3236 3244 3284 3276
rect 3316 3244 3364 3276
rect 3396 3244 3444 3276
rect 3476 3244 3524 3276
rect 3556 3244 3604 3276
rect 3636 3244 3684 3276
rect 3716 3244 3764 3276
rect 3796 3244 3844 3276
rect 3876 3244 3924 3276
rect 3956 3244 4004 3276
rect 4036 3244 4084 3276
rect 4116 3244 4164 3276
rect 4196 3244 4244 3276
rect 4276 3244 4324 3276
rect 4356 3244 4404 3276
rect 4436 3244 4484 3276
rect 4516 3244 4564 3276
rect 4596 3244 4644 3276
rect 4676 3244 4724 3276
rect 4756 3244 4804 3276
rect 4836 3244 4840 3276
rect -800 3240 4840 3244
rect 4880 3276 5720 3280
rect 4880 3244 4884 3276
rect 4916 3244 5044 3276
rect 5076 3244 5204 3276
rect 5236 3244 5364 3276
rect 5396 3244 5524 3276
rect 5556 3244 5684 3276
rect 5716 3244 5720 3276
rect 4880 3240 5720 3244
rect -1520 3196 -840 3200
rect -1520 3164 -1516 3196
rect -1484 3164 -1356 3196
rect -1324 3164 -1196 3196
rect -1164 3164 -1036 3196
rect -1004 3164 -876 3196
rect -844 3164 -840 3196
rect -1520 3160 -840 3164
rect -800 3196 4840 3200
rect -800 3164 -796 3196
rect -764 3164 -716 3196
rect -684 3164 -636 3196
rect -604 3164 -556 3196
rect -524 3164 -476 3196
rect -444 3164 -396 3196
rect -364 3164 -316 3196
rect -284 3164 -236 3196
rect -204 3164 -156 3196
rect -124 3164 -76 3196
rect -44 3164 4 3196
rect 36 3164 84 3196
rect 116 3164 164 3196
rect 196 3164 244 3196
rect 276 3164 324 3196
rect 356 3164 404 3196
rect 436 3164 484 3196
rect 516 3164 564 3196
rect 596 3164 644 3196
rect 676 3164 724 3196
rect 756 3164 804 3196
rect 836 3164 884 3196
rect 916 3164 964 3196
rect 996 3164 1044 3196
rect 1076 3164 1124 3196
rect 1156 3164 1204 3196
rect 1236 3164 1284 3196
rect 1316 3164 1364 3196
rect 1396 3164 1444 3196
rect 1476 3164 1524 3196
rect 1556 3164 1604 3196
rect 1636 3164 1684 3196
rect 1716 3164 1764 3196
rect 1796 3164 1844 3196
rect 1876 3164 1924 3196
rect 1956 3164 2004 3196
rect 2036 3164 2084 3196
rect 2116 3164 2164 3196
rect 2196 3164 2244 3196
rect 2276 3164 2324 3196
rect 2356 3164 2404 3196
rect 2436 3164 2484 3196
rect 2516 3164 2564 3196
rect 2596 3164 2644 3196
rect 2676 3164 2724 3196
rect 2756 3164 2804 3196
rect 2836 3164 2884 3196
rect 2916 3164 2964 3196
rect 2996 3164 3044 3196
rect 3076 3164 3124 3196
rect 3156 3164 3204 3196
rect 3236 3164 3284 3196
rect 3316 3164 3364 3196
rect 3396 3164 3444 3196
rect 3476 3164 3524 3196
rect 3556 3164 3604 3196
rect 3636 3164 3684 3196
rect 3716 3164 3764 3196
rect 3796 3164 3844 3196
rect 3876 3164 3924 3196
rect 3956 3164 4004 3196
rect 4036 3164 4084 3196
rect 4116 3164 4164 3196
rect 4196 3164 4244 3196
rect 4276 3164 4324 3196
rect 4356 3164 4404 3196
rect 4436 3164 4484 3196
rect 4516 3164 4564 3196
rect 4596 3164 4644 3196
rect 4676 3164 4724 3196
rect 4756 3164 4804 3196
rect 4836 3164 4840 3196
rect -800 3160 4840 3164
rect 4880 3196 5720 3200
rect 4880 3164 4884 3196
rect 4916 3164 5044 3196
rect 5076 3164 5204 3196
rect 5236 3164 5364 3196
rect 5396 3164 5524 3196
rect 5556 3164 5684 3196
rect 5716 3164 5720 3196
rect 4880 3160 5720 3164
rect -1520 3116 -840 3120
rect -1520 3084 -1516 3116
rect -1484 3084 -1356 3116
rect -1324 3084 -1196 3116
rect -1164 3084 -1036 3116
rect -1004 3084 -876 3116
rect -844 3084 -840 3116
rect -1520 3080 -840 3084
rect -800 3116 4840 3120
rect -800 3084 -796 3116
rect -764 3084 -716 3116
rect -684 3084 -636 3116
rect -604 3084 -556 3116
rect -524 3084 -476 3116
rect -444 3084 -396 3116
rect -364 3084 -316 3116
rect -284 3084 -236 3116
rect -204 3084 -156 3116
rect -124 3084 -76 3116
rect -44 3084 4 3116
rect 36 3084 84 3116
rect 116 3084 164 3116
rect 196 3084 244 3116
rect 276 3084 324 3116
rect 356 3084 404 3116
rect 436 3084 484 3116
rect 516 3084 564 3116
rect 596 3084 644 3116
rect 676 3084 724 3116
rect 756 3084 804 3116
rect 836 3084 884 3116
rect 916 3084 964 3116
rect 996 3084 1044 3116
rect 1076 3084 1124 3116
rect 1156 3084 1204 3116
rect 1236 3084 1284 3116
rect 1316 3084 1364 3116
rect 1396 3084 1444 3116
rect 1476 3084 1524 3116
rect 1556 3084 1604 3116
rect 1636 3084 1684 3116
rect 1716 3084 1764 3116
rect 1796 3084 1844 3116
rect 1876 3084 1924 3116
rect 1956 3084 2004 3116
rect 2036 3084 2084 3116
rect 2116 3084 2164 3116
rect 2196 3084 2244 3116
rect 2276 3084 2324 3116
rect 2356 3084 2404 3116
rect 2436 3084 2484 3116
rect 2516 3084 2564 3116
rect 2596 3084 2644 3116
rect 2676 3084 2724 3116
rect 2756 3084 2804 3116
rect 2836 3084 2884 3116
rect 2916 3084 2964 3116
rect 2996 3084 3044 3116
rect 3076 3084 3124 3116
rect 3156 3084 3204 3116
rect 3236 3084 3284 3116
rect 3316 3084 3364 3116
rect 3396 3084 3444 3116
rect 3476 3084 3524 3116
rect 3556 3084 3604 3116
rect 3636 3084 3684 3116
rect 3716 3084 3764 3116
rect 3796 3084 3844 3116
rect 3876 3084 3924 3116
rect 3956 3084 4004 3116
rect 4036 3084 4084 3116
rect 4116 3084 4164 3116
rect 4196 3084 4244 3116
rect 4276 3084 4324 3116
rect 4356 3084 4404 3116
rect 4436 3084 4484 3116
rect 4516 3084 4564 3116
rect 4596 3084 4644 3116
rect 4676 3084 4724 3116
rect 4756 3084 4804 3116
rect 4836 3084 4840 3116
rect -800 3080 4840 3084
rect 4880 3116 5720 3120
rect 4880 3084 4884 3116
rect 4916 3084 5044 3116
rect 5076 3084 5204 3116
rect 5236 3084 5364 3116
rect 5396 3084 5524 3116
rect 5556 3084 5684 3116
rect 5716 3084 5720 3116
rect 4880 3080 5720 3084
rect -1520 3036 -840 3040
rect -1520 3004 -1516 3036
rect -1484 3004 -1356 3036
rect -1324 3004 -1196 3036
rect -1164 3004 -1036 3036
rect -1004 3004 -876 3036
rect -844 3004 -840 3036
rect -1520 3000 -840 3004
rect -800 3036 4840 3040
rect -800 3004 -796 3036
rect -764 3004 -716 3036
rect -684 3004 -636 3036
rect -604 3004 -556 3036
rect -524 3004 -476 3036
rect -444 3004 -396 3036
rect -364 3004 -316 3036
rect -284 3004 -236 3036
rect -204 3004 -156 3036
rect -124 3004 -76 3036
rect -44 3004 4 3036
rect 36 3004 84 3036
rect 116 3004 164 3036
rect 196 3004 244 3036
rect 276 3004 324 3036
rect 356 3004 404 3036
rect 436 3004 484 3036
rect 516 3004 564 3036
rect 596 3004 644 3036
rect 676 3004 724 3036
rect 756 3004 804 3036
rect 836 3004 884 3036
rect 916 3004 964 3036
rect 996 3004 1044 3036
rect 1076 3004 1124 3036
rect 1156 3004 1204 3036
rect 1236 3004 1284 3036
rect 1316 3004 1364 3036
rect 1396 3004 1444 3036
rect 1476 3004 1524 3036
rect 1556 3004 1604 3036
rect 1636 3004 1684 3036
rect 1716 3004 1764 3036
rect 1796 3004 1844 3036
rect 1876 3004 1924 3036
rect 1956 3004 2004 3036
rect 2036 3004 2084 3036
rect 2116 3004 2164 3036
rect 2196 3004 2244 3036
rect 2276 3004 2324 3036
rect 2356 3004 2404 3036
rect 2436 3004 2484 3036
rect 2516 3004 2564 3036
rect 2596 3004 2644 3036
rect 2676 3004 2724 3036
rect 2756 3004 2804 3036
rect 2836 3004 2884 3036
rect 2916 3004 2964 3036
rect 2996 3004 3044 3036
rect 3076 3004 3124 3036
rect 3156 3004 3204 3036
rect 3236 3004 3284 3036
rect 3316 3004 3364 3036
rect 3396 3004 3444 3036
rect 3476 3004 3524 3036
rect 3556 3004 3604 3036
rect 3636 3004 3684 3036
rect 3716 3004 3764 3036
rect 3796 3004 3844 3036
rect 3876 3004 3924 3036
rect 3956 3004 4004 3036
rect 4036 3004 4084 3036
rect 4116 3004 4164 3036
rect 4196 3004 4244 3036
rect 4276 3004 4324 3036
rect 4356 3004 4404 3036
rect 4436 3004 4484 3036
rect 4516 3004 4564 3036
rect 4596 3004 4644 3036
rect 4676 3004 4724 3036
rect 4756 3004 4804 3036
rect 4836 3004 4840 3036
rect -800 3000 4840 3004
rect 4880 3036 5720 3040
rect 4880 3004 4884 3036
rect 4916 3004 5044 3036
rect 5076 3004 5204 3036
rect 5236 3004 5364 3036
rect 5396 3004 5524 3036
rect 5556 3004 5684 3036
rect 5716 3004 5720 3036
rect 4880 3000 5720 3004
rect -1520 2956 -840 2960
rect -1520 2924 -1516 2956
rect -1484 2924 -1356 2956
rect -1324 2924 -1196 2956
rect -1164 2924 -1036 2956
rect -1004 2924 -876 2956
rect -844 2924 -840 2956
rect -1520 2920 -840 2924
rect -800 2956 4840 2960
rect -800 2924 -796 2956
rect -764 2924 -716 2956
rect -684 2924 -636 2956
rect -604 2924 -556 2956
rect -524 2924 -476 2956
rect -444 2924 -396 2956
rect -364 2924 -316 2956
rect -284 2924 -236 2956
rect -204 2924 -156 2956
rect -124 2924 -76 2956
rect -44 2924 4 2956
rect 36 2924 84 2956
rect 116 2924 164 2956
rect 196 2924 244 2956
rect 276 2924 324 2956
rect 356 2924 404 2956
rect 436 2924 484 2956
rect 516 2924 564 2956
rect 596 2924 644 2956
rect 676 2924 724 2956
rect 756 2924 804 2956
rect 836 2924 884 2956
rect 916 2924 964 2956
rect 996 2924 1044 2956
rect 1076 2924 1124 2956
rect 1156 2924 1204 2956
rect 1236 2924 1284 2956
rect 1316 2924 1364 2956
rect 1396 2924 1444 2956
rect 1476 2924 1524 2956
rect 1556 2924 1604 2956
rect 1636 2924 1684 2956
rect 1716 2924 1764 2956
rect 1796 2924 1844 2956
rect 1876 2924 1924 2956
rect 1956 2924 2004 2956
rect 2036 2924 2084 2956
rect 2116 2924 2164 2956
rect 2196 2924 2244 2956
rect 2276 2924 2324 2956
rect 2356 2924 2404 2956
rect 2436 2924 2484 2956
rect 2516 2924 2564 2956
rect 2596 2924 2644 2956
rect 2676 2924 2724 2956
rect 2756 2924 2804 2956
rect 2836 2924 2884 2956
rect 2916 2924 2964 2956
rect 2996 2924 3044 2956
rect 3076 2924 3124 2956
rect 3156 2924 3204 2956
rect 3236 2924 3284 2956
rect 3316 2924 3364 2956
rect 3396 2924 3444 2956
rect 3476 2924 3524 2956
rect 3556 2924 3604 2956
rect 3636 2924 3684 2956
rect 3716 2924 3764 2956
rect 3796 2924 3844 2956
rect 3876 2924 3924 2956
rect 3956 2924 4004 2956
rect 4036 2924 4084 2956
rect 4116 2924 4164 2956
rect 4196 2924 4244 2956
rect 4276 2924 4324 2956
rect 4356 2924 4404 2956
rect 4436 2924 4484 2956
rect 4516 2924 4564 2956
rect 4596 2924 4644 2956
rect 4676 2924 4724 2956
rect 4756 2924 4804 2956
rect 4836 2924 4840 2956
rect -800 2920 4840 2924
rect 4880 2956 5720 2960
rect 4880 2924 4884 2956
rect 4916 2924 5044 2956
rect 5076 2924 5204 2956
rect 5236 2924 5364 2956
rect 5396 2924 5524 2956
rect 5556 2924 5684 2956
rect 5716 2924 5720 2956
rect 4880 2920 5720 2924
rect -1520 2876 -840 2880
rect -1520 2844 -1516 2876
rect -1484 2844 -1356 2876
rect -1324 2844 -1196 2876
rect -1164 2844 -1036 2876
rect -1004 2844 -876 2876
rect -844 2844 -840 2876
rect -1520 2840 -840 2844
rect -800 2876 4840 2880
rect -800 2844 -796 2876
rect -764 2844 -716 2876
rect -684 2844 -636 2876
rect -604 2844 -556 2876
rect -524 2844 -476 2876
rect -444 2844 -396 2876
rect -364 2844 -316 2876
rect -284 2844 -236 2876
rect -204 2844 -156 2876
rect -124 2844 -76 2876
rect -44 2844 4 2876
rect 36 2844 84 2876
rect 116 2844 164 2876
rect 196 2844 244 2876
rect 276 2844 324 2876
rect 356 2844 404 2876
rect 436 2844 484 2876
rect 516 2844 564 2876
rect 596 2844 644 2876
rect 676 2844 724 2876
rect 756 2844 804 2876
rect 836 2844 884 2876
rect 916 2844 964 2876
rect 996 2844 1044 2876
rect 1076 2844 1124 2876
rect 1156 2844 1204 2876
rect 1236 2844 1284 2876
rect 1316 2844 1364 2876
rect 1396 2844 1444 2876
rect 1476 2844 1524 2876
rect 1556 2844 1604 2876
rect 1636 2844 1684 2876
rect 1716 2844 1764 2876
rect 1796 2844 1844 2876
rect 1876 2844 1924 2876
rect 1956 2844 2004 2876
rect 2036 2844 2084 2876
rect 2116 2844 2164 2876
rect 2196 2844 2244 2876
rect 2276 2844 2324 2876
rect 2356 2844 2404 2876
rect 2436 2844 2484 2876
rect 2516 2844 2564 2876
rect 2596 2844 2644 2876
rect 2676 2844 2724 2876
rect 2756 2844 2804 2876
rect 2836 2844 2884 2876
rect 2916 2844 2964 2876
rect 2996 2844 3044 2876
rect 3076 2844 3124 2876
rect 3156 2844 3204 2876
rect 3236 2844 3284 2876
rect 3316 2844 3364 2876
rect 3396 2844 3444 2876
rect 3476 2844 3524 2876
rect 3556 2844 3604 2876
rect 3636 2844 3684 2876
rect 3716 2844 3764 2876
rect 3796 2844 3844 2876
rect 3876 2844 3924 2876
rect 3956 2844 4004 2876
rect 4036 2844 4084 2876
rect 4116 2844 4164 2876
rect 4196 2844 4244 2876
rect 4276 2844 4324 2876
rect 4356 2844 4404 2876
rect 4436 2844 4484 2876
rect 4516 2844 4564 2876
rect 4596 2844 4644 2876
rect 4676 2844 4724 2876
rect 4756 2844 4804 2876
rect 4836 2844 4840 2876
rect -800 2840 4840 2844
rect 4880 2876 5720 2880
rect 4880 2844 4884 2876
rect 4916 2844 5044 2876
rect 5076 2844 5204 2876
rect 5236 2844 5364 2876
rect 5396 2844 5524 2876
rect 5556 2844 5684 2876
rect 5716 2844 5720 2876
rect 4880 2840 5720 2844
rect -1520 2796 -840 2800
rect -1520 2764 -1516 2796
rect -1484 2764 -1356 2796
rect -1324 2764 -1196 2796
rect -1164 2764 -1036 2796
rect -1004 2764 -876 2796
rect -844 2764 -840 2796
rect -1520 2760 -840 2764
rect -800 2796 4840 2800
rect -800 2764 -796 2796
rect -764 2764 -716 2796
rect -684 2764 -636 2796
rect -604 2764 -556 2796
rect -524 2764 -476 2796
rect -444 2764 -396 2796
rect -364 2764 -316 2796
rect -284 2764 -236 2796
rect -204 2764 -156 2796
rect -124 2764 -76 2796
rect -44 2764 4 2796
rect 36 2764 84 2796
rect 116 2764 164 2796
rect 196 2764 244 2796
rect 276 2764 324 2796
rect 356 2764 404 2796
rect 436 2764 484 2796
rect 516 2764 564 2796
rect 596 2764 644 2796
rect 676 2764 724 2796
rect 756 2764 804 2796
rect 836 2764 884 2796
rect 916 2764 964 2796
rect 996 2764 1044 2796
rect 1076 2764 1124 2796
rect 1156 2764 1204 2796
rect 1236 2764 1284 2796
rect 1316 2764 1364 2796
rect 1396 2764 1444 2796
rect 1476 2764 1524 2796
rect 1556 2764 1604 2796
rect 1636 2764 1684 2796
rect 1716 2764 1764 2796
rect 1796 2764 1844 2796
rect 1876 2764 1924 2796
rect 1956 2764 2004 2796
rect 2036 2764 2084 2796
rect 2116 2764 2164 2796
rect 2196 2764 2244 2796
rect 2276 2764 2324 2796
rect 2356 2764 2404 2796
rect 2436 2764 2484 2796
rect 2516 2764 2564 2796
rect 2596 2764 2644 2796
rect 2676 2764 2724 2796
rect 2756 2764 2804 2796
rect 2836 2764 2884 2796
rect 2916 2764 2964 2796
rect 2996 2764 3044 2796
rect 3076 2764 3124 2796
rect 3156 2764 3204 2796
rect 3236 2764 3284 2796
rect 3316 2764 3364 2796
rect 3396 2764 3444 2796
rect 3476 2764 3524 2796
rect 3556 2764 3604 2796
rect 3636 2764 3684 2796
rect 3716 2764 3764 2796
rect 3796 2764 3844 2796
rect 3876 2764 3924 2796
rect 3956 2764 4004 2796
rect 4036 2764 4084 2796
rect 4116 2764 4164 2796
rect 4196 2764 4244 2796
rect 4276 2764 4324 2796
rect 4356 2764 4404 2796
rect 4436 2764 4484 2796
rect 4516 2764 4564 2796
rect 4596 2764 4644 2796
rect 4676 2764 4724 2796
rect 4756 2764 4804 2796
rect 4836 2764 4840 2796
rect -800 2760 4840 2764
rect 4880 2796 5720 2800
rect 4880 2764 4884 2796
rect 4916 2764 5044 2796
rect 5076 2764 5204 2796
rect 5236 2764 5364 2796
rect 5396 2764 5524 2796
rect 5556 2764 5684 2796
rect 5716 2764 5720 2796
rect 4880 2760 5720 2764
rect -1520 2716 -840 2720
rect -1520 2684 -1516 2716
rect -1484 2684 -1356 2716
rect -1324 2684 -1196 2716
rect -1164 2684 -1036 2716
rect -1004 2684 -876 2716
rect -844 2684 -840 2716
rect -1520 2680 -840 2684
rect -800 2716 4840 2720
rect -800 2684 -796 2716
rect -764 2684 -716 2716
rect -684 2684 -636 2716
rect -604 2684 -556 2716
rect -524 2684 -476 2716
rect -444 2684 -396 2716
rect -364 2684 -316 2716
rect -284 2684 -236 2716
rect -204 2684 -156 2716
rect -124 2684 -76 2716
rect -44 2684 4 2716
rect 36 2684 84 2716
rect 116 2684 164 2716
rect 196 2684 244 2716
rect 276 2684 324 2716
rect 356 2684 404 2716
rect 436 2684 484 2716
rect 516 2684 564 2716
rect 596 2684 644 2716
rect 676 2684 724 2716
rect 756 2684 804 2716
rect 836 2684 884 2716
rect 916 2684 964 2716
rect 996 2684 1044 2716
rect 1076 2684 1124 2716
rect 1156 2684 1204 2716
rect 1236 2684 1284 2716
rect 1316 2684 1364 2716
rect 1396 2684 1444 2716
rect 1476 2684 1524 2716
rect 1556 2684 1604 2716
rect 1636 2684 1684 2716
rect 1716 2684 1764 2716
rect 1796 2684 1844 2716
rect 1876 2684 1924 2716
rect 1956 2684 2004 2716
rect 2036 2684 2084 2716
rect 2116 2684 2164 2716
rect 2196 2684 2244 2716
rect 2276 2684 2324 2716
rect 2356 2684 2404 2716
rect 2436 2684 2484 2716
rect 2516 2684 2564 2716
rect 2596 2684 2644 2716
rect 2676 2684 2724 2716
rect 2756 2684 2804 2716
rect 2836 2684 2884 2716
rect 2916 2684 2964 2716
rect 2996 2684 3044 2716
rect 3076 2684 3124 2716
rect 3156 2684 3204 2716
rect 3236 2684 3284 2716
rect 3316 2684 3364 2716
rect 3396 2684 3444 2716
rect 3476 2684 3524 2716
rect 3556 2684 3604 2716
rect 3636 2684 3684 2716
rect 3716 2684 3764 2716
rect 3796 2684 3844 2716
rect 3876 2684 3924 2716
rect 3956 2684 4004 2716
rect 4036 2684 4084 2716
rect 4116 2684 4164 2716
rect 4196 2684 4244 2716
rect 4276 2684 4324 2716
rect 4356 2684 4404 2716
rect 4436 2684 4484 2716
rect 4516 2684 4564 2716
rect 4596 2684 4644 2716
rect 4676 2684 4724 2716
rect 4756 2684 4804 2716
rect 4836 2684 4840 2716
rect -800 2680 4840 2684
rect 4880 2716 5720 2720
rect 4880 2684 4884 2716
rect 4916 2684 5044 2716
rect 5076 2684 5204 2716
rect 5236 2684 5364 2716
rect 5396 2684 5524 2716
rect 5556 2684 5684 2716
rect 5716 2684 5720 2716
rect 4880 2680 5720 2684
rect -1520 2636 -840 2640
rect -1520 2604 -1516 2636
rect -1484 2604 -1356 2636
rect -1324 2604 -1196 2636
rect -1164 2604 -1036 2636
rect -1004 2604 -876 2636
rect -844 2604 -840 2636
rect -1520 2600 -840 2604
rect -800 2636 4840 2640
rect -800 2604 -796 2636
rect -764 2604 -716 2636
rect -684 2604 -636 2636
rect -604 2604 -556 2636
rect -524 2604 -476 2636
rect -444 2604 -396 2636
rect -364 2604 -316 2636
rect -284 2604 -236 2636
rect -204 2604 -156 2636
rect -124 2604 -76 2636
rect -44 2604 4 2636
rect 36 2604 84 2636
rect 116 2604 164 2636
rect 196 2604 244 2636
rect 276 2604 324 2636
rect 356 2604 404 2636
rect 436 2604 484 2636
rect 516 2604 564 2636
rect 596 2604 644 2636
rect 676 2604 724 2636
rect 756 2604 804 2636
rect 836 2604 884 2636
rect 916 2604 964 2636
rect 996 2604 1044 2636
rect 1076 2604 1124 2636
rect 1156 2604 1204 2636
rect 1236 2604 1284 2636
rect 1316 2604 1364 2636
rect 1396 2604 1444 2636
rect 1476 2604 1524 2636
rect 1556 2604 1604 2636
rect 1636 2604 1684 2636
rect 1716 2604 1764 2636
rect 1796 2604 1844 2636
rect 1876 2604 1924 2636
rect 1956 2604 2004 2636
rect 2036 2604 2084 2636
rect 2116 2604 2164 2636
rect 2196 2604 2244 2636
rect 2276 2604 2324 2636
rect 2356 2604 2404 2636
rect 2436 2604 2484 2636
rect 2516 2604 2564 2636
rect 2596 2604 2644 2636
rect 2676 2604 2724 2636
rect 2756 2604 2804 2636
rect 2836 2604 2884 2636
rect 2916 2604 2964 2636
rect 2996 2604 3044 2636
rect 3076 2604 3124 2636
rect 3156 2604 3204 2636
rect 3236 2604 3284 2636
rect 3316 2604 3364 2636
rect 3396 2604 3444 2636
rect 3476 2604 3524 2636
rect 3556 2604 3604 2636
rect 3636 2604 3684 2636
rect 3716 2604 3764 2636
rect 3796 2604 3844 2636
rect 3876 2604 3924 2636
rect 3956 2604 4004 2636
rect 4036 2604 4084 2636
rect 4116 2604 4164 2636
rect 4196 2604 4244 2636
rect 4276 2604 4324 2636
rect 4356 2604 4404 2636
rect 4436 2604 4484 2636
rect 4516 2604 4564 2636
rect 4596 2604 4644 2636
rect 4676 2604 4724 2636
rect 4756 2604 4804 2636
rect 4836 2604 4840 2636
rect -800 2600 4840 2604
rect 4880 2636 5720 2640
rect 4880 2604 4884 2636
rect 4916 2604 5044 2636
rect 5076 2604 5204 2636
rect 5236 2604 5364 2636
rect 5396 2604 5524 2636
rect 5556 2604 5684 2636
rect 5716 2604 5720 2636
rect 4880 2600 5720 2604
rect -1520 2556 -840 2560
rect -1520 2524 -1516 2556
rect -1484 2524 -1356 2556
rect -1324 2524 -1196 2556
rect -1164 2524 -1036 2556
rect -1004 2524 -876 2556
rect -844 2524 -840 2556
rect -1520 2520 -840 2524
rect -800 2556 4840 2560
rect -800 2524 -796 2556
rect -764 2524 -716 2556
rect -684 2524 -636 2556
rect -604 2524 -556 2556
rect -524 2524 -476 2556
rect -444 2524 -396 2556
rect -364 2524 -316 2556
rect -284 2524 -236 2556
rect -204 2524 -156 2556
rect -124 2524 -76 2556
rect -44 2524 4 2556
rect 36 2524 84 2556
rect 116 2524 164 2556
rect 196 2524 244 2556
rect 276 2524 324 2556
rect 356 2524 404 2556
rect 436 2524 484 2556
rect 516 2524 564 2556
rect 596 2524 644 2556
rect 676 2524 724 2556
rect 756 2524 804 2556
rect 836 2524 884 2556
rect 916 2524 964 2556
rect 996 2524 1044 2556
rect 1076 2524 1124 2556
rect 1156 2524 1204 2556
rect 1236 2524 1284 2556
rect 1316 2524 1364 2556
rect 1396 2524 1444 2556
rect 1476 2524 1524 2556
rect 1556 2524 1604 2556
rect 1636 2524 1684 2556
rect 1716 2524 1764 2556
rect 1796 2524 1844 2556
rect 1876 2524 1924 2556
rect 1956 2524 2004 2556
rect 2036 2524 2084 2556
rect 2116 2524 2164 2556
rect 2196 2524 2244 2556
rect 2276 2524 2324 2556
rect 2356 2524 2404 2556
rect 2436 2524 2484 2556
rect 2516 2524 2564 2556
rect 2596 2524 2644 2556
rect 2676 2524 2724 2556
rect 2756 2524 2804 2556
rect 2836 2524 2884 2556
rect 2916 2524 2964 2556
rect 2996 2524 3044 2556
rect 3076 2524 3124 2556
rect 3156 2524 3204 2556
rect 3236 2524 3284 2556
rect 3316 2524 3364 2556
rect 3396 2524 3444 2556
rect 3476 2524 3524 2556
rect 3556 2524 3604 2556
rect 3636 2524 3684 2556
rect 3716 2524 3764 2556
rect 3796 2524 3844 2556
rect 3876 2524 3924 2556
rect 3956 2524 4004 2556
rect 4036 2524 4084 2556
rect 4116 2524 4164 2556
rect 4196 2524 4244 2556
rect 4276 2524 4324 2556
rect 4356 2524 4404 2556
rect 4436 2524 4484 2556
rect 4516 2524 4564 2556
rect 4596 2524 4644 2556
rect 4676 2524 4724 2556
rect 4756 2524 4804 2556
rect 4836 2524 4840 2556
rect -800 2520 4840 2524
rect 4880 2556 5720 2560
rect 4880 2524 4884 2556
rect 4916 2524 5044 2556
rect 5076 2524 5204 2556
rect 5236 2524 5364 2556
rect 5396 2524 5524 2556
rect 5556 2524 5684 2556
rect 5716 2524 5720 2556
rect 4880 2520 5720 2524
rect -1520 2476 -840 2480
rect -1520 2444 -1516 2476
rect -1484 2444 -1356 2476
rect -1324 2444 -1196 2476
rect -1164 2444 -1036 2476
rect -1004 2444 -876 2476
rect -844 2444 -840 2476
rect -1520 2440 -840 2444
rect -800 2476 4840 2480
rect -800 2444 -796 2476
rect -764 2444 -716 2476
rect -684 2444 -636 2476
rect -604 2444 -556 2476
rect -524 2444 -476 2476
rect -444 2444 -396 2476
rect -364 2444 -316 2476
rect -284 2444 -236 2476
rect -204 2444 -156 2476
rect -124 2444 -76 2476
rect -44 2444 4 2476
rect 36 2444 84 2476
rect 116 2444 164 2476
rect 196 2444 244 2476
rect 276 2444 324 2476
rect 356 2444 404 2476
rect 436 2444 484 2476
rect 516 2444 564 2476
rect 596 2444 644 2476
rect 676 2444 724 2476
rect 756 2444 804 2476
rect 836 2444 884 2476
rect 916 2444 964 2476
rect 996 2444 1044 2476
rect 1076 2444 1124 2476
rect 1156 2444 1204 2476
rect 1236 2444 1284 2476
rect 1316 2444 1364 2476
rect 1396 2444 1444 2476
rect 1476 2444 1524 2476
rect 1556 2444 1604 2476
rect 1636 2444 1684 2476
rect 1716 2444 1764 2476
rect 1796 2444 1844 2476
rect 1876 2444 1924 2476
rect 1956 2444 2004 2476
rect 2036 2444 2084 2476
rect 2116 2444 2164 2476
rect 2196 2444 2244 2476
rect 2276 2444 2324 2476
rect 2356 2444 2404 2476
rect 2436 2444 2484 2476
rect 2516 2444 2564 2476
rect 2596 2444 2644 2476
rect 2676 2444 2724 2476
rect 2756 2444 2804 2476
rect 2836 2444 2884 2476
rect 2916 2444 2964 2476
rect 2996 2444 3044 2476
rect 3076 2444 3124 2476
rect 3156 2444 3204 2476
rect 3236 2444 3284 2476
rect 3316 2444 3364 2476
rect 3396 2444 3444 2476
rect 3476 2444 3524 2476
rect 3556 2444 3604 2476
rect 3636 2444 3684 2476
rect 3716 2444 3764 2476
rect 3796 2444 3844 2476
rect 3876 2444 3924 2476
rect 3956 2444 4004 2476
rect 4036 2444 4084 2476
rect 4116 2444 4164 2476
rect 4196 2444 4244 2476
rect 4276 2444 4324 2476
rect 4356 2444 4404 2476
rect 4436 2444 4484 2476
rect 4516 2444 4564 2476
rect 4596 2444 4644 2476
rect 4676 2444 4724 2476
rect 4756 2444 4804 2476
rect 4836 2444 4840 2476
rect -800 2440 4840 2444
rect 4880 2476 5720 2480
rect 4880 2444 4884 2476
rect 4916 2444 5044 2476
rect 5076 2444 5204 2476
rect 5236 2444 5364 2476
rect 5396 2444 5524 2476
rect 5556 2444 5684 2476
rect 5716 2444 5720 2476
rect 4880 2440 5720 2444
rect -1520 2396 -840 2400
rect -1520 2364 -1516 2396
rect -1484 2364 -1356 2396
rect -1324 2364 -1196 2396
rect -1164 2364 -1036 2396
rect -1004 2364 -876 2396
rect -844 2364 -840 2396
rect -1520 2360 -840 2364
rect -800 2396 4840 2400
rect -800 2364 -796 2396
rect -764 2364 -716 2396
rect -684 2364 -636 2396
rect -604 2364 -556 2396
rect -524 2364 -476 2396
rect -444 2364 -396 2396
rect -364 2364 -316 2396
rect -284 2364 -236 2396
rect -204 2364 -156 2396
rect -124 2364 -76 2396
rect -44 2364 4 2396
rect 36 2364 84 2396
rect 116 2364 164 2396
rect 196 2364 244 2396
rect 276 2364 324 2396
rect 356 2364 404 2396
rect 436 2364 484 2396
rect 516 2364 564 2396
rect 596 2364 644 2396
rect 676 2364 724 2396
rect 756 2364 804 2396
rect 836 2364 884 2396
rect 916 2364 964 2396
rect 996 2364 1044 2396
rect 1076 2364 1124 2396
rect 1156 2364 1204 2396
rect 1236 2364 1284 2396
rect 1316 2364 1364 2396
rect 1396 2364 1444 2396
rect 1476 2364 1524 2396
rect 1556 2364 1604 2396
rect 1636 2364 1684 2396
rect 1716 2364 1764 2396
rect 1796 2364 1844 2396
rect 1876 2364 1924 2396
rect 1956 2364 2004 2396
rect 2036 2364 2084 2396
rect 2116 2364 2164 2396
rect 2196 2364 2244 2396
rect 2276 2364 2324 2396
rect 2356 2364 2404 2396
rect 2436 2364 2484 2396
rect 2516 2364 2564 2396
rect 2596 2364 2644 2396
rect 2676 2364 2724 2396
rect 2756 2364 2804 2396
rect 2836 2364 2884 2396
rect 2916 2364 2964 2396
rect 2996 2364 3044 2396
rect 3076 2364 3124 2396
rect 3156 2364 3204 2396
rect 3236 2364 3284 2396
rect 3316 2364 3364 2396
rect 3396 2364 3444 2396
rect 3476 2364 3524 2396
rect 3556 2364 3604 2396
rect 3636 2364 3684 2396
rect 3716 2364 3764 2396
rect 3796 2364 3844 2396
rect 3876 2364 3924 2396
rect 3956 2364 4004 2396
rect 4036 2364 4084 2396
rect 4116 2364 4164 2396
rect 4196 2364 4244 2396
rect 4276 2364 4324 2396
rect 4356 2364 4404 2396
rect 4436 2364 4484 2396
rect 4516 2364 4564 2396
rect 4596 2364 4644 2396
rect 4676 2364 4724 2396
rect 4756 2364 4804 2396
rect 4836 2364 4840 2396
rect -800 2360 4840 2364
rect 4880 2396 5720 2400
rect 4880 2364 4884 2396
rect 4916 2364 5044 2396
rect 5076 2364 5204 2396
rect 5236 2364 5364 2396
rect 5396 2364 5524 2396
rect 5556 2364 5684 2396
rect 5716 2364 5720 2396
rect 4880 2360 5720 2364
rect -1520 2316 -840 2320
rect -1520 2284 -1516 2316
rect -1484 2284 -1356 2316
rect -1324 2284 -1196 2316
rect -1164 2284 -1036 2316
rect -1004 2284 -876 2316
rect -844 2284 -840 2316
rect -1520 2280 -840 2284
rect -800 2316 4840 2320
rect -800 2284 -796 2316
rect -764 2284 -716 2316
rect -684 2284 -636 2316
rect -604 2284 -556 2316
rect -524 2284 -476 2316
rect -444 2284 -396 2316
rect -364 2284 -316 2316
rect -284 2284 -236 2316
rect -204 2284 -156 2316
rect -124 2284 -76 2316
rect -44 2284 4 2316
rect 36 2284 84 2316
rect 116 2284 164 2316
rect 196 2284 244 2316
rect 276 2284 324 2316
rect 356 2284 404 2316
rect 436 2284 484 2316
rect 516 2284 564 2316
rect 596 2284 644 2316
rect 676 2284 724 2316
rect 756 2284 804 2316
rect 836 2284 884 2316
rect 916 2284 964 2316
rect 996 2284 1044 2316
rect 1076 2284 1124 2316
rect 1156 2284 1204 2316
rect 1236 2284 1284 2316
rect 1316 2284 1364 2316
rect 1396 2284 1444 2316
rect 1476 2284 1524 2316
rect 1556 2284 1604 2316
rect 1636 2284 1684 2316
rect 1716 2284 1764 2316
rect 1796 2284 1844 2316
rect 1876 2284 1924 2316
rect 1956 2284 2004 2316
rect 2036 2284 2084 2316
rect 2116 2284 2164 2316
rect 2196 2284 2244 2316
rect 2276 2284 2324 2316
rect 2356 2284 2404 2316
rect 2436 2284 2484 2316
rect 2516 2284 2564 2316
rect 2596 2284 2644 2316
rect 2676 2284 2724 2316
rect 2756 2284 2804 2316
rect 2836 2284 2884 2316
rect 2916 2284 2964 2316
rect 2996 2284 3044 2316
rect 3076 2284 3124 2316
rect 3156 2284 3204 2316
rect 3236 2284 3284 2316
rect 3316 2284 3364 2316
rect 3396 2284 3444 2316
rect 3476 2284 3524 2316
rect 3556 2284 3604 2316
rect 3636 2284 3684 2316
rect 3716 2284 3764 2316
rect 3796 2284 3844 2316
rect 3876 2284 3924 2316
rect 3956 2284 4004 2316
rect 4036 2284 4084 2316
rect 4116 2284 4164 2316
rect 4196 2284 4244 2316
rect 4276 2284 4324 2316
rect 4356 2284 4404 2316
rect 4436 2284 4484 2316
rect 4516 2284 4564 2316
rect 4596 2284 4644 2316
rect 4676 2284 4724 2316
rect 4756 2284 4804 2316
rect 4836 2284 4840 2316
rect -800 2280 4840 2284
rect 4880 2316 5720 2320
rect 4880 2284 4884 2316
rect 4916 2284 5044 2316
rect 5076 2284 5204 2316
rect 5236 2284 5364 2316
rect 5396 2284 5524 2316
rect 5556 2284 5684 2316
rect 5716 2284 5720 2316
rect 4880 2280 5720 2284
rect -1520 2236 -840 2240
rect -1520 2204 -1516 2236
rect -1484 2204 -1356 2236
rect -1324 2204 -1196 2236
rect -1164 2204 -1036 2236
rect -1004 2204 -876 2236
rect -844 2204 -840 2236
rect -1520 2200 -840 2204
rect -800 2236 4840 2240
rect -800 2204 -796 2236
rect -764 2204 -716 2236
rect -684 2204 -636 2236
rect -604 2204 -556 2236
rect -524 2204 -476 2236
rect -444 2204 -396 2236
rect -364 2204 -316 2236
rect -284 2204 -236 2236
rect -204 2204 -156 2236
rect -124 2204 -76 2236
rect -44 2204 4 2236
rect 36 2204 84 2236
rect 116 2204 164 2236
rect 196 2204 244 2236
rect 276 2204 324 2236
rect 356 2204 404 2236
rect 436 2204 484 2236
rect 516 2204 564 2236
rect 596 2204 644 2236
rect 676 2204 724 2236
rect 756 2204 804 2236
rect 836 2204 884 2236
rect 916 2204 964 2236
rect 996 2204 1044 2236
rect 1076 2204 1124 2236
rect 1156 2204 1204 2236
rect 1236 2204 1284 2236
rect 1316 2204 1364 2236
rect 1396 2204 1444 2236
rect 1476 2204 1524 2236
rect 1556 2204 1604 2236
rect 1636 2204 1684 2236
rect 1716 2204 1764 2236
rect 1796 2204 1844 2236
rect 1876 2204 1924 2236
rect 1956 2204 2004 2236
rect 2036 2204 2084 2236
rect 2116 2204 2164 2236
rect 2196 2204 2244 2236
rect 2276 2204 2324 2236
rect 2356 2204 2404 2236
rect 2436 2204 2484 2236
rect 2516 2204 2564 2236
rect 2596 2204 2644 2236
rect 2676 2204 2724 2236
rect 2756 2204 2804 2236
rect 2836 2204 2884 2236
rect 2916 2204 2964 2236
rect 2996 2204 3044 2236
rect 3076 2204 3124 2236
rect 3156 2204 3204 2236
rect 3236 2204 3284 2236
rect 3316 2204 3364 2236
rect 3396 2204 3444 2236
rect 3476 2204 3524 2236
rect 3556 2204 3604 2236
rect 3636 2204 3684 2236
rect 3716 2204 3764 2236
rect 3796 2204 3844 2236
rect 3876 2204 3924 2236
rect 3956 2204 4004 2236
rect 4036 2204 4084 2236
rect 4116 2204 4164 2236
rect 4196 2204 4244 2236
rect 4276 2204 4324 2236
rect 4356 2204 4404 2236
rect 4436 2204 4484 2236
rect 4516 2204 4564 2236
rect 4596 2204 4644 2236
rect 4676 2204 4724 2236
rect 4756 2204 4804 2236
rect 4836 2204 4840 2236
rect -800 2200 4840 2204
rect 4880 2236 5720 2240
rect 4880 2204 4884 2236
rect 4916 2204 5044 2236
rect 5076 2204 5204 2236
rect 5236 2204 5364 2236
rect 5396 2204 5524 2236
rect 5556 2204 5684 2236
rect 5716 2204 5720 2236
rect 4880 2200 5720 2204
rect -1520 2156 -840 2160
rect -1520 2124 -1516 2156
rect -1484 2124 -1356 2156
rect -1324 2124 -1196 2156
rect -1164 2124 -1036 2156
rect -1004 2124 -876 2156
rect -844 2124 -840 2156
rect -1520 2120 -840 2124
rect -800 2156 4840 2160
rect -800 2124 -796 2156
rect -764 2124 -716 2156
rect -684 2124 -636 2156
rect -604 2124 -556 2156
rect -524 2124 -476 2156
rect -444 2124 -396 2156
rect -364 2124 -316 2156
rect -284 2124 -236 2156
rect -204 2124 -156 2156
rect -124 2124 -76 2156
rect -44 2124 4 2156
rect 36 2124 84 2156
rect 116 2124 164 2156
rect 196 2124 244 2156
rect 276 2124 324 2156
rect 356 2124 404 2156
rect 436 2124 484 2156
rect 516 2124 564 2156
rect 596 2124 644 2156
rect 676 2124 724 2156
rect 756 2124 804 2156
rect 836 2124 884 2156
rect 916 2124 964 2156
rect 996 2124 1044 2156
rect 1076 2124 1124 2156
rect 1156 2124 1204 2156
rect 1236 2124 1284 2156
rect 1316 2124 1364 2156
rect 1396 2124 1444 2156
rect 1476 2124 1524 2156
rect 1556 2124 1604 2156
rect 1636 2124 1684 2156
rect 1716 2124 1764 2156
rect 1796 2124 1844 2156
rect 1876 2124 1924 2156
rect 1956 2124 2004 2156
rect 2036 2124 2084 2156
rect 2116 2124 2164 2156
rect 2196 2124 2244 2156
rect 2276 2124 2324 2156
rect 2356 2124 2404 2156
rect 2436 2124 2484 2156
rect 2516 2124 2564 2156
rect 2596 2124 2644 2156
rect 2676 2124 2724 2156
rect 2756 2124 2804 2156
rect 2836 2124 2884 2156
rect 2916 2124 2964 2156
rect 2996 2124 3044 2156
rect 3076 2124 3124 2156
rect 3156 2124 3204 2156
rect 3236 2124 3284 2156
rect 3316 2124 3364 2156
rect 3396 2124 3444 2156
rect 3476 2124 3524 2156
rect 3556 2124 3604 2156
rect 3636 2124 3684 2156
rect 3716 2124 3764 2156
rect 3796 2124 3844 2156
rect 3876 2124 3924 2156
rect 3956 2124 4004 2156
rect 4036 2124 4084 2156
rect 4116 2124 4164 2156
rect 4196 2124 4244 2156
rect 4276 2124 4324 2156
rect 4356 2124 4404 2156
rect 4436 2124 4484 2156
rect 4516 2124 4564 2156
rect 4596 2124 4644 2156
rect 4676 2124 4724 2156
rect 4756 2124 4804 2156
rect 4836 2124 4840 2156
rect -800 2120 4840 2124
rect 4880 2156 5720 2160
rect 4880 2124 4884 2156
rect 4916 2124 5044 2156
rect 5076 2124 5204 2156
rect 5236 2124 5364 2156
rect 5396 2124 5524 2156
rect 5556 2124 5684 2156
rect 5716 2124 5720 2156
rect 4880 2120 5720 2124
rect -1520 2076 -840 2080
rect -1520 2044 -1516 2076
rect -1484 2044 -1356 2076
rect -1324 2044 -1196 2076
rect -1164 2044 -1036 2076
rect -1004 2044 -876 2076
rect -844 2044 -840 2076
rect -1520 2040 -840 2044
rect -800 2076 4840 2080
rect -800 2044 -796 2076
rect -764 2044 -716 2076
rect -684 2044 -636 2076
rect -604 2044 -556 2076
rect -524 2044 -476 2076
rect -444 2044 -396 2076
rect -364 2044 -316 2076
rect -284 2044 -236 2076
rect -204 2044 -156 2076
rect -124 2044 -76 2076
rect -44 2044 4 2076
rect 36 2044 84 2076
rect 116 2044 164 2076
rect 196 2044 244 2076
rect 276 2044 324 2076
rect 356 2044 404 2076
rect 436 2044 484 2076
rect 516 2044 564 2076
rect 596 2044 644 2076
rect 676 2044 724 2076
rect 756 2044 804 2076
rect 836 2044 884 2076
rect 916 2044 964 2076
rect 996 2044 1044 2076
rect 1076 2044 1124 2076
rect 1156 2044 1204 2076
rect 1236 2044 1284 2076
rect 1316 2044 1364 2076
rect 1396 2044 1444 2076
rect 1476 2044 1524 2076
rect 1556 2044 1604 2076
rect 1636 2044 1684 2076
rect 1716 2044 1764 2076
rect 1796 2044 1844 2076
rect 1876 2044 1924 2076
rect 1956 2044 2004 2076
rect 2036 2044 2084 2076
rect 2116 2044 2164 2076
rect 2196 2044 2244 2076
rect 2276 2044 2324 2076
rect 2356 2044 2404 2076
rect 2436 2044 2484 2076
rect 2516 2044 2564 2076
rect 2596 2044 2644 2076
rect 2676 2044 2724 2076
rect 2756 2044 2804 2076
rect 2836 2044 2884 2076
rect 2916 2044 2964 2076
rect 2996 2044 3044 2076
rect 3076 2044 3124 2076
rect 3156 2044 3204 2076
rect 3236 2044 3284 2076
rect 3316 2044 3364 2076
rect 3396 2044 3444 2076
rect 3476 2044 3524 2076
rect 3556 2044 3604 2076
rect 3636 2044 3684 2076
rect 3716 2044 3764 2076
rect 3796 2044 3844 2076
rect 3876 2044 3924 2076
rect 3956 2044 4004 2076
rect 4036 2044 4084 2076
rect 4116 2044 4164 2076
rect 4196 2044 4244 2076
rect 4276 2044 4324 2076
rect 4356 2044 4404 2076
rect 4436 2044 4484 2076
rect 4516 2044 4564 2076
rect 4596 2044 4644 2076
rect 4676 2044 4724 2076
rect 4756 2044 4804 2076
rect 4836 2044 4840 2076
rect -800 2040 4840 2044
rect 4880 2076 5720 2080
rect 4880 2044 4884 2076
rect 4916 2044 5044 2076
rect 5076 2044 5204 2076
rect 5236 2044 5364 2076
rect 5396 2044 5524 2076
rect 5556 2044 5684 2076
rect 5716 2044 5720 2076
rect 4880 2040 5720 2044
rect -1520 1996 -840 2000
rect -1520 1964 -1516 1996
rect -1484 1964 -1356 1996
rect -1324 1964 -1196 1996
rect -1164 1964 -1036 1996
rect -1004 1964 -876 1996
rect -844 1964 -840 1996
rect -1520 1960 -840 1964
rect -800 1996 4840 2000
rect -800 1964 -796 1996
rect -764 1964 -716 1996
rect -684 1964 -636 1996
rect -604 1964 -556 1996
rect -524 1964 -476 1996
rect -444 1964 -396 1996
rect -364 1964 -316 1996
rect -284 1964 -236 1996
rect -204 1964 -156 1996
rect -124 1964 -76 1996
rect -44 1964 4 1996
rect 36 1964 84 1996
rect 116 1964 164 1996
rect 196 1964 244 1996
rect 276 1964 324 1996
rect 356 1964 404 1996
rect 436 1964 484 1996
rect 516 1964 564 1996
rect 596 1964 644 1996
rect 676 1964 724 1996
rect 756 1964 804 1996
rect 836 1964 884 1996
rect 916 1964 964 1996
rect 996 1964 1044 1996
rect 1076 1964 1124 1996
rect 1156 1964 1204 1996
rect 1236 1964 1284 1996
rect 1316 1964 1364 1996
rect 1396 1964 1444 1996
rect 1476 1964 1524 1996
rect 1556 1964 1604 1996
rect 1636 1964 1684 1996
rect 1716 1964 1764 1996
rect 1796 1964 1844 1996
rect 1876 1964 1924 1996
rect 1956 1964 2004 1996
rect 2036 1964 2084 1996
rect 2116 1964 2164 1996
rect 2196 1964 2244 1996
rect 2276 1964 2324 1996
rect 2356 1964 2404 1996
rect 2436 1964 2484 1996
rect 2516 1964 2564 1996
rect 2596 1964 2644 1996
rect 2676 1964 2724 1996
rect 2756 1964 2804 1996
rect 2836 1964 2884 1996
rect 2916 1964 2964 1996
rect 2996 1964 3044 1996
rect 3076 1964 3124 1996
rect 3156 1964 3204 1996
rect 3236 1964 3284 1996
rect 3316 1964 3364 1996
rect 3396 1964 3444 1996
rect 3476 1964 3524 1996
rect 3556 1964 3604 1996
rect 3636 1964 3684 1996
rect 3716 1964 3764 1996
rect 3796 1964 3844 1996
rect 3876 1964 3924 1996
rect 3956 1964 4004 1996
rect 4036 1964 4084 1996
rect 4116 1964 4164 1996
rect 4196 1964 4244 1996
rect 4276 1964 4324 1996
rect 4356 1964 4404 1996
rect 4436 1964 4484 1996
rect 4516 1964 4564 1996
rect 4596 1964 4644 1996
rect 4676 1964 4724 1996
rect 4756 1964 4804 1996
rect 4836 1964 4840 1996
rect -800 1960 4840 1964
rect 4880 1996 5720 2000
rect 4880 1964 4884 1996
rect 4916 1964 5044 1996
rect 5076 1964 5204 1996
rect 5236 1964 5364 1996
rect 5396 1964 5524 1996
rect 5556 1964 5684 1996
rect 5716 1964 5720 1996
rect 4880 1960 5720 1964
rect -1520 1916 -840 1920
rect -1520 1884 -1516 1916
rect -1484 1884 -1356 1916
rect -1324 1884 -1196 1916
rect -1164 1884 -1036 1916
rect -1004 1884 -876 1916
rect -844 1884 -840 1916
rect -1520 1880 -840 1884
rect -800 1916 4840 1920
rect -800 1884 -796 1916
rect -764 1884 -716 1916
rect -684 1884 -636 1916
rect -604 1884 -556 1916
rect -524 1884 -476 1916
rect -444 1884 -396 1916
rect -364 1884 -316 1916
rect -284 1884 -236 1916
rect -204 1884 -156 1916
rect -124 1884 -76 1916
rect -44 1884 4 1916
rect 36 1884 84 1916
rect 116 1884 164 1916
rect 196 1884 244 1916
rect 276 1884 324 1916
rect 356 1884 404 1916
rect 436 1884 484 1916
rect 516 1884 564 1916
rect 596 1884 644 1916
rect 676 1884 724 1916
rect 756 1884 804 1916
rect 836 1884 884 1916
rect 916 1884 964 1916
rect 996 1884 1044 1916
rect 1076 1884 1124 1916
rect 1156 1884 1204 1916
rect 1236 1884 1284 1916
rect 1316 1884 1364 1916
rect 1396 1884 1444 1916
rect 1476 1884 1524 1916
rect 1556 1884 1604 1916
rect 1636 1884 1684 1916
rect 1716 1884 1764 1916
rect 1796 1884 1844 1916
rect 1876 1884 1924 1916
rect 1956 1884 2004 1916
rect 2036 1884 2084 1916
rect 2116 1884 2164 1916
rect 2196 1884 2244 1916
rect 2276 1884 2324 1916
rect 2356 1884 2404 1916
rect 2436 1884 2484 1916
rect 2516 1884 2564 1916
rect 2596 1884 2644 1916
rect 2676 1884 2724 1916
rect 2756 1884 2804 1916
rect 2836 1884 2884 1916
rect 2916 1884 2964 1916
rect 2996 1884 3044 1916
rect 3076 1884 3124 1916
rect 3156 1884 3204 1916
rect 3236 1884 3284 1916
rect 3316 1884 3364 1916
rect 3396 1884 3444 1916
rect 3476 1884 3524 1916
rect 3556 1884 3604 1916
rect 3636 1884 3684 1916
rect 3716 1884 3764 1916
rect 3796 1884 3844 1916
rect 3876 1884 3924 1916
rect 3956 1884 4004 1916
rect 4036 1884 4084 1916
rect 4116 1884 4164 1916
rect 4196 1884 4244 1916
rect 4276 1884 4324 1916
rect 4356 1884 4404 1916
rect 4436 1884 4484 1916
rect 4516 1884 4564 1916
rect 4596 1884 4644 1916
rect 4676 1884 4724 1916
rect 4756 1884 4804 1916
rect 4836 1884 4840 1916
rect -800 1880 4840 1884
rect 4880 1916 5720 1920
rect 4880 1884 4884 1916
rect 4916 1884 5044 1916
rect 5076 1884 5204 1916
rect 5236 1884 5364 1916
rect 5396 1884 5524 1916
rect 5556 1884 5684 1916
rect 5716 1884 5720 1916
rect 4880 1880 5720 1884
rect -1520 1836 -840 1840
rect -1520 1804 -1516 1836
rect -1484 1804 -1356 1836
rect -1324 1804 -1196 1836
rect -1164 1804 -1036 1836
rect -1004 1804 -876 1836
rect -844 1804 -840 1836
rect -1520 1800 -840 1804
rect -800 1836 4840 1840
rect -800 1804 -796 1836
rect -764 1804 -716 1836
rect -684 1804 -636 1836
rect -604 1804 -556 1836
rect -524 1804 -476 1836
rect -444 1804 -396 1836
rect -364 1804 -316 1836
rect -284 1804 -236 1836
rect -204 1804 -156 1836
rect -124 1804 -76 1836
rect -44 1804 4 1836
rect 36 1804 84 1836
rect 116 1804 164 1836
rect 196 1804 244 1836
rect 276 1804 324 1836
rect 356 1804 404 1836
rect 436 1804 484 1836
rect 516 1804 564 1836
rect 596 1804 644 1836
rect 676 1804 724 1836
rect 756 1804 804 1836
rect 836 1804 884 1836
rect 916 1804 964 1836
rect 996 1804 1044 1836
rect 1076 1804 1124 1836
rect 1156 1804 1204 1836
rect 1236 1804 1284 1836
rect 1316 1804 1364 1836
rect 1396 1804 1444 1836
rect 1476 1804 1524 1836
rect 1556 1804 1604 1836
rect 1636 1804 1684 1836
rect 1716 1804 1764 1836
rect 1796 1804 1844 1836
rect 1876 1804 1924 1836
rect 1956 1804 2004 1836
rect 2036 1804 2084 1836
rect 2116 1804 2164 1836
rect 2196 1804 2244 1836
rect 2276 1804 2324 1836
rect 2356 1804 2404 1836
rect 2436 1804 2484 1836
rect 2516 1804 2564 1836
rect 2596 1804 2644 1836
rect 2676 1804 2724 1836
rect 2756 1804 2804 1836
rect 2836 1804 2884 1836
rect 2916 1804 2964 1836
rect 2996 1804 3044 1836
rect 3076 1804 3124 1836
rect 3156 1804 3204 1836
rect 3236 1804 3284 1836
rect 3316 1804 3364 1836
rect 3396 1804 3444 1836
rect 3476 1804 3524 1836
rect 3556 1804 3604 1836
rect 3636 1804 3684 1836
rect 3716 1804 3764 1836
rect 3796 1804 3844 1836
rect 3876 1804 3924 1836
rect 3956 1804 4004 1836
rect 4036 1804 4084 1836
rect 4116 1804 4164 1836
rect 4196 1804 4244 1836
rect 4276 1804 4324 1836
rect 4356 1804 4404 1836
rect 4436 1804 4484 1836
rect 4516 1804 4564 1836
rect 4596 1804 4644 1836
rect 4676 1804 4724 1836
rect 4756 1804 4804 1836
rect 4836 1804 4840 1836
rect -800 1800 4840 1804
rect 4880 1836 5720 1840
rect 4880 1804 4884 1836
rect 4916 1804 5044 1836
rect 5076 1804 5204 1836
rect 5236 1804 5364 1836
rect 5396 1804 5524 1836
rect 5556 1804 5684 1836
rect 5716 1804 5720 1836
rect 4880 1800 5720 1804
rect -1520 1756 -840 1760
rect -1520 1724 -1516 1756
rect -1484 1724 -1356 1756
rect -1324 1724 -1196 1756
rect -1164 1724 -1036 1756
rect -1004 1724 -876 1756
rect -844 1724 -840 1756
rect -1520 1720 -840 1724
rect -800 1756 4840 1760
rect -800 1724 -796 1756
rect -764 1724 -716 1756
rect -684 1724 -636 1756
rect -604 1724 -556 1756
rect -524 1724 -476 1756
rect -444 1724 -396 1756
rect -364 1724 -316 1756
rect -284 1724 -236 1756
rect -204 1724 -156 1756
rect -124 1724 -76 1756
rect -44 1724 4 1756
rect 36 1724 84 1756
rect 116 1724 164 1756
rect 196 1724 244 1756
rect 276 1724 324 1756
rect 356 1724 404 1756
rect 436 1724 484 1756
rect 516 1724 564 1756
rect 596 1724 644 1756
rect 676 1724 724 1756
rect 756 1724 804 1756
rect 836 1724 884 1756
rect 916 1724 964 1756
rect 996 1724 1044 1756
rect 1076 1724 1124 1756
rect 1156 1724 1204 1756
rect 1236 1724 1284 1756
rect 1316 1724 1364 1756
rect 1396 1724 1444 1756
rect 1476 1724 1524 1756
rect 1556 1724 1604 1756
rect 1636 1724 1684 1756
rect 1716 1724 1764 1756
rect 1796 1724 1844 1756
rect 1876 1724 1924 1756
rect 1956 1724 2004 1756
rect 2036 1724 2084 1756
rect 2116 1724 2164 1756
rect 2196 1724 2244 1756
rect 2276 1724 2324 1756
rect 2356 1724 2404 1756
rect 2436 1724 2484 1756
rect 2516 1724 2564 1756
rect 2596 1724 2644 1756
rect 2676 1724 2724 1756
rect 2756 1724 2804 1756
rect 2836 1724 2884 1756
rect 2916 1724 2964 1756
rect 2996 1724 3044 1756
rect 3076 1724 3124 1756
rect 3156 1724 3204 1756
rect 3236 1724 3284 1756
rect 3316 1724 3364 1756
rect 3396 1724 3444 1756
rect 3476 1724 3524 1756
rect 3556 1724 3604 1756
rect 3636 1724 3684 1756
rect 3716 1724 3764 1756
rect 3796 1724 3844 1756
rect 3876 1724 3924 1756
rect 3956 1724 4004 1756
rect 4036 1724 4084 1756
rect 4116 1724 4164 1756
rect 4196 1724 4244 1756
rect 4276 1724 4324 1756
rect 4356 1724 4404 1756
rect 4436 1724 4484 1756
rect 4516 1724 4564 1756
rect 4596 1724 4644 1756
rect 4676 1724 4724 1756
rect 4756 1724 4804 1756
rect 4836 1724 4840 1756
rect -800 1720 4840 1724
rect 4880 1756 5720 1760
rect 4880 1724 4884 1756
rect 4916 1724 5044 1756
rect 5076 1724 5204 1756
rect 5236 1724 5364 1756
rect 5396 1724 5524 1756
rect 5556 1724 5684 1756
rect 5716 1724 5720 1756
rect 4880 1720 5720 1724
rect -1520 1676 -840 1680
rect -1520 1644 -1516 1676
rect -1484 1644 -1356 1676
rect -1324 1644 -1196 1676
rect -1164 1644 -1036 1676
rect -1004 1644 -876 1676
rect -844 1644 -840 1676
rect -1520 1640 -840 1644
rect -800 1676 4840 1680
rect -800 1644 -796 1676
rect -764 1644 -716 1676
rect -684 1644 -636 1676
rect -604 1644 -556 1676
rect -524 1644 -476 1676
rect -444 1644 -396 1676
rect -364 1644 -316 1676
rect -284 1644 -236 1676
rect -204 1644 -156 1676
rect -124 1644 -76 1676
rect -44 1644 4 1676
rect 36 1644 84 1676
rect 116 1644 164 1676
rect 196 1644 244 1676
rect 276 1644 324 1676
rect 356 1644 404 1676
rect 436 1644 484 1676
rect 516 1644 564 1676
rect 596 1644 644 1676
rect 676 1644 724 1676
rect 756 1644 804 1676
rect 836 1644 884 1676
rect 916 1644 964 1676
rect 996 1644 1044 1676
rect 1076 1644 1124 1676
rect 1156 1644 1204 1676
rect 1236 1644 1284 1676
rect 1316 1644 1364 1676
rect 1396 1644 1444 1676
rect 1476 1644 1524 1676
rect 1556 1644 1604 1676
rect 1636 1644 1684 1676
rect 1716 1644 1764 1676
rect 1796 1644 1844 1676
rect 1876 1644 1924 1676
rect 1956 1644 2004 1676
rect 2036 1644 2084 1676
rect 2116 1644 2164 1676
rect 2196 1644 2244 1676
rect 2276 1644 2324 1676
rect 2356 1644 2404 1676
rect 2436 1644 2484 1676
rect 2516 1644 2564 1676
rect 2596 1644 2644 1676
rect 2676 1644 2724 1676
rect 2756 1644 2804 1676
rect 2836 1644 2884 1676
rect 2916 1644 2964 1676
rect 2996 1644 3044 1676
rect 3076 1644 3124 1676
rect 3156 1644 3204 1676
rect 3236 1644 3284 1676
rect 3316 1644 3364 1676
rect 3396 1644 3444 1676
rect 3476 1644 3524 1676
rect 3556 1644 3604 1676
rect 3636 1644 3684 1676
rect 3716 1644 3764 1676
rect 3796 1644 3844 1676
rect 3876 1644 3924 1676
rect 3956 1644 4004 1676
rect 4036 1644 4084 1676
rect 4116 1644 4164 1676
rect 4196 1644 4244 1676
rect 4276 1644 4324 1676
rect 4356 1644 4404 1676
rect 4436 1644 4484 1676
rect 4516 1644 4564 1676
rect 4596 1644 4644 1676
rect 4676 1644 4724 1676
rect 4756 1644 4804 1676
rect 4836 1644 4840 1676
rect -800 1640 4840 1644
rect 4880 1676 5720 1680
rect 4880 1644 4884 1676
rect 4916 1644 5044 1676
rect 5076 1644 5204 1676
rect 5236 1644 5364 1676
rect 5396 1644 5524 1676
rect 5556 1644 5684 1676
rect 5716 1644 5720 1676
rect 4880 1640 5720 1644
rect -1520 1596 -840 1600
rect -1520 1564 -1516 1596
rect -1484 1564 -1356 1596
rect -1324 1564 -1196 1596
rect -1164 1564 -1036 1596
rect -1004 1564 -876 1596
rect -844 1564 -840 1596
rect -1520 1560 -840 1564
rect -800 1596 4840 1600
rect -800 1564 -796 1596
rect -764 1564 -716 1596
rect -684 1564 -636 1596
rect -604 1564 -556 1596
rect -524 1564 -476 1596
rect -444 1564 -396 1596
rect -364 1564 -316 1596
rect -284 1564 -236 1596
rect -204 1564 -156 1596
rect -124 1564 -76 1596
rect -44 1564 4 1596
rect 36 1564 84 1596
rect 116 1564 164 1596
rect 196 1564 244 1596
rect 276 1564 324 1596
rect 356 1564 404 1596
rect 436 1564 484 1596
rect 516 1564 564 1596
rect 596 1564 644 1596
rect 676 1564 724 1596
rect 756 1564 804 1596
rect 836 1564 884 1596
rect 916 1564 964 1596
rect 996 1564 1044 1596
rect 1076 1564 1124 1596
rect 1156 1564 1204 1596
rect 1236 1564 1284 1596
rect 1316 1564 1364 1596
rect 1396 1564 1444 1596
rect 1476 1564 1524 1596
rect 1556 1564 1604 1596
rect 1636 1564 1684 1596
rect 1716 1564 1764 1596
rect 1796 1564 1844 1596
rect 1876 1564 1924 1596
rect 1956 1564 2004 1596
rect 2036 1564 2084 1596
rect 2116 1564 2164 1596
rect 2196 1564 2244 1596
rect 2276 1564 2324 1596
rect 2356 1564 2404 1596
rect 2436 1564 2484 1596
rect 2516 1564 2564 1596
rect 2596 1564 2644 1596
rect 2676 1564 2724 1596
rect 2756 1564 2804 1596
rect 2836 1564 2884 1596
rect 2916 1564 2964 1596
rect 2996 1564 3044 1596
rect 3076 1564 3124 1596
rect 3156 1564 3204 1596
rect 3236 1564 3284 1596
rect 3316 1564 3364 1596
rect 3396 1564 3444 1596
rect 3476 1564 3524 1596
rect 3556 1564 3604 1596
rect 3636 1564 3684 1596
rect 3716 1564 3764 1596
rect 3796 1564 3844 1596
rect 3876 1564 3924 1596
rect 3956 1564 4004 1596
rect 4036 1564 4084 1596
rect 4116 1564 4164 1596
rect 4196 1564 4244 1596
rect 4276 1564 4324 1596
rect 4356 1564 4404 1596
rect 4436 1564 4484 1596
rect 4516 1564 4564 1596
rect 4596 1564 4644 1596
rect 4676 1564 4724 1596
rect 4756 1564 4804 1596
rect 4836 1564 4840 1596
rect -800 1560 4840 1564
rect 4880 1596 5720 1600
rect 4880 1564 4884 1596
rect 4916 1564 5044 1596
rect 5076 1564 5204 1596
rect 5236 1564 5364 1596
rect 5396 1564 5524 1596
rect 5556 1564 5684 1596
rect 5716 1564 5720 1596
rect 4880 1560 5720 1564
rect -1520 1516 -840 1520
rect -1520 1484 -1516 1516
rect -1484 1484 -1356 1516
rect -1324 1484 -1196 1516
rect -1164 1484 -1036 1516
rect -1004 1484 -876 1516
rect -844 1484 -840 1516
rect -1520 1480 -840 1484
rect -800 1516 4840 1520
rect -800 1484 -796 1516
rect -764 1484 -716 1516
rect -684 1484 -636 1516
rect -604 1484 -556 1516
rect -524 1484 -476 1516
rect -444 1484 -396 1516
rect -364 1484 -316 1516
rect -284 1484 -236 1516
rect -204 1484 -156 1516
rect -124 1484 -76 1516
rect -44 1484 4 1516
rect 36 1484 84 1516
rect 116 1484 164 1516
rect 196 1484 244 1516
rect 276 1484 324 1516
rect 356 1484 404 1516
rect 436 1484 484 1516
rect 516 1484 564 1516
rect 596 1484 644 1516
rect 676 1484 724 1516
rect 756 1484 804 1516
rect 836 1484 884 1516
rect 916 1484 964 1516
rect 996 1484 1044 1516
rect 1076 1484 1124 1516
rect 1156 1484 1204 1516
rect 1236 1484 1284 1516
rect 1316 1484 1364 1516
rect 1396 1484 1444 1516
rect 1476 1484 1524 1516
rect 1556 1484 1604 1516
rect 1636 1484 1684 1516
rect 1716 1484 1764 1516
rect 1796 1484 1844 1516
rect 1876 1484 1924 1516
rect 1956 1484 2004 1516
rect 2036 1484 2084 1516
rect 2116 1484 2164 1516
rect 2196 1484 2244 1516
rect 2276 1484 2324 1516
rect 2356 1484 2404 1516
rect 2436 1484 2484 1516
rect 2516 1484 2564 1516
rect 2596 1484 2644 1516
rect 2676 1484 2724 1516
rect 2756 1484 2804 1516
rect 2836 1484 2884 1516
rect 2916 1484 2964 1516
rect 2996 1484 3044 1516
rect 3076 1484 3124 1516
rect 3156 1484 3204 1516
rect 3236 1484 3284 1516
rect 3316 1484 3364 1516
rect 3396 1484 3444 1516
rect 3476 1484 3524 1516
rect 3556 1484 3604 1516
rect 3636 1484 3684 1516
rect 3716 1484 3764 1516
rect 3796 1484 3844 1516
rect 3876 1484 3924 1516
rect 3956 1484 4004 1516
rect 4036 1484 4084 1516
rect 4116 1484 4164 1516
rect 4196 1484 4244 1516
rect 4276 1484 4324 1516
rect 4356 1484 4404 1516
rect 4436 1484 4484 1516
rect 4516 1484 4564 1516
rect 4596 1484 4644 1516
rect 4676 1484 4724 1516
rect 4756 1484 4804 1516
rect 4836 1484 4840 1516
rect -800 1480 4840 1484
rect 4880 1516 5720 1520
rect 4880 1484 4884 1516
rect 4916 1484 5044 1516
rect 5076 1484 5204 1516
rect 5236 1484 5364 1516
rect 5396 1484 5524 1516
rect 5556 1484 5684 1516
rect 5716 1484 5720 1516
rect 4880 1480 5720 1484
rect -1520 1436 -840 1440
rect -1520 1404 -1516 1436
rect -1484 1404 -1356 1436
rect -1324 1404 -1196 1436
rect -1164 1404 -1036 1436
rect -1004 1404 -876 1436
rect -844 1404 -840 1436
rect -1520 1400 -840 1404
rect -800 1436 4840 1440
rect -800 1404 -796 1436
rect -764 1404 -716 1436
rect -684 1404 -636 1436
rect -604 1404 -556 1436
rect -524 1404 -476 1436
rect -444 1404 -396 1436
rect -364 1404 -316 1436
rect -284 1404 -236 1436
rect -204 1404 -156 1436
rect -124 1404 -76 1436
rect -44 1404 4 1436
rect 36 1404 84 1436
rect 116 1404 164 1436
rect 196 1404 244 1436
rect 276 1404 324 1436
rect 356 1404 404 1436
rect 436 1404 484 1436
rect 516 1404 564 1436
rect 596 1404 644 1436
rect 676 1404 724 1436
rect 756 1404 804 1436
rect 836 1404 884 1436
rect 916 1404 964 1436
rect 996 1404 1044 1436
rect 1076 1404 1124 1436
rect 1156 1404 1204 1436
rect 1236 1404 1284 1436
rect 1316 1404 1364 1436
rect 1396 1404 1444 1436
rect 1476 1404 1524 1436
rect 1556 1404 1604 1436
rect 1636 1404 1684 1436
rect 1716 1404 1764 1436
rect 1796 1404 1844 1436
rect 1876 1404 1924 1436
rect 1956 1404 2004 1436
rect 2036 1404 2084 1436
rect 2116 1404 2164 1436
rect 2196 1404 2244 1436
rect 2276 1404 2324 1436
rect 2356 1404 2404 1436
rect 2436 1404 2484 1436
rect 2516 1404 2564 1436
rect 2596 1404 2644 1436
rect 2676 1404 2724 1436
rect 2756 1404 2804 1436
rect 2836 1404 2884 1436
rect 2916 1404 2964 1436
rect 2996 1404 3044 1436
rect 3076 1404 3124 1436
rect 3156 1404 3204 1436
rect 3236 1404 3284 1436
rect 3316 1404 3364 1436
rect 3396 1404 3444 1436
rect 3476 1404 3524 1436
rect 3556 1404 3604 1436
rect 3636 1404 3684 1436
rect 3716 1404 3764 1436
rect 3796 1404 3844 1436
rect 3876 1404 3924 1436
rect 3956 1404 4004 1436
rect 4036 1404 4084 1436
rect 4116 1404 4164 1436
rect 4196 1404 4244 1436
rect 4276 1404 4324 1436
rect 4356 1404 4404 1436
rect 4436 1404 4484 1436
rect 4516 1404 4564 1436
rect 4596 1404 4644 1436
rect 4676 1404 4724 1436
rect 4756 1404 4804 1436
rect 4836 1404 4840 1436
rect -800 1400 4840 1404
rect 4880 1436 5720 1440
rect 4880 1404 4884 1436
rect 4916 1404 5044 1436
rect 5076 1404 5204 1436
rect 5236 1404 5364 1436
rect 5396 1404 5524 1436
rect 5556 1404 5684 1436
rect 5716 1404 5720 1436
rect 4880 1400 5720 1404
rect -1520 1356 -840 1360
rect -1520 1324 -1516 1356
rect -1484 1324 -1356 1356
rect -1324 1324 -1196 1356
rect -1164 1324 -1036 1356
rect -1004 1324 -876 1356
rect -844 1324 -840 1356
rect -1520 1320 -840 1324
rect -800 1356 4840 1360
rect -800 1324 -796 1356
rect -764 1324 -716 1356
rect -684 1324 -636 1356
rect -604 1324 -556 1356
rect -524 1324 -476 1356
rect -444 1324 -396 1356
rect -364 1324 -316 1356
rect -284 1324 -236 1356
rect -204 1324 -156 1356
rect -124 1324 -76 1356
rect -44 1324 4 1356
rect 36 1324 84 1356
rect 116 1324 164 1356
rect 196 1324 244 1356
rect 276 1324 324 1356
rect 356 1324 404 1356
rect 436 1324 484 1356
rect 516 1324 564 1356
rect 596 1324 644 1356
rect 676 1324 724 1356
rect 756 1324 804 1356
rect 836 1324 884 1356
rect 916 1324 964 1356
rect 996 1324 1044 1356
rect 1076 1324 1124 1356
rect 1156 1324 1204 1356
rect 1236 1324 1284 1356
rect 1316 1324 1364 1356
rect 1396 1324 1444 1356
rect 1476 1324 1524 1356
rect 1556 1324 1604 1356
rect 1636 1324 1684 1356
rect 1716 1324 1764 1356
rect 1796 1324 1844 1356
rect 1876 1324 1924 1356
rect 1956 1324 2004 1356
rect 2036 1324 2084 1356
rect 2116 1324 2164 1356
rect 2196 1324 2244 1356
rect 2276 1324 2324 1356
rect 2356 1324 2404 1356
rect 2436 1324 2484 1356
rect 2516 1324 2564 1356
rect 2596 1324 2644 1356
rect 2676 1324 2724 1356
rect 2756 1324 2804 1356
rect 2836 1324 2884 1356
rect 2916 1324 2964 1356
rect 2996 1324 3044 1356
rect 3076 1324 3124 1356
rect 3156 1324 3204 1356
rect 3236 1324 3284 1356
rect 3316 1324 3364 1356
rect 3396 1324 3444 1356
rect 3476 1324 3524 1356
rect 3556 1324 3604 1356
rect 3636 1324 3684 1356
rect 3716 1324 3764 1356
rect 3796 1324 3844 1356
rect 3876 1324 3924 1356
rect 3956 1324 4004 1356
rect 4036 1324 4084 1356
rect 4116 1324 4164 1356
rect 4196 1324 4244 1356
rect 4276 1324 4324 1356
rect 4356 1324 4404 1356
rect 4436 1324 4484 1356
rect 4516 1324 4564 1356
rect 4596 1324 4644 1356
rect 4676 1324 4724 1356
rect 4756 1324 4804 1356
rect 4836 1324 4840 1356
rect -800 1320 4840 1324
rect 4880 1356 5720 1360
rect 4880 1324 4884 1356
rect 4916 1324 5044 1356
rect 5076 1324 5204 1356
rect 5236 1324 5364 1356
rect 5396 1324 5524 1356
rect 5556 1324 5684 1356
rect 5716 1324 5720 1356
rect 4880 1320 5720 1324
rect -1520 1276 -840 1280
rect -1520 1244 -1516 1276
rect -1484 1244 -1356 1276
rect -1324 1244 -1196 1276
rect -1164 1244 -1036 1276
rect -1004 1244 -876 1276
rect -844 1244 -840 1276
rect -1520 1240 -840 1244
rect -800 1276 4840 1280
rect -800 1244 -796 1276
rect -764 1244 -716 1276
rect -684 1244 -636 1276
rect -604 1244 -556 1276
rect -524 1244 -476 1276
rect -444 1244 -396 1276
rect -364 1244 -316 1276
rect -284 1244 -236 1276
rect -204 1244 -156 1276
rect -124 1244 -76 1276
rect -44 1244 4 1276
rect 36 1244 84 1276
rect 116 1244 164 1276
rect 196 1244 244 1276
rect 276 1244 324 1276
rect 356 1244 404 1276
rect 436 1244 484 1276
rect 516 1244 564 1276
rect 596 1244 644 1276
rect 676 1244 724 1276
rect 756 1244 804 1276
rect 836 1244 884 1276
rect 916 1244 964 1276
rect 996 1244 1044 1276
rect 1076 1244 1124 1276
rect 1156 1244 1204 1276
rect 1236 1244 1284 1276
rect 1316 1244 1364 1276
rect 1396 1244 1444 1276
rect 1476 1244 1524 1276
rect 1556 1244 1604 1276
rect 1636 1244 1684 1276
rect 1716 1244 1764 1276
rect 1796 1244 1844 1276
rect 1876 1244 1924 1276
rect 1956 1244 2004 1276
rect 2036 1244 2084 1276
rect 2116 1244 2164 1276
rect 2196 1244 2244 1276
rect 2276 1244 2324 1276
rect 2356 1244 2404 1276
rect 2436 1244 2484 1276
rect 2516 1244 2564 1276
rect 2596 1244 2644 1276
rect 2676 1244 2724 1276
rect 2756 1244 2804 1276
rect 2836 1244 2884 1276
rect 2916 1244 2964 1276
rect 2996 1244 3044 1276
rect 3076 1244 3124 1276
rect 3156 1244 3204 1276
rect 3236 1244 3284 1276
rect 3316 1244 3364 1276
rect 3396 1244 3444 1276
rect 3476 1244 3524 1276
rect 3556 1244 3604 1276
rect 3636 1244 3684 1276
rect 3716 1244 3764 1276
rect 3796 1244 3844 1276
rect 3876 1244 3924 1276
rect 3956 1244 4004 1276
rect 4036 1244 4084 1276
rect 4116 1244 4164 1276
rect 4196 1244 4244 1276
rect 4276 1244 4324 1276
rect 4356 1244 4404 1276
rect 4436 1244 4484 1276
rect 4516 1244 4564 1276
rect 4596 1244 4644 1276
rect 4676 1244 4724 1276
rect 4756 1244 4804 1276
rect 4836 1244 4840 1276
rect -800 1240 4840 1244
rect 4880 1276 5720 1280
rect 4880 1244 4884 1276
rect 4916 1244 5044 1276
rect 5076 1244 5204 1276
rect 5236 1244 5364 1276
rect 5396 1244 5524 1276
rect 5556 1244 5684 1276
rect 5716 1244 5720 1276
rect 4880 1240 5720 1244
rect -1520 1196 -840 1200
rect -1520 1164 -1516 1196
rect -1484 1164 -1356 1196
rect -1324 1164 -1196 1196
rect -1164 1164 -1036 1196
rect -1004 1164 -876 1196
rect -844 1164 -840 1196
rect -1520 1160 -840 1164
rect -800 1196 4840 1200
rect -800 1164 -796 1196
rect -764 1164 -716 1196
rect -684 1164 -636 1196
rect -604 1164 -556 1196
rect -524 1164 -476 1196
rect -444 1164 -396 1196
rect -364 1164 -316 1196
rect -284 1164 -236 1196
rect -204 1164 -156 1196
rect -124 1164 -76 1196
rect -44 1164 4 1196
rect 36 1164 84 1196
rect 116 1164 164 1196
rect 196 1164 244 1196
rect 276 1164 324 1196
rect 356 1164 404 1196
rect 436 1164 484 1196
rect 516 1164 564 1196
rect 596 1164 644 1196
rect 676 1164 724 1196
rect 756 1164 804 1196
rect 836 1164 884 1196
rect 916 1164 964 1196
rect 996 1164 1044 1196
rect 1076 1164 1124 1196
rect 1156 1164 1204 1196
rect 1236 1164 1284 1196
rect 1316 1164 1364 1196
rect 1396 1164 1444 1196
rect 1476 1164 1524 1196
rect 1556 1164 1604 1196
rect 1636 1164 1684 1196
rect 1716 1164 1764 1196
rect 1796 1164 1844 1196
rect 1876 1164 1924 1196
rect 1956 1164 2004 1196
rect 2036 1164 2084 1196
rect 2116 1164 2164 1196
rect 2196 1164 2244 1196
rect 2276 1164 2324 1196
rect 2356 1164 2404 1196
rect 2436 1164 2484 1196
rect 2516 1164 2564 1196
rect 2596 1164 2644 1196
rect 2676 1164 2724 1196
rect 2756 1164 2804 1196
rect 2836 1164 2884 1196
rect 2916 1164 2964 1196
rect 2996 1164 3044 1196
rect 3076 1164 3124 1196
rect 3156 1164 3204 1196
rect 3236 1164 3284 1196
rect 3316 1164 3364 1196
rect 3396 1164 3444 1196
rect 3476 1164 3524 1196
rect 3556 1164 3604 1196
rect 3636 1164 3684 1196
rect 3716 1164 3764 1196
rect 3796 1164 3844 1196
rect 3876 1164 3924 1196
rect 3956 1164 4004 1196
rect 4036 1164 4084 1196
rect 4116 1164 4164 1196
rect 4196 1164 4244 1196
rect 4276 1164 4324 1196
rect 4356 1164 4404 1196
rect 4436 1164 4484 1196
rect 4516 1164 4564 1196
rect 4596 1164 4644 1196
rect 4676 1164 4724 1196
rect 4756 1164 4804 1196
rect 4836 1164 4840 1196
rect -800 1160 4840 1164
rect 4880 1196 5720 1200
rect 4880 1164 4884 1196
rect 4916 1164 5044 1196
rect 5076 1164 5204 1196
rect 5236 1164 5364 1196
rect 5396 1164 5524 1196
rect 5556 1164 5684 1196
rect 5716 1164 5720 1196
rect 4880 1160 5720 1164
rect -1520 1116 -840 1120
rect -1520 1084 -1516 1116
rect -1484 1084 -1356 1116
rect -1324 1084 -1196 1116
rect -1164 1084 -1036 1116
rect -1004 1084 -876 1116
rect -844 1084 -840 1116
rect -1520 1080 -840 1084
rect -800 1116 4840 1120
rect -800 1084 -796 1116
rect -764 1084 -716 1116
rect -684 1084 -636 1116
rect -604 1084 -556 1116
rect -524 1084 -476 1116
rect -444 1084 -396 1116
rect -364 1084 -316 1116
rect -284 1084 -236 1116
rect -204 1084 -156 1116
rect -124 1084 -76 1116
rect -44 1084 4 1116
rect 36 1084 84 1116
rect 116 1084 164 1116
rect 196 1084 244 1116
rect 276 1084 324 1116
rect 356 1084 404 1116
rect 436 1084 484 1116
rect 516 1084 564 1116
rect 596 1084 644 1116
rect 676 1084 724 1116
rect 756 1084 804 1116
rect 836 1084 884 1116
rect 916 1084 964 1116
rect 996 1084 1044 1116
rect 1076 1084 1124 1116
rect 1156 1084 1204 1116
rect 1236 1084 1284 1116
rect 1316 1084 1364 1116
rect 1396 1084 1444 1116
rect 1476 1084 1524 1116
rect 1556 1084 1604 1116
rect 1636 1084 1684 1116
rect 1716 1084 1764 1116
rect 1796 1084 1844 1116
rect 1876 1084 1924 1116
rect 1956 1084 2004 1116
rect 2036 1084 2084 1116
rect 2116 1084 2164 1116
rect 2196 1084 2244 1116
rect 2276 1084 2324 1116
rect 2356 1084 2404 1116
rect 2436 1084 2484 1116
rect 2516 1084 2564 1116
rect 2596 1084 2644 1116
rect 2676 1084 2724 1116
rect 2756 1084 2804 1116
rect 2836 1084 2884 1116
rect 2916 1084 2964 1116
rect 2996 1084 3044 1116
rect 3076 1084 3124 1116
rect 3156 1084 3204 1116
rect 3236 1084 3284 1116
rect 3316 1084 3364 1116
rect 3396 1084 3444 1116
rect 3476 1084 3524 1116
rect 3556 1084 3604 1116
rect 3636 1084 3684 1116
rect 3716 1084 3764 1116
rect 3796 1084 3844 1116
rect 3876 1084 3924 1116
rect 3956 1084 4004 1116
rect 4036 1084 4084 1116
rect 4116 1084 4164 1116
rect 4196 1084 4244 1116
rect 4276 1084 4324 1116
rect 4356 1084 4404 1116
rect 4436 1084 4484 1116
rect 4516 1084 4564 1116
rect 4596 1084 4644 1116
rect 4676 1084 4724 1116
rect 4756 1084 4804 1116
rect 4836 1084 4840 1116
rect -800 1080 4840 1084
rect 4880 1116 5720 1120
rect 4880 1084 4884 1116
rect 4916 1084 5044 1116
rect 5076 1084 5204 1116
rect 5236 1084 5364 1116
rect 5396 1084 5524 1116
rect 5556 1084 5684 1116
rect 5716 1084 5720 1116
rect 4880 1080 5720 1084
rect -1520 1036 -840 1040
rect -1520 1004 -1516 1036
rect -1484 1004 -1356 1036
rect -1324 1004 -1196 1036
rect -1164 1004 -1036 1036
rect -1004 1004 -876 1036
rect -844 1004 -840 1036
rect -1520 1000 -840 1004
rect -800 1036 4840 1040
rect -800 1004 -796 1036
rect -764 1004 -716 1036
rect -684 1004 -636 1036
rect -604 1004 -556 1036
rect -524 1004 -476 1036
rect -444 1004 -396 1036
rect -364 1004 -316 1036
rect -284 1004 -236 1036
rect -204 1004 -156 1036
rect -124 1004 -76 1036
rect -44 1004 4 1036
rect 36 1004 84 1036
rect 116 1004 164 1036
rect 196 1004 244 1036
rect 276 1004 324 1036
rect 356 1004 404 1036
rect 436 1004 484 1036
rect 516 1004 564 1036
rect 596 1004 644 1036
rect 676 1004 724 1036
rect 756 1004 804 1036
rect 836 1004 884 1036
rect 916 1004 964 1036
rect 996 1004 1044 1036
rect 1076 1004 1124 1036
rect 1156 1004 1204 1036
rect 1236 1004 1284 1036
rect 1316 1004 1364 1036
rect 1396 1004 1444 1036
rect 1476 1004 1524 1036
rect 1556 1004 1604 1036
rect 1636 1004 1684 1036
rect 1716 1004 1764 1036
rect 1796 1004 1844 1036
rect 1876 1004 1924 1036
rect 1956 1004 2004 1036
rect 2036 1004 2084 1036
rect 2116 1004 2164 1036
rect 2196 1004 2244 1036
rect 2276 1004 2324 1036
rect 2356 1004 2404 1036
rect 2436 1004 2484 1036
rect 2516 1004 2564 1036
rect 2596 1004 2644 1036
rect 2676 1004 2724 1036
rect 2756 1004 2804 1036
rect 2836 1004 2884 1036
rect 2916 1004 2964 1036
rect 2996 1004 3044 1036
rect 3076 1004 3124 1036
rect 3156 1004 3204 1036
rect 3236 1004 3284 1036
rect 3316 1004 3364 1036
rect 3396 1004 3444 1036
rect 3476 1004 3524 1036
rect 3556 1004 3604 1036
rect 3636 1004 3684 1036
rect 3716 1004 3764 1036
rect 3796 1004 3844 1036
rect 3876 1004 3924 1036
rect 3956 1004 4004 1036
rect 4036 1004 4084 1036
rect 4116 1004 4164 1036
rect 4196 1004 4244 1036
rect 4276 1004 4324 1036
rect 4356 1004 4404 1036
rect 4436 1004 4484 1036
rect 4516 1004 4564 1036
rect 4596 1004 4644 1036
rect 4676 1004 4724 1036
rect 4756 1004 4804 1036
rect 4836 1004 4840 1036
rect -800 1000 4840 1004
rect 4880 1036 5720 1040
rect 4880 1004 4884 1036
rect 4916 1004 5044 1036
rect 5076 1004 5204 1036
rect 5236 1004 5364 1036
rect 5396 1004 5524 1036
rect 5556 1004 5684 1036
rect 5716 1004 5720 1036
rect 4880 1000 5720 1004
rect -1520 956 -840 960
rect -1520 924 -1516 956
rect -1484 924 -1356 956
rect -1324 924 -1196 956
rect -1164 924 -1036 956
rect -1004 924 -876 956
rect -844 924 -840 956
rect -1520 920 -840 924
rect -800 956 4840 960
rect -800 924 -796 956
rect -764 924 -716 956
rect -684 924 -636 956
rect -604 924 -556 956
rect -524 924 -476 956
rect -444 924 -396 956
rect -364 924 -316 956
rect -284 924 -236 956
rect -204 924 -156 956
rect -124 924 -76 956
rect -44 924 4 956
rect 36 924 84 956
rect 116 924 164 956
rect 196 924 244 956
rect 276 924 324 956
rect 356 924 404 956
rect 436 924 484 956
rect 516 924 564 956
rect 596 924 644 956
rect 676 924 724 956
rect 756 924 804 956
rect 836 924 884 956
rect 916 924 964 956
rect 996 924 1044 956
rect 1076 924 1124 956
rect 1156 924 1204 956
rect 1236 924 1284 956
rect 1316 924 1364 956
rect 1396 924 1444 956
rect 1476 924 1524 956
rect 1556 924 1604 956
rect 1636 924 1684 956
rect 1716 924 1764 956
rect 1796 924 1844 956
rect 1876 924 1924 956
rect 1956 924 2004 956
rect 2036 924 2084 956
rect 2116 924 2164 956
rect 2196 924 2244 956
rect 2276 924 2324 956
rect 2356 924 2404 956
rect 2436 924 2484 956
rect 2516 924 2564 956
rect 2596 924 2644 956
rect 2676 924 2724 956
rect 2756 924 2804 956
rect 2836 924 2884 956
rect 2916 924 2964 956
rect 2996 924 3044 956
rect 3076 924 3124 956
rect 3156 924 3204 956
rect 3236 924 3284 956
rect 3316 924 3364 956
rect 3396 924 3444 956
rect 3476 924 3524 956
rect 3556 924 3604 956
rect 3636 924 3684 956
rect 3716 924 3764 956
rect 3796 924 3844 956
rect 3876 924 3924 956
rect 3956 924 4004 956
rect 4036 924 4084 956
rect 4116 924 4164 956
rect 4196 924 4244 956
rect 4276 924 4324 956
rect 4356 924 4404 956
rect 4436 924 4484 956
rect 4516 924 4564 956
rect 4596 924 4644 956
rect 4676 924 4724 956
rect 4756 924 4804 956
rect 4836 924 4840 956
rect -800 920 4840 924
rect 4880 956 5720 960
rect 4880 924 4884 956
rect 4916 924 5044 956
rect 5076 924 5204 956
rect 5236 924 5364 956
rect 5396 924 5524 956
rect 5556 924 5684 956
rect 5716 924 5720 956
rect 4880 920 5720 924
rect -1520 876 -840 880
rect -1520 844 -1516 876
rect -1484 844 -1356 876
rect -1324 844 -1196 876
rect -1164 844 -1036 876
rect -1004 844 -876 876
rect -844 844 -840 876
rect -1520 840 -840 844
rect -800 876 4840 880
rect -800 844 -796 876
rect -764 844 -716 876
rect -684 844 -636 876
rect -604 844 -556 876
rect -524 844 -476 876
rect -444 844 -396 876
rect -364 844 -316 876
rect -284 844 -236 876
rect -204 844 -156 876
rect -124 844 -76 876
rect -44 844 4 876
rect 36 844 84 876
rect 116 844 164 876
rect 196 844 244 876
rect 276 844 324 876
rect 356 844 404 876
rect 436 844 484 876
rect 516 844 564 876
rect 596 844 644 876
rect 676 844 724 876
rect 756 844 804 876
rect 836 844 884 876
rect 916 844 964 876
rect 996 844 1044 876
rect 1076 844 1124 876
rect 1156 844 1204 876
rect 1236 844 1284 876
rect 1316 844 1364 876
rect 1396 844 1444 876
rect 1476 844 1524 876
rect 1556 844 1604 876
rect 1636 844 1684 876
rect 1716 844 1764 876
rect 1796 844 1844 876
rect 1876 844 1924 876
rect 1956 844 2004 876
rect 2036 844 2084 876
rect 2116 844 2164 876
rect 2196 844 2244 876
rect 2276 844 2324 876
rect 2356 844 2404 876
rect 2436 844 2484 876
rect 2516 844 2564 876
rect 2596 844 2644 876
rect 2676 844 2724 876
rect 2756 844 2804 876
rect 2836 844 2884 876
rect 2916 844 2964 876
rect 2996 844 3044 876
rect 3076 844 3124 876
rect 3156 844 3204 876
rect 3236 844 3284 876
rect 3316 844 3364 876
rect 3396 844 3444 876
rect 3476 844 3524 876
rect 3556 844 3604 876
rect 3636 844 3684 876
rect 3716 844 3764 876
rect 3796 844 3844 876
rect 3876 844 3924 876
rect 3956 844 4004 876
rect 4036 844 4084 876
rect 4116 844 4164 876
rect 4196 844 4244 876
rect 4276 844 4324 876
rect 4356 844 4404 876
rect 4436 844 4484 876
rect 4516 844 4564 876
rect 4596 844 4644 876
rect 4676 844 4724 876
rect 4756 844 4804 876
rect 4836 844 4840 876
rect -800 840 4840 844
rect 4880 876 5720 880
rect 4880 844 4884 876
rect 4916 844 5044 876
rect 5076 844 5204 876
rect 5236 844 5364 876
rect 5396 844 5524 876
rect 5556 844 5684 876
rect 5716 844 5720 876
rect 4880 840 5720 844
rect -1520 796 -840 800
rect -1520 764 -1516 796
rect -1484 764 -1356 796
rect -1324 764 -1196 796
rect -1164 764 -1036 796
rect -1004 764 -876 796
rect -844 764 -840 796
rect -1520 760 -840 764
rect -800 796 4840 800
rect -800 764 -796 796
rect -764 764 -716 796
rect -684 764 -636 796
rect -604 764 -556 796
rect -524 764 -476 796
rect -444 764 -396 796
rect -364 764 -316 796
rect -284 764 -236 796
rect -204 764 -156 796
rect -124 764 -76 796
rect -44 764 4 796
rect 36 764 84 796
rect 116 764 164 796
rect 196 764 244 796
rect 276 764 324 796
rect 356 764 404 796
rect 436 764 484 796
rect 516 764 564 796
rect 596 764 644 796
rect 676 764 724 796
rect 756 764 804 796
rect 836 764 884 796
rect 916 764 964 796
rect 996 764 1044 796
rect 1076 764 1124 796
rect 1156 764 1204 796
rect 1236 764 1284 796
rect 1316 764 1364 796
rect 1396 764 1444 796
rect 1476 764 1524 796
rect 1556 764 1604 796
rect 1636 764 1684 796
rect 1716 764 1764 796
rect 1796 764 1844 796
rect 1876 764 1924 796
rect 1956 764 2004 796
rect 2036 764 2084 796
rect 2116 764 2164 796
rect 2196 764 2244 796
rect 2276 764 2324 796
rect 2356 764 2404 796
rect 2436 764 2484 796
rect 2516 764 2564 796
rect 2596 764 2644 796
rect 2676 764 2724 796
rect 2756 764 2804 796
rect 2836 764 2884 796
rect 2916 764 2964 796
rect 2996 764 3044 796
rect 3076 764 3124 796
rect 3156 764 3204 796
rect 3236 764 3284 796
rect 3316 764 3364 796
rect 3396 764 3444 796
rect 3476 764 3524 796
rect 3556 764 3604 796
rect 3636 764 3684 796
rect 3716 764 3764 796
rect 3796 764 3844 796
rect 3876 764 3924 796
rect 3956 764 4004 796
rect 4036 764 4084 796
rect 4116 764 4164 796
rect 4196 764 4244 796
rect 4276 764 4324 796
rect 4356 764 4404 796
rect 4436 764 4484 796
rect 4516 764 4564 796
rect 4596 764 4644 796
rect 4676 764 4724 796
rect 4756 764 4804 796
rect 4836 764 4840 796
rect -800 760 4840 764
rect 4880 796 5720 800
rect 4880 764 4884 796
rect 4916 764 5044 796
rect 5076 764 5204 796
rect 5236 764 5364 796
rect 5396 764 5524 796
rect 5556 764 5684 796
rect 5716 764 5720 796
rect 4880 760 5720 764
rect -1520 716 -840 720
rect -1520 684 -1516 716
rect -1484 684 -1356 716
rect -1324 684 -1196 716
rect -1164 684 -1036 716
rect -1004 684 -876 716
rect -844 684 -840 716
rect -1520 680 -840 684
rect -800 716 4840 720
rect -800 684 -796 716
rect -764 684 -716 716
rect -684 684 -636 716
rect -604 684 -556 716
rect -524 684 -476 716
rect -444 684 -396 716
rect -364 684 -316 716
rect -284 684 -236 716
rect -204 684 -156 716
rect -124 684 -76 716
rect -44 684 4 716
rect 36 684 84 716
rect 116 684 164 716
rect 196 684 244 716
rect 276 684 324 716
rect 356 684 404 716
rect 436 684 484 716
rect 516 684 564 716
rect 596 684 644 716
rect 676 684 724 716
rect 756 684 804 716
rect 836 684 884 716
rect 916 684 964 716
rect 996 684 1044 716
rect 1076 684 1124 716
rect 1156 684 1204 716
rect 1236 684 1284 716
rect 1316 684 1364 716
rect 1396 684 1444 716
rect 1476 684 1524 716
rect 1556 684 1604 716
rect 1636 684 1684 716
rect 1716 684 1764 716
rect 1796 684 1844 716
rect 1876 684 1924 716
rect 1956 684 2004 716
rect 2036 684 2084 716
rect 2116 684 2164 716
rect 2196 684 2244 716
rect 2276 684 2324 716
rect 2356 684 2404 716
rect 2436 684 2484 716
rect 2516 684 2564 716
rect 2596 684 2644 716
rect 2676 684 2724 716
rect 2756 684 2804 716
rect 2836 684 2884 716
rect 2916 684 2964 716
rect 2996 684 3044 716
rect 3076 684 3124 716
rect 3156 684 3204 716
rect 3236 684 3284 716
rect 3316 684 3364 716
rect 3396 684 3444 716
rect 3476 684 3524 716
rect 3556 684 3604 716
rect 3636 684 3684 716
rect 3716 684 3764 716
rect 3796 684 3844 716
rect 3876 684 3924 716
rect 3956 684 4004 716
rect 4036 684 4084 716
rect 4116 684 4164 716
rect 4196 684 4244 716
rect 4276 684 4324 716
rect 4356 684 4404 716
rect 4436 684 4484 716
rect 4516 684 4564 716
rect 4596 684 4644 716
rect 4676 684 4724 716
rect 4756 684 4804 716
rect 4836 684 4840 716
rect -800 680 4840 684
rect 4880 716 5720 720
rect 4880 684 4884 716
rect 4916 684 5044 716
rect 5076 684 5204 716
rect 5236 684 5364 716
rect 5396 684 5524 716
rect 5556 684 5684 716
rect 5716 684 5720 716
rect 4880 680 5720 684
rect -1520 636 -840 640
rect -1520 604 -1516 636
rect -1484 604 -1356 636
rect -1324 604 -1196 636
rect -1164 604 -1036 636
rect -1004 604 -876 636
rect -844 604 -840 636
rect -1520 600 -840 604
rect -800 636 4840 640
rect -800 604 -796 636
rect -764 604 -716 636
rect -684 604 -636 636
rect -604 604 -556 636
rect -524 604 -476 636
rect -444 604 -396 636
rect -364 604 -316 636
rect -284 604 -236 636
rect -204 604 -156 636
rect -124 604 -76 636
rect -44 604 4 636
rect 36 604 84 636
rect 116 604 164 636
rect 196 604 244 636
rect 276 604 324 636
rect 356 604 404 636
rect 436 604 484 636
rect 516 604 564 636
rect 596 604 644 636
rect 676 604 724 636
rect 756 604 804 636
rect 836 604 884 636
rect 916 604 964 636
rect 996 604 1044 636
rect 1076 604 1124 636
rect 1156 604 1204 636
rect 1236 604 1284 636
rect 1316 604 1364 636
rect 1396 604 1444 636
rect 1476 604 1524 636
rect 1556 604 1604 636
rect 1636 604 1684 636
rect 1716 604 1764 636
rect 1796 604 1844 636
rect 1876 604 1924 636
rect 1956 604 2004 636
rect 2036 604 2084 636
rect 2116 604 2164 636
rect 2196 604 2244 636
rect 2276 604 2324 636
rect 2356 604 2404 636
rect 2436 604 2484 636
rect 2516 604 2564 636
rect 2596 604 2644 636
rect 2676 604 2724 636
rect 2756 604 2804 636
rect 2836 604 2884 636
rect 2916 604 2964 636
rect 2996 604 3044 636
rect 3076 604 3124 636
rect 3156 604 3204 636
rect 3236 604 3284 636
rect 3316 604 3364 636
rect 3396 604 3444 636
rect 3476 604 3524 636
rect 3556 604 3604 636
rect 3636 604 3684 636
rect 3716 604 3764 636
rect 3796 604 3844 636
rect 3876 604 3924 636
rect 3956 604 4004 636
rect 4036 604 4084 636
rect 4116 604 4164 636
rect 4196 604 4244 636
rect 4276 604 4324 636
rect 4356 604 4404 636
rect 4436 604 4484 636
rect 4516 604 4564 636
rect 4596 604 4644 636
rect 4676 604 4724 636
rect 4756 604 4804 636
rect 4836 604 4840 636
rect -800 600 4840 604
rect 4880 636 5720 640
rect 4880 604 4884 636
rect 4916 604 5044 636
rect 5076 604 5204 636
rect 5236 604 5364 636
rect 5396 604 5524 636
rect 5556 604 5684 636
rect 5716 604 5720 636
rect 4880 600 5720 604
rect -1520 556 -840 560
rect -1520 524 -1516 556
rect -1484 524 -1356 556
rect -1324 524 -1196 556
rect -1164 524 -1036 556
rect -1004 524 -876 556
rect -844 524 -840 556
rect -1520 520 -840 524
rect -800 556 4840 560
rect -800 524 -796 556
rect -764 524 -716 556
rect -684 524 -636 556
rect -604 524 -556 556
rect -524 524 -476 556
rect -444 524 -396 556
rect -364 524 -316 556
rect -284 524 -236 556
rect -204 524 -156 556
rect -124 524 -76 556
rect -44 524 4 556
rect 36 524 84 556
rect 116 524 164 556
rect 196 524 244 556
rect 276 524 324 556
rect 356 524 404 556
rect 436 524 484 556
rect 516 524 564 556
rect 596 524 644 556
rect 676 524 724 556
rect 756 524 804 556
rect 836 524 884 556
rect 916 524 964 556
rect 996 524 1044 556
rect 1076 524 1124 556
rect 1156 524 1204 556
rect 1236 524 1284 556
rect 1316 524 1364 556
rect 1396 524 1444 556
rect 1476 524 1524 556
rect 1556 524 1604 556
rect 1636 524 1684 556
rect 1716 524 1764 556
rect 1796 524 1844 556
rect 1876 524 1924 556
rect 1956 524 2004 556
rect 2036 524 2084 556
rect 2116 524 2164 556
rect 2196 524 2244 556
rect 2276 524 2324 556
rect 2356 524 2404 556
rect 2436 524 2484 556
rect 2516 524 2564 556
rect 2596 524 2644 556
rect 2676 524 2724 556
rect 2756 524 2804 556
rect 2836 524 2884 556
rect 2916 524 2964 556
rect 2996 524 3044 556
rect 3076 524 3124 556
rect 3156 524 3204 556
rect 3236 524 3284 556
rect 3316 524 3364 556
rect 3396 524 3444 556
rect 3476 524 3524 556
rect 3556 524 3604 556
rect 3636 524 3684 556
rect 3716 524 3764 556
rect 3796 524 3844 556
rect 3876 524 3924 556
rect 3956 524 4004 556
rect 4036 524 4084 556
rect 4116 524 4164 556
rect 4196 524 4244 556
rect 4276 524 4324 556
rect 4356 524 4404 556
rect 4436 524 4484 556
rect 4516 524 4564 556
rect 4596 524 4644 556
rect 4676 524 4724 556
rect 4756 524 4804 556
rect 4836 524 4840 556
rect -800 520 4840 524
rect 4880 556 5720 560
rect 4880 524 4884 556
rect 4916 524 5044 556
rect 5076 524 5204 556
rect 5236 524 5364 556
rect 5396 524 5524 556
rect 5556 524 5684 556
rect 5716 524 5720 556
rect 4880 520 5720 524
rect -1520 476 -840 480
rect -1520 444 -1516 476
rect -1484 444 -1356 476
rect -1324 444 -1196 476
rect -1164 444 -1036 476
rect -1004 444 -876 476
rect -844 444 -840 476
rect -1520 440 -840 444
rect -800 476 4840 480
rect -800 444 -796 476
rect -764 444 -716 476
rect -684 444 -636 476
rect -604 444 -556 476
rect -524 444 -476 476
rect -444 444 -396 476
rect -364 444 -316 476
rect -284 444 -236 476
rect -204 444 -156 476
rect -124 444 -76 476
rect -44 444 4 476
rect 36 444 84 476
rect 116 444 164 476
rect 196 444 244 476
rect 276 444 324 476
rect 356 444 404 476
rect 436 444 484 476
rect 516 444 564 476
rect 596 444 644 476
rect 676 444 724 476
rect 756 444 804 476
rect 836 444 884 476
rect 916 444 964 476
rect 996 444 1044 476
rect 1076 444 1124 476
rect 1156 444 1204 476
rect 1236 444 1284 476
rect 1316 444 1364 476
rect 1396 444 1444 476
rect 1476 444 1524 476
rect 1556 444 1604 476
rect 1636 444 1684 476
rect 1716 444 1764 476
rect 1796 444 1844 476
rect 1876 444 1924 476
rect 1956 444 2004 476
rect 2036 444 2084 476
rect 2116 444 2164 476
rect 2196 444 2244 476
rect 2276 444 2324 476
rect 2356 444 2404 476
rect 2436 444 2484 476
rect 2516 444 2564 476
rect 2596 444 2644 476
rect 2676 444 2724 476
rect 2756 444 2804 476
rect 2836 444 2884 476
rect 2916 444 2964 476
rect 2996 444 3044 476
rect 3076 444 3124 476
rect 3156 444 3204 476
rect 3236 444 3284 476
rect 3316 444 3364 476
rect 3396 444 3444 476
rect 3476 444 3524 476
rect 3556 444 3604 476
rect 3636 444 3684 476
rect 3716 444 3764 476
rect 3796 444 3844 476
rect 3876 444 3924 476
rect 3956 444 4004 476
rect 4036 444 4084 476
rect 4116 444 4164 476
rect 4196 444 4244 476
rect 4276 444 4324 476
rect 4356 444 4404 476
rect 4436 444 4484 476
rect 4516 444 4564 476
rect 4596 444 4644 476
rect 4676 444 4724 476
rect 4756 444 4804 476
rect 4836 444 4840 476
rect -800 440 4840 444
rect 4880 476 5720 480
rect 4880 444 4884 476
rect 4916 444 5044 476
rect 5076 444 5204 476
rect 5236 444 5364 476
rect 5396 444 5524 476
rect 5556 444 5684 476
rect 5716 444 5720 476
rect 4880 440 5720 444
rect -1520 396 -840 400
rect -1520 364 -1516 396
rect -1484 364 -1356 396
rect -1324 364 -1196 396
rect -1164 364 -1036 396
rect -1004 364 -876 396
rect -844 364 -840 396
rect -1520 360 -840 364
rect -800 396 4840 400
rect -800 364 -796 396
rect -764 364 -716 396
rect -684 364 -636 396
rect -604 364 -556 396
rect -524 364 -476 396
rect -444 364 -396 396
rect -364 364 -316 396
rect -284 364 -236 396
rect -204 364 -156 396
rect -124 364 -76 396
rect -44 364 4 396
rect 36 364 84 396
rect 116 364 164 396
rect 196 364 244 396
rect 276 364 324 396
rect 356 364 404 396
rect 436 364 484 396
rect 516 364 564 396
rect 596 364 644 396
rect 676 364 724 396
rect 756 364 804 396
rect 836 364 884 396
rect 916 364 964 396
rect 996 364 1044 396
rect 1076 364 1124 396
rect 1156 364 1204 396
rect 1236 364 1284 396
rect 1316 364 1364 396
rect 1396 364 1444 396
rect 1476 364 1524 396
rect 1556 364 1604 396
rect 1636 364 1684 396
rect 1716 364 1764 396
rect 1796 364 1844 396
rect 1876 364 1924 396
rect 1956 364 2004 396
rect 2036 364 2084 396
rect 2116 364 2164 396
rect 2196 364 2244 396
rect 2276 364 2324 396
rect 2356 364 2404 396
rect 2436 364 2484 396
rect 2516 364 2564 396
rect 2596 364 2644 396
rect 2676 364 2724 396
rect 2756 364 2804 396
rect 2836 364 2884 396
rect 2916 364 2964 396
rect 2996 364 3044 396
rect 3076 364 3124 396
rect 3156 364 3204 396
rect 3236 364 3284 396
rect 3316 364 3364 396
rect 3396 364 3444 396
rect 3476 364 3524 396
rect 3556 364 3604 396
rect 3636 364 3684 396
rect 3716 364 3764 396
rect 3796 364 3844 396
rect 3876 364 3924 396
rect 3956 364 4004 396
rect 4036 364 4084 396
rect 4116 364 4164 396
rect 4196 364 4244 396
rect 4276 364 4324 396
rect 4356 364 4404 396
rect 4436 364 4484 396
rect 4516 364 4564 396
rect 4596 364 4644 396
rect 4676 364 4724 396
rect 4756 364 4804 396
rect 4836 364 4840 396
rect -800 360 4840 364
rect 4880 396 5720 400
rect 4880 364 4884 396
rect 4916 364 5044 396
rect 5076 364 5204 396
rect 5236 364 5364 396
rect 5396 364 5524 396
rect 5556 364 5684 396
rect 5716 364 5720 396
rect 4880 360 5720 364
rect -1520 316 -840 320
rect -1520 284 -1516 316
rect -1484 284 -1356 316
rect -1324 284 -1196 316
rect -1164 284 -1036 316
rect -1004 284 -876 316
rect -844 284 -840 316
rect -1520 280 -840 284
rect -800 316 4840 320
rect -800 284 -796 316
rect -764 284 -716 316
rect -684 284 -636 316
rect -604 284 -556 316
rect -524 284 -476 316
rect -444 284 -396 316
rect -364 284 -316 316
rect -284 284 -236 316
rect -204 284 -156 316
rect -124 284 -76 316
rect -44 284 4 316
rect 36 284 84 316
rect 116 284 164 316
rect 196 284 244 316
rect 276 284 324 316
rect 356 284 404 316
rect 436 284 484 316
rect 516 284 564 316
rect 596 284 644 316
rect 676 284 724 316
rect 756 284 804 316
rect 836 284 884 316
rect 916 284 964 316
rect 996 284 1044 316
rect 1076 284 1124 316
rect 1156 284 1204 316
rect 1236 284 1284 316
rect 1316 284 1364 316
rect 1396 284 1444 316
rect 1476 284 1524 316
rect 1556 284 1604 316
rect 1636 284 1684 316
rect 1716 284 1764 316
rect 1796 284 1844 316
rect 1876 284 1924 316
rect 1956 284 2004 316
rect 2036 284 2084 316
rect 2116 284 2164 316
rect 2196 284 2244 316
rect 2276 284 2324 316
rect 2356 284 2404 316
rect 2436 284 2484 316
rect 2516 284 2564 316
rect 2596 284 2644 316
rect 2676 284 2724 316
rect 2756 284 2804 316
rect 2836 284 2884 316
rect 2916 284 2964 316
rect 2996 284 3044 316
rect 3076 284 3124 316
rect 3156 284 3204 316
rect 3236 284 3284 316
rect 3316 284 3364 316
rect 3396 284 3444 316
rect 3476 284 3524 316
rect 3556 284 3604 316
rect 3636 284 3684 316
rect 3716 284 3764 316
rect 3796 284 3844 316
rect 3876 284 3924 316
rect 3956 284 4004 316
rect 4036 284 4084 316
rect 4116 284 4164 316
rect 4196 284 4244 316
rect 4276 284 4324 316
rect 4356 284 4404 316
rect 4436 284 4484 316
rect 4516 284 4564 316
rect 4596 284 4644 316
rect 4676 284 4724 316
rect 4756 284 4804 316
rect 4836 284 4840 316
rect -800 280 4840 284
rect 4880 316 5720 320
rect 4880 284 4884 316
rect 4916 284 5044 316
rect 5076 284 5204 316
rect 5236 284 5364 316
rect 5396 284 5524 316
rect 5556 284 5684 316
rect 5716 284 5720 316
rect 4880 280 5720 284
rect -1520 236 -840 240
rect -1520 204 -1516 236
rect -1484 204 -1356 236
rect -1324 204 -1196 236
rect -1164 204 -1036 236
rect -1004 204 -876 236
rect -844 204 -840 236
rect -1520 200 -840 204
rect -800 236 4840 240
rect -800 204 -796 236
rect -764 204 -716 236
rect -684 204 -636 236
rect -604 204 -556 236
rect -524 204 -476 236
rect -444 204 -396 236
rect -364 204 -316 236
rect -284 204 -236 236
rect -204 204 -156 236
rect -124 204 -76 236
rect -44 204 4 236
rect 36 204 84 236
rect 116 204 164 236
rect 196 204 244 236
rect 276 204 324 236
rect 356 204 404 236
rect 436 204 484 236
rect 516 204 564 236
rect 596 204 644 236
rect 676 204 724 236
rect 756 204 804 236
rect 836 204 884 236
rect 916 204 964 236
rect 996 204 1044 236
rect 1076 204 1124 236
rect 1156 204 1204 236
rect 1236 204 1284 236
rect 1316 204 1364 236
rect 1396 204 1444 236
rect 1476 204 1524 236
rect 1556 204 1604 236
rect 1636 204 1684 236
rect 1716 204 1764 236
rect 1796 204 1844 236
rect 1876 204 1924 236
rect 1956 204 2004 236
rect 2036 204 2084 236
rect 2116 204 2164 236
rect 2196 204 2244 236
rect 2276 204 2324 236
rect 2356 204 2404 236
rect 2436 204 2484 236
rect 2516 204 2564 236
rect 2596 204 2644 236
rect 2676 204 2724 236
rect 2756 204 2804 236
rect 2836 204 2884 236
rect 2916 204 2964 236
rect 2996 204 3044 236
rect 3076 204 3124 236
rect 3156 204 3204 236
rect 3236 204 3284 236
rect 3316 204 3364 236
rect 3396 204 3444 236
rect 3476 204 3524 236
rect 3556 204 3604 236
rect 3636 204 3684 236
rect 3716 204 3764 236
rect 3796 204 3844 236
rect 3876 204 3924 236
rect 3956 204 4004 236
rect 4036 204 4084 236
rect 4116 204 4164 236
rect 4196 204 4244 236
rect 4276 204 4324 236
rect 4356 204 4404 236
rect 4436 204 4484 236
rect 4516 204 4564 236
rect 4596 204 4644 236
rect 4676 204 4724 236
rect 4756 204 4804 236
rect 4836 204 4840 236
rect -800 200 4840 204
rect 4880 236 5720 240
rect 4880 204 4884 236
rect 4916 204 5044 236
rect 5076 204 5204 236
rect 5236 204 5364 236
rect 5396 204 5524 236
rect 5556 204 5684 236
rect 5716 204 5720 236
rect 4880 200 5720 204
rect -1520 156 -840 160
rect -1520 124 -1516 156
rect -1484 124 -1356 156
rect -1324 124 -1196 156
rect -1164 124 -1036 156
rect -1004 124 -876 156
rect -844 124 -840 156
rect -1520 120 -840 124
rect -800 156 4840 160
rect -800 124 -796 156
rect -764 124 -716 156
rect -684 124 -636 156
rect -604 124 -556 156
rect -524 124 -476 156
rect -444 124 -396 156
rect -364 124 -316 156
rect -284 124 -236 156
rect -204 124 -156 156
rect -124 124 -76 156
rect -44 124 4 156
rect 36 124 84 156
rect 116 124 164 156
rect 196 124 244 156
rect 276 124 324 156
rect 356 124 404 156
rect 436 124 484 156
rect 516 124 564 156
rect 596 124 644 156
rect 676 124 724 156
rect 756 124 804 156
rect 836 124 884 156
rect 916 124 964 156
rect 996 124 1044 156
rect 1076 124 1124 156
rect 1156 124 1204 156
rect 1236 124 1284 156
rect 1316 124 1364 156
rect 1396 124 1444 156
rect 1476 124 1524 156
rect 1556 124 1604 156
rect 1636 124 1684 156
rect 1716 124 1764 156
rect 1796 124 1844 156
rect 1876 124 1924 156
rect 1956 124 2004 156
rect 2036 124 2084 156
rect 2116 124 2164 156
rect 2196 124 2244 156
rect 2276 124 2324 156
rect 2356 124 2404 156
rect 2436 124 2484 156
rect 2516 124 2564 156
rect 2596 124 2644 156
rect 2676 124 2724 156
rect 2756 124 2804 156
rect 2836 124 2884 156
rect 2916 124 2964 156
rect 2996 124 3044 156
rect 3076 124 3124 156
rect 3156 124 3204 156
rect 3236 124 3284 156
rect 3316 124 3364 156
rect 3396 124 3444 156
rect 3476 124 3524 156
rect 3556 124 3604 156
rect 3636 124 3684 156
rect 3716 124 3764 156
rect 3796 124 3844 156
rect 3876 124 3924 156
rect 3956 124 4004 156
rect 4036 124 4084 156
rect 4116 124 4164 156
rect 4196 124 4244 156
rect 4276 124 4324 156
rect 4356 124 4404 156
rect 4436 124 4484 156
rect 4516 124 4564 156
rect 4596 124 4644 156
rect 4676 124 4724 156
rect 4756 124 4804 156
rect 4836 124 4840 156
rect -800 120 4840 124
rect 4880 156 5720 160
rect 4880 124 4884 156
rect 4916 124 5044 156
rect 5076 124 5204 156
rect 5236 124 5364 156
rect 5396 124 5524 156
rect 5556 124 5684 156
rect 5716 124 5720 156
rect 4880 120 5720 124
rect -1520 76 -840 80
rect -1520 44 -1516 76
rect -1484 44 -1356 76
rect -1324 44 -1196 76
rect -1164 44 -1036 76
rect -1004 44 -876 76
rect -844 44 -840 76
rect -1520 40 -840 44
rect -800 76 4840 80
rect -800 44 -796 76
rect -764 44 -716 76
rect -684 44 -636 76
rect -604 44 -556 76
rect -524 44 -476 76
rect -444 44 -396 76
rect -364 44 -316 76
rect -284 44 -236 76
rect -204 44 -156 76
rect -124 44 -76 76
rect -44 44 4 76
rect 36 44 84 76
rect 116 44 164 76
rect 196 44 244 76
rect 276 44 324 76
rect 356 44 404 76
rect 436 44 484 76
rect 516 44 564 76
rect 596 44 644 76
rect 676 44 724 76
rect 756 44 804 76
rect 836 44 884 76
rect 916 44 964 76
rect 996 44 1044 76
rect 1076 44 1124 76
rect 1156 44 1204 76
rect 1236 44 1284 76
rect 1316 44 1364 76
rect 1396 44 1444 76
rect 1476 44 1524 76
rect 1556 44 1604 76
rect 1636 44 1684 76
rect 1716 44 1764 76
rect 1796 44 1844 76
rect 1876 44 1924 76
rect 1956 44 2004 76
rect 2036 44 2084 76
rect 2116 44 2164 76
rect 2196 44 2244 76
rect 2276 44 2324 76
rect 2356 44 2404 76
rect 2436 44 2484 76
rect 2516 44 2564 76
rect 2596 44 2644 76
rect 2676 44 2724 76
rect 2756 44 2804 76
rect 2836 44 2884 76
rect 2916 44 2964 76
rect 2996 44 3044 76
rect 3076 44 3124 76
rect 3156 44 3204 76
rect 3236 44 3284 76
rect 3316 44 3364 76
rect 3396 44 3444 76
rect 3476 44 3524 76
rect 3556 44 3604 76
rect 3636 44 3684 76
rect 3716 44 3764 76
rect 3796 44 3844 76
rect 3876 44 3924 76
rect 3956 44 4004 76
rect 4036 44 4084 76
rect 4116 44 4164 76
rect 4196 44 4244 76
rect 4276 44 4324 76
rect 4356 44 4404 76
rect 4436 44 4484 76
rect 4516 44 4564 76
rect 4596 44 4644 76
rect 4676 44 4724 76
rect 4756 44 4804 76
rect 4836 44 4840 76
rect -800 40 4840 44
rect 4880 76 5720 80
rect 4880 44 4884 76
rect 4916 44 5044 76
rect 5076 44 5204 76
rect 5236 44 5364 76
rect 5396 44 5524 76
rect 5556 44 5684 76
rect 5716 44 5720 76
rect 4880 40 5720 44
rect -1520 -4 -840 0
rect -1520 -36 -1516 -4
rect -1484 -36 -1356 -4
rect -1324 -36 -1196 -4
rect -1164 -36 -1036 -4
rect -1004 -36 -876 -4
rect -844 -36 -840 -4
rect -1520 -40 -840 -36
rect -800 -4 4840 0
rect -800 -36 -796 -4
rect -764 -36 -716 -4
rect -684 -36 -636 -4
rect -604 -36 -556 -4
rect -524 -36 -476 -4
rect -444 -36 -396 -4
rect -364 -36 -316 -4
rect -284 -36 -236 -4
rect -204 -36 -156 -4
rect -124 -36 -76 -4
rect -44 -36 4 -4
rect 36 -36 84 -4
rect 116 -36 164 -4
rect 196 -36 244 -4
rect 276 -36 324 -4
rect 356 -36 404 -4
rect 436 -36 484 -4
rect 516 -36 564 -4
rect 596 -36 644 -4
rect 676 -36 724 -4
rect 756 -36 804 -4
rect 836 -36 884 -4
rect 916 -36 964 -4
rect 996 -36 1044 -4
rect 1076 -36 1124 -4
rect 1156 -36 1204 -4
rect 1236 -36 1284 -4
rect 1316 -36 1364 -4
rect 1396 -36 1444 -4
rect 1476 -36 1524 -4
rect 1556 -36 1604 -4
rect 1636 -36 1684 -4
rect 1716 -36 1764 -4
rect 1796 -36 1844 -4
rect 1876 -36 1924 -4
rect 1956 -36 2004 -4
rect 2036 -36 2084 -4
rect 2116 -36 2164 -4
rect 2196 -36 2244 -4
rect 2276 -36 2324 -4
rect 2356 -36 2404 -4
rect 2436 -36 2484 -4
rect 2516 -36 2564 -4
rect 2596 -36 2644 -4
rect 2676 -36 2724 -4
rect 2756 -36 2804 -4
rect 2836 -36 2884 -4
rect 2916 -36 2964 -4
rect 2996 -36 3044 -4
rect 3076 -36 3124 -4
rect 3156 -36 3204 -4
rect 3236 -36 3284 -4
rect 3316 -36 3364 -4
rect 3396 -36 3444 -4
rect 3476 -36 3524 -4
rect 3556 -36 3604 -4
rect 3636 -36 3684 -4
rect 3716 -36 3764 -4
rect 3796 -36 3844 -4
rect 3876 -36 3924 -4
rect 3956 -36 4004 -4
rect 4036 -36 4084 -4
rect 4116 -36 4164 -4
rect 4196 -36 4244 -4
rect 4276 -36 4324 -4
rect 4356 -36 4404 -4
rect 4436 -36 4484 -4
rect 4516 -36 4564 -4
rect 4596 -36 4644 -4
rect 4676 -36 4724 -4
rect 4756 -36 4804 -4
rect 4836 -36 4840 -4
rect -800 -40 4840 -36
rect 4880 -4 5720 0
rect 4880 -36 4884 -4
rect 4916 -36 5044 -4
rect 5076 -36 5204 -4
rect 5236 -36 5364 -4
rect 5396 -36 5524 -4
rect 5556 -36 5684 -4
rect 5716 -36 5720 -4
rect 4880 -40 5720 -36
rect -1520 -84 -840 -80
rect -1520 -116 -1516 -84
rect -1484 -116 -1356 -84
rect -1324 -116 -1196 -84
rect -1164 -116 -1036 -84
rect -1004 -116 -876 -84
rect -844 -116 -840 -84
rect -1520 -120 -840 -116
rect -800 -84 4840 -80
rect -800 -116 -796 -84
rect -764 -116 -716 -84
rect -684 -116 -636 -84
rect -604 -116 -556 -84
rect -524 -116 -476 -84
rect -444 -116 -396 -84
rect -364 -116 -316 -84
rect -284 -116 -236 -84
rect -204 -116 -156 -84
rect -124 -116 -76 -84
rect -44 -116 4 -84
rect 36 -116 84 -84
rect 116 -116 164 -84
rect 196 -116 244 -84
rect 276 -116 324 -84
rect 356 -116 404 -84
rect 436 -116 484 -84
rect 516 -116 564 -84
rect 596 -116 644 -84
rect 676 -116 724 -84
rect 756 -116 804 -84
rect 836 -116 884 -84
rect 916 -116 964 -84
rect 996 -116 1044 -84
rect 1076 -116 1124 -84
rect 1156 -116 1204 -84
rect 1236 -116 1284 -84
rect 1316 -116 1364 -84
rect 1396 -116 1444 -84
rect 1476 -116 1524 -84
rect 1556 -116 1604 -84
rect 1636 -116 1684 -84
rect 1716 -116 1764 -84
rect 1796 -116 1844 -84
rect 1876 -116 1924 -84
rect 1956 -116 2004 -84
rect 2036 -116 2084 -84
rect 2116 -116 2164 -84
rect 2196 -116 2244 -84
rect 2276 -116 2324 -84
rect 2356 -116 2404 -84
rect 2436 -116 2484 -84
rect 2516 -116 2564 -84
rect 2596 -116 2644 -84
rect 2676 -116 2724 -84
rect 2756 -116 2804 -84
rect 2836 -116 2884 -84
rect 2916 -116 2964 -84
rect 2996 -116 3044 -84
rect 3076 -116 3124 -84
rect 3156 -116 3204 -84
rect 3236 -116 3284 -84
rect 3316 -116 3364 -84
rect 3396 -116 3444 -84
rect 3476 -116 3524 -84
rect 3556 -116 3604 -84
rect 3636 -116 3684 -84
rect 3716 -116 3764 -84
rect 3796 -116 3844 -84
rect 3876 -116 3924 -84
rect 3956 -116 4004 -84
rect 4036 -116 4084 -84
rect 4116 -116 4164 -84
rect 4196 -116 4244 -84
rect 4276 -116 4324 -84
rect 4356 -116 4404 -84
rect 4436 -116 4484 -84
rect 4516 -116 4564 -84
rect 4596 -116 4644 -84
rect 4676 -116 4724 -84
rect 4756 -116 4804 -84
rect 4836 -116 4840 -84
rect -800 -120 4840 -116
rect 4880 -84 5720 -80
rect 4880 -116 4884 -84
rect 4916 -116 5044 -84
rect 5076 -116 5204 -84
rect 5236 -116 5364 -84
rect 5396 -116 5524 -84
rect 5556 -116 5684 -84
rect 5716 -116 5720 -84
rect 4880 -120 5720 -116
<< labels >>
rlabel metal3 -960 5600 -920 5640 0 p1
rlabel metal3 -1120 5600 -1080 5640 0 p2
rlabel metal3 -1280 5600 -1240 5640 0 p0
rlabel metal3 -1440 5600 -1400 5640 0 s
rlabel metal3 -1520 5600 -1480 5640 0 vdda
port 2 nsew
rlabel metal3 4960 5600 5000 5640 0 n
rlabel metal3 5120 5600 5160 5640 0 z
rlabel metal3 5280 5600 5320 5640 0 y
rlabel metal3 5440 5600 5480 5640 0 x
port 4 nsew
rlabel metal3 5600 5600 5640 5640 0 io
port 1 nsew
rlabel metal3 5680 5600 5720 5640 0 vssa
port 3 nsew
<< end >>
