magic
tech sky130A
timestamp 1640965787
<< metal1 >>
rect 10720 351395 10760 351400
rect 10720 351365 10725 351395
rect 10755 351365 10760 351395
rect 10720 351360 10760 351365
rect 10800 351395 10840 351400
rect 10800 351365 10805 351395
rect 10835 351365 10840 351395
rect 10800 351360 10840 351365
rect 10880 351395 10920 351400
rect 10880 351365 10885 351395
rect 10915 351365 10920 351395
rect 10880 351360 10920 351365
rect 10960 351395 11000 351400
rect 10960 351365 10965 351395
rect 10995 351365 11000 351395
rect 10960 351360 11000 351365
rect 11040 351395 11080 351400
rect 11040 351365 11045 351395
rect 11075 351365 11080 351395
rect 11040 351360 11080 351365
rect 11120 351395 11160 351400
rect 11120 351365 11125 351395
rect 11155 351365 11160 351395
rect 11120 351360 11160 351365
rect 11200 351395 11240 351400
rect 11200 351365 11205 351395
rect 11235 351365 11240 351395
rect 11200 351360 11240 351365
rect 11280 351395 11320 351400
rect 11280 351365 11285 351395
rect 11315 351365 11320 351395
rect 11280 351360 11320 351365
rect 11360 351395 11400 351400
rect 11360 351365 11365 351395
rect 11395 351365 11400 351395
rect 11360 351360 11400 351365
rect 11440 351395 11480 351400
rect 11440 351365 11445 351395
rect 11475 351365 11480 351395
rect 11440 351360 11480 351365
rect 11520 351395 11560 351400
rect 11520 351365 11525 351395
rect 11555 351365 11560 351395
rect 11520 351360 11560 351365
rect 11600 351395 11640 351400
rect 11600 351365 11605 351395
rect 11635 351365 11640 351395
rect 11600 351360 11640 351365
rect 11680 351395 11720 351400
rect 11680 351365 11685 351395
rect 11715 351365 11720 351395
rect 11680 351360 11720 351365
rect 11760 351395 11800 351400
rect 11760 351365 11765 351395
rect 11795 351365 11800 351395
rect 11760 351360 11800 351365
rect 11840 351395 11880 351400
rect 11840 351365 11845 351395
rect 11875 351365 11880 351395
rect 11840 351360 11880 351365
rect 11920 351395 11960 351400
rect 11920 351365 11925 351395
rect 11955 351365 11960 351395
rect 11920 351360 11960 351365
rect 12000 351395 12040 351400
rect 12000 351365 12005 351395
rect 12035 351365 12040 351395
rect 12000 351360 12040 351365
rect 12080 351395 12120 351400
rect 12080 351365 12085 351395
rect 12115 351365 12120 351395
rect 12080 351360 12120 351365
rect 12160 351395 12200 351400
rect 12160 351365 12165 351395
rect 12195 351365 12200 351395
rect 12160 351360 12200 351365
rect 12240 351395 12280 351400
rect 12240 351365 12245 351395
rect 12275 351365 12280 351395
rect 12240 351360 12280 351365
rect 12320 351395 12360 351400
rect 12320 351365 12325 351395
rect 12355 351365 12360 351395
rect 12320 351360 12360 351365
rect 12400 351395 12440 351400
rect 12400 351365 12405 351395
rect 12435 351365 12440 351395
rect 12400 351360 12440 351365
rect 12480 351395 12520 351400
rect 12480 351365 12485 351395
rect 12515 351365 12520 351395
rect 12480 351360 12520 351365
rect 12560 351395 12600 351400
rect 12560 351365 12565 351395
rect 12595 351365 12600 351395
rect 12560 351360 12600 351365
rect 12640 351395 12680 351400
rect 12640 351365 12645 351395
rect 12675 351365 12680 351395
rect 12640 351360 12680 351365
rect 12720 351395 12760 351400
rect 12720 351365 12725 351395
rect 12755 351365 12760 351395
rect 12720 351360 12760 351365
rect 12800 351395 12840 351400
rect 12800 351365 12805 351395
rect 12835 351365 12840 351395
rect 12800 351360 12840 351365
rect 12880 351395 12920 351400
rect 12880 351365 12885 351395
rect 12915 351365 12920 351395
rect 12880 351360 12920 351365
rect 12960 351395 13000 351400
rect 12960 351365 12965 351395
rect 12995 351365 13000 351395
rect 12960 351360 13000 351365
rect 13040 351395 13080 351400
rect 13040 351365 13045 351395
rect 13075 351365 13080 351395
rect 13040 351360 13080 351365
rect 13120 351395 13160 351400
rect 13120 351365 13125 351395
rect 13155 351365 13160 351395
rect 13120 351360 13160 351365
rect 13200 351395 13240 351400
rect 13200 351365 13205 351395
rect 13235 351365 13240 351395
rect 13200 351360 13240 351365
rect 13280 351395 13320 351400
rect 13280 351365 13285 351395
rect 13315 351365 13320 351395
rect 13280 351360 13320 351365
rect 13360 351395 13400 351400
rect 13360 351365 13365 351395
rect 13395 351365 13400 351395
rect 13360 351360 13400 351365
rect 13440 351395 13480 351400
rect 13440 351365 13445 351395
rect 13475 351365 13480 351395
rect 13440 351360 13480 351365
rect 13520 351395 13560 351400
rect 13520 351365 13525 351395
rect 13555 351365 13560 351395
rect 13520 351360 13560 351365
rect 13600 351395 13640 351400
rect 13600 351365 13605 351395
rect 13635 351365 13640 351395
rect 13600 351360 13640 351365
rect 13680 351395 13720 351400
rect 13680 351365 13685 351395
rect 13715 351365 13720 351395
rect 13680 351360 13720 351365
rect 13760 351395 13800 351400
rect 13760 351365 13765 351395
rect 13795 351365 13800 351395
rect 13760 351360 13800 351365
rect 13840 351395 13880 351400
rect 13840 351365 13845 351395
rect 13875 351365 13880 351395
rect 13840 351360 13880 351365
rect 13920 351395 13960 351400
rect 13920 351365 13925 351395
rect 13955 351365 13960 351395
rect 13920 351360 13960 351365
rect 14000 351395 14040 351400
rect 14000 351365 14005 351395
rect 14035 351365 14040 351395
rect 14000 351360 14040 351365
rect 14080 351395 14120 351400
rect 14080 351365 14085 351395
rect 14115 351365 14120 351395
rect 14080 351360 14120 351365
rect 14160 351395 14200 351400
rect 14160 351365 14165 351395
rect 14195 351365 14200 351395
rect 14160 351360 14200 351365
rect 14240 351395 14280 351400
rect 14240 351365 14245 351395
rect 14275 351365 14280 351395
rect 14240 351360 14280 351365
rect 14320 351395 14360 351400
rect 14320 351365 14325 351395
rect 14355 351365 14360 351395
rect 14320 351360 14360 351365
rect 14400 351395 14440 351400
rect 14400 351365 14405 351395
rect 14435 351365 14440 351395
rect 14400 351360 14440 351365
rect 14480 351395 14520 351400
rect 14480 351365 14485 351395
rect 14515 351365 14520 351395
rect 14480 351360 14520 351365
rect 14560 351395 14600 351400
rect 14560 351365 14565 351395
rect 14595 351365 14600 351395
rect 14560 351360 14600 351365
rect 14640 351395 14680 351400
rect 14640 351365 14645 351395
rect 14675 351365 14680 351395
rect 14640 351360 14680 351365
rect 14720 351395 14760 351400
rect 14720 351365 14725 351395
rect 14755 351365 14760 351395
rect 14720 351360 14760 351365
rect 14800 351395 14840 351400
rect 14800 351365 14805 351395
rect 14835 351365 14840 351395
rect 14800 351360 14840 351365
rect 14880 351395 14920 351400
rect 14880 351365 14885 351395
rect 14915 351365 14920 351395
rect 14880 351360 14920 351365
rect 14960 351395 15000 351400
rect 14960 351365 14965 351395
rect 14995 351365 15000 351395
rect 14960 351360 15000 351365
rect 15040 351395 15080 351400
rect 15040 351365 15045 351395
rect 15075 351365 15080 351395
rect 15040 351360 15080 351365
rect 15120 351395 15160 351400
rect 15120 351365 15125 351395
rect 15155 351365 15160 351395
rect 15120 351360 15160 351365
rect 15200 351395 15240 351400
rect 15200 351365 15205 351395
rect 15235 351365 15240 351395
rect 15200 351360 15240 351365
rect 15280 351395 15320 351400
rect 15280 351365 15285 351395
rect 15315 351365 15320 351395
rect 15280 351360 15320 351365
rect 15360 351395 15400 351400
rect 15360 351365 15365 351395
rect 15395 351365 15400 351395
rect 15360 351360 15400 351365
rect 15440 351395 15480 351400
rect 15440 351365 15445 351395
rect 15475 351365 15480 351395
rect 15440 351360 15480 351365
rect 15520 351395 15560 351400
rect 15520 351365 15525 351395
rect 15555 351365 15560 351395
rect 15520 351360 15560 351365
rect 15600 351395 15640 351400
rect 15600 351365 15605 351395
rect 15635 351365 15640 351395
rect 15600 351360 15640 351365
rect 15680 351395 15720 351400
rect 15680 351365 15685 351395
rect 15715 351365 15720 351395
rect 15680 351360 15720 351365
rect 15760 351395 15800 351400
rect 15760 351365 15765 351395
rect 15795 351365 15800 351395
rect 15760 351360 15800 351365
rect 15840 351395 15880 351400
rect 15840 351365 15845 351395
rect 15875 351365 15880 351395
rect 15840 351360 15880 351365
rect 15920 351395 15960 351400
rect 15920 351365 15925 351395
rect 15955 351365 15960 351395
rect 15920 351360 15960 351365
rect 16000 351395 16040 351400
rect 16000 351365 16005 351395
rect 16035 351365 16040 351395
rect 16000 351360 16040 351365
rect 16080 351395 16120 351400
rect 16080 351365 16085 351395
rect 16115 351365 16120 351395
rect 16080 351360 16120 351365
rect 16160 351395 16200 351400
rect 16160 351365 16165 351395
rect 16195 351365 16200 351395
rect 16160 351360 16200 351365
rect 16240 351395 16280 351400
rect 16240 351365 16245 351395
rect 16275 351365 16280 351395
rect 16240 351360 16280 351365
rect 16320 351395 16360 351400
rect 16320 351365 16325 351395
rect 16355 351365 16360 351395
rect 16320 351360 16360 351365
rect 16400 351395 16440 351400
rect 16400 351365 16405 351395
rect 16435 351365 16440 351395
rect 16400 351360 16440 351365
rect 16480 351395 16520 351400
rect 16480 351365 16485 351395
rect 16515 351365 16520 351395
rect 16480 351360 16520 351365
rect 16560 351395 16600 351400
rect 16560 351365 16565 351395
rect 16595 351365 16600 351395
rect 16560 351360 16600 351365
rect 16640 351395 16680 351400
rect 16640 351365 16645 351395
rect 16675 351365 16680 351395
rect 16640 351360 16680 351365
rect 16720 351395 16760 351400
rect 16720 351365 16725 351395
rect 16755 351365 16760 351395
rect 16720 351360 16760 351365
rect 16800 351395 16840 351400
rect 16800 351365 16805 351395
rect 16835 351365 16840 351395
rect 16800 351360 16840 351365
rect 16880 351395 16920 351400
rect 16880 351365 16885 351395
rect 16915 351365 16920 351395
rect 16880 351360 16920 351365
rect 16960 351395 17000 351400
rect 16960 351365 16965 351395
rect 16995 351365 17000 351395
rect 16960 351360 17000 351365
rect 17040 351395 17080 351400
rect 17040 351365 17045 351395
rect 17075 351365 17080 351395
rect 17040 351360 17080 351365
rect 17120 351395 17160 351400
rect 17120 351365 17125 351395
rect 17155 351365 17160 351395
rect 17120 351360 17160 351365
rect 17200 351395 17240 351400
rect 17200 351365 17205 351395
rect 17235 351365 17240 351395
rect 17200 351360 17240 351365
rect 17280 351395 17320 351400
rect 17280 351365 17285 351395
rect 17315 351365 17320 351395
rect 17280 351360 17320 351365
rect 17360 351395 17400 351400
rect 17360 351365 17365 351395
rect 17395 351365 17400 351395
rect 17360 351360 17400 351365
rect 17440 351395 17480 351400
rect 17440 351365 17445 351395
rect 17475 351365 17480 351395
rect 17440 351360 17480 351365
rect 17520 351395 17560 351400
rect 17520 351365 17525 351395
rect 17555 351365 17560 351395
rect 17520 351360 17560 351365
rect 17600 351395 17640 351400
rect 17600 351365 17605 351395
rect 17635 351365 17640 351395
rect 17600 351360 17640 351365
rect 17680 351395 17720 351400
rect 17680 351365 17685 351395
rect 17715 351365 17720 351395
rect 17680 351360 17720 351365
rect 17760 351395 17800 351400
rect 17760 351365 17765 351395
rect 17795 351365 17800 351395
rect 17760 351360 17800 351365
rect 17840 351395 17880 351400
rect 17840 351365 17845 351395
rect 17875 351365 17880 351395
rect 17840 351360 17880 351365
rect 17920 351395 17960 351400
rect 17920 351365 17925 351395
rect 17955 351365 17960 351395
rect 17920 351360 17960 351365
rect 18000 351395 18040 351400
rect 18000 351365 18005 351395
rect 18035 351365 18040 351395
rect 18000 351360 18040 351365
rect 18080 351395 18120 351400
rect 18080 351365 18085 351395
rect 18115 351365 18120 351395
rect 18080 351360 18120 351365
rect 18160 351395 18200 351400
rect 18160 351365 18165 351395
rect 18195 351365 18200 351395
rect 18160 351360 18200 351365
rect 18240 351395 18280 351400
rect 18240 351365 18245 351395
rect 18275 351365 18280 351395
rect 18240 351360 18280 351365
rect 18320 351395 18360 351400
rect 18320 351365 18325 351395
rect 18355 351365 18360 351395
rect 18320 351360 18360 351365
rect 18400 351395 18440 351400
rect 18400 351365 18405 351395
rect 18435 351365 18440 351395
rect 18400 351360 18440 351365
rect 18480 351395 18520 351400
rect 18480 351365 18485 351395
rect 18515 351365 18520 351395
rect 18480 351360 18520 351365
rect 18560 351395 18600 351400
rect 18560 351365 18565 351395
rect 18595 351365 18600 351395
rect 18560 351360 18600 351365
rect 18640 351395 18680 351400
rect 18640 351365 18645 351395
rect 18675 351365 18680 351395
rect 18640 351360 18680 351365
rect 18720 351395 18760 351400
rect 18720 351365 18725 351395
rect 18755 351365 18760 351395
rect 18720 351360 18760 351365
rect 18800 351395 18840 351400
rect 18800 351365 18805 351395
rect 18835 351365 18840 351395
rect 18800 351360 18840 351365
rect 18880 351395 18920 351400
rect 18880 351365 18885 351395
rect 18915 351365 18920 351395
rect 18880 351360 18920 351365
rect 18960 351395 19000 351400
rect 18960 351365 18965 351395
rect 18995 351365 19000 351395
rect 18960 351360 19000 351365
rect 19040 351395 19080 351400
rect 19040 351365 19045 351395
rect 19075 351365 19080 351395
rect 19040 351360 19080 351365
rect 19120 351395 19160 351400
rect 19120 351365 19125 351395
rect 19155 351365 19160 351395
rect 19120 351360 19160 351365
rect 19200 351395 19240 351400
rect 19200 351365 19205 351395
rect 19235 351365 19240 351395
rect 19200 351360 19240 351365
rect 19280 351395 19320 351400
rect 19280 351365 19285 351395
rect 19315 351365 19320 351395
rect 19280 351360 19320 351365
rect 19360 351395 19400 351400
rect 19360 351365 19365 351395
rect 19395 351365 19400 351395
rect 19360 351360 19400 351365
rect 19440 351395 19480 351400
rect 19440 351365 19445 351395
rect 19475 351365 19480 351395
rect 19440 351360 19480 351365
rect 19520 351395 19560 351400
rect 19520 351365 19525 351395
rect 19555 351365 19560 351395
rect 19520 351360 19560 351365
rect 19600 351395 19640 351400
rect 19600 351365 19605 351395
rect 19635 351365 19640 351395
rect 19600 351360 19640 351365
rect 19680 351395 19720 351400
rect 19680 351365 19685 351395
rect 19715 351365 19720 351395
rect 19680 351360 19720 351365
rect 19840 351395 19880 351400
rect 19840 351365 19845 351395
rect 19875 351365 19880 351395
rect 19840 351360 19880 351365
rect 10720 351235 10760 351240
rect 10720 351205 10725 351235
rect 10755 351205 10760 351235
rect 10720 351200 10760 351205
rect 10800 351235 10840 351240
rect 10800 351205 10805 351235
rect 10835 351205 10840 351235
rect 10800 351200 10840 351205
rect 10880 351235 10920 351240
rect 10880 351205 10885 351235
rect 10915 351205 10920 351235
rect 10880 351200 10920 351205
rect 10960 351235 11000 351240
rect 10960 351205 10965 351235
rect 10995 351205 11000 351235
rect 10960 351200 11000 351205
rect 11040 351235 11080 351240
rect 11040 351205 11045 351235
rect 11075 351205 11080 351235
rect 11040 351200 11080 351205
rect 11120 351235 11160 351240
rect 11120 351205 11125 351235
rect 11155 351205 11160 351235
rect 11120 351200 11160 351205
rect 11200 351235 11240 351240
rect 11200 351205 11205 351235
rect 11235 351205 11240 351235
rect 11200 351200 11240 351205
rect 11280 351235 11320 351240
rect 11280 351205 11285 351235
rect 11315 351205 11320 351235
rect 11280 351200 11320 351205
rect 11360 351235 11400 351240
rect 11360 351205 11365 351235
rect 11395 351205 11400 351235
rect 11360 351200 11400 351205
rect 11440 351235 11480 351240
rect 11440 351205 11445 351235
rect 11475 351205 11480 351235
rect 11440 351200 11480 351205
rect 11520 351235 11560 351240
rect 11520 351205 11525 351235
rect 11555 351205 11560 351235
rect 11520 351200 11560 351205
rect 11600 351235 11640 351240
rect 11600 351205 11605 351235
rect 11635 351205 11640 351235
rect 11600 351200 11640 351205
rect 11680 351235 11720 351240
rect 11680 351205 11685 351235
rect 11715 351205 11720 351235
rect 11680 351200 11720 351205
rect 11760 351235 11800 351240
rect 11760 351205 11765 351235
rect 11795 351205 11800 351235
rect 11760 351200 11800 351205
rect 11840 351235 11880 351240
rect 11840 351205 11845 351235
rect 11875 351205 11880 351235
rect 11840 351200 11880 351205
rect 11920 351235 11960 351240
rect 11920 351205 11925 351235
rect 11955 351205 11960 351235
rect 11920 351200 11960 351205
rect 12000 351235 12040 351240
rect 12000 351205 12005 351235
rect 12035 351205 12040 351235
rect 12000 351200 12040 351205
rect 12080 351235 12120 351240
rect 12080 351205 12085 351235
rect 12115 351205 12120 351235
rect 12080 351200 12120 351205
rect 12160 351235 12200 351240
rect 12160 351205 12165 351235
rect 12195 351205 12200 351235
rect 12160 351200 12200 351205
rect 12240 351235 12280 351240
rect 12240 351205 12245 351235
rect 12275 351205 12280 351235
rect 12240 351200 12280 351205
rect 12320 351235 12360 351240
rect 12320 351205 12325 351235
rect 12355 351205 12360 351235
rect 12320 351200 12360 351205
rect 12400 351235 12440 351240
rect 12400 351205 12405 351235
rect 12435 351205 12440 351235
rect 12400 351200 12440 351205
rect 12480 351235 12520 351240
rect 12480 351205 12485 351235
rect 12515 351205 12520 351235
rect 12480 351200 12520 351205
rect 12560 351235 12600 351240
rect 12560 351205 12565 351235
rect 12595 351205 12600 351235
rect 12560 351200 12600 351205
rect 12640 351235 12680 351240
rect 12640 351205 12645 351235
rect 12675 351205 12680 351235
rect 12640 351200 12680 351205
rect 12720 351235 12760 351240
rect 12720 351205 12725 351235
rect 12755 351205 12760 351235
rect 12720 351200 12760 351205
rect 12800 351235 12840 351240
rect 12800 351205 12805 351235
rect 12835 351205 12840 351235
rect 12800 351200 12840 351205
rect 12880 351235 12920 351240
rect 12880 351205 12885 351235
rect 12915 351205 12920 351235
rect 12880 351200 12920 351205
rect 12960 351235 13000 351240
rect 12960 351205 12965 351235
rect 12995 351205 13000 351235
rect 12960 351200 13000 351205
rect 13040 351235 13080 351240
rect 13040 351205 13045 351235
rect 13075 351205 13080 351235
rect 13040 351200 13080 351205
rect 13120 351235 13160 351240
rect 13120 351205 13125 351235
rect 13155 351205 13160 351235
rect 13120 351200 13160 351205
rect 13200 351235 13240 351240
rect 13200 351205 13205 351235
rect 13235 351205 13240 351235
rect 13200 351200 13240 351205
rect 13280 351235 13320 351240
rect 13280 351205 13285 351235
rect 13315 351205 13320 351235
rect 13280 351200 13320 351205
rect 13360 351235 13400 351240
rect 13360 351205 13365 351235
rect 13395 351205 13400 351235
rect 13360 351200 13400 351205
rect 13440 351235 13480 351240
rect 13440 351205 13445 351235
rect 13475 351205 13480 351235
rect 13440 351200 13480 351205
rect 13520 351235 13560 351240
rect 13520 351205 13525 351235
rect 13555 351205 13560 351235
rect 13520 351200 13560 351205
rect 13600 351235 13640 351240
rect 13600 351205 13605 351235
rect 13635 351205 13640 351235
rect 13600 351200 13640 351205
rect 13680 351235 13720 351240
rect 13680 351205 13685 351235
rect 13715 351205 13720 351235
rect 13680 351200 13720 351205
rect 13760 351235 13800 351240
rect 13760 351205 13765 351235
rect 13795 351205 13800 351235
rect 13760 351200 13800 351205
rect 13840 351235 13880 351240
rect 13840 351205 13845 351235
rect 13875 351205 13880 351235
rect 13840 351200 13880 351205
rect 13920 351235 13960 351240
rect 13920 351205 13925 351235
rect 13955 351205 13960 351235
rect 13920 351200 13960 351205
rect 14000 351235 14040 351240
rect 14000 351205 14005 351235
rect 14035 351205 14040 351235
rect 14000 351200 14040 351205
rect 14080 351235 14120 351240
rect 14080 351205 14085 351235
rect 14115 351205 14120 351235
rect 14080 351200 14120 351205
rect 14160 351235 14200 351240
rect 14160 351205 14165 351235
rect 14195 351205 14200 351235
rect 14160 351200 14200 351205
rect 14240 351235 14280 351240
rect 14240 351205 14245 351235
rect 14275 351205 14280 351235
rect 14240 351200 14280 351205
rect 14320 351235 14360 351240
rect 14320 351205 14325 351235
rect 14355 351205 14360 351235
rect 14320 351200 14360 351205
rect 14400 351235 14440 351240
rect 14400 351205 14405 351235
rect 14435 351205 14440 351235
rect 14400 351200 14440 351205
rect 14480 351235 14520 351240
rect 14480 351205 14485 351235
rect 14515 351205 14520 351235
rect 14480 351200 14520 351205
rect 14560 351235 14600 351240
rect 14560 351205 14565 351235
rect 14595 351205 14600 351235
rect 14560 351200 14600 351205
rect 14640 351235 14680 351240
rect 14640 351205 14645 351235
rect 14675 351205 14680 351235
rect 14640 351200 14680 351205
rect 14720 351235 14760 351240
rect 14720 351205 14725 351235
rect 14755 351205 14760 351235
rect 14720 351200 14760 351205
rect 14800 351235 14840 351240
rect 14800 351205 14805 351235
rect 14835 351205 14840 351235
rect 14800 351200 14840 351205
rect 14880 351235 14920 351240
rect 14880 351205 14885 351235
rect 14915 351205 14920 351235
rect 14880 351200 14920 351205
rect 14960 351235 15000 351240
rect 14960 351205 14965 351235
rect 14995 351205 15000 351235
rect 14960 351200 15000 351205
rect 15040 351235 15080 351240
rect 15040 351205 15045 351235
rect 15075 351205 15080 351235
rect 15040 351200 15080 351205
rect 15120 351235 15160 351240
rect 15120 351205 15125 351235
rect 15155 351205 15160 351235
rect 15120 351200 15160 351205
rect 15200 351235 15240 351240
rect 15200 351205 15205 351235
rect 15235 351205 15240 351235
rect 15200 351200 15240 351205
rect 15280 351235 15320 351240
rect 15280 351205 15285 351235
rect 15315 351205 15320 351235
rect 15280 351200 15320 351205
rect 15360 351235 15400 351240
rect 15360 351205 15365 351235
rect 15395 351205 15400 351235
rect 15360 351200 15400 351205
rect 15440 351235 15480 351240
rect 15440 351205 15445 351235
rect 15475 351205 15480 351235
rect 15440 351200 15480 351205
rect 15520 351235 15560 351240
rect 15520 351205 15525 351235
rect 15555 351205 15560 351235
rect 15520 351200 15560 351205
rect 15600 351235 15640 351240
rect 15600 351205 15605 351235
rect 15635 351205 15640 351235
rect 15600 351200 15640 351205
rect 15680 351235 15720 351240
rect 15680 351205 15685 351235
rect 15715 351205 15720 351235
rect 15680 351200 15720 351205
rect 15760 351235 15800 351240
rect 15760 351205 15765 351235
rect 15795 351205 15800 351235
rect 15760 351200 15800 351205
rect 15840 351235 15880 351240
rect 15840 351205 15845 351235
rect 15875 351205 15880 351235
rect 15840 351200 15880 351205
rect 15920 351235 15960 351240
rect 15920 351205 15925 351235
rect 15955 351205 15960 351235
rect 15920 351200 15960 351205
rect 16000 351235 16040 351240
rect 16000 351205 16005 351235
rect 16035 351205 16040 351235
rect 16000 351200 16040 351205
rect 16080 351235 16120 351240
rect 16080 351205 16085 351235
rect 16115 351205 16120 351235
rect 16080 351200 16120 351205
rect 16160 351235 16200 351240
rect 16160 351205 16165 351235
rect 16195 351205 16200 351235
rect 16160 351200 16200 351205
rect 16240 351235 16280 351240
rect 16240 351205 16245 351235
rect 16275 351205 16280 351235
rect 16240 351200 16280 351205
rect 16320 351235 16360 351240
rect 16320 351205 16325 351235
rect 16355 351205 16360 351235
rect 16320 351200 16360 351205
rect 16400 351235 16440 351240
rect 16400 351205 16405 351235
rect 16435 351205 16440 351235
rect 16400 351200 16440 351205
rect 16480 351235 16520 351240
rect 16480 351205 16485 351235
rect 16515 351205 16520 351235
rect 16480 351200 16520 351205
rect 16560 351235 16600 351240
rect 16560 351205 16565 351235
rect 16595 351205 16600 351235
rect 16560 351200 16600 351205
rect 16640 351235 16680 351240
rect 16640 351205 16645 351235
rect 16675 351205 16680 351235
rect 16640 351200 16680 351205
rect 16720 351235 16760 351240
rect 16720 351205 16725 351235
rect 16755 351205 16760 351235
rect 16720 351200 16760 351205
rect 16800 351235 16840 351240
rect 16800 351205 16805 351235
rect 16835 351205 16840 351235
rect 16800 351200 16840 351205
rect 16880 351235 16920 351240
rect 16880 351205 16885 351235
rect 16915 351205 16920 351235
rect 16880 351200 16920 351205
rect 16960 351235 17000 351240
rect 16960 351205 16965 351235
rect 16995 351205 17000 351235
rect 16960 351200 17000 351205
rect 17040 351235 17080 351240
rect 17040 351205 17045 351235
rect 17075 351205 17080 351235
rect 17040 351200 17080 351205
rect 17120 351235 17160 351240
rect 17120 351205 17125 351235
rect 17155 351205 17160 351235
rect 17120 351200 17160 351205
rect 17200 351235 17240 351240
rect 17200 351205 17205 351235
rect 17235 351205 17240 351235
rect 17200 351200 17240 351205
rect 17280 351235 17320 351240
rect 17280 351205 17285 351235
rect 17315 351205 17320 351235
rect 17280 351200 17320 351205
rect 17360 351235 17400 351240
rect 17360 351205 17365 351235
rect 17395 351205 17400 351235
rect 17360 351200 17400 351205
rect 17440 351235 17480 351240
rect 17440 351205 17445 351235
rect 17475 351205 17480 351235
rect 17440 351200 17480 351205
rect 17520 351235 17560 351240
rect 17520 351205 17525 351235
rect 17555 351205 17560 351235
rect 17520 351200 17560 351205
rect 17600 351235 17640 351240
rect 17600 351205 17605 351235
rect 17635 351205 17640 351235
rect 17600 351200 17640 351205
rect 17680 351235 17720 351240
rect 17680 351205 17685 351235
rect 17715 351205 17720 351235
rect 17680 351200 17720 351205
rect 17760 351235 17800 351240
rect 17760 351205 17765 351235
rect 17795 351205 17800 351235
rect 17760 351200 17800 351205
rect 17840 351235 17880 351240
rect 17840 351205 17845 351235
rect 17875 351205 17880 351235
rect 17840 351200 17880 351205
rect 17920 351235 17960 351240
rect 17920 351205 17925 351235
rect 17955 351205 17960 351235
rect 17920 351200 17960 351205
rect 18000 351235 18040 351240
rect 18000 351205 18005 351235
rect 18035 351205 18040 351235
rect 18000 351200 18040 351205
rect 18080 351235 18120 351240
rect 18080 351205 18085 351235
rect 18115 351205 18120 351235
rect 18080 351200 18120 351205
rect 18160 351235 18200 351240
rect 18160 351205 18165 351235
rect 18195 351205 18200 351235
rect 18160 351200 18200 351205
rect 18240 351235 18280 351240
rect 18240 351205 18245 351235
rect 18275 351205 18280 351235
rect 18240 351200 18280 351205
rect 18320 351235 18360 351240
rect 18320 351205 18325 351235
rect 18355 351205 18360 351235
rect 18320 351200 18360 351205
rect 18400 351235 18440 351240
rect 18400 351205 18405 351235
rect 18435 351205 18440 351235
rect 18400 351200 18440 351205
rect 18480 351235 18520 351240
rect 18480 351205 18485 351235
rect 18515 351205 18520 351235
rect 18480 351200 18520 351205
rect 18560 351235 18600 351240
rect 18560 351205 18565 351235
rect 18595 351205 18600 351235
rect 18560 351200 18600 351205
rect 18640 351235 18680 351240
rect 18640 351205 18645 351235
rect 18675 351205 18680 351235
rect 18640 351200 18680 351205
rect 18720 351235 18760 351240
rect 18720 351205 18725 351235
rect 18755 351205 18760 351235
rect 18720 351200 18760 351205
rect 18800 351235 18840 351240
rect 18800 351205 18805 351235
rect 18835 351205 18840 351235
rect 18800 351200 18840 351205
rect 18880 351235 18920 351240
rect 18880 351205 18885 351235
rect 18915 351205 18920 351235
rect 18880 351200 18920 351205
rect 18960 351235 19000 351240
rect 18960 351205 18965 351235
rect 18995 351205 19000 351235
rect 18960 351200 19000 351205
rect 19040 351235 19080 351240
rect 19040 351205 19045 351235
rect 19075 351205 19080 351235
rect 19040 351200 19080 351205
rect 19120 351235 19160 351240
rect 19120 351205 19125 351235
rect 19155 351205 19160 351235
rect 19120 351200 19160 351205
rect 19200 351235 19240 351240
rect 19200 351205 19205 351235
rect 19235 351205 19240 351235
rect 19200 351200 19240 351205
rect 19280 351235 19320 351240
rect 19280 351205 19285 351235
rect 19315 351205 19320 351235
rect 19280 351200 19320 351205
rect 19360 351235 19400 351240
rect 19360 351205 19365 351235
rect 19395 351205 19400 351235
rect 19360 351200 19400 351205
rect 19440 351235 19480 351240
rect 19440 351205 19445 351235
rect 19475 351205 19480 351235
rect 19440 351200 19480 351205
rect 19520 351235 19560 351240
rect 19520 351205 19525 351235
rect 19555 351205 19560 351235
rect 19520 351200 19560 351205
rect 19600 351235 19640 351240
rect 19600 351205 19605 351235
rect 19635 351205 19640 351235
rect 19600 351200 19640 351205
rect 19680 351235 19720 351240
rect 19680 351205 19685 351235
rect 19715 351205 19720 351235
rect 19680 351200 19720 351205
rect 19840 351235 19880 351240
rect 19840 351205 19845 351235
rect 19875 351205 19880 351235
rect 19840 351200 19880 351205
rect 19680 351155 19720 351160
rect 19680 351125 19685 351155
rect 19715 351125 19720 351155
rect 19680 351120 19720 351125
rect 19840 351155 19880 351160
rect 19840 351125 19845 351155
rect 19875 351125 19880 351155
rect 19840 351120 19880 351125
rect 19680 351075 19720 351080
rect 19680 351045 19685 351075
rect 19715 351045 19720 351075
rect 19680 351040 19720 351045
rect 19840 351075 19880 351080
rect 19840 351045 19845 351075
rect 19875 351045 19880 351075
rect 19840 351040 19880 351045
rect 19680 350995 19720 351000
rect 19680 350965 19685 350995
rect 19715 350965 19720 350995
rect 19680 350960 19720 350965
rect 19840 350995 19880 351000
rect 19840 350965 19845 350995
rect 19875 350965 19880 350995
rect 19840 350960 19880 350965
rect 19680 350915 19720 350920
rect 19680 350885 19685 350915
rect 19715 350885 19720 350915
rect 19680 350880 19720 350885
rect 19840 350915 19880 350920
rect 19840 350885 19845 350915
rect 19875 350885 19880 350915
rect 19840 350880 19880 350885
rect 19680 350835 19720 350840
rect 19680 350805 19685 350835
rect 19715 350805 19720 350835
rect 19680 350800 19720 350805
rect 19840 350835 19880 350840
rect 19840 350805 19845 350835
rect 19875 350805 19880 350835
rect 19840 350800 19880 350805
rect 19680 350755 19720 350760
rect 19680 350725 19685 350755
rect 19715 350725 19720 350755
rect 19680 350720 19720 350725
rect 19840 350755 19880 350760
rect 19840 350725 19845 350755
rect 19875 350725 19880 350755
rect 19840 350720 19880 350725
rect 19680 350675 19720 350680
rect 19680 350645 19685 350675
rect 19715 350645 19720 350675
rect 19680 350640 19720 350645
rect 19840 350675 19880 350680
rect 19840 350645 19845 350675
rect 19875 350645 19880 350675
rect 19840 350640 19880 350645
rect 19680 350595 19720 350600
rect 19680 350565 19685 350595
rect 19715 350565 19720 350595
rect 19680 350560 19720 350565
rect 19840 350595 19880 350600
rect 19840 350565 19845 350595
rect 19875 350565 19880 350595
rect 19840 350560 19880 350565
rect 19680 350515 19720 350520
rect 19680 350485 19685 350515
rect 19715 350485 19720 350515
rect 19680 350480 19720 350485
rect 19840 350515 19880 350520
rect 19840 350485 19845 350515
rect 19875 350485 19880 350515
rect 19840 350480 19880 350485
rect 19680 350435 19720 350440
rect 19680 350405 19685 350435
rect 19715 350405 19720 350435
rect 19680 350400 19720 350405
rect 19840 350435 19880 350440
rect 19840 350405 19845 350435
rect 19875 350405 19880 350435
rect 19840 350400 19880 350405
rect 19680 350355 19720 350360
rect 19680 350325 19685 350355
rect 19715 350325 19720 350355
rect 19680 350320 19720 350325
rect 19840 350355 19880 350360
rect 19840 350325 19845 350355
rect 19875 350325 19880 350355
rect 19840 350320 19880 350325
rect 19680 350275 19720 350280
rect 19680 350245 19685 350275
rect 19715 350245 19720 350275
rect 19680 350240 19720 350245
rect 19840 350275 19880 350280
rect 19840 350245 19845 350275
rect 19875 350245 19880 350275
rect 19840 350240 19880 350245
rect 19680 350195 19720 350200
rect 19680 350165 19685 350195
rect 19715 350165 19720 350195
rect 19680 350160 19720 350165
rect 19840 350195 19880 350200
rect 19840 350165 19845 350195
rect 19875 350165 19880 350195
rect 19840 350160 19880 350165
rect 19680 350115 19720 350120
rect 19680 350085 19685 350115
rect 19715 350085 19720 350115
rect 19680 350080 19720 350085
rect 19840 350115 19880 350120
rect 19840 350085 19845 350115
rect 19875 350085 19880 350115
rect 19840 350080 19880 350085
rect 19680 350035 19720 350040
rect 19680 350005 19685 350035
rect 19715 350005 19720 350035
rect 19680 350000 19720 350005
rect 19840 350035 19880 350040
rect 19840 350005 19845 350035
rect 19875 350005 19880 350035
rect 19840 350000 19880 350005
rect 19680 349955 19720 349960
rect 19680 349925 19685 349955
rect 19715 349925 19720 349955
rect 19680 349920 19720 349925
rect 19840 349955 19880 349960
rect 19840 349925 19845 349955
rect 19875 349925 19880 349955
rect 19840 349920 19880 349925
rect 19680 349875 19720 349880
rect 19680 349845 19685 349875
rect 19715 349845 19720 349875
rect 19680 349840 19720 349845
rect 19840 349875 19880 349880
rect 19840 349845 19845 349875
rect 19875 349845 19880 349875
rect 19840 349840 19880 349845
rect 19680 349795 19720 349800
rect 19680 349765 19685 349795
rect 19715 349765 19720 349795
rect 19680 349760 19720 349765
rect 19840 349795 19880 349800
rect 19840 349765 19845 349795
rect 19875 349765 19880 349795
rect 19840 349760 19880 349765
rect 19680 349715 19720 349720
rect 19680 349685 19685 349715
rect 19715 349685 19720 349715
rect 19680 349680 19720 349685
rect 19840 349715 19880 349720
rect 19840 349685 19845 349715
rect 19875 349685 19880 349715
rect 19840 349680 19880 349685
rect 19680 349635 19720 349640
rect 19680 349605 19685 349635
rect 19715 349605 19720 349635
rect 19680 349600 19720 349605
rect 19840 349635 19880 349640
rect 19840 349605 19845 349635
rect 19875 349605 19880 349635
rect 19840 349600 19880 349605
rect 19680 349555 19720 349560
rect 19680 349525 19685 349555
rect 19715 349525 19720 349555
rect 19680 349520 19720 349525
rect 19840 349555 19880 349560
rect 19840 349525 19845 349555
rect 19875 349525 19880 349555
rect 19840 349520 19880 349525
rect 19680 349475 19720 349480
rect 19680 349445 19685 349475
rect 19715 349445 19720 349475
rect 19680 349440 19720 349445
rect 19840 349475 19880 349480
rect 19840 349445 19845 349475
rect 19875 349445 19880 349475
rect 19840 349440 19880 349445
rect 19680 349395 19720 349400
rect 19680 349365 19685 349395
rect 19715 349365 19720 349395
rect 19680 349360 19720 349365
rect 19840 349395 19880 349400
rect 19840 349365 19845 349395
rect 19875 349365 19880 349395
rect 19840 349360 19880 349365
rect 19680 349315 19720 349320
rect 19680 349285 19685 349315
rect 19715 349285 19720 349315
rect 19680 349280 19720 349285
rect 19840 349315 19880 349320
rect 19840 349285 19845 349315
rect 19875 349285 19880 349315
rect 19840 349280 19880 349285
rect 19680 349235 19720 349240
rect 19680 349205 19685 349235
rect 19715 349205 19720 349235
rect 19680 349200 19720 349205
rect 19840 349235 19880 349240
rect 19840 349205 19845 349235
rect 19875 349205 19880 349235
rect 19840 349200 19880 349205
rect 19680 349155 19720 349160
rect 19680 349125 19685 349155
rect 19715 349125 19720 349155
rect 19680 349120 19720 349125
rect 19840 349155 19880 349160
rect 19840 349125 19845 349155
rect 19875 349125 19880 349155
rect 19840 349120 19880 349125
rect 19680 349075 19720 349080
rect 19680 349045 19685 349075
rect 19715 349045 19720 349075
rect 19680 349040 19720 349045
rect 19840 349075 19880 349080
rect 19840 349045 19845 349075
rect 19875 349045 19880 349075
rect 19840 349040 19880 349045
rect 19680 348995 19720 349000
rect 19680 348965 19685 348995
rect 19715 348965 19720 348995
rect 19680 348960 19720 348965
rect 19840 348995 19880 349000
rect 19840 348965 19845 348995
rect 19875 348965 19880 348995
rect 19840 348960 19880 348965
rect 19680 348915 19720 348920
rect 19680 348885 19685 348915
rect 19715 348885 19720 348915
rect 19680 348880 19720 348885
rect 19840 348915 19880 348920
rect 19840 348885 19845 348915
rect 19875 348885 19880 348915
rect 19840 348880 19880 348885
rect 19680 348835 19720 348840
rect 19680 348805 19685 348835
rect 19715 348805 19720 348835
rect 19680 348800 19720 348805
rect 19840 348835 19880 348840
rect 19840 348805 19845 348835
rect 19875 348805 19880 348835
rect 19840 348800 19880 348805
rect 19680 348755 19720 348760
rect 19680 348725 19685 348755
rect 19715 348725 19720 348755
rect 19680 348720 19720 348725
rect 19840 348755 19880 348760
rect 19840 348725 19845 348755
rect 19875 348725 19880 348755
rect 19840 348720 19880 348725
rect 19680 348675 19720 348680
rect 19680 348645 19685 348675
rect 19715 348645 19720 348675
rect 19680 348640 19720 348645
rect 19840 348675 19880 348680
rect 19840 348645 19845 348675
rect 19875 348645 19880 348675
rect 19840 348640 19880 348645
rect 19680 348595 19720 348600
rect 19680 348565 19685 348595
rect 19715 348565 19720 348595
rect 19680 348560 19720 348565
rect 19840 348595 19880 348600
rect 19840 348565 19845 348595
rect 19875 348565 19880 348595
rect 19840 348560 19880 348565
rect 19680 348515 19720 348520
rect 19680 348485 19685 348515
rect 19715 348485 19720 348515
rect 19680 348480 19720 348485
rect 19840 348515 19880 348520
rect 19840 348485 19845 348515
rect 19875 348485 19880 348515
rect 19840 348480 19880 348485
rect 19680 348435 19720 348440
rect 19680 348405 19685 348435
rect 19715 348405 19720 348435
rect 19680 348400 19720 348405
rect 19840 348435 19880 348440
rect 19840 348405 19845 348435
rect 19875 348405 19880 348435
rect 19840 348400 19880 348405
rect 19680 348355 19720 348360
rect 19680 348325 19685 348355
rect 19715 348325 19720 348355
rect 19680 348320 19720 348325
rect 19840 348355 19880 348360
rect 19840 348325 19845 348355
rect 19875 348325 19880 348355
rect 19840 348320 19880 348325
rect 19680 348275 19720 348280
rect 19680 348245 19685 348275
rect 19715 348245 19720 348275
rect 19680 348240 19720 348245
rect 19840 348275 19880 348280
rect 19840 348245 19845 348275
rect 19875 348245 19880 348275
rect 19840 348240 19880 348245
rect 19680 348195 19720 348200
rect 19680 348165 19685 348195
rect 19715 348165 19720 348195
rect 19680 348160 19720 348165
rect 19840 348195 19880 348200
rect 19840 348165 19845 348195
rect 19875 348165 19880 348195
rect 19840 348160 19880 348165
rect 19680 348115 19720 348120
rect 19680 348085 19685 348115
rect 19715 348085 19720 348115
rect 19680 348080 19720 348085
rect 19840 348115 19880 348120
rect 19840 348085 19845 348115
rect 19875 348085 19880 348115
rect 19840 348080 19880 348085
rect 19680 348035 19720 348040
rect 19680 348005 19685 348035
rect 19715 348005 19720 348035
rect 19680 348000 19720 348005
rect 19840 348035 19880 348040
rect 19840 348005 19845 348035
rect 19875 348005 19880 348035
rect 19840 348000 19880 348005
rect 19680 347955 19720 347960
rect 19680 347925 19685 347955
rect 19715 347925 19720 347955
rect 19680 347920 19720 347925
rect 19840 347955 19880 347960
rect 19840 347925 19845 347955
rect 19875 347925 19880 347955
rect 19840 347920 19880 347925
rect 19680 347875 19720 347880
rect 19680 347845 19685 347875
rect 19715 347845 19720 347875
rect 19680 347840 19720 347845
rect 19840 347875 19880 347880
rect 19840 347845 19845 347875
rect 19875 347845 19880 347875
rect 19840 347840 19880 347845
rect 19680 347795 19720 347800
rect 19680 347765 19685 347795
rect 19715 347765 19720 347795
rect 19680 347760 19720 347765
rect 19840 347795 19880 347800
rect 19840 347765 19845 347795
rect 19875 347765 19880 347795
rect 19840 347760 19880 347765
rect 19680 347715 19720 347720
rect 19680 347685 19685 347715
rect 19715 347685 19720 347715
rect 19680 347680 19720 347685
rect 19840 347715 19880 347720
rect 19840 347685 19845 347715
rect 19875 347685 19880 347715
rect 19840 347680 19880 347685
rect 19680 347635 19720 347640
rect 19680 347605 19685 347635
rect 19715 347605 19720 347635
rect 19680 347600 19720 347605
rect 19840 347635 19880 347640
rect 19840 347605 19845 347635
rect 19875 347605 19880 347635
rect 19840 347600 19880 347605
rect 19680 347555 19720 347560
rect 19680 347525 19685 347555
rect 19715 347525 19720 347555
rect 19680 347520 19720 347525
rect 19840 347555 19880 347560
rect 19840 347525 19845 347555
rect 19875 347525 19880 347555
rect 19840 347520 19880 347525
rect 19680 347475 19720 347480
rect 19680 347445 19685 347475
rect 19715 347445 19720 347475
rect 19680 347440 19720 347445
rect 19840 347475 19880 347480
rect 19840 347445 19845 347475
rect 19875 347445 19880 347475
rect 19840 347440 19880 347445
rect 19680 347395 19720 347400
rect 19680 347365 19685 347395
rect 19715 347365 19720 347395
rect 19680 347360 19720 347365
rect 19840 347395 19880 347400
rect 19840 347365 19845 347395
rect 19875 347365 19880 347395
rect 19840 347360 19880 347365
rect 19680 347315 19720 347320
rect 19680 347285 19685 347315
rect 19715 347285 19720 347315
rect 19680 347280 19720 347285
rect 19840 347315 19880 347320
rect 19840 347285 19845 347315
rect 19875 347285 19880 347315
rect 19840 347280 19880 347285
rect 19680 347235 19720 347240
rect 19680 347205 19685 347235
rect 19715 347205 19720 347235
rect 19680 347200 19720 347205
rect 19840 347235 19880 347240
rect 19840 347205 19845 347235
rect 19875 347205 19880 347235
rect 19840 347200 19880 347205
rect 19680 347155 19720 347160
rect 19680 347125 19685 347155
rect 19715 347125 19720 347155
rect 19680 347120 19720 347125
rect 19840 347155 19880 347160
rect 19840 347125 19845 347155
rect 19875 347125 19880 347155
rect 19840 347120 19880 347125
rect 19680 347075 19720 347080
rect 19680 347045 19685 347075
rect 19715 347045 19720 347075
rect 19680 347040 19720 347045
rect 19840 347075 19880 347080
rect 19840 347045 19845 347075
rect 19875 347045 19880 347075
rect 19840 347040 19880 347045
rect 19680 346995 19720 347000
rect 19680 346965 19685 346995
rect 19715 346965 19720 346995
rect 19680 346960 19720 346965
rect 19840 346995 19880 347000
rect 19840 346965 19845 346995
rect 19875 346965 19880 346995
rect 19840 346960 19880 346965
rect 19680 346915 19720 346920
rect 19680 346885 19685 346915
rect 19715 346885 19720 346915
rect 19680 346880 19720 346885
rect 19840 346915 19880 346920
rect 19840 346885 19845 346915
rect 19875 346885 19880 346915
rect 19840 346880 19880 346885
rect 19680 346835 19720 346840
rect 19680 346805 19685 346835
rect 19715 346805 19720 346835
rect 19680 346800 19720 346805
rect 19840 346835 19880 346840
rect 19840 346805 19845 346835
rect 19875 346805 19880 346835
rect 19840 346800 19880 346805
rect 19680 346755 19720 346760
rect 19680 346725 19685 346755
rect 19715 346725 19720 346755
rect 19680 346720 19720 346725
rect 19840 346755 19880 346760
rect 19840 346725 19845 346755
rect 19875 346725 19880 346755
rect 19840 346720 19880 346725
rect 19680 346675 19720 346680
rect 19680 346645 19685 346675
rect 19715 346645 19720 346675
rect 19680 346640 19720 346645
rect 19840 346675 19880 346680
rect 19840 346645 19845 346675
rect 19875 346645 19880 346675
rect 19840 346640 19880 346645
rect 19680 346595 19720 346600
rect 19680 346565 19685 346595
rect 19715 346565 19720 346595
rect 19680 346560 19720 346565
rect 19840 346595 19880 346600
rect 19840 346565 19845 346595
rect 19875 346565 19880 346595
rect 19840 346560 19880 346565
rect 19680 346515 19720 346520
rect 19680 346485 19685 346515
rect 19715 346485 19720 346515
rect 19680 346480 19720 346485
rect 19840 346515 19880 346520
rect 19840 346485 19845 346515
rect 19875 346485 19880 346515
rect 19840 346480 19880 346485
rect 19680 346435 19720 346440
rect 19680 346405 19685 346435
rect 19715 346405 19720 346435
rect 19680 346400 19720 346405
rect 19840 346435 19880 346440
rect 19840 346405 19845 346435
rect 19875 346405 19880 346435
rect 19840 346400 19880 346405
rect 19680 346355 19720 346360
rect 19680 346325 19685 346355
rect 19715 346325 19720 346355
rect 19680 346320 19720 346325
rect 19840 346355 19880 346360
rect 19840 346325 19845 346355
rect 19875 346325 19880 346355
rect 19840 346320 19880 346325
rect 19680 346275 19720 346280
rect 19680 346245 19685 346275
rect 19715 346245 19720 346275
rect 19680 346240 19720 346245
rect 19840 346275 19880 346280
rect 19840 346245 19845 346275
rect 19875 346245 19880 346275
rect 19840 346240 19880 346245
rect 19680 346195 19720 346200
rect 19680 346165 19685 346195
rect 19715 346165 19720 346195
rect 19680 346160 19720 346165
rect 19840 346195 19880 346200
rect 19840 346165 19845 346195
rect 19875 346165 19880 346195
rect 19840 346160 19880 346165
rect 19680 346115 19720 346120
rect 19680 346085 19685 346115
rect 19715 346085 19720 346115
rect 19680 346080 19720 346085
rect 19840 346115 19880 346120
rect 19840 346085 19845 346115
rect 19875 346085 19880 346115
rect 19840 346080 19880 346085
rect 19680 346035 19720 346040
rect 19680 346005 19685 346035
rect 19715 346005 19720 346035
rect 19680 346000 19720 346005
rect 19840 346035 19880 346040
rect 19840 346005 19845 346035
rect 19875 346005 19880 346035
rect 19840 346000 19880 346005
rect 19680 345955 19720 345960
rect 19680 345925 19685 345955
rect 19715 345925 19720 345955
rect 19680 345920 19720 345925
rect 19840 345955 19880 345960
rect 19840 345925 19845 345955
rect 19875 345925 19880 345955
rect 19840 345920 19880 345925
rect 19680 345875 19720 345880
rect 19680 345845 19685 345875
rect 19715 345845 19720 345875
rect 19680 345840 19720 345845
rect 19840 345875 19880 345880
rect 19840 345845 19845 345875
rect 19875 345845 19880 345875
rect 19840 345840 19880 345845
rect 19680 345795 19720 345800
rect 19680 345765 19685 345795
rect 19715 345765 19720 345795
rect 19680 345760 19720 345765
rect 19840 345795 19880 345800
rect 19840 345765 19845 345795
rect 19875 345765 19880 345795
rect 19840 345760 19880 345765
rect 19680 345715 19720 345720
rect 19680 345685 19685 345715
rect 19715 345685 19720 345715
rect 19680 345680 19720 345685
rect 19840 345715 19880 345720
rect 19840 345685 19845 345715
rect 19875 345685 19880 345715
rect 19840 345680 19880 345685
rect 19680 345635 19720 345640
rect 19680 345605 19685 345635
rect 19715 345605 19720 345635
rect 19680 345600 19720 345605
rect 19840 345635 19880 345640
rect 19840 345605 19845 345635
rect 19875 345605 19880 345635
rect 19840 345600 19880 345605
rect 19680 345555 19720 345560
rect 19680 345525 19685 345555
rect 19715 345525 19720 345555
rect 19680 345520 19720 345525
rect 19840 345555 19880 345560
rect 19840 345525 19845 345555
rect 19875 345525 19880 345555
rect 19840 345520 19880 345525
rect 19680 345475 19720 345480
rect 19680 345445 19685 345475
rect 19715 345445 19720 345475
rect 19680 345440 19720 345445
rect 19840 345475 19880 345480
rect 19840 345445 19845 345475
rect 19875 345445 19880 345475
rect 19840 345440 19880 345445
rect 19680 345395 19720 345400
rect 19680 345365 19685 345395
rect 19715 345365 19720 345395
rect 19680 345360 19720 345365
rect 19840 345395 19880 345400
rect 19840 345365 19845 345395
rect 19875 345365 19880 345395
rect 19840 345360 19880 345365
rect 19680 345315 19720 345320
rect 19680 345285 19685 345315
rect 19715 345285 19720 345315
rect 19680 345280 19720 345285
rect 19840 345315 19880 345320
rect 19840 345285 19845 345315
rect 19875 345285 19880 345315
rect 19840 345280 19880 345285
rect 19680 345235 19720 345240
rect 19680 345205 19685 345235
rect 19715 345205 19720 345235
rect 19680 345200 19720 345205
rect 19840 345235 19880 345240
rect 19840 345205 19845 345235
rect 19875 345205 19880 345235
rect 19840 345200 19880 345205
rect 19680 345155 19720 345160
rect 19680 345125 19685 345155
rect 19715 345125 19720 345155
rect 19680 345120 19720 345125
rect 19840 345155 19880 345160
rect 19840 345125 19845 345155
rect 19875 345125 19880 345155
rect 19840 345120 19880 345125
rect 19680 345075 19720 345080
rect 19680 345045 19685 345075
rect 19715 345045 19720 345075
rect 19680 345040 19720 345045
rect 19840 345075 19880 345080
rect 19840 345045 19845 345075
rect 19875 345045 19880 345075
rect 19840 345040 19880 345045
rect 19680 344995 19720 345000
rect 19680 344965 19685 344995
rect 19715 344965 19720 344995
rect 19680 344960 19720 344965
rect 19840 344995 19880 345000
rect 19840 344965 19845 344995
rect 19875 344965 19880 344995
rect 19840 344960 19880 344965
rect 19680 344915 19720 344920
rect 19680 344885 19685 344915
rect 19715 344885 19720 344915
rect 19680 344880 19720 344885
rect 19840 344915 19880 344920
rect 19840 344885 19845 344915
rect 19875 344885 19880 344915
rect 19840 344880 19880 344885
rect 19680 344835 19720 344840
rect 19680 344805 19685 344835
rect 19715 344805 19720 344835
rect 19680 344800 19720 344805
rect 19840 344835 19880 344840
rect 19840 344805 19845 344835
rect 19875 344805 19880 344835
rect 19840 344800 19880 344805
rect 19680 344755 19720 344760
rect 19680 344725 19685 344755
rect 19715 344725 19720 344755
rect 19680 344720 19720 344725
rect 19840 344755 19880 344760
rect 19840 344725 19845 344755
rect 19875 344725 19880 344755
rect 19840 344720 19880 344725
rect 19680 344675 19720 344680
rect 19680 344645 19685 344675
rect 19715 344645 19720 344675
rect 19680 344640 19720 344645
rect 19840 344675 19880 344680
rect 19840 344645 19845 344675
rect 19875 344645 19880 344675
rect 19840 344640 19880 344645
rect 19680 344595 19720 344600
rect 19680 344565 19685 344595
rect 19715 344565 19720 344595
rect 19680 344560 19720 344565
rect 19840 344595 19880 344600
rect 19840 344565 19845 344595
rect 19875 344565 19880 344595
rect 19840 344560 19880 344565
rect 19680 344515 19720 344520
rect 19680 344485 19685 344515
rect 19715 344485 19720 344515
rect 19680 344480 19720 344485
rect 19840 344515 19880 344520
rect 19840 344485 19845 344515
rect 19875 344485 19880 344515
rect 19840 344480 19880 344485
rect 19680 344435 19720 344440
rect 19680 344405 19685 344435
rect 19715 344405 19720 344435
rect 19680 344400 19720 344405
rect 19840 344435 19880 344440
rect 19840 344405 19845 344435
rect 19875 344405 19880 344435
rect 19840 344400 19880 344405
rect 19680 344355 19720 344360
rect 19680 344325 19685 344355
rect 19715 344325 19720 344355
rect 19680 344320 19720 344325
rect 19840 344355 19880 344360
rect 19840 344325 19845 344355
rect 19875 344325 19880 344355
rect 19840 344320 19880 344325
rect 19680 344275 19720 344280
rect 19680 344245 19685 344275
rect 19715 344245 19720 344275
rect 19680 344240 19720 344245
rect 19840 344275 19880 344280
rect 19840 344245 19845 344275
rect 19875 344245 19880 344275
rect 19840 344240 19880 344245
rect 19680 344195 19720 344200
rect 19680 344165 19685 344195
rect 19715 344165 19720 344195
rect 19680 344160 19720 344165
rect 19840 344195 19880 344200
rect 19840 344165 19845 344195
rect 19875 344165 19880 344195
rect 19840 344160 19880 344165
rect 19680 344115 19720 344120
rect 19680 344085 19685 344115
rect 19715 344085 19720 344115
rect 19680 344080 19720 344085
rect 19840 344115 19880 344120
rect 19840 344085 19845 344115
rect 19875 344085 19880 344115
rect 19840 344080 19880 344085
rect 19680 344035 19720 344040
rect 19680 344005 19685 344035
rect 19715 344005 19720 344035
rect 19680 344000 19720 344005
rect 19840 344035 19880 344040
rect 19840 344005 19845 344035
rect 19875 344005 19880 344035
rect 19840 344000 19880 344005
rect 19680 343955 19720 343960
rect 19680 343925 19685 343955
rect 19715 343925 19720 343955
rect 19680 343920 19720 343925
rect 19840 343955 19880 343960
rect 19840 343925 19845 343955
rect 19875 343925 19880 343955
rect 19840 343920 19880 343925
rect 19680 343875 19720 343880
rect 19680 343845 19685 343875
rect 19715 343845 19720 343875
rect 19680 343840 19720 343845
rect 19840 343875 19880 343880
rect 19840 343845 19845 343875
rect 19875 343845 19880 343875
rect 19840 343840 19880 343845
rect 19680 343795 19720 343800
rect 19680 343765 19685 343795
rect 19715 343765 19720 343795
rect 19680 343760 19720 343765
rect 19840 343795 19880 343800
rect 19840 343765 19845 343795
rect 19875 343765 19880 343795
rect 19840 343760 19880 343765
rect 19680 343715 19720 343720
rect 19680 343685 19685 343715
rect 19715 343685 19720 343715
rect 19680 343680 19720 343685
rect 19840 343715 19880 343720
rect 19840 343685 19845 343715
rect 19875 343685 19880 343715
rect 19840 343680 19880 343685
rect 19680 343635 19720 343640
rect 19680 343605 19685 343635
rect 19715 343605 19720 343635
rect 19680 343600 19720 343605
rect 19840 343635 19880 343640
rect 19840 343605 19845 343635
rect 19875 343605 19880 343635
rect 19840 343600 19880 343605
rect 19680 343555 19720 343560
rect 19680 343525 19685 343555
rect 19715 343525 19720 343555
rect 19680 343520 19720 343525
rect 19840 343555 19880 343560
rect 19840 343525 19845 343555
rect 19875 343525 19880 343555
rect 19840 343520 19880 343525
rect 19680 343475 19720 343480
rect 19680 343445 19685 343475
rect 19715 343445 19720 343475
rect 19680 343440 19720 343445
rect 19840 343475 19880 343480
rect 19840 343445 19845 343475
rect 19875 343445 19880 343475
rect 19840 343440 19880 343445
rect 19680 343395 19720 343400
rect 19680 343365 19685 343395
rect 19715 343365 19720 343395
rect 19680 343360 19720 343365
rect 19840 343395 19880 343400
rect 19840 343365 19845 343395
rect 19875 343365 19880 343395
rect 19840 343360 19880 343365
rect 19680 343315 19720 343320
rect 19680 343285 19685 343315
rect 19715 343285 19720 343315
rect 19680 343280 19720 343285
rect 19840 343315 19880 343320
rect 19840 343285 19845 343315
rect 19875 343285 19880 343315
rect 19840 343280 19880 343285
rect 19680 343235 19720 343240
rect 19680 343205 19685 343235
rect 19715 343205 19720 343235
rect 19680 343200 19720 343205
rect 19840 343235 19880 343240
rect 19840 343205 19845 343235
rect 19875 343205 19880 343235
rect 19840 343200 19880 343205
rect 19680 343155 19720 343160
rect 19680 343125 19685 343155
rect 19715 343125 19720 343155
rect 19680 343120 19720 343125
rect 19840 343155 19880 343160
rect 19840 343125 19845 343155
rect 19875 343125 19880 343155
rect 19840 343120 19880 343125
rect 19680 343075 19720 343080
rect 19680 343045 19685 343075
rect 19715 343045 19720 343075
rect 19680 343040 19720 343045
rect 19840 343075 19880 343080
rect 19840 343045 19845 343075
rect 19875 343045 19880 343075
rect 19840 343040 19880 343045
rect 19680 342995 19720 343000
rect 19680 342965 19685 342995
rect 19715 342965 19720 342995
rect 19680 342960 19720 342965
rect 19840 342995 19880 343000
rect 19840 342965 19845 342995
rect 19875 342965 19880 342995
rect 19840 342960 19880 342965
rect 19680 342915 19720 342920
rect 19680 342885 19685 342915
rect 19715 342885 19720 342915
rect 19680 342880 19720 342885
rect 19840 342915 19880 342920
rect 19840 342885 19845 342915
rect 19875 342885 19880 342915
rect 19840 342880 19880 342885
rect 19680 342835 19720 342840
rect 19680 342805 19685 342835
rect 19715 342805 19720 342835
rect 19680 342800 19720 342805
rect 19840 342835 19880 342840
rect 19840 342805 19845 342835
rect 19875 342805 19880 342835
rect 19840 342800 19880 342805
rect 19680 342755 19720 342760
rect 19680 342725 19685 342755
rect 19715 342725 19720 342755
rect 19680 342720 19720 342725
rect 19840 342755 19880 342760
rect 19840 342725 19845 342755
rect 19875 342725 19880 342755
rect 19840 342720 19880 342725
rect 19680 342675 19720 342680
rect 19680 342645 19685 342675
rect 19715 342645 19720 342675
rect 19680 342640 19720 342645
rect 19840 342675 19880 342680
rect 19840 342645 19845 342675
rect 19875 342645 19880 342675
rect 19840 342640 19880 342645
rect 19680 342595 19720 342600
rect 19680 342565 19685 342595
rect 19715 342565 19720 342595
rect 19680 342560 19720 342565
rect 19840 342595 19880 342600
rect 19840 342565 19845 342595
rect 19875 342565 19880 342595
rect 19840 342560 19880 342565
rect 19680 342515 19720 342520
rect 19680 342485 19685 342515
rect 19715 342485 19720 342515
rect 19680 342480 19720 342485
rect 19840 342515 19880 342520
rect 19840 342485 19845 342515
rect 19875 342485 19880 342515
rect 19840 342480 19880 342485
rect 19680 342435 19720 342440
rect 19680 342405 19685 342435
rect 19715 342405 19720 342435
rect 19680 342400 19720 342405
rect 19840 342435 19880 342440
rect 19840 342405 19845 342435
rect 19875 342405 19880 342435
rect 19840 342400 19880 342405
rect 19680 342355 19720 342360
rect 19680 342325 19685 342355
rect 19715 342325 19720 342355
rect 19680 342320 19720 342325
rect 19840 342355 19880 342360
rect 19840 342325 19845 342355
rect 19875 342325 19880 342355
rect 19840 342320 19880 342325
rect 19680 342275 19720 342280
rect 19680 342245 19685 342275
rect 19715 342245 19720 342275
rect 19680 342240 19720 342245
rect 19840 342275 19880 342280
rect 19840 342245 19845 342275
rect 19875 342245 19880 342275
rect 19840 342240 19880 342245
rect 19680 342195 19720 342200
rect 19680 342165 19685 342195
rect 19715 342165 19720 342195
rect 19680 342160 19720 342165
rect 19840 342195 19880 342200
rect 19840 342165 19845 342195
rect 19875 342165 19880 342195
rect 19840 342160 19880 342165
rect 19680 342115 19720 342120
rect 19680 342085 19685 342115
rect 19715 342085 19720 342115
rect 19680 342080 19720 342085
rect 19840 342115 19880 342120
rect 19840 342085 19845 342115
rect 19875 342085 19880 342115
rect 19840 342080 19880 342085
rect 19680 342035 19720 342040
rect 19680 342005 19685 342035
rect 19715 342005 19720 342035
rect 19680 342000 19720 342005
rect 19840 342035 19880 342040
rect 19840 342005 19845 342035
rect 19875 342005 19880 342035
rect 19840 342000 19880 342005
rect 19680 341955 19720 341960
rect 19680 341925 19685 341955
rect 19715 341925 19720 341955
rect 19680 341920 19720 341925
rect 19840 341955 19880 341960
rect 19840 341925 19845 341955
rect 19875 341925 19880 341955
rect 19840 341920 19880 341925
rect 19680 341875 19720 341880
rect 19680 341845 19685 341875
rect 19715 341845 19720 341875
rect 19680 341840 19720 341845
rect 19840 341875 19880 341880
rect 19840 341845 19845 341875
rect 19875 341845 19880 341875
rect 19840 341840 19880 341845
rect 19680 341795 19720 341800
rect 19680 341765 19685 341795
rect 19715 341765 19720 341795
rect 19680 341760 19720 341765
rect 19840 341795 19880 341800
rect 19840 341765 19845 341795
rect 19875 341765 19880 341795
rect 19840 341760 19880 341765
rect 19680 341715 19720 341720
rect 19680 341685 19685 341715
rect 19715 341685 19720 341715
rect 19680 341680 19720 341685
rect 19840 341715 19880 341720
rect 19840 341685 19845 341715
rect 19875 341685 19880 341715
rect 19840 341680 19880 341685
rect 19680 341635 19720 341640
rect 19680 341605 19685 341635
rect 19715 341605 19720 341635
rect 19680 341600 19720 341605
rect 19840 341635 19880 341640
rect 19840 341605 19845 341635
rect 19875 341605 19880 341635
rect 19840 341600 19880 341605
rect 19680 341555 19720 341560
rect 19680 341525 19685 341555
rect 19715 341525 19720 341555
rect 19680 341520 19720 341525
rect 19840 341555 19880 341560
rect 19840 341525 19845 341555
rect 19875 341525 19880 341555
rect 19840 341520 19880 341525
rect 19680 341475 19720 341480
rect 19680 341445 19685 341475
rect 19715 341445 19720 341475
rect 19680 341440 19720 341445
rect 19840 341475 19880 341480
rect 19840 341445 19845 341475
rect 19875 341445 19880 341475
rect 19840 341440 19880 341445
rect 19680 341395 19720 341400
rect 19680 341365 19685 341395
rect 19715 341365 19720 341395
rect 19680 341360 19720 341365
rect 19840 341395 19880 341400
rect 19840 341365 19845 341395
rect 19875 341365 19880 341395
rect 19840 341360 19880 341365
rect 19680 341315 19720 341320
rect 19680 341285 19685 341315
rect 19715 341285 19720 341315
rect 19680 341280 19720 341285
rect 19840 341315 19880 341320
rect 19840 341285 19845 341315
rect 19875 341285 19880 341315
rect 19840 341280 19880 341285
rect 19680 341235 19720 341240
rect 19680 341205 19685 341235
rect 19715 341205 19720 341235
rect 19680 341200 19720 341205
rect 19840 341235 19880 341240
rect 19840 341205 19845 341235
rect 19875 341205 19880 341235
rect 19840 341200 19880 341205
rect 19680 341155 19720 341160
rect 19680 341125 19685 341155
rect 19715 341125 19720 341155
rect 19680 341120 19720 341125
rect 19840 341155 19880 341160
rect 19840 341125 19845 341155
rect 19875 341125 19880 341155
rect 19840 341120 19880 341125
rect 19680 341075 19720 341080
rect 19680 341045 19685 341075
rect 19715 341045 19720 341075
rect 19680 341040 19720 341045
rect 19840 341075 19880 341080
rect 19840 341045 19845 341075
rect 19875 341045 19880 341075
rect 19840 341040 19880 341045
rect 19680 340995 19720 341000
rect 19680 340965 19685 340995
rect 19715 340965 19720 340995
rect 19680 340960 19720 340965
rect 19840 340995 19880 341000
rect 19840 340965 19845 340995
rect 19875 340965 19880 340995
rect 19840 340960 19880 340965
rect 19680 340915 19720 340920
rect 19680 340885 19685 340915
rect 19715 340885 19720 340915
rect 19680 340880 19720 340885
rect 19840 340915 19880 340920
rect 19840 340885 19845 340915
rect 19875 340885 19880 340915
rect 19840 340880 19880 340885
rect 19680 340835 19720 340840
rect 19680 340805 19685 340835
rect 19715 340805 19720 340835
rect 19680 340800 19720 340805
rect 19840 340835 19880 340840
rect 19840 340805 19845 340835
rect 19875 340805 19880 340835
rect 19840 340800 19880 340805
rect 19680 340755 19720 340760
rect 19680 340725 19685 340755
rect 19715 340725 19720 340755
rect 19680 340720 19720 340725
rect 19840 340755 19880 340760
rect 19840 340725 19845 340755
rect 19875 340725 19880 340755
rect 19840 340720 19880 340725
rect 19680 340675 19720 340680
rect 19680 340645 19685 340675
rect 19715 340645 19720 340675
rect 19680 340640 19720 340645
rect 19840 340675 19880 340680
rect 19840 340645 19845 340675
rect 19875 340645 19880 340675
rect 19840 340640 19880 340645
rect 19680 340595 19720 340600
rect 19680 340565 19685 340595
rect 19715 340565 19720 340595
rect 19680 340560 19720 340565
rect 19840 340595 19880 340600
rect 19840 340565 19845 340595
rect 19875 340565 19880 340595
rect 19840 340560 19880 340565
rect 19680 340515 19720 340520
rect 19680 340485 19685 340515
rect 19715 340485 19720 340515
rect 19680 340480 19720 340485
rect 19840 340515 19880 340520
rect 19840 340485 19845 340515
rect 19875 340485 19880 340515
rect 19840 340480 19880 340485
rect 19680 340435 19720 340440
rect 19680 340405 19685 340435
rect 19715 340405 19720 340435
rect 19680 340400 19720 340405
rect 19840 340435 19880 340440
rect 19840 340405 19845 340435
rect 19875 340405 19880 340435
rect 19840 340400 19880 340405
rect 19680 340355 19720 340360
rect 19680 340325 19685 340355
rect 19715 340325 19720 340355
rect 19680 340320 19720 340325
rect 19840 340355 19880 340360
rect 19840 340325 19845 340355
rect 19875 340325 19880 340355
rect 19840 340320 19880 340325
rect 19680 340275 19720 340280
rect 19680 340245 19685 340275
rect 19715 340245 19720 340275
rect 19680 340240 19720 340245
rect 19840 340275 19880 340280
rect 19840 340245 19845 340275
rect 19875 340245 19880 340275
rect 19840 340240 19880 340245
rect 19680 340195 19720 340200
rect 19680 340165 19685 340195
rect 19715 340165 19720 340195
rect 19680 340160 19720 340165
rect 19840 340195 19880 340200
rect 19840 340165 19845 340195
rect 19875 340165 19880 340195
rect 19840 340160 19880 340165
rect 19680 340115 19720 340120
rect 19680 340085 19685 340115
rect 19715 340085 19720 340115
rect 19680 340080 19720 340085
rect 19840 340115 19880 340120
rect 19840 340085 19845 340115
rect 19875 340085 19880 340115
rect 19840 340080 19880 340085
rect 19680 340035 19720 340040
rect 19680 340005 19685 340035
rect 19715 340005 19720 340035
rect 19680 340000 19720 340005
rect 19840 340035 19880 340040
rect 19840 340005 19845 340035
rect 19875 340005 19880 340035
rect 19840 340000 19880 340005
rect 19680 339955 19720 339960
rect 19680 339925 19685 339955
rect 19715 339925 19720 339955
rect 19680 339920 19720 339925
rect 19840 339955 19880 339960
rect 19840 339925 19845 339955
rect 19875 339925 19880 339955
rect 19840 339920 19880 339925
rect 19680 339875 19720 339880
rect 19680 339845 19685 339875
rect 19715 339845 19720 339875
rect 19680 339840 19720 339845
rect 19840 339875 19880 339880
rect 19840 339845 19845 339875
rect 19875 339845 19880 339875
rect 19840 339840 19880 339845
rect 19680 339795 19720 339800
rect 19680 339765 19685 339795
rect 19715 339765 19720 339795
rect 19680 339760 19720 339765
rect 19840 339795 19880 339800
rect 19840 339765 19845 339795
rect 19875 339765 19880 339795
rect 19840 339760 19880 339765
rect 19680 339715 19720 339720
rect 19680 339685 19685 339715
rect 19715 339685 19720 339715
rect 19680 339680 19720 339685
rect 19840 339715 19880 339720
rect 19840 339685 19845 339715
rect 19875 339685 19880 339715
rect 19840 339680 19880 339685
rect 19680 339635 19720 339640
rect 19680 339605 19685 339635
rect 19715 339605 19720 339635
rect 19680 339600 19720 339605
rect 19840 339635 19880 339640
rect 19840 339605 19845 339635
rect 19875 339605 19880 339635
rect 19840 339600 19880 339605
rect 19680 339555 19720 339560
rect 19680 339525 19685 339555
rect 19715 339525 19720 339555
rect 19680 339520 19720 339525
rect 19840 339555 19880 339560
rect 19840 339525 19845 339555
rect 19875 339525 19880 339555
rect 19840 339520 19880 339525
rect 19680 339475 19720 339480
rect 19680 339445 19685 339475
rect 19715 339445 19720 339475
rect 19680 339440 19720 339445
rect 19840 339475 19880 339480
rect 19840 339445 19845 339475
rect 19875 339445 19880 339475
rect 19840 339440 19880 339445
rect 19680 339395 19720 339400
rect 19680 339365 19685 339395
rect 19715 339365 19720 339395
rect 19680 339360 19720 339365
rect 19840 339395 19880 339400
rect 19840 339365 19845 339395
rect 19875 339365 19880 339395
rect 19840 339360 19880 339365
rect 19680 339315 19720 339320
rect 19680 339285 19685 339315
rect 19715 339285 19720 339315
rect 19680 339280 19720 339285
rect 19840 339315 19880 339320
rect 19840 339285 19845 339315
rect 19875 339285 19880 339315
rect 19840 339280 19880 339285
rect 19680 339235 19720 339240
rect 19680 339205 19685 339235
rect 19715 339205 19720 339235
rect 19680 339200 19720 339205
rect 19840 339235 19880 339240
rect 19840 339205 19845 339235
rect 19875 339205 19880 339235
rect 19840 339200 19880 339205
rect 19680 339155 19720 339160
rect 19680 339125 19685 339155
rect 19715 339125 19720 339155
rect 19680 339120 19720 339125
rect 19840 339155 19880 339160
rect 19840 339125 19845 339155
rect 19875 339125 19880 339155
rect 19840 339120 19880 339125
rect 19680 339075 19720 339080
rect 19680 339045 19685 339075
rect 19715 339045 19720 339075
rect 19680 339040 19720 339045
rect 19840 339075 19880 339080
rect 19840 339045 19845 339075
rect 19875 339045 19880 339075
rect 19840 339040 19880 339045
rect 19680 338995 19720 339000
rect 19680 338965 19685 338995
rect 19715 338965 19720 338995
rect 19680 338960 19720 338965
rect 19840 338995 19880 339000
rect 19840 338965 19845 338995
rect 19875 338965 19880 338995
rect 19840 338960 19880 338965
rect 19680 338915 19720 338920
rect 19680 338885 19685 338915
rect 19715 338885 19720 338915
rect 19680 338880 19720 338885
rect 19840 338915 19880 338920
rect 19840 338885 19845 338915
rect 19875 338885 19880 338915
rect 19840 338880 19880 338885
rect 19680 338835 19720 338840
rect 19680 338805 19685 338835
rect 19715 338805 19720 338835
rect 19680 338800 19720 338805
rect 19840 338835 19880 338840
rect 19840 338805 19845 338835
rect 19875 338805 19880 338835
rect 19840 338800 19880 338805
rect 19680 338755 19720 338760
rect 19680 338725 19685 338755
rect 19715 338725 19720 338755
rect 19680 338720 19720 338725
rect 19840 338755 19880 338760
rect 19840 338725 19845 338755
rect 19875 338725 19880 338755
rect 19840 338720 19880 338725
rect 19680 338675 19720 338680
rect 19680 338645 19685 338675
rect 19715 338645 19720 338675
rect 19680 338640 19720 338645
rect 19840 338675 19880 338680
rect 19840 338645 19845 338675
rect 19875 338645 19880 338675
rect 19840 338640 19880 338645
rect 19680 338595 19720 338600
rect 19680 338565 19685 338595
rect 19715 338565 19720 338595
rect 19680 338560 19720 338565
rect 19840 338595 19880 338600
rect 19840 338565 19845 338595
rect 19875 338565 19880 338595
rect 19840 338560 19880 338565
rect 19680 338515 19720 338520
rect 19680 338485 19685 338515
rect 19715 338485 19720 338515
rect 19680 338480 19720 338485
rect 19840 338515 19880 338520
rect 19840 338485 19845 338515
rect 19875 338485 19880 338515
rect 19840 338480 19880 338485
rect 19680 338435 19720 338440
rect 19680 338405 19685 338435
rect 19715 338405 19720 338435
rect 19680 338400 19720 338405
rect 19840 338435 19880 338440
rect 19840 338405 19845 338435
rect 19875 338405 19880 338435
rect 19840 338400 19880 338405
rect 19680 338355 19720 338360
rect 19680 338325 19685 338355
rect 19715 338325 19720 338355
rect 19680 338320 19720 338325
rect 19840 338355 19880 338360
rect 19840 338325 19845 338355
rect 19875 338325 19880 338355
rect 19840 338320 19880 338325
rect 19680 338275 19720 338280
rect 19680 338245 19685 338275
rect 19715 338245 19720 338275
rect 19680 338240 19720 338245
rect 19840 338275 19880 338280
rect 19840 338245 19845 338275
rect 19875 338245 19880 338275
rect 19840 338240 19880 338245
rect 19680 338195 19720 338200
rect 19680 338165 19685 338195
rect 19715 338165 19720 338195
rect 19680 338160 19720 338165
rect 19840 338195 19880 338200
rect 19840 338165 19845 338195
rect 19875 338165 19880 338195
rect 19840 338160 19880 338165
rect 19680 338115 19720 338120
rect 19680 338085 19685 338115
rect 19715 338085 19720 338115
rect 19680 338080 19720 338085
rect 19840 338115 19880 338120
rect 19840 338085 19845 338115
rect 19875 338085 19880 338115
rect 19840 338080 19880 338085
rect 19680 338035 19720 338040
rect 19680 338005 19685 338035
rect 19715 338005 19720 338035
rect 19680 338000 19720 338005
rect 19840 338035 19880 338040
rect 19840 338005 19845 338035
rect 19875 338005 19880 338035
rect 19840 338000 19880 338005
rect 19680 337955 19720 337960
rect 19680 337925 19685 337955
rect 19715 337925 19720 337955
rect 19680 337920 19720 337925
rect 19840 337955 19880 337960
rect 19840 337925 19845 337955
rect 19875 337925 19880 337955
rect 19840 337920 19880 337925
rect 19680 337875 19720 337880
rect 19680 337845 19685 337875
rect 19715 337845 19720 337875
rect 19680 337840 19720 337845
rect 19840 337875 19880 337880
rect 19840 337845 19845 337875
rect 19875 337845 19880 337875
rect 19840 337840 19880 337845
rect 19680 337795 19720 337800
rect 19680 337765 19685 337795
rect 19715 337765 19720 337795
rect 19680 337760 19720 337765
rect 19840 337795 19880 337800
rect 19840 337765 19845 337795
rect 19875 337765 19880 337795
rect 19840 337760 19880 337765
rect 19680 337715 19720 337720
rect 19680 337685 19685 337715
rect 19715 337685 19720 337715
rect 19680 337680 19720 337685
rect 19840 337715 19880 337720
rect 19840 337685 19845 337715
rect 19875 337685 19880 337715
rect 19840 337680 19880 337685
rect 19680 337635 19720 337640
rect 19680 337605 19685 337635
rect 19715 337605 19720 337635
rect 19680 337600 19720 337605
rect 19840 337635 19880 337640
rect 19840 337605 19845 337635
rect 19875 337605 19880 337635
rect 19840 337600 19880 337605
rect 19680 337555 19720 337560
rect 19680 337525 19685 337555
rect 19715 337525 19720 337555
rect 19680 337520 19720 337525
rect 19840 337555 19880 337560
rect 19840 337525 19845 337555
rect 19875 337525 19880 337555
rect 19840 337520 19880 337525
rect 19680 337475 19720 337480
rect 19680 337445 19685 337475
rect 19715 337445 19720 337475
rect 19680 337440 19720 337445
rect 19840 337475 19880 337480
rect 19840 337445 19845 337475
rect 19875 337445 19880 337475
rect 19840 337440 19880 337445
rect 19680 337395 19720 337400
rect 19680 337365 19685 337395
rect 19715 337365 19720 337395
rect 19680 337360 19720 337365
rect 19840 337395 19880 337400
rect 19840 337365 19845 337395
rect 19875 337365 19880 337395
rect 19840 337360 19880 337365
rect 19680 337315 19720 337320
rect 19680 337285 19685 337315
rect 19715 337285 19720 337315
rect 19680 337280 19720 337285
rect 19840 337315 19880 337320
rect 19840 337285 19845 337315
rect 19875 337285 19880 337315
rect 19840 337280 19880 337285
rect 19680 337235 19720 337240
rect 19680 337205 19685 337235
rect 19715 337205 19720 337235
rect 19680 337200 19720 337205
rect 19840 337235 19880 337240
rect 19840 337205 19845 337235
rect 19875 337205 19880 337235
rect 19840 337200 19880 337205
rect 19680 337155 19720 337160
rect 19680 337125 19685 337155
rect 19715 337125 19720 337155
rect 19680 337120 19720 337125
rect 19840 337155 19880 337160
rect 19840 337125 19845 337155
rect 19875 337125 19880 337155
rect 19840 337120 19880 337125
rect 19680 337075 19720 337080
rect 19680 337045 19685 337075
rect 19715 337045 19720 337075
rect 19680 337040 19720 337045
rect 19840 337075 19880 337080
rect 19840 337045 19845 337075
rect 19875 337045 19880 337075
rect 19840 337040 19880 337045
rect 19680 336995 19720 337000
rect 19680 336965 19685 336995
rect 19715 336965 19720 336995
rect 19680 336960 19720 336965
rect 19840 336995 19880 337000
rect 19840 336965 19845 336995
rect 19875 336965 19880 336995
rect 19840 336960 19880 336965
rect 19680 336915 19720 336920
rect 19680 336885 19685 336915
rect 19715 336885 19720 336915
rect 19680 336880 19720 336885
rect 19840 336915 19880 336920
rect 19840 336885 19845 336915
rect 19875 336885 19880 336915
rect 19840 336880 19880 336885
rect 19680 336835 19720 336840
rect 19680 336805 19685 336835
rect 19715 336805 19720 336835
rect 19680 336800 19720 336805
rect 19840 336835 19880 336840
rect 19840 336805 19845 336835
rect 19875 336805 19880 336835
rect 19840 336800 19880 336805
rect 19680 336755 19720 336760
rect 19680 336725 19685 336755
rect 19715 336725 19720 336755
rect 19680 336720 19720 336725
rect 19840 336755 19880 336760
rect 19840 336725 19845 336755
rect 19875 336725 19880 336755
rect 19840 336720 19880 336725
rect 19680 336675 19720 336680
rect 19680 336645 19685 336675
rect 19715 336645 19720 336675
rect 19680 336640 19720 336645
rect 19840 336675 19880 336680
rect 19840 336645 19845 336675
rect 19875 336645 19880 336675
rect 19840 336640 19880 336645
rect 19680 336595 19720 336600
rect 19680 336565 19685 336595
rect 19715 336565 19720 336595
rect 19680 336560 19720 336565
rect 19840 336595 19880 336600
rect 19840 336565 19845 336595
rect 19875 336565 19880 336595
rect 19840 336560 19880 336565
rect 19680 336515 19720 336520
rect 19680 336485 19685 336515
rect 19715 336485 19720 336515
rect 19680 336480 19720 336485
rect 19840 336515 19880 336520
rect 19840 336485 19845 336515
rect 19875 336485 19880 336515
rect 19840 336480 19880 336485
rect 19680 336435 19720 336440
rect 19680 336405 19685 336435
rect 19715 336405 19720 336435
rect 19680 336400 19720 336405
rect 19840 336435 19880 336440
rect 19840 336405 19845 336435
rect 19875 336405 19880 336435
rect 19840 336400 19880 336405
rect 19680 336355 19720 336360
rect 19680 336325 19685 336355
rect 19715 336325 19720 336355
rect 19680 336320 19720 336325
rect 19840 336355 19880 336360
rect 19840 336325 19845 336355
rect 19875 336325 19880 336355
rect 19840 336320 19880 336325
rect 19680 336275 19720 336280
rect 19680 336245 19685 336275
rect 19715 336245 19720 336275
rect 19680 336240 19720 336245
rect 19840 336275 19880 336280
rect 19840 336245 19845 336275
rect 19875 336245 19880 336275
rect 19840 336240 19880 336245
rect 19680 336195 19720 336200
rect 19680 336165 19685 336195
rect 19715 336165 19720 336195
rect 19680 336160 19720 336165
rect 19840 336195 19880 336200
rect 19840 336165 19845 336195
rect 19875 336165 19880 336195
rect 19840 336160 19880 336165
rect 19680 336115 19720 336120
rect 19680 336085 19685 336115
rect 19715 336085 19720 336115
rect 19680 336080 19720 336085
rect 19840 336115 19880 336120
rect 19840 336085 19845 336115
rect 19875 336085 19880 336115
rect 19840 336080 19880 336085
rect 19680 336035 19720 336040
rect 19680 336005 19685 336035
rect 19715 336005 19720 336035
rect 19680 336000 19720 336005
rect 19840 336035 19880 336040
rect 19840 336005 19845 336035
rect 19875 336005 19880 336035
rect 19840 336000 19880 336005
rect 19680 335955 19720 335960
rect 19680 335925 19685 335955
rect 19715 335925 19720 335955
rect 19680 335920 19720 335925
rect 19840 335955 19880 335960
rect 19840 335925 19845 335955
rect 19875 335925 19880 335955
rect 19840 335920 19880 335925
rect 19680 335875 19720 335880
rect 19680 335845 19685 335875
rect 19715 335845 19720 335875
rect 19680 335840 19720 335845
rect 19840 335875 19880 335880
rect 19840 335845 19845 335875
rect 19875 335845 19880 335875
rect 19840 335840 19880 335845
rect 19680 335795 19720 335800
rect 19680 335765 19685 335795
rect 19715 335765 19720 335795
rect 19680 335760 19720 335765
rect 19840 335795 19880 335800
rect 19840 335765 19845 335795
rect 19875 335765 19880 335795
rect 19840 335760 19880 335765
rect 19680 335715 19720 335720
rect 19680 335685 19685 335715
rect 19715 335685 19720 335715
rect 19680 335680 19720 335685
rect 19840 335715 19880 335720
rect 19840 335685 19845 335715
rect 19875 335685 19880 335715
rect 19840 335680 19880 335685
rect 19680 335635 19720 335640
rect 19680 335605 19685 335635
rect 19715 335605 19720 335635
rect 19680 335600 19720 335605
rect 19840 335635 19880 335640
rect 19840 335605 19845 335635
rect 19875 335605 19880 335635
rect 19840 335600 19880 335605
rect 19680 335555 19720 335560
rect 19680 335525 19685 335555
rect 19715 335525 19720 335555
rect 19680 335520 19720 335525
rect 19840 335555 19880 335560
rect 19840 335525 19845 335555
rect 19875 335525 19880 335555
rect 19840 335520 19880 335525
rect 19680 335475 19720 335480
rect 19680 335445 19685 335475
rect 19715 335445 19720 335475
rect 19680 335440 19720 335445
rect 19840 335475 19880 335480
rect 19840 335445 19845 335475
rect 19875 335445 19880 335475
rect 19840 335440 19880 335445
rect 19680 335395 19720 335400
rect 19680 335365 19685 335395
rect 19715 335365 19720 335395
rect 19680 335360 19720 335365
rect 19840 335395 19880 335400
rect 19840 335365 19845 335395
rect 19875 335365 19880 335395
rect 19840 335360 19880 335365
rect 19680 335315 19720 335320
rect 19680 335285 19685 335315
rect 19715 335285 19720 335315
rect 19680 335280 19720 335285
rect 19840 335315 19880 335320
rect 19840 335285 19845 335315
rect 19875 335285 19880 335315
rect 19840 335280 19880 335285
rect 19680 335235 19720 335240
rect 19680 335205 19685 335235
rect 19715 335205 19720 335235
rect 19680 335200 19720 335205
rect 19840 335235 19880 335240
rect 19840 335205 19845 335235
rect 19875 335205 19880 335235
rect 19840 335200 19880 335205
rect 19680 335155 19720 335160
rect 19680 335125 19685 335155
rect 19715 335125 19720 335155
rect 19680 335120 19720 335125
rect 19840 335155 19880 335160
rect 19840 335125 19845 335155
rect 19875 335125 19880 335155
rect 19840 335120 19880 335125
rect 19680 335075 19720 335080
rect 19680 335045 19685 335075
rect 19715 335045 19720 335075
rect 19680 335040 19720 335045
rect 19840 335075 19880 335080
rect 19840 335045 19845 335075
rect 19875 335045 19880 335075
rect 19840 335040 19880 335045
rect 19680 334995 19720 335000
rect 19680 334965 19685 334995
rect 19715 334965 19720 334995
rect 19680 334960 19720 334965
rect 19840 334995 19880 335000
rect 19840 334965 19845 334995
rect 19875 334965 19880 334995
rect 19840 334960 19880 334965
rect 19680 334915 19720 334920
rect 19680 334885 19685 334915
rect 19715 334885 19720 334915
rect 19680 334880 19720 334885
rect 19840 334915 19880 334920
rect 19840 334885 19845 334915
rect 19875 334885 19880 334915
rect 19840 334880 19880 334885
rect 19680 334835 19720 334840
rect 19680 334805 19685 334835
rect 19715 334805 19720 334835
rect 19680 334800 19720 334805
rect 19840 334835 19880 334840
rect 19840 334805 19845 334835
rect 19875 334805 19880 334835
rect 19840 334800 19880 334805
rect 19680 334755 19720 334760
rect 19680 334725 19685 334755
rect 19715 334725 19720 334755
rect 19680 334720 19720 334725
rect 19840 334755 19880 334760
rect 19840 334725 19845 334755
rect 19875 334725 19880 334755
rect 19840 334720 19880 334725
rect 19680 334675 19720 334680
rect 19680 334645 19685 334675
rect 19715 334645 19720 334675
rect 19680 334640 19720 334645
rect 19840 334675 19880 334680
rect 19840 334645 19845 334675
rect 19875 334645 19880 334675
rect 19840 334640 19880 334645
rect 19680 334595 19720 334600
rect 19680 334565 19685 334595
rect 19715 334565 19720 334595
rect 19680 334560 19720 334565
rect 19840 334595 19880 334600
rect 19840 334565 19845 334595
rect 19875 334565 19880 334595
rect 19840 334560 19880 334565
rect 19680 334515 19720 334520
rect 19680 334485 19685 334515
rect 19715 334485 19720 334515
rect 19680 334480 19720 334485
rect 19840 334515 19880 334520
rect 19840 334485 19845 334515
rect 19875 334485 19880 334515
rect 19840 334480 19880 334485
rect 19680 334435 19720 334440
rect 19680 334405 19685 334435
rect 19715 334405 19720 334435
rect 19680 334400 19720 334405
rect 19840 334435 19880 334440
rect 19840 334405 19845 334435
rect 19875 334405 19880 334435
rect 19840 334400 19880 334405
rect 19680 334355 19720 334360
rect 19680 334325 19685 334355
rect 19715 334325 19720 334355
rect 19680 334320 19720 334325
rect 19840 334355 19880 334360
rect 19840 334325 19845 334355
rect 19875 334325 19880 334355
rect 19840 334320 19880 334325
rect 19680 334275 19720 334280
rect 19680 334245 19685 334275
rect 19715 334245 19720 334275
rect 19680 334240 19720 334245
rect 19840 334275 19880 334280
rect 19840 334245 19845 334275
rect 19875 334245 19880 334275
rect 19840 334240 19880 334245
rect 19680 334195 19720 334200
rect 19680 334165 19685 334195
rect 19715 334165 19720 334195
rect 19680 334160 19720 334165
rect 19840 334195 19880 334200
rect 19840 334165 19845 334195
rect 19875 334165 19880 334195
rect 19840 334160 19880 334165
rect 19680 334115 19720 334120
rect 19680 334085 19685 334115
rect 19715 334085 19720 334115
rect 19680 334080 19720 334085
rect 19840 334115 19880 334120
rect 19840 334085 19845 334115
rect 19875 334085 19880 334115
rect 19840 334080 19880 334085
rect 19680 334035 19720 334040
rect 19680 334005 19685 334035
rect 19715 334005 19720 334035
rect 19680 334000 19720 334005
rect 19840 334035 19880 334040
rect 19840 334005 19845 334035
rect 19875 334005 19880 334035
rect 19840 334000 19880 334005
rect 19680 333955 19720 333960
rect 19680 333925 19685 333955
rect 19715 333925 19720 333955
rect 19680 333920 19720 333925
rect 19840 333955 19880 333960
rect 19840 333925 19845 333955
rect 19875 333925 19880 333955
rect 19840 333920 19880 333925
rect 19680 333875 19720 333880
rect 19680 333845 19685 333875
rect 19715 333845 19720 333875
rect 19680 333840 19720 333845
rect 19840 333875 19880 333880
rect 19840 333845 19845 333875
rect 19875 333845 19880 333875
rect 19840 333840 19880 333845
rect 19680 333795 19720 333800
rect 19680 333765 19685 333795
rect 19715 333765 19720 333795
rect 19680 333760 19720 333765
rect 19840 333795 19880 333800
rect 19840 333765 19845 333795
rect 19875 333765 19880 333795
rect 19840 333760 19880 333765
rect 19680 333715 19720 333720
rect 19680 333685 19685 333715
rect 19715 333685 19720 333715
rect 19680 333680 19720 333685
rect 19840 333715 19880 333720
rect 19840 333685 19845 333715
rect 19875 333685 19880 333715
rect 19840 333680 19880 333685
rect 19680 333635 19720 333640
rect 19680 333605 19685 333635
rect 19715 333605 19720 333635
rect 19680 333600 19720 333605
rect 19840 333635 19880 333640
rect 19840 333605 19845 333635
rect 19875 333605 19880 333635
rect 19840 333600 19880 333605
rect 19680 333555 19720 333560
rect 19680 333525 19685 333555
rect 19715 333525 19720 333555
rect 19680 333520 19720 333525
rect 19840 333555 19880 333560
rect 19840 333525 19845 333555
rect 19875 333525 19880 333555
rect 19840 333520 19880 333525
rect 19680 333475 19720 333480
rect 19680 333445 19685 333475
rect 19715 333445 19720 333475
rect 19680 333440 19720 333445
rect 19840 333475 19880 333480
rect 19840 333445 19845 333475
rect 19875 333445 19880 333475
rect 19840 333440 19880 333445
rect 19680 333395 19720 333400
rect 19680 333365 19685 333395
rect 19715 333365 19720 333395
rect 19680 333360 19720 333365
rect 19840 333395 19880 333400
rect 19840 333365 19845 333395
rect 19875 333365 19880 333395
rect 19840 333360 19880 333365
rect 19680 333315 19720 333320
rect 19680 333285 19685 333315
rect 19715 333285 19720 333315
rect 19680 333280 19720 333285
rect 19840 333315 19880 333320
rect 19840 333285 19845 333315
rect 19875 333285 19880 333315
rect 19840 333280 19880 333285
rect 19680 333235 19720 333240
rect 19680 333205 19685 333235
rect 19715 333205 19720 333235
rect 19680 333200 19720 333205
rect 19840 333235 19880 333240
rect 19840 333205 19845 333235
rect 19875 333205 19880 333235
rect 19840 333200 19880 333205
rect 19680 333155 19720 333160
rect 19680 333125 19685 333155
rect 19715 333125 19720 333155
rect 19680 333120 19720 333125
rect 19840 333155 19880 333160
rect 19840 333125 19845 333155
rect 19875 333125 19880 333155
rect 19840 333120 19880 333125
rect 19680 333075 19720 333080
rect 19680 333045 19685 333075
rect 19715 333045 19720 333075
rect 19680 333040 19720 333045
rect 19840 333075 19880 333080
rect 19840 333045 19845 333075
rect 19875 333045 19880 333075
rect 19840 333040 19880 333045
rect 19680 332995 19720 333000
rect 19680 332965 19685 332995
rect 19715 332965 19720 332995
rect 19680 332960 19720 332965
rect 19840 332995 19880 333000
rect 19840 332965 19845 332995
rect 19875 332965 19880 332995
rect 19840 332960 19880 332965
rect 19680 332915 19720 332920
rect 19680 332885 19685 332915
rect 19715 332885 19720 332915
rect 19680 332880 19720 332885
rect 19840 332915 19880 332920
rect 19840 332885 19845 332915
rect 19875 332885 19880 332915
rect 19840 332880 19880 332885
rect 19680 332835 19720 332840
rect 19680 332805 19685 332835
rect 19715 332805 19720 332835
rect 19680 332800 19720 332805
rect 19840 332835 19880 332840
rect 19840 332805 19845 332835
rect 19875 332805 19880 332835
rect 19840 332800 19880 332805
rect 19680 332755 19720 332760
rect 19680 332725 19685 332755
rect 19715 332725 19720 332755
rect 19680 332720 19720 332725
rect 19840 332755 19880 332760
rect 19840 332725 19845 332755
rect 19875 332725 19880 332755
rect 19840 332720 19880 332725
rect 19680 332675 19720 332680
rect 19680 332645 19685 332675
rect 19715 332645 19720 332675
rect 19680 332640 19720 332645
rect 19840 332675 19880 332680
rect 19840 332645 19845 332675
rect 19875 332645 19880 332675
rect 19840 332640 19880 332645
rect 19680 332595 19720 332600
rect 19680 332565 19685 332595
rect 19715 332565 19720 332595
rect 19680 332560 19720 332565
rect 19840 332595 19880 332600
rect 19840 332565 19845 332595
rect 19875 332565 19880 332595
rect 19840 332560 19880 332565
rect 19680 332515 19720 332520
rect 19680 332485 19685 332515
rect 19715 332485 19720 332515
rect 19680 332480 19720 332485
rect 19840 332515 19880 332520
rect 19840 332485 19845 332515
rect 19875 332485 19880 332515
rect 19840 332480 19880 332485
rect 19680 332435 19720 332440
rect 19680 332405 19685 332435
rect 19715 332405 19720 332435
rect 19680 332400 19720 332405
rect 19840 332435 19880 332440
rect 19840 332405 19845 332435
rect 19875 332405 19880 332435
rect 19840 332400 19880 332405
rect 19680 332355 19720 332360
rect 19680 332325 19685 332355
rect 19715 332325 19720 332355
rect 19680 332320 19720 332325
rect 19840 332355 19880 332360
rect 19840 332325 19845 332355
rect 19875 332325 19880 332355
rect 19840 332320 19880 332325
rect 19680 332275 19720 332280
rect 19680 332245 19685 332275
rect 19715 332245 19720 332275
rect 19680 332240 19720 332245
rect 19840 332275 19880 332280
rect 19840 332245 19845 332275
rect 19875 332245 19880 332275
rect 19840 332240 19880 332245
rect 19680 332195 19720 332200
rect 19680 332165 19685 332195
rect 19715 332165 19720 332195
rect 19680 332160 19720 332165
rect 19840 332195 19880 332200
rect 19840 332165 19845 332195
rect 19875 332165 19880 332195
rect 19840 332160 19880 332165
rect 19680 332115 19720 332120
rect 19680 332085 19685 332115
rect 19715 332085 19720 332115
rect 19680 332080 19720 332085
rect 19840 332115 19880 332120
rect 19840 332085 19845 332115
rect 19875 332085 19880 332115
rect 19840 332080 19880 332085
rect 19680 332035 19720 332040
rect 19680 332005 19685 332035
rect 19715 332005 19720 332035
rect 19680 332000 19720 332005
rect 19840 332035 19880 332040
rect 19840 332005 19845 332035
rect 19875 332005 19880 332035
rect 19840 332000 19880 332005
rect 19680 331955 19720 331960
rect 19680 331925 19685 331955
rect 19715 331925 19720 331955
rect 19680 331920 19720 331925
rect 19840 331955 19880 331960
rect 19840 331925 19845 331955
rect 19875 331925 19880 331955
rect 19840 331920 19880 331925
rect 19680 331875 19720 331880
rect 19680 331845 19685 331875
rect 19715 331845 19720 331875
rect 19680 331840 19720 331845
rect 19840 331875 19880 331880
rect 19840 331845 19845 331875
rect 19875 331845 19880 331875
rect 19840 331840 19880 331845
rect 19680 331795 19720 331800
rect 19680 331765 19685 331795
rect 19715 331765 19720 331795
rect 19680 331760 19720 331765
rect 19840 331795 19880 331800
rect 19840 331765 19845 331795
rect 19875 331765 19880 331795
rect 19840 331760 19880 331765
rect 19680 331715 19720 331720
rect 19680 331685 19685 331715
rect 19715 331685 19720 331715
rect 19680 331680 19720 331685
rect 19840 331715 19880 331720
rect 19840 331685 19845 331715
rect 19875 331685 19880 331715
rect 19840 331680 19880 331685
rect 19680 331635 19720 331640
rect 19680 331605 19685 331635
rect 19715 331605 19720 331635
rect 19680 331600 19720 331605
rect 19840 331635 19880 331640
rect 19840 331605 19845 331635
rect 19875 331605 19880 331635
rect 19840 331600 19880 331605
rect 19680 331555 19720 331560
rect 19680 331525 19685 331555
rect 19715 331525 19720 331555
rect 19680 331520 19720 331525
rect 19840 331555 19880 331560
rect 19840 331525 19845 331555
rect 19875 331525 19880 331555
rect 19840 331520 19880 331525
rect 19680 331475 19720 331480
rect 19680 331445 19685 331475
rect 19715 331445 19720 331475
rect 19680 331440 19720 331445
rect 19840 331475 19880 331480
rect 19840 331445 19845 331475
rect 19875 331445 19880 331475
rect 19840 331440 19880 331445
rect 19680 331395 19720 331400
rect 19680 331365 19685 331395
rect 19715 331365 19720 331395
rect 19680 331360 19720 331365
rect 19840 331395 19880 331400
rect 19840 331365 19845 331395
rect 19875 331365 19880 331395
rect 19840 331360 19880 331365
rect 19680 331315 19720 331320
rect 19680 331285 19685 331315
rect 19715 331285 19720 331315
rect 19680 331280 19720 331285
rect 19840 331315 19880 331320
rect 19840 331285 19845 331315
rect 19875 331285 19880 331315
rect 19840 331280 19880 331285
rect 19680 331235 19720 331240
rect 19680 331205 19685 331235
rect 19715 331205 19720 331235
rect 19680 331200 19720 331205
rect 19840 331235 19880 331240
rect 19840 331205 19845 331235
rect 19875 331205 19880 331235
rect 19840 331200 19880 331205
rect 19680 331155 19720 331160
rect 19680 331125 19685 331155
rect 19715 331125 19720 331155
rect 19680 331120 19720 331125
rect 19840 331155 19880 331160
rect 19840 331125 19845 331155
rect 19875 331125 19880 331155
rect 19840 331120 19880 331125
rect 19680 331075 19720 331080
rect 19680 331045 19685 331075
rect 19715 331045 19720 331075
rect 19680 331040 19720 331045
rect 19840 331075 19880 331080
rect 19840 331045 19845 331075
rect 19875 331045 19880 331075
rect 19840 331040 19880 331045
rect 19680 330995 19720 331000
rect 19680 330965 19685 330995
rect 19715 330965 19720 330995
rect 19680 330960 19720 330965
rect 19840 330995 19880 331000
rect 19840 330965 19845 330995
rect 19875 330965 19880 330995
rect 19840 330960 19880 330965
rect 19680 330915 19720 330920
rect 19680 330885 19685 330915
rect 19715 330885 19720 330915
rect 19680 330880 19720 330885
rect 19840 330915 19880 330920
rect 19840 330885 19845 330915
rect 19875 330885 19880 330915
rect 19840 330880 19880 330885
rect 19680 330835 19720 330840
rect 19680 330805 19685 330835
rect 19715 330805 19720 330835
rect 19680 330800 19720 330805
rect 19840 330835 19880 330840
rect 19840 330805 19845 330835
rect 19875 330805 19880 330835
rect 19840 330800 19880 330805
rect 19680 330755 19720 330760
rect 19680 330725 19685 330755
rect 19715 330725 19720 330755
rect 19680 330720 19720 330725
rect 19840 330755 19880 330760
rect 19840 330725 19845 330755
rect 19875 330725 19880 330755
rect 19840 330720 19880 330725
rect 19680 330675 19720 330680
rect 19680 330645 19685 330675
rect 19715 330645 19720 330675
rect 19680 330640 19720 330645
rect 19840 330675 19880 330680
rect 19840 330645 19845 330675
rect 19875 330645 19880 330675
rect 19840 330640 19880 330645
rect 19680 330595 19720 330600
rect 19680 330565 19685 330595
rect 19715 330565 19720 330595
rect 19680 330560 19720 330565
rect 19840 330595 19880 330600
rect 19840 330565 19845 330595
rect 19875 330565 19880 330595
rect 19840 330560 19880 330565
rect 19680 330515 19720 330520
rect 19680 330485 19685 330515
rect 19715 330485 19720 330515
rect 19680 330480 19720 330485
rect 19840 330515 19880 330520
rect 19840 330485 19845 330515
rect 19875 330485 19880 330515
rect 19840 330480 19880 330485
rect 19680 330435 19720 330440
rect 19680 330405 19685 330435
rect 19715 330405 19720 330435
rect 19680 330400 19720 330405
rect 19840 330435 19880 330440
rect 19840 330405 19845 330435
rect 19875 330405 19880 330435
rect 19840 330400 19880 330405
rect 19680 330355 19720 330360
rect 19680 330325 19685 330355
rect 19715 330325 19720 330355
rect 19680 330320 19720 330325
rect 19840 330355 19880 330360
rect 19840 330325 19845 330355
rect 19875 330325 19880 330355
rect 19840 330320 19880 330325
rect 19680 330275 19720 330280
rect 19680 330245 19685 330275
rect 19715 330245 19720 330275
rect 19680 330240 19720 330245
rect 19840 330275 19880 330280
rect 19840 330245 19845 330275
rect 19875 330245 19880 330275
rect 19840 330240 19880 330245
rect 19680 330195 19720 330200
rect 19680 330165 19685 330195
rect 19715 330165 19720 330195
rect 19680 330160 19720 330165
rect 19840 330195 19880 330200
rect 19840 330165 19845 330195
rect 19875 330165 19880 330195
rect 19840 330160 19880 330165
rect 19680 330115 19720 330120
rect 19680 330085 19685 330115
rect 19715 330085 19720 330115
rect 19680 330080 19720 330085
rect 19840 330115 19880 330120
rect 19840 330085 19845 330115
rect 19875 330085 19880 330115
rect 19840 330080 19880 330085
rect 19680 330035 19720 330040
rect 19680 330005 19685 330035
rect 19715 330005 19720 330035
rect 19680 330000 19720 330005
rect 19840 330035 19880 330040
rect 19840 330005 19845 330035
rect 19875 330005 19880 330035
rect 19840 330000 19880 330005
rect 19680 329955 19720 329960
rect 19680 329925 19685 329955
rect 19715 329925 19720 329955
rect 19680 329920 19720 329925
rect 19840 329955 19880 329960
rect 19840 329925 19845 329955
rect 19875 329925 19880 329955
rect 19840 329920 19880 329925
rect 19680 329875 19720 329880
rect 19680 329845 19685 329875
rect 19715 329845 19720 329875
rect 19680 329840 19720 329845
rect 19840 329875 19880 329880
rect 19840 329845 19845 329875
rect 19875 329845 19880 329875
rect 19840 329840 19880 329845
rect 19680 329795 19720 329800
rect 19680 329765 19685 329795
rect 19715 329765 19720 329795
rect 19680 329760 19720 329765
rect 19840 329795 19880 329800
rect 19840 329765 19845 329795
rect 19875 329765 19880 329795
rect 19840 329760 19880 329765
rect 19680 329715 19720 329720
rect 19680 329685 19685 329715
rect 19715 329685 19720 329715
rect 19680 329680 19720 329685
rect 19840 329715 19880 329720
rect 19840 329685 19845 329715
rect 19875 329685 19880 329715
rect 19840 329680 19880 329685
rect 19680 329635 19720 329640
rect 19680 329605 19685 329635
rect 19715 329605 19720 329635
rect 19680 329600 19720 329605
rect 19840 329635 19880 329640
rect 19840 329605 19845 329635
rect 19875 329605 19880 329635
rect 19840 329600 19880 329605
rect 19680 329555 19720 329560
rect 19680 329525 19685 329555
rect 19715 329525 19720 329555
rect 19680 329520 19720 329525
rect 19840 329555 19880 329560
rect 19840 329525 19845 329555
rect 19875 329525 19880 329555
rect 19840 329520 19880 329525
rect 19680 329475 19720 329480
rect 19680 329445 19685 329475
rect 19715 329445 19720 329475
rect 19680 329440 19720 329445
rect 19840 329475 19880 329480
rect 19840 329445 19845 329475
rect 19875 329445 19880 329475
rect 19840 329440 19880 329445
rect 19680 329395 19720 329400
rect 19680 329365 19685 329395
rect 19715 329365 19720 329395
rect 19680 329360 19720 329365
rect 19840 329395 19880 329400
rect 19840 329365 19845 329395
rect 19875 329365 19880 329395
rect 19840 329360 19880 329365
rect 19680 329315 19720 329320
rect 19680 329285 19685 329315
rect 19715 329285 19720 329315
rect 19680 329280 19720 329285
rect 19840 329315 19880 329320
rect 19840 329285 19845 329315
rect 19875 329285 19880 329315
rect 19840 329280 19880 329285
rect 19680 329235 19720 329240
rect 19680 329205 19685 329235
rect 19715 329205 19720 329235
rect 19680 329200 19720 329205
rect 19840 329235 19880 329240
rect 19840 329205 19845 329235
rect 19875 329205 19880 329235
rect 19840 329200 19880 329205
rect 19680 329155 19720 329160
rect 19680 329125 19685 329155
rect 19715 329125 19720 329155
rect 19680 329120 19720 329125
rect 19840 329155 19880 329160
rect 19840 329125 19845 329155
rect 19875 329125 19880 329155
rect 19840 329120 19880 329125
rect 19680 329075 19720 329080
rect 19680 329045 19685 329075
rect 19715 329045 19720 329075
rect 19680 329040 19720 329045
rect 19840 329075 19880 329080
rect 19840 329045 19845 329075
rect 19875 329045 19880 329075
rect 19840 329040 19880 329045
rect 19680 328995 19720 329000
rect 19680 328965 19685 328995
rect 19715 328965 19720 328995
rect 19680 328960 19720 328965
rect 19840 328995 19880 329000
rect 19840 328965 19845 328995
rect 19875 328965 19880 328995
rect 19840 328960 19880 328965
rect 19680 328915 19720 328920
rect 19680 328885 19685 328915
rect 19715 328885 19720 328915
rect 19680 328880 19720 328885
rect 19840 328915 19880 328920
rect 19840 328885 19845 328915
rect 19875 328885 19880 328915
rect 19840 328880 19880 328885
rect 19680 328835 19720 328840
rect 19680 328805 19685 328835
rect 19715 328805 19720 328835
rect 19680 328800 19720 328805
rect 19840 328835 19880 328840
rect 19840 328805 19845 328835
rect 19875 328805 19880 328835
rect 19840 328800 19880 328805
rect 19680 328755 19720 328760
rect 19680 328725 19685 328755
rect 19715 328725 19720 328755
rect 19680 328720 19720 328725
rect 19840 328755 19880 328760
rect 19840 328725 19845 328755
rect 19875 328725 19880 328755
rect 19840 328720 19880 328725
rect 19680 328675 19720 328680
rect 19680 328645 19685 328675
rect 19715 328645 19720 328675
rect 19680 328640 19720 328645
rect 19840 328675 19880 328680
rect 19840 328645 19845 328675
rect 19875 328645 19880 328675
rect 19840 328640 19880 328645
rect 19680 328595 19720 328600
rect 19680 328565 19685 328595
rect 19715 328565 19720 328595
rect 19680 328560 19720 328565
rect 19840 328595 19880 328600
rect 19840 328565 19845 328595
rect 19875 328565 19880 328595
rect 19840 328560 19880 328565
rect 19680 328515 19720 328520
rect 19680 328485 19685 328515
rect 19715 328485 19720 328515
rect 19680 328480 19720 328485
rect 19840 328515 19880 328520
rect 19840 328485 19845 328515
rect 19875 328485 19880 328515
rect 19840 328480 19880 328485
rect 19680 328435 19720 328440
rect 19680 328405 19685 328435
rect 19715 328405 19720 328435
rect 19680 328400 19720 328405
rect 19840 328435 19880 328440
rect 19840 328405 19845 328435
rect 19875 328405 19880 328435
rect 19840 328400 19880 328405
rect 19680 328355 19720 328360
rect 19680 328325 19685 328355
rect 19715 328325 19720 328355
rect 19680 328320 19720 328325
rect 19840 328355 19880 328360
rect 19840 328325 19845 328355
rect 19875 328325 19880 328355
rect 19840 328320 19880 328325
rect 19680 328275 19720 328280
rect 19680 328245 19685 328275
rect 19715 328245 19720 328275
rect 19680 328240 19720 328245
rect 19840 328275 19880 328280
rect 19840 328245 19845 328275
rect 19875 328245 19880 328275
rect 19840 328240 19880 328245
rect 19680 328195 19720 328200
rect 19680 328165 19685 328195
rect 19715 328165 19720 328195
rect 19680 328160 19720 328165
rect 19840 328195 19880 328200
rect 19840 328165 19845 328195
rect 19875 328165 19880 328195
rect 19840 328160 19880 328165
rect 19680 328115 19720 328120
rect 19680 328085 19685 328115
rect 19715 328085 19720 328115
rect 19680 328080 19720 328085
rect 19840 328115 19880 328120
rect 19840 328085 19845 328115
rect 19875 328085 19880 328115
rect 19840 328080 19880 328085
rect 19680 328035 19720 328040
rect 19680 328005 19685 328035
rect 19715 328005 19720 328035
rect 19680 328000 19720 328005
rect 19840 328035 19880 328040
rect 19840 328005 19845 328035
rect 19875 328005 19880 328035
rect 19840 328000 19880 328005
rect 19680 327955 19720 327960
rect 19680 327925 19685 327955
rect 19715 327925 19720 327955
rect 19680 327920 19720 327925
rect 19840 327955 19880 327960
rect 19840 327925 19845 327955
rect 19875 327925 19880 327955
rect 19840 327920 19880 327925
rect 19680 327875 19720 327880
rect 19680 327845 19685 327875
rect 19715 327845 19720 327875
rect 19680 327840 19720 327845
rect 19840 327875 19880 327880
rect 19840 327845 19845 327875
rect 19875 327845 19880 327875
rect 19840 327840 19880 327845
rect 19680 327795 19720 327800
rect 19680 327765 19685 327795
rect 19715 327765 19720 327795
rect 19680 327760 19720 327765
rect 19840 327795 19880 327800
rect 19840 327765 19845 327795
rect 19875 327765 19880 327795
rect 19840 327760 19880 327765
rect 19680 327715 19720 327720
rect 19680 327685 19685 327715
rect 19715 327685 19720 327715
rect 19680 327680 19720 327685
rect 19840 327715 19880 327720
rect 19840 327685 19845 327715
rect 19875 327685 19880 327715
rect 19840 327680 19880 327685
rect 19680 327635 19720 327640
rect 19680 327605 19685 327635
rect 19715 327605 19720 327635
rect 19680 327600 19720 327605
rect 19840 327635 19880 327640
rect 19840 327605 19845 327635
rect 19875 327605 19880 327635
rect 19840 327600 19880 327605
rect 19680 327555 19720 327560
rect 19680 327525 19685 327555
rect 19715 327525 19720 327555
rect 19680 327520 19720 327525
rect 19840 327555 19880 327560
rect 19840 327525 19845 327555
rect 19875 327525 19880 327555
rect 19840 327520 19880 327525
rect 19680 327475 19720 327480
rect 19680 327445 19685 327475
rect 19715 327445 19720 327475
rect 19680 327440 19720 327445
rect 19840 327475 19880 327480
rect 19840 327445 19845 327475
rect 19875 327445 19880 327475
rect 19840 327440 19880 327445
rect 19680 327395 19720 327400
rect 19680 327365 19685 327395
rect 19715 327365 19720 327395
rect 19680 327360 19720 327365
rect 19840 327395 19880 327400
rect 19840 327365 19845 327395
rect 19875 327365 19880 327395
rect 19840 327360 19880 327365
rect 19680 327315 19720 327320
rect 19680 327285 19685 327315
rect 19715 327285 19720 327315
rect 19680 327280 19720 327285
rect 19840 327315 19880 327320
rect 19840 327285 19845 327315
rect 19875 327285 19880 327315
rect 19840 327280 19880 327285
rect 19680 327235 19720 327240
rect 19680 327205 19685 327235
rect 19715 327205 19720 327235
rect 19680 327200 19720 327205
rect 19840 327235 19880 327240
rect 19840 327205 19845 327235
rect 19875 327205 19880 327235
rect 19840 327200 19880 327205
rect 19680 327155 19720 327160
rect 19680 327125 19685 327155
rect 19715 327125 19720 327155
rect 19680 327120 19720 327125
rect 19840 327155 19880 327160
rect 19840 327125 19845 327155
rect 19875 327125 19880 327155
rect 19840 327120 19880 327125
rect 19680 327075 19720 327080
rect 19680 327045 19685 327075
rect 19715 327045 19720 327075
rect 19680 327040 19720 327045
rect 19840 327075 19880 327080
rect 19840 327045 19845 327075
rect 19875 327045 19880 327075
rect 19840 327040 19880 327045
rect 19680 326995 19720 327000
rect 19680 326965 19685 326995
rect 19715 326965 19720 326995
rect 19680 326960 19720 326965
rect 19840 326995 19880 327000
rect 19840 326965 19845 326995
rect 19875 326965 19880 326995
rect 19840 326960 19880 326965
rect 19680 326915 19720 326920
rect 19680 326885 19685 326915
rect 19715 326885 19720 326915
rect 19680 326880 19720 326885
rect 19840 326915 19880 326920
rect 19840 326885 19845 326915
rect 19875 326885 19880 326915
rect 19840 326880 19880 326885
rect 19680 326835 19720 326840
rect 19680 326805 19685 326835
rect 19715 326805 19720 326835
rect 19680 326800 19720 326805
rect 19840 326835 19880 326840
rect 19840 326805 19845 326835
rect 19875 326805 19880 326835
rect 19840 326800 19880 326805
rect 19680 326755 19720 326760
rect 19680 326725 19685 326755
rect 19715 326725 19720 326755
rect 19680 326720 19720 326725
rect 19840 326755 19880 326760
rect 19840 326725 19845 326755
rect 19875 326725 19880 326755
rect 19840 326720 19880 326725
rect 19680 326675 19720 326680
rect 19680 326645 19685 326675
rect 19715 326645 19720 326675
rect 19680 326640 19720 326645
rect 19840 326675 19880 326680
rect 19840 326645 19845 326675
rect 19875 326645 19880 326675
rect 19840 326640 19880 326645
rect 19680 326595 19720 326600
rect 19680 326565 19685 326595
rect 19715 326565 19720 326595
rect 19680 326560 19720 326565
rect 19840 326595 19880 326600
rect 19840 326565 19845 326595
rect 19875 326565 19880 326595
rect 19840 326560 19880 326565
rect 19680 326515 19720 326520
rect 19680 326485 19685 326515
rect 19715 326485 19720 326515
rect 19680 326480 19720 326485
rect 19840 326515 19880 326520
rect 19840 326485 19845 326515
rect 19875 326485 19880 326515
rect 19840 326480 19880 326485
rect 19680 326435 19720 326440
rect 19680 326405 19685 326435
rect 19715 326405 19720 326435
rect 19680 326400 19720 326405
rect 19840 326435 19880 326440
rect 19840 326405 19845 326435
rect 19875 326405 19880 326435
rect 19840 326400 19880 326405
rect 19680 326355 19720 326360
rect 19680 326325 19685 326355
rect 19715 326325 19720 326355
rect 19680 326320 19720 326325
rect 19840 326355 19880 326360
rect 19840 326325 19845 326355
rect 19875 326325 19880 326355
rect 19840 326320 19880 326325
rect 19680 326275 19720 326280
rect 19680 326245 19685 326275
rect 19715 326245 19720 326275
rect 19680 326240 19720 326245
rect 19840 326275 19880 326280
rect 19840 326245 19845 326275
rect 19875 326245 19880 326275
rect 19840 326240 19880 326245
rect 19680 326195 19720 326200
rect 19680 326165 19685 326195
rect 19715 326165 19720 326195
rect 19680 326160 19720 326165
rect 19840 326195 19880 326200
rect 19840 326165 19845 326195
rect 19875 326165 19880 326195
rect 19840 326160 19880 326165
rect 19680 326115 19720 326120
rect 19680 326085 19685 326115
rect 19715 326085 19720 326115
rect 19680 326080 19720 326085
rect 19840 326115 19880 326120
rect 19840 326085 19845 326115
rect 19875 326085 19880 326115
rect 19840 326080 19880 326085
rect 19680 326035 19720 326040
rect 19680 326005 19685 326035
rect 19715 326005 19720 326035
rect 19680 326000 19720 326005
rect 19840 326035 19880 326040
rect 19840 326005 19845 326035
rect 19875 326005 19880 326035
rect 19840 326000 19880 326005
rect 19680 325955 19720 325960
rect 19680 325925 19685 325955
rect 19715 325925 19720 325955
rect 19680 325920 19720 325925
rect 19840 325955 19880 325960
rect 19840 325925 19845 325955
rect 19875 325925 19880 325955
rect 19840 325920 19880 325925
rect 19680 325875 19720 325880
rect 19680 325845 19685 325875
rect 19715 325845 19720 325875
rect 19680 325840 19720 325845
rect 19840 325875 19880 325880
rect 19840 325845 19845 325875
rect 19875 325845 19880 325875
rect 19840 325840 19880 325845
rect 19680 325795 19720 325800
rect 19680 325765 19685 325795
rect 19715 325765 19720 325795
rect 19680 325760 19720 325765
rect 19840 325795 19880 325800
rect 19840 325765 19845 325795
rect 19875 325765 19880 325795
rect 19840 325760 19880 325765
rect 19680 325715 19720 325720
rect 19680 325685 19685 325715
rect 19715 325685 19720 325715
rect 19680 325680 19720 325685
rect 19840 325715 19880 325720
rect 19840 325685 19845 325715
rect 19875 325685 19880 325715
rect 19840 325680 19880 325685
rect 19680 325635 19720 325640
rect 19680 325605 19685 325635
rect 19715 325605 19720 325635
rect 19680 325600 19720 325605
rect 19840 325635 19880 325640
rect 19840 325605 19845 325635
rect 19875 325605 19880 325635
rect 19840 325600 19880 325605
rect 19680 325555 19720 325560
rect 19680 325525 19685 325555
rect 19715 325525 19720 325555
rect 19680 325520 19720 325525
rect 19840 325555 19880 325560
rect 19840 325525 19845 325555
rect 19875 325525 19880 325555
rect 19840 325520 19880 325525
rect 19680 325475 19720 325480
rect 19680 325445 19685 325475
rect 19715 325445 19720 325475
rect 19680 325440 19720 325445
rect 19840 325475 19880 325480
rect 19840 325445 19845 325475
rect 19875 325445 19880 325475
rect 19840 325440 19880 325445
rect 19680 325395 19720 325400
rect 19680 325365 19685 325395
rect 19715 325365 19720 325395
rect 19680 325360 19720 325365
rect 19840 325395 19880 325400
rect 19840 325365 19845 325395
rect 19875 325365 19880 325395
rect 19840 325360 19880 325365
rect 19680 325315 19720 325320
rect 19680 325285 19685 325315
rect 19715 325285 19720 325315
rect 19680 325280 19720 325285
rect 19840 325315 19880 325320
rect 19840 325285 19845 325315
rect 19875 325285 19880 325315
rect 19840 325280 19880 325285
rect 19680 325235 19720 325240
rect 19680 325205 19685 325235
rect 19715 325205 19720 325235
rect 19680 325200 19720 325205
rect 19840 325235 19880 325240
rect 19840 325205 19845 325235
rect 19875 325205 19880 325235
rect 19840 325200 19880 325205
rect 19680 325155 19720 325160
rect 19680 325125 19685 325155
rect 19715 325125 19720 325155
rect 19680 325120 19720 325125
rect 19840 325155 19880 325160
rect 19840 325125 19845 325155
rect 19875 325125 19880 325155
rect 19840 325120 19880 325125
rect 19680 325075 19720 325080
rect 19680 325045 19685 325075
rect 19715 325045 19720 325075
rect 19680 325040 19720 325045
rect 19840 325075 19880 325080
rect 19840 325045 19845 325075
rect 19875 325045 19880 325075
rect 19840 325040 19880 325045
rect 19680 324995 19720 325000
rect 19680 324965 19685 324995
rect 19715 324965 19720 324995
rect 19680 324960 19720 324965
rect 19840 324995 19880 325000
rect 19840 324965 19845 324995
rect 19875 324965 19880 324995
rect 19840 324960 19880 324965
rect 19680 324915 19720 324920
rect 19680 324885 19685 324915
rect 19715 324885 19720 324915
rect 19680 324880 19720 324885
rect 19840 324915 19880 324920
rect 19840 324885 19845 324915
rect 19875 324885 19880 324915
rect 19840 324880 19880 324885
rect 19680 324835 19720 324840
rect 19680 324805 19685 324835
rect 19715 324805 19720 324835
rect 19680 324800 19720 324805
rect 19840 324835 19880 324840
rect 19840 324805 19845 324835
rect 19875 324805 19880 324835
rect 19840 324800 19880 324805
rect 19680 324755 19720 324760
rect 19680 324725 19685 324755
rect 19715 324725 19720 324755
rect 19680 324720 19720 324725
rect 19840 324755 19880 324760
rect 19840 324725 19845 324755
rect 19875 324725 19880 324755
rect 19840 324720 19880 324725
rect 19680 324675 19720 324680
rect 19680 324645 19685 324675
rect 19715 324645 19720 324675
rect 19680 324640 19720 324645
rect 19840 324675 19880 324680
rect 19840 324645 19845 324675
rect 19875 324645 19880 324675
rect 19840 324640 19880 324645
rect 19680 324595 19720 324600
rect 19680 324565 19685 324595
rect 19715 324565 19720 324595
rect 19680 324560 19720 324565
rect 19840 324595 19880 324600
rect 19840 324565 19845 324595
rect 19875 324565 19880 324595
rect 19840 324560 19880 324565
rect 19680 324515 19720 324520
rect 19680 324485 19685 324515
rect 19715 324485 19720 324515
rect 19680 324480 19720 324485
rect 19840 324515 19880 324520
rect 19840 324485 19845 324515
rect 19875 324485 19880 324515
rect 19840 324480 19880 324485
rect 19680 324435 19720 324440
rect 19680 324405 19685 324435
rect 19715 324405 19720 324435
rect 19680 324400 19720 324405
rect 19840 324435 19880 324440
rect 19840 324405 19845 324435
rect 19875 324405 19880 324435
rect 19840 324400 19880 324405
rect 19680 324355 19720 324360
rect 19680 324325 19685 324355
rect 19715 324325 19720 324355
rect 19680 324320 19720 324325
rect 19840 324355 19880 324360
rect 19840 324325 19845 324355
rect 19875 324325 19880 324355
rect 19840 324320 19880 324325
rect 19680 324275 19720 324280
rect 19680 324245 19685 324275
rect 19715 324245 19720 324275
rect 19680 324240 19720 324245
rect 19840 324275 19880 324280
rect 19840 324245 19845 324275
rect 19875 324245 19880 324275
rect 19840 324240 19880 324245
rect 19680 324195 19720 324200
rect 19680 324165 19685 324195
rect 19715 324165 19720 324195
rect 19680 324160 19720 324165
rect 19840 324195 19880 324200
rect 19840 324165 19845 324195
rect 19875 324165 19880 324195
rect 19840 324160 19880 324165
rect 19680 324115 19720 324120
rect 19680 324085 19685 324115
rect 19715 324085 19720 324115
rect 19680 324080 19720 324085
rect 19840 324115 19880 324120
rect 19840 324085 19845 324115
rect 19875 324085 19880 324115
rect 19840 324080 19880 324085
rect 19680 324035 19720 324040
rect 19680 324005 19685 324035
rect 19715 324005 19720 324035
rect 19680 324000 19720 324005
rect 19840 324035 19880 324040
rect 19840 324005 19845 324035
rect 19875 324005 19880 324035
rect 19840 324000 19880 324005
rect 19680 323955 19720 323960
rect 19680 323925 19685 323955
rect 19715 323925 19720 323955
rect 19680 323920 19720 323925
rect 19840 323955 19880 323960
rect 19840 323925 19845 323955
rect 19875 323925 19880 323955
rect 19840 323920 19880 323925
rect 19680 323875 19720 323880
rect 19680 323845 19685 323875
rect 19715 323845 19720 323875
rect 19680 323840 19720 323845
rect 19840 323875 19880 323880
rect 19840 323845 19845 323875
rect 19875 323845 19880 323875
rect 19840 323840 19880 323845
rect 19680 323795 19720 323800
rect 19680 323765 19685 323795
rect 19715 323765 19720 323795
rect 19680 323760 19720 323765
rect 19840 323795 19880 323800
rect 19840 323765 19845 323795
rect 19875 323765 19880 323795
rect 19840 323760 19880 323765
rect 19680 323715 19720 323720
rect 19680 323685 19685 323715
rect 19715 323685 19720 323715
rect 19680 323680 19720 323685
rect 19840 323715 19880 323720
rect 19840 323685 19845 323715
rect 19875 323685 19880 323715
rect 19840 323680 19880 323685
rect 19680 323635 19720 323640
rect 19680 323605 19685 323635
rect 19715 323605 19720 323635
rect 19680 323600 19720 323605
rect 19840 323635 19880 323640
rect 19840 323605 19845 323635
rect 19875 323605 19880 323635
rect 19840 323600 19880 323605
rect 19680 323555 19720 323560
rect 19680 323525 19685 323555
rect 19715 323525 19720 323555
rect 19680 323520 19720 323525
rect 19840 323555 19880 323560
rect 19840 323525 19845 323555
rect 19875 323525 19880 323555
rect 19840 323520 19880 323525
rect 19680 323475 19720 323480
rect 19680 323445 19685 323475
rect 19715 323445 19720 323475
rect 19680 323440 19720 323445
rect 19840 323475 19880 323480
rect 19840 323445 19845 323475
rect 19875 323445 19880 323475
rect 19840 323440 19880 323445
rect 19680 323395 19720 323400
rect 19680 323365 19685 323395
rect 19715 323365 19720 323395
rect 19680 323360 19720 323365
rect 19840 323395 19880 323400
rect 19840 323365 19845 323395
rect 19875 323365 19880 323395
rect 19840 323360 19880 323365
rect 19680 323315 19720 323320
rect 19680 323285 19685 323315
rect 19715 323285 19720 323315
rect 19680 323280 19720 323285
rect 19840 323315 19880 323320
rect 19840 323285 19845 323315
rect 19875 323285 19880 323315
rect 19840 323280 19880 323285
rect 19680 323235 19720 323240
rect 19680 323205 19685 323235
rect 19715 323205 19720 323235
rect 19680 323200 19720 323205
rect 19840 323235 19880 323240
rect 19840 323205 19845 323235
rect 19875 323205 19880 323235
rect 19840 323200 19880 323205
rect 19680 323155 19720 323160
rect 19680 323125 19685 323155
rect 19715 323125 19720 323155
rect 19680 323120 19720 323125
rect 19840 323155 19880 323160
rect 19840 323125 19845 323155
rect 19875 323125 19880 323155
rect 19840 323120 19880 323125
rect 19680 323075 19720 323080
rect 19680 323045 19685 323075
rect 19715 323045 19720 323075
rect 19680 323040 19720 323045
rect 19840 323075 19880 323080
rect 19840 323045 19845 323075
rect 19875 323045 19880 323075
rect 19840 323040 19880 323045
rect 19680 322995 19720 323000
rect 19680 322965 19685 322995
rect 19715 322965 19720 322995
rect 19680 322960 19720 322965
rect 19840 322995 19880 323000
rect 19840 322965 19845 322995
rect 19875 322965 19880 322995
rect 19840 322960 19880 322965
rect 19680 322915 19720 322920
rect 19680 322885 19685 322915
rect 19715 322885 19720 322915
rect 19680 322880 19720 322885
rect 19840 322915 19880 322920
rect 19840 322885 19845 322915
rect 19875 322885 19880 322915
rect 19840 322880 19880 322885
rect 19680 322835 19720 322840
rect 19680 322805 19685 322835
rect 19715 322805 19720 322835
rect 19680 322800 19720 322805
rect 19840 322835 19880 322840
rect 19840 322805 19845 322835
rect 19875 322805 19880 322835
rect 19840 322800 19880 322805
rect 19680 322755 19720 322760
rect 19680 322725 19685 322755
rect 19715 322725 19720 322755
rect 19680 322720 19720 322725
rect 19840 322755 19880 322760
rect 19840 322725 19845 322755
rect 19875 322725 19880 322755
rect 19840 322720 19880 322725
rect 19680 322675 19720 322680
rect 19680 322645 19685 322675
rect 19715 322645 19720 322675
rect 19680 322640 19720 322645
rect 19840 322675 19880 322680
rect 19840 322645 19845 322675
rect 19875 322645 19880 322675
rect 19840 322640 19880 322645
rect 19680 322595 19720 322600
rect 19680 322565 19685 322595
rect 19715 322565 19720 322595
rect 19680 322560 19720 322565
rect 19840 322595 19880 322600
rect 19840 322565 19845 322595
rect 19875 322565 19880 322595
rect 19840 322560 19880 322565
rect 19680 322515 19720 322520
rect 19680 322485 19685 322515
rect 19715 322485 19720 322515
rect 19680 322480 19720 322485
rect 19840 322515 19880 322520
rect 19840 322485 19845 322515
rect 19875 322485 19880 322515
rect 19840 322480 19880 322485
rect 19680 322435 19720 322440
rect 19680 322405 19685 322435
rect 19715 322405 19720 322435
rect 19680 322400 19720 322405
rect 19840 322435 19880 322440
rect 19840 322405 19845 322435
rect 19875 322405 19880 322435
rect 19840 322400 19880 322405
rect 19680 322355 19720 322360
rect 19680 322325 19685 322355
rect 19715 322325 19720 322355
rect 19680 322320 19720 322325
rect 19840 322355 19880 322360
rect 19840 322325 19845 322355
rect 19875 322325 19880 322355
rect 19840 322320 19880 322325
rect 19680 322275 19720 322280
rect 19680 322245 19685 322275
rect 19715 322245 19720 322275
rect 19680 322240 19720 322245
rect 19840 322275 19880 322280
rect 19840 322245 19845 322275
rect 19875 322245 19880 322275
rect 19840 322240 19880 322245
rect 19680 322195 19720 322200
rect 19680 322165 19685 322195
rect 19715 322165 19720 322195
rect 19680 322160 19720 322165
rect 19840 322195 19880 322200
rect 19840 322165 19845 322195
rect 19875 322165 19880 322195
rect 19840 322160 19880 322165
rect 19680 322115 19720 322120
rect 19680 322085 19685 322115
rect 19715 322085 19720 322115
rect 19680 322080 19720 322085
rect 19840 322115 19880 322120
rect 19840 322085 19845 322115
rect 19875 322085 19880 322115
rect 19840 322080 19880 322085
rect 19680 322035 19720 322040
rect 19680 322005 19685 322035
rect 19715 322005 19720 322035
rect 19680 322000 19720 322005
rect 19840 322035 19880 322040
rect 19840 322005 19845 322035
rect 19875 322005 19880 322035
rect 19840 322000 19880 322005
rect 19680 321955 19720 321960
rect 19680 321925 19685 321955
rect 19715 321925 19720 321955
rect 19680 321920 19720 321925
rect 19840 321955 19880 321960
rect 19840 321925 19845 321955
rect 19875 321925 19880 321955
rect 19840 321920 19880 321925
rect 19680 321875 19720 321880
rect 19680 321845 19685 321875
rect 19715 321845 19720 321875
rect 19680 321840 19720 321845
rect 19840 321875 19880 321880
rect 19840 321845 19845 321875
rect 19875 321845 19880 321875
rect 19840 321840 19880 321845
rect 19680 321795 19720 321800
rect 19680 321765 19685 321795
rect 19715 321765 19720 321795
rect 19680 321760 19720 321765
rect 19840 321795 19880 321800
rect 19840 321765 19845 321795
rect 19875 321765 19880 321795
rect 19840 321760 19880 321765
rect 19680 321715 19720 321720
rect 19680 321685 19685 321715
rect 19715 321685 19720 321715
rect 19680 321680 19720 321685
rect 19840 321715 19880 321720
rect 19840 321685 19845 321715
rect 19875 321685 19880 321715
rect 19840 321680 19880 321685
rect 19680 321635 19720 321640
rect 19680 321605 19685 321635
rect 19715 321605 19720 321635
rect 19680 321600 19720 321605
rect 19840 321635 19880 321640
rect 19840 321605 19845 321635
rect 19875 321605 19880 321635
rect 19840 321600 19880 321605
rect 19680 321555 19720 321560
rect 19680 321525 19685 321555
rect 19715 321525 19720 321555
rect 19680 321520 19720 321525
rect 19840 321555 19880 321560
rect 19840 321525 19845 321555
rect 19875 321525 19880 321555
rect 19840 321520 19880 321525
rect 19680 321475 19720 321480
rect 19680 321445 19685 321475
rect 19715 321445 19720 321475
rect 19680 321440 19720 321445
rect 19840 321475 19880 321480
rect 19840 321445 19845 321475
rect 19875 321445 19880 321475
rect 19840 321440 19880 321445
rect 19680 321395 19720 321400
rect 19680 321365 19685 321395
rect 19715 321365 19720 321395
rect 19680 321360 19720 321365
rect 19840 321395 19880 321400
rect 19840 321365 19845 321395
rect 19875 321365 19880 321395
rect 19840 321360 19880 321365
rect 19680 321315 19720 321320
rect 19680 321285 19685 321315
rect 19715 321285 19720 321315
rect 19680 321280 19720 321285
rect 19840 321315 19880 321320
rect 19840 321285 19845 321315
rect 19875 321285 19880 321315
rect 19840 321280 19880 321285
rect 19680 321235 19720 321240
rect 19680 321205 19685 321235
rect 19715 321205 19720 321235
rect 19680 321200 19720 321205
rect 19840 321235 19880 321240
rect 19840 321205 19845 321235
rect 19875 321205 19880 321235
rect 19840 321200 19880 321205
rect 19680 321155 19720 321160
rect 19680 321125 19685 321155
rect 19715 321125 19720 321155
rect 19680 321120 19720 321125
rect 19840 321155 19880 321160
rect 19840 321125 19845 321155
rect 19875 321125 19880 321155
rect 19840 321120 19880 321125
rect 19680 321075 19720 321080
rect 19680 321045 19685 321075
rect 19715 321045 19720 321075
rect 19680 321040 19720 321045
rect 19840 321075 19880 321080
rect 19840 321045 19845 321075
rect 19875 321045 19880 321075
rect 19840 321040 19880 321045
rect 19680 320995 19720 321000
rect 19680 320965 19685 320995
rect 19715 320965 19720 320995
rect 19680 320960 19720 320965
rect 19840 320995 19880 321000
rect 19840 320965 19845 320995
rect 19875 320965 19880 320995
rect 19840 320960 19880 320965
rect 19680 320915 19720 320920
rect 19680 320885 19685 320915
rect 19715 320885 19720 320915
rect 19680 320880 19720 320885
rect 19840 320915 19880 320920
rect 19840 320885 19845 320915
rect 19875 320885 19880 320915
rect 19840 320880 19880 320885
rect 19680 320835 19720 320840
rect 19680 320805 19685 320835
rect 19715 320805 19720 320835
rect 19680 320800 19720 320805
rect 19840 320835 19880 320840
rect 19840 320805 19845 320835
rect 19875 320805 19880 320835
rect 19840 320800 19880 320805
rect 19680 320755 19720 320760
rect 19680 320725 19685 320755
rect 19715 320725 19720 320755
rect 19680 320720 19720 320725
rect 19840 320755 19880 320760
rect 19840 320725 19845 320755
rect 19875 320725 19880 320755
rect 19840 320720 19880 320725
rect 19680 320675 19720 320680
rect 19680 320645 19685 320675
rect 19715 320645 19720 320675
rect 19680 320640 19720 320645
rect 19840 320675 19880 320680
rect 19840 320645 19845 320675
rect 19875 320645 19880 320675
rect 19840 320640 19880 320645
rect 19680 320595 19720 320600
rect 19680 320565 19685 320595
rect 19715 320565 19720 320595
rect 19680 320560 19720 320565
rect 19840 320595 19880 320600
rect 19840 320565 19845 320595
rect 19875 320565 19880 320595
rect 19840 320560 19880 320565
rect 19680 320515 19720 320520
rect 19680 320485 19685 320515
rect 19715 320485 19720 320515
rect 19680 320480 19720 320485
rect 19840 320515 19880 320520
rect 19840 320485 19845 320515
rect 19875 320485 19880 320515
rect 19840 320480 19880 320485
rect 19680 320435 19720 320440
rect 19680 320405 19685 320435
rect 19715 320405 19720 320435
rect 19680 320400 19720 320405
rect 19840 320435 19880 320440
rect 19840 320405 19845 320435
rect 19875 320405 19880 320435
rect 19840 320400 19880 320405
rect 19680 320355 19720 320360
rect 19680 320325 19685 320355
rect 19715 320325 19720 320355
rect 19680 320320 19720 320325
rect 19840 320355 19880 320360
rect 19840 320325 19845 320355
rect 19875 320325 19880 320355
rect 19840 320320 19880 320325
rect 19680 320275 19720 320280
rect 19680 320245 19685 320275
rect 19715 320245 19720 320275
rect 19680 320240 19720 320245
rect 19840 320275 19880 320280
rect 19840 320245 19845 320275
rect 19875 320245 19880 320275
rect 19840 320240 19880 320245
rect 19680 320195 19720 320200
rect 19680 320165 19685 320195
rect 19715 320165 19720 320195
rect 19680 320160 19720 320165
rect 19840 320195 19880 320200
rect 19840 320165 19845 320195
rect 19875 320165 19880 320195
rect 19840 320160 19880 320165
rect 19680 320115 19720 320120
rect 19680 320085 19685 320115
rect 19715 320085 19720 320115
rect 19680 320080 19720 320085
rect 19840 320115 19880 320120
rect 19840 320085 19845 320115
rect 19875 320085 19880 320115
rect 19840 320080 19880 320085
rect 19680 320035 19720 320040
rect 19680 320005 19685 320035
rect 19715 320005 19720 320035
rect 19680 320000 19720 320005
rect 19840 320035 19880 320040
rect 19840 320005 19845 320035
rect 19875 320005 19880 320035
rect 19840 320000 19880 320005
rect 19680 319955 19720 319960
rect 19680 319925 19685 319955
rect 19715 319925 19720 319955
rect 19680 319920 19720 319925
rect 19840 319955 19880 319960
rect 19840 319925 19845 319955
rect 19875 319925 19880 319955
rect 19840 319920 19880 319925
rect 19680 319875 19720 319880
rect 19680 319845 19685 319875
rect 19715 319845 19720 319875
rect 19680 319840 19720 319845
rect 19840 319875 19880 319880
rect 19840 319845 19845 319875
rect 19875 319845 19880 319875
rect 19840 319840 19880 319845
rect 19680 319795 19720 319800
rect 19680 319765 19685 319795
rect 19715 319765 19720 319795
rect 19680 319760 19720 319765
rect 19840 319795 19880 319800
rect 19840 319765 19845 319795
rect 19875 319765 19880 319795
rect 19840 319760 19880 319765
rect 19680 319715 19720 319720
rect 19680 319685 19685 319715
rect 19715 319685 19720 319715
rect 19680 319680 19720 319685
rect 19840 319715 19880 319720
rect 19840 319685 19845 319715
rect 19875 319685 19880 319715
rect 19840 319680 19880 319685
rect 19680 319635 19720 319640
rect 19680 319605 19685 319635
rect 19715 319605 19720 319635
rect 19680 319600 19720 319605
rect 19840 319635 19880 319640
rect 19840 319605 19845 319635
rect 19875 319605 19880 319635
rect 19840 319600 19880 319605
rect 19680 319555 19720 319560
rect 19680 319525 19685 319555
rect 19715 319525 19720 319555
rect 19680 319520 19720 319525
rect 19840 319555 19880 319560
rect 19840 319525 19845 319555
rect 19875 319525 19880 319555
rect 19840 319520 19880 319525
rect 19680 319475 19720 319480
rect 19680 319445 19685 319475
rect 19715 319445 19720 319475
rect 19680 319440 19720 319445
rect 19840 319475 19880 319480
rect 19840 319445 19845 319475
rect 19875 319445 19880 319475
rect 19840 319440 19880 319445
rect 19680 319395 19720 319400
rect 19680 319365 19685 319395
rect 19715 319365 19720 319395
rect 19680 319360 19720 319365
rect 19840 319395 19880 319400
rect 19840 319365 19845 319395
rect 19875 319365 19880 319395
rect 19840 319360 19880 319365
rect 19680 319315 19720 319320
rect 19680 319285 19685 319315
rect 19715 319285 19720 319315
rect 19680 319280 19720 319285
rect 19840 319315 19880 319320
rect 19840 319285 19845 319315
rect 19875 319285 19880 319315
rect 19840 319280 19880 319285
rect 19680 319235 19720 319240
rect 19680 319205 19685 319235
rect 19715 319205 19720 319235
rect 19680 319200 19720 319205
rect 19840 319235 19880 319240
rect 19840 319205 19845 319235
rect 19875 319205 19880 319235
rect 19840 319200 19880 319205
rect 19680 319155 19720 319160
rect 19680 319125 19685 319155
rect 19715 319125 19720 319155
rect 19680 319120 19720 319125
rect 19840 319155 19880 319160
rect 19840 319125 19845 319155
rect 19875 319125 19880 319155
rect 19840 319120 19880 319125
rect 19680 319075 19720 319080
rect 19680 319045 19685 319075
rect 19715 319045 19720 319075
rect 19680 319040 19720 319045
rect 19840 319075 19880 319080
rect 19840 319045 19845 319075
rect 19875 319045 19880 319075
rect 19840 319040 19880 319045
rect 19680 318995 19720 319000
rect 19680 318965 19685 318995
rect 19715 318965 19720 318995
rect 19680 318960 19720 318965
rect 19840 318995 19880 319000
rect 19840 318965 19845 318995
rect 19875 318965 19880 318995
rect 19840 318960 19880 318965
rect 19680 318915 19720 318920
rect 19680 318885 19685 318915
rect 19715 318885 19720 318915
rect 19680 318880 19720 318885
rect 19840 318915 19880 318920
rect 19840 318885 19845 318915
rect 19875 318885 19880 318915
rect 19840 318880 19880 318885
rect 19680 318835 19720 318840
rect 19680 318805 19685 318835
rect 19715 318805 19720 318835
rect 19680 318800 19720 318805
rect 19840 318835 19880 318840
rect 19840 318805 19845 318835
rect 19875 318805 19880 318835
rect 19840 318800 19880 318805
rect 19680 318755 19720 318760
rect 19680 318725 19685 318755
rect 19715 318725 19720 318755
rect 19680 318720 19720 318725
rect 19840 318755 19880 318760
rect 19840 318725 19845 318755
rect 19875 318725 19880 318755
rect 19840 318720 19880 318725
rect 19680 318675 19720 318680
rect 19680 318645 19685 318675
rect 19715 318645 19720 318675
rect 19680 318640 19720 318645
rect 19840 318675 19880 318680
rect 19840 318645 19845 318675
rect 19875 318645 19880 318675
rect 19840 318640 19880 318645
rect 19680 318595 19720 318600
rect 19680 318565 19685 318595
rect 19715 318565 19720 318595
rect 19680 318560 19720 318565
rect 19840 318595 19880 318600
rect 19840 318565 19845 318595
rect 19875 318565 19880 318595
rect 19840 318560 19880 318565
rect 19680 318515 19720 318520
rect 19680 318485 19685 318515
rect 19715 318485 19720 318515
rect 19680 318480 19720 318485
rect 19840 318515 19880 318520
rect 19840 318485 19845 318515
rect 19875 318485 19880 318515
rect 19840 318480 19880 318485
rect 19680 318435 19720 318440
rect 19680 318405 19685 318435
rect 19715 318405 19720 318435
rect 19680 318400 19720 318405
rect 19840 318435 19880 318440
rect 19840 318405 19845 318435
rect 19875 318405 19880 318435
rect 19840 318400 19880 318405
rect 19680 318355 19720 318360
rect 19680 318325 19685 318355
rect 19715 318325 19720 318355
rect 19680 318320 19720 318325
rect 19840 318355 19880 318360
rect 19840 318325 19845 318355
rect 19875 318325 19880 318355
rect 19840 318320 19880 318325
rect 19680 318275 19720 318280
rect 19680 318245 19685 318275
rect 19715 318245 19720 318275
rect 19680 318240 19720 318245
rect 19840 318275 19880 318280
rect 19840 318245 19845 318275
rect 19875 318245 19880 318275
rect 19840 318240 19880 318245
rect 19680 318195 19720 318200
rect 19680 318165 19685 318195
rect 19715 318165 19720 318195
rect 19680 318160 19720 318165
rect 19840 318195 19880 318200
rect 19840 318165 19845 318195
rect 19875 318165 19880 318195
rect 19840 318160 19880 318165
rect 19680 318115 19720 318120
rect 19680 318085 19685 318115
rect 19715 318085 19720 318115
rect 19680 318080 19720 318085
rect 19840 318115 19880 318120
rect 19840 318085 19845 318115
rect 19875 318085 19880 318115
rect 19840 318080 19880 318085
rect 19680 318035 19720 318040
rect 19680 318005 19685 318035
rect 19715 318005 19720 318035
rect 19680 318000 19720 318005
rect 19840 318035 19880 318040
rect 19840 318005 19845 318035
rect 19875 318005 19880 318035
rect 19840 318000 19880 318005
rect 19680 317955 19720 317960
rect 19680 317925 19685 317955
rect 19715 317925 19720 317955
rect 19680 317920 19720 317925
rect 19840 317955 19880 317960
rect 19840 317925 19845 317955
rect 19875 317925 19880 317955
rect 19840 317920 19880 317925
rect 19680 317875 19720 317880
rect 19680 317845 19685 317875
rect 19715 317845 19720 317875
rect 19680 317840 19720 317845
rect 19840 317875 19880 317880
rect 19840 317845 19845 317875
rect 19875 317845 19880 317875
rect 19840 317840 19880 317845
rect 19680 317795 19720 317800
rect 19680 317765 19685 317795
rect 19715 317765 19720 317795
rect 19680 317760 19720 317765
rect 19840 317795 19880 317800
rect 19840 317765 19845 317795
rect 19875 317765 19880 317795
rect 19840 317760 19880 317765
rect 19680 317715 19720 317720
rect 19680 317685 19685 317715
rect 19715 317685 19720 317715
rect 19680 317680 19720 317685
rect 19840 317715 19880 317720
rect 19840 317685 19845 317715
rect 19875 317685 19880 317715
rect 19840 317680 19880 317685
rect 19680 317635 19720 317640
rect 19680 317605 19685 317635
rect 19715 317605 19720 317635
rect 19680 317600 19720 317605
rect 19840 317635 19880 317640
rect 19840 317605 19845 317635
rect 19875 317605 19880 317635
rect 19840 317600 19880 317605
rect 19680 317555 19720 317560
rect 19680 317525 19685 317555
rect 19715 317525 19720 317555
rect 19680 317520 19720 317525
rect 19840 317555 19880 317560
rect 19840 317525 19845 317555
rect 19875 317525 19880 317555
rect 19840 317520 19880 317525
rect 19680 317475 19720 317480
rect 19680 317445 19685 317475
rect 19715 317445 19720 317475
rect 19680 317440 19720 317445
rect 19840 317475 19880 317480
rect 19840 317445 19845 317475
rect 19875 317445 19880 317475
rect 19840 317440 19880 317445
rect 19680 317395 19720 317400
rect 19680 317365 19685 317395
rect 19715 317365 19720 317395
rect 19680 317360 19720 317365
rect 19840 317395 19880 317400
rect 19840 317365 19845 317395
rect 19875 317365 19880 317395
rect 19840 317360 19880 317365
rect 19680 317315 19720 317320
rect 19680 317285 19685 317315
rect 19715 317285 19720 317315
rect 19680 317280 19720 317285
rect 19840 317315 19880 317320
rect 19840 317285 19845 317315
rect 19875 317285 19880 317315
rect 19840 317280 19880 317285
rect 19680 317235 19720 317240
rect 19680 317205 19685 317235
rect 19715 317205 19720 317235
rect 19680 317200 19720 317205
rect 19840 317235 19880 317240
rect 19840 317205 19845 317235
rect 19875 317205 19880 317235
rect 19840 317200 19880 317205
rect 19680 317155 19720 317160
rect 19680 317125 19685 317155
rect 19715 317125 19720 317155
rect 19680 317120 19720 317125
rect 19840 317155 19880 317160
rect 19840 317125 19845 317155
rect 19875 317125 19880 317155
rect 19840 317120 19880 317125
rect 19680 317075 19720 317080
rect 19680 317045 19685 317075
rect 19715 317045 19720 317075
rect 19680 317040 19720 317045
rect 19840 317075 19880 317080
rect 19840 317045 19845 317075
rect 19875 317045 19880 317075
rect 19840 317040 19880 317045
rect 19680 316995 19720 317000
rect 19680 316965 19685 316995
rect 19715 316965 19720 316995
rect 19680 316960 19720 316965
rect 19840 316995 19880 317000
rect 19840 316965 19845 316995
rect 19875 316965 19880 316995
rect 19840 316960 19880 316965
rect 19680 316915 19720 316920
rect 19680 316885 19685 316915
rect 19715 316885 19720 316915
rect 19680 316880 19720 316885
rect 19840 316915 19880 316920
rect 19840 316885 19845 316915
rect 19875 316885 19880 316915
rect 19840 316880 19880 316885
rect 19680 316835 19720 316840
rect 19680 316805 19685 316835
rect 19715 316805 19720 316835
rect 19680 316800 19720 316805
rect 19840 316835 19880 316840
rect 19840 316805 19845 316835
rect 19875 316805 19880 316835
rect 19840 316800 19880 316805
rect 19680 316755 19720 316760
rect 19680 316725 19685 316755
rect 19715 316725 19720 316755
rect 19680 316720 19720 316725
rect 19840 316755 19880 316760
rect 19840 316725 19845 316755
rect 19875 316725 19880 316755
rect 19840 316720 19880 316725
rect 19680 316675 19720 316680
rect 19680 316645 19685 316675
rect 19715 316645 19720 316675
rect 19680 316640 19720 316645
rect 19840 316675 19880 316680
rect 19840 316645 19845 316675
rect 19875 316645 19880 316675
rect 19840 316640 19880 316645
rect 19680 316595 19720 316600
rect 19680 316565 19685 316595
rect 19715 316565 19720 316595
rect 19680 316560 19720 316565
rect 19840 316595 19880 316600
rect 19840 316565 19845 316595
rect 19875 316565 19880 316595
rect 19840 316560 19880 316565
rect 19680 316515 19720 316520
rect 19680 316485 19685 316515
rect 19715 316485 19720 316515
rect 19680 316480 19720 316485
rect 19840 316515 19880 316520
rect 19840 316485 19845 316515
rect 19875 316485 19880 316515
rect 19840 316480 19880 316485
rect 19680 316435 19720 316440
rect 19680 316405 19685 316435
rect 19715 316405 19720 316435
rect 19680 316400 19720 316405
rect 19840 316435 19880 316440
rect 19840 316405 19845 316435
rect 19875 316405 19880 316435
rect 19840 316400 19880 316405
rect 19680 316355 19720 316360
rect 19680 316325 19685 316355
rect 19715 316325 19720 316355
rect 19680 316320 19720 316325
rect 19840 316355 19880 316360
rect 19840 316325 19845 316355
rect 19875 316325 19880 316355
rect 19840 316320 19880 316325
rect 19680 316275 19720 316280
rect 19680 316245 19685 316275
rect 19715 316245 19720 316275
rect 19680 316240 19720 316245
rect 19840 316275 19880 316280
rect 19840 316245 19845 316275
rect 19875 316245 19880 316275
rect 19840 316240 19880 316245
rect 19680 316195 19720 316200
rect 19680 316165 19685 316195
rect 19715 316165 19720 316195
rect 19680 316160 19720 316165
rect 19840 316195 19880 316200
rect 19840 316165 19845 316195
rect 19875 316165 19880 316195
rect 19840 316160 19880 316165
rect 19680 316115 19720 316120
rect 19680 316085 19685 316115
rect 19715 316085 19720 316115
rect 19680 316080 19720 316085
rect 19840 316115 19880 316120
rect 19840 316085 19845 316115
rect 19875 316085 19880 316115
rect 19840 316080 19880 316085
rect 19680 316035 19720 316040
rect 19680 316005 19685 316035
rect 19715 316005 19720 316035
rect 19680 316000 19720 316005
rect 19840 316035 19880 316040
rect 19840 316005 19845 316035
rect 19875 316005 19880 316035
rect 19840 316000 19880 316005
rect 19680 315955 19720 315960
rect 19680 315925 19685 315955
rect 19715 315925 19720 315955
rect 19680 315920 19720 315925
rect 19840 315955 19880 315960
rect 19840 315925 19845 315955
rect 19875 315925 19880 315955
rect 19840 315920 19880 315925
rect 19680 315875 19720 315880
rect 19680 315845 19685 315875
rect 19715 315845 19720 315875
rect 19680 315840 19720 315845
rect 19840 315875 19880 315880
rect 19840 315845 19845 315875
rect 19875 315845 19880 315875
rect 19840 315840 19880 315845
rect 19680 315795 19720 315800
rect 19680 315765 19685 315795
rect 19715 315765 19720 315795
rect 19680 315760 19720 315765
rect 19840 315795 19880 315800
rect 19840 315765 19845 315795
rect 19875 315765 19880 315795
rect 19840 315760 19880 315765
rect 19680 315715 19720 315720
rect 19680 315685 19685 315715
rect 19715 315685 19720 315715
rect 19680 315680 19720 315685
rect 19840 315715 19880 315720
rect 19840 315685 19845 315715
rect 19875 315685 19880 315715
rect 19840 315680 19880 315685
rect 19680 315635 19720 315640
rect 19680 315605 19685 315635
rect 19715 315605 19720 315635
rect 19680 315600 19720 315605
rect 19840 315635 19880 315640
rect 19840 315605 19845 315635
rect 19875 315605 19880 315635
rect 19840 315600 19880 315605
rect 19680 315555 19720 315560
rect 19680 315525 19685 315555
rect 19715 315525 19720 315555
rect 19680 315520 19720 315525
rect 19840 315555 19880 315560
rect 19840 315525 19845 315555
rect 19875 315525 19880 315555
rect 19840 315520 19880 315525
rect 19680 315475 19720 315480
rect 19680 315445 19685 315475
rect 19715 315445 19720 315475
rect 19680 315440 19720 315445
rect 19840 315475 19880 315480
rect 19840 315445 19845 315475
rect 19875 315445 19880 315475
rect 19840 315440 19880 315445
rect 19680 315395 19720 315400
rect 19680 315365 19685 315395
rect 19715 315365 19720 315395
rect 19680 315360 19720 315365
rect 19840 315395 19880 315400
rect 19840 315365 19845 315395
rect 19875 315365 19880 315395
rect 19840 315360 19880 315365
rect 19680 315315 19720 315320
rect 19680 315285 19685 315315
rect 19715 315285 19720 315315
rect 19680 315280 19720 315285
rect 19840 315315 19880 315320
rect 19840 315285 19845 315315
rect 19875 315285 19880 315315
rect 19840 315280 19880 315285
rect 19680 315235 19720 315240
rect 19680 315205 19685 315235
rect 19715 315205 19720 315235
rect 19680 315200 19720 315205
rect 19840 315235 19880 315240
rect 19840 315205 19845 315235
rect 19875 315205 19880 315235
rect 19840 315200 19880 315205
rect 19680 315155 19720 315160
rect 19680 315125 19685 315155
rect 19715 315125 19720 315155
rect 19680 315120 19720 315125
rect 19840 315155 19880 315160
rect 19840 315125 19845 315155
rect 19875 315125 19880 315155
rect 19840 315120 19880 315125
rect 19680 315075 19720 315080
rect 19680 315045 19685 315075
rect 19715 315045 19720 315075
rect 19680 315040 19720 315045
rect 19840 315075 19880 315080
rect 19840 315045 19845 315075
rect 19875 315045 19880 315075
rect 19840 315040 19880 315045
rect 19680 314995 19720 315000
rect 19680 314965 19685 314995
rect 19715 314965 19720 314995
rect 19680 314960 19720 314965
rect 19840 314995 19880 315000
rect 19840 314965 19845 314995
rect 19875 314965 19880 314995
rect 19840 314960 19880 314965
rect 19680 314915 19720 314920
rect 19680 314885 19685 314915
rect 19715 314885 19720 314915
rect 19680 314880 19720 314885
rect 19840 314915 19880 314920
rect 19840 314885 19845 314915
rect 19875 314885 19880 314915
rect 19840 314880 19880 314885
rect 19680 314835 19720 314840
rect 19680 314805 19685 314835
rect 19715 314805 19720 314835
rect 19680 314800 19720 314805
rect 19840 314835 19880 314840
rect 19840 314805 19845 314835
rect 19875 314805 19880 314835
rect 19840 314800 19880 314805
rect 19680 314755 19720 314760
rect 19680 314725 19685 314755
rect 19715 314725 19720 314755
rect 19680 314720 19720 314725
rect 19840 314755 19880 314760
rect 19840 314725 19845 314755
rect 19875 314725 19880 314755
rect 19840 314720 19880 314725
rect 19680 314675 19720 314680
rect 19680 314645 19685 314675
rect 19715 314645 19720 314675
rect 19680 314640 19720 314645
rect 19840 314675 19880 314680
rect 19840 314645 19845 314675
rect 19875 314645 19880 314675
rect 19840 314640 19880 314645
rect 19680 314595 19720 314600
rect 19680 314565 19685 314595
rect 19715 314565 19720 314595
rect 19680 314560 19720 314565
rect 19840 314595 19880 314600
rect 19840 314565 19845 314595
rect 19875 314565 19880 314595
rect 19840 314560 19880 314565
rect 19680 314515 19720 314520
rect 19680 314485 19685 314515
rect 19715 314485 19720 314515
rect 19680 314480 19720 314485
rect 19840 314515 19880 314520
rect 19840 314485 19845 314515
rect 19875 314485 19880 314515
rect 19840 314480 19880 314485
rect 19680 314435 19720 314440
rect 19680 314405 19685 314435
rect 19715 314405 19720 314435
rect 19680 314400 19720 314405
rect 19840 314435 19880 314440
rect 19840 314405 19845 314435
rect 19875 314405 19880 314435
rect 19840 314400 19880 314405
rect 19680 314355 19720 314360
rect 19680 314325 19685 314355
rect 19715 314325 19720 314355
rect 19680 314320 19720 314325
rect 19840 314355 19880 314360
rect 19840 314325 19845 314355
rect 19875 314325 19880 314355
rect 19840 314320 19880 314325
rect 19680 314275 19720 314280
rect 19680 314245 19685 314275
rect 19715 314245 19720 314275
rect 19680 314240 19720 314245
rect 19840 314275 19880 314280
rect 19840 314245 19845 314275
rect 19875 314245 19880 314275
rect 19840 314240 19880 314245
rect 19680 314195 19720 314200
rect 19680 314165 19685 314195
rect 19715 314165 19720 314195
rect 19680 314160 19720 314165
rect 19840 314195 19880 314200
rect 19840 314165 19845 314195
rect 19875 314165 19880 314195
rect 19840 314160 19880 314165
rect 19680 314115 19720 314120
rect 19680 314085 19685 314115
rect 19715 314085 19720 314115
rect 19680 314080 19720 314085
rect 19840 314115 19880 314120
rect 19840 314085 19845 314115
rect 19875 314085 19880 314115
rect 19840 314080 19880 314085
rect 19680 314035 19720 314040
rect 19680 314005 19685 314035
rect 19715 314005 19720 314035
rect 19680 314000 19720 314005
rect 19840 314035 19880 314040
rect 19840 314005 19845 314035
rect 19875 314005 19880 314035
rect 19840 314000 19880 314005
rect 19680 313955 19720 313960
rect 19680 313925 19685 313955
rect 19715 313925 19720 313955
rect 19680 313920 19720 313925
rect 19840 313955 19880 313960
rect 19840 313925 19845 313955
rect 19875 313925 19880 313955
rect 19840 313920 19880 313925
rect 19680 313875 19720 313880
rect 19680 313845 19685 313875
rect 19715 313845 19720 313875
rect 19680 313840 19720 313845
rect 19840 313875 19880 313880
rect 19840 313845 19845 313875
rect 19875 313845 19880 313875
rect 19840 313840 19880 313845
rect 19680 313795 19720 313800
rect 19680 313765 19685 313795
rect 19715 313765 19720 313795
rect 19680 313760 19720 313765
rect 19840 313795 19880 313800
rect 19840 313765 19845 313795
rect 19875 313765 19880 313795
rect 19840 313760 19880 313765
rect 19680 313715 19720 313720
rect 19680 313685 19685 313715
rect 19715 313685 19720 313715
rect 19680 313680 19720 313685
rect 19840 313715 19880 313720
rect 19840 313685 19845 313715
rect 19875 313685 19880 313715
rect 19840 313680 19880 313685
rect 19680 313635 19720 313640
rect 19680 313605 19685 313635
rect 19715 313605 19720 313635
rect 19680 313600 19720 313605
rect 19840 313635 19880 313640
rect 19840 313605 19845 313635
rect 19875 313605 19880 313635
rect 19840 313600 19880 313605
rect 19680 313555 19720 313560
rect 19680 313525 19685 313555
rect 19715 313525 19720 313555
rect 19680 313520 19720 313525
rect 19840 313555 19880 313560
rect 19840 313525 19845 313555
rect 19875 313525 19880 313555
rect 19840 313520 19880 313525
rect 19680 313475 19720 313480
rect 19680 313445 19685 313475
rect 19715 313445 19720 313475
rect 19680 313440 19720 313445
rect 19840 313475 19880 313480
rect 19840 313445 19845 313475
rect 19875 313445 19880 313475
rect 19840 313440 19880 313445
rect 19680 313395 19720 313400
rect 19680 313365 19685 313395
rect 19715 313365 19720 313395
rect 19680 313360 19720 313365
rect 19840 313395 19880 313400
rect 19840 313365 19845 313395
rect 19875 313365 19880 313395
rect 19840 313360 19880 313365
rect 19680 313315 19720 313320
rect 19680 313285 19685 313315
rect 19715 313285 19720 313315
rect 19680 313280 19720 313285
rect 19840 313315 19880 313320
rect 19840 313285 19845 313315
rect 19875 313285 19880 313315
rect 19840 313280 19880 313285
rect 19680 313235 19720 313240
rect 19680 313205 19685 313235
rect 19715 313205 19720 313235
rect 19680 313200 19720 313205
rect 19840 313235 19880 313240
rect 19840 313205 19845 313235
rect 19875 313205 19880 313235
rect 19840 313200 19880 313205
rect 19680 313155 19720 313160
rect 19680 313125 19685 313155
rect 19715 313125 19720 313155
rect 19680 313120 19720 313125
rect 19840 313155 19880 313160
rect 19840 313125 19845 313155
rect 19875 313125 19880 313155
rect 19840 313120 19880 313125
rect 19680 313075 19720 313080
rect 19680 313045 19685 313075
rect 19715 313045 19720 313075
rect 19680 313040 19720 313045
rect 19840 313075 19880 313080
rect 19840 313045 19845 313075
rect 19875 313045 19880 313075
rect 19840 313040 19880 313045
rect 19680 312995 19720 313000
rect 19680 312965 19685 312995
rect 19715 312965 19720 312995
rect 19680 312960 19720 312965
rect 19840 312995 19880 313000
rect 19840 312965 19845 312995
rect 19875 312965 19880 312995
rect 19840 312960 19880 312965
rect 19680 312915 19720 312920
rect 19680 312885 19685 312915
rect 19715 312885 19720 312915
rect 19680 312880 19720 312885
rect 19840 312915 19880 312920
rect 19840 312885 19845 312915
rect 19875 312885 19880 312915
rect 19840 312880 19880 312885
rect 19680 312835 19720 312840
rect 19680 312805 19685 312835
rect 19715 312805 19720 312835
rect 19680 312800 19720 312805
rect 19840 312835 19880 312840
rect 19840 312805 19845 312835
rect 19875 312805 19880 312835
rect 19840 312800 19880 312805
rect 19680 312755 19720 312760
rect 19680 312725 19685 312755
rect 19715 312725 19720 312755
rect 19680 312720 19720 312725
rect 19840 312755 19880 312760
rect 19840 312725 19845 312755
rect 19875 312725 19880 312755
rect 19840 312720 19880 312725
rect 19680 312675 19720 312680
rect 19680 312645 19685 312675
rect 19715 312645 19720 312675
rect 19680 312640 19720 312645
rect 19840 312675 19880 312680
rect 19840 312645 19845 312675
rect 19875 312645 19880 312675
rect 19840 312640 19880 312645
rect 19680 312595 19720 312600
rect 19680 312565 19685 312595
rect 19715 312565 19720 312595
rect 19680 312560 19720 312565
rect 19840 312595 19880 312600
rect 19840 312565 19845 312595
rect 19875 312565 19880 312595
rect 19840 312560 19880 312565
rect 19680 312515 19720 312520
rect 19680 312485 19685 312515
rect 19715 312485 19720 312515
rect 19680 312480 19720 312485
rect 19840 312515 19880 312520
rect 19840 312485 19845 312515
rect 19875 312485 19880 312515
rect 19840 312480 19880 312485
rect 19680 312435 19720 312440
rect 19680 312405 19685 312435
rect 19715 312405 19720 312435
rect 19680 312400 19720 312405
rect 19840 312435 19880 312440
rect 19840 312405 19845 312435
rect 19875 312405 19880 312435
rect 19840 312400 19880 312405
rect 19680 312355 19720 312360
rect 19680 312325 19685 312355
rect 19715 312325 19720 312355
rect 19680 312320 19720 312325
rect 19840 312355 19880 312360
rect 19840 312325 19845 312355
rect 19875 312325 19880 312355
rect 19840 312320 19880 312325
rect 19680 312275 19720 312280
rect 19680 312245 19685 312275
rect 19715 312245 19720 312275
rect 19680 312240 19720 312245
rect 19840 312275 19880 312280
rect 19840 312245 19845 312275
rect 19875 312245 19880 312275
rect 19840 312240 19880 312245
rect 19680 312195 19720 312200
rect 19680 312165 19685 312195
rect 19715 312165 19720 312195
rect 19680 312160 19720 312165
rect 19840 312195 19880 312200
rect 19840 312165 19845 312195
rect 19875 312165 19880 312195
rect 19840 312160 19880 312165
rect 19680 312115 19720 312120
rect 19680 312085 19685 312115
rect 19715 312085 19720 312115
rect 19680 312080 19720 312085
rect 19840 312115 19880 312120
rect 19840 312085 19845 312115
rect 19875 312085 19880 312115
rect 19840 312080 19880 312085
rect 19680 312035 19720 312040
rect 19680 312005 19685 312035
rect 19715 312005 19720 312035
rect 19680 312000 19720 312005
rect 19840 312035 19880 312040
rect 19840 312005 19845 312035
rect 19875 312005 19880 312035
rect 19840 312000 19880 312005
rect 19680 311955 19720 311960
rect 19680 311925 19685 311955
rect 19715 311925 19720 311955
rect 19680 311920 19720 311925
rect 19840 311955 19880 311960
rect 19840 311925 19845 311955
rect 19875 311925 19880 311955
rect 19840 311920 19880 311925
rect 19680 311875 19720 311880
rect 19680 311845 19685 311875
rect 19715 311845 19720 311875
rect 19680 311840 19720 311845
rect 19840 311875 19880 311880
rect 19840 311845 19845 311875
rect 19875 311845 19880 311875
rect 19840 311840 19880 311845
rect 19680 311795 19720 311800
rect 19680 311765 19685 311795
rect 19715 311765 19720 311795
rect 19680 311760 19720 311765
rect 19840 311795 19880 311800
rect 19840 311765 19845 311795
rect 19875 311765 19880 311795
rect 19840 311760 19880 311765
rect 19680 311715 19720 311720
rect 19680 311685 19685 311715
rect 19715 311685 19720 311715
rect 19680 311680 19720 311685
rect 19840 311715 19880 311720
rect 19840 311685 19845 311715
rect 19875 311685 19880 311715
rect 19840 311680 19880 311685
rect 19680 311635 19720 311640
rect 19680 311605 19685 311635
rect 19715 311605 19720 311635
rect 19680 311600 19720 311605
rect 19840 311635 19880 311640
rect 19840 311605 19845 311635
rect 19875 311605 19880 311635
rect 19840 311600 19880 311605
rect 19680 311555 19720 311560
rect 19680 311525 19685 311555
rect 19715 311525 19720 311555
rect 19680 311520 19720 311525
rect 19840 311555 19880 311560
rect 19840 311525 19845 311555
rect 19875 311525 19880 311555
rect 19840 311520 19880 311525
rect 19680 311475 19720 311480
rect 19680 311445 19685 311475
rect 19715 311445 19720 311475
rect 19680 311440 19720 311445
rect 19840 311475 19880 311480
rect 19840 311445 19845 311475
rect 19875 311445 19880 311475
rect 19840 311440 19880 311445
rect 19680 311395 19720 311400
rect 19680 311365 19685 311395
rect 19715 311365 19720 311395
rect 19680 311360 19720 311365
rect 19840 311395 19880 311400
rect 19840 311365 19845 311395
rect 19875 311365 19880 311395
rect 19840 311360 19880 311365
rect 19680 311315 19720 311320
rect 19680 311285 19685 311315
rect 19715 311285 19720 311315
rect 19680 311280 19720 311285
rect 19840 311315 19880 311320
rect 19840 311285 19845 311315
rect 19875 311285 19880 311315
rect 19840 311280 19880 311285
rect 19680 311235 19720 311240
rect 19680 311205 19685 311235
rect 19715 311205 19720 311235
rect 19680 311200 19720 311205
rect 19840 311235 19880 311240
rect 19840 311205 19845 311235
rect 19875 311205 19880 311235
rect 19840 311200 19880 311205
rect 19680 311155 19720 311160
rect 19680 311125 19685 311155
rect 19715 311125 19720 311155
rect 19680 311120 19720 311125
rect 19840 311155 19880 311160
rect 19840 311125 19845 311155
rect 19875 311125 19880 311155
rect 19840 311120 19880 311125
rect 19680 311075 19720 311080
rect 19680 311045 19685 311075
rect 19715 311045 19720 311075
rect 19680 311040 19720 311045
rect 19840 311075 19880 311080
rect 19840 311045 19845 311075
rect 19875 311045 19880 311075
rect 19840 311040 19880 311045
rect 19680 310995 19720 311000
rect 19680 310965 19685 310995
rect 19715 310965 19720 310995
rect 19680 310960 19720 310965
rect 19840 310995 19880 311000
rect 19840 310965 19845 310995
rect 19875 310965 19880 310995
rect 19840 310960 19880 310965
rect 19680 310915 19720 310920
rect 19680 310885 19685 310915
rect 19715 310885 19720 310915
rect 19680 310880 19720 310885
rect 19840 310915 19880 310920
rect 19840 310885 19845 310915
rect 19875 310885 19880 310915
rect 19840 310880 19880 310885
rect 19680 310835 19720 310840
rect 19680 310805 19685 310835
rect 19715 310805 19720 310835
rect 19680 310800 19720 310805
rect 19840 310835 19880 310840
rect 19840 310805 19845 310835
rect 19875 310805 19880 310835
rect 19840 310800 19880 310805
rect 19680 310755 19720 310760
rect 19680 310725 19685 310755
rect 19715 310725 19720 310755
rect 19680 310720 19720 310725
rect 19840 310755 19880 310760
rect 19840 310725 19845 310755
rect 19875 310725 19880 310755
rect 19840 310720 19880 310725
rect 19680 310675 19720 310680
rect 19680 310645 19685 310675
rect 19715 310645 19720 310675
rect 19680 310640 19720 310645
rect 19840 310675 19880 310680
rect 19840 310645 19845 310675
rect 19875 310645 19880 310675
rect 19840 310640 19880 310645
rect 19680 310595 19720 310600
rect 19680 310565 19685 310595
rect 19715 310565 19720 310595
rect 19680 310560 19720 310565
rect 19840 310595 19880 310600
rect 19840 310565 19845 310595
rect 19875 310565 19880 310595
rect 19840 310560 19880 310565
rect 19680 310515 19720 310520
rect 19680 310485 19685 310515
rect 19715 310485 19720 310515
rect 19680 310480 19720 310485
rect 19840 310515 19880 310520
rect 19840 310485 19845 310515
rect 19875 310485 19880 310515
rect 19840 310480 19880 310485
rect 19680 310435 19720 310440
rect 19680 310405 19685 310435
rect 19715 310405 19720 310435
rect 19680 310400 19720 310405
rect 19840 310435 19880 310440
rect 19840 310405 19845 310435
rect 19875 310405 19880 310435
rect 19840 310400 19880 310405
rect 19680 310355 19720 310360
rect 19680 310325 19685 310355
rect 19715 310325 19720 310355
rect 19680 310320 19720 310325
rect 19840 310355 19880 310360
rect 19840 310325 19845 310355
rect 19875 310325 19880 310355
rect 19840 310320 19880 310325
rect 19680 310275 19720 310280
rect 19680 310245 19685 310275
rect 19715 310245 19720 310275
rect 19680 310240 19720 310245
rect 19840 310275 19880 310280
rect 19840 310245 19845 310275
rect 19875 310245 19880 310275
rect 19840 310240 19880 310245
rect 19680 310195 19720 310200
rect 19680 310165 19685 310195
rect 19715 310165 19720 310195
rect 19680 310160 19720 310165
rect 19840 310195 19880 310200
rect 19840 310165 19845 310195
rect 19875 310165 19880 310195
rect 19840 310160 19880 310165
rect 19680 310115 19720 310120
rect 19680 310085 19685 310115
rect 19715 310085 19720 310115
rect 19680 310080 19720 310085
rect 19840 310115 19880 310120
rect 19840 310085 19845 310115
rect 19875 310085 19880 310115
rect 19840 310080 19880 310085
rect 19680 310035 19720 310040
rect 19680 310005 19685 310035
rect 19715 310005 19720 310035
rect 19680 310000 19720 310005
rect 19840 310035 19880 310040
rect 19840 310005 19845 310035
rect 19875 310005 19880 310035
rect 19840 310000 19880 310005
rect 19680 309955 19720 309960
rect 19680 309925 19685 309955
rect 19715 309925 19720 309955
rect 19680 309920 19720 309925
rect 19840 309955 19880 309960
rect 19840 309925 19845 309955
rect 19875 309925 19880 309955
rect 19840 309920 19880 309925
rect 19680 309875 19720 309880
rect 19680 309845 19685 309875
rect 19715 309845 19720 309875
rect 19680 309840 19720 309845
rect 19840 309875 19880 309880
rect 19840 309845 19845 309875
rect 19875 309845 19880 309875
rect 19840 309840 19880 309845
rect 19680 309795 19720 309800
rect 19680 309765 19685 309795
rect 19715 309765 19720 309795
rect 19680 309760 19720 309765
rect 19840 309795 19880 309800
rect 19840 309765 19845 309795
rect 19875 309765 19880 309795
rect 19840 309760 19880 309765
rect 19680 309715 19720 309720
rect 19680 309685 19685 309715
rect 19715 309685 19720 309715
rect 19680 309680 19720 309685
rect 19840 309715 19880 309720
rect 19840 309685 19845 309715
rect 19875 309685 19880 309715
rect 19840 309680 19880 309685
rect 19680 309635 19720 309640
rect 19680 309605 19685 309635
rect 19715 309605 19720 309635
rect 19680 309600 19720 309605
rect 19840 309635 19880 309640
rect 19840 309605 19845 309635
rect 19875 309605 19880 309635
rect 19840 309600 19880 309605
rect 19680 309555 19720 309560
rect 19680 309525 19685 309555
rect 19715 309525 19720 309555
rect 19680 309520 19720 309525
rect 19840 309555 19880 309560
rect 19840 309525 19845 309555
rect 19875 309525 19880 309555
rect 19840 309520 19880 309525
rect 19680 309475 19720 309480
rect 19680 309445 19685 309475
rect 19715 309445 19720 309475
rect 19680 309440 19720 309445
rect 19840 309475 19880 309480
rect 19840 309445 19845 309475
rect 19875 309445 19880 309475
rect 19840 309440 19880 309445
rect 19680 309395 19720 309400
rect 19680 309365 19685 309395
rect 19715 309365 19720 309395
rect 19680 309360 19720 309365
rect 19840 309395 19880 309400
rect 19840 309365 19845 309395
rect 19875 309365 19880 309395
rect 19840 309360 19880 309365
rect 19680 309315 19720 309320
rect 19680 309285 19685 309315
rect 19715 309285 19720 309315
rect 19680 309280 19720 309285
rect 19840 309315 19880 309320
rect 19840 309285 19845 309315
rect 19875 309285 19880 309315
rect 19840 309280 19880 309285
rect 19680 309235 19720 309240
rect 19680 309205 19685 309235
rect 19715 309205 19720 309235
rect 19680 309200 19720 309205
rect 19840 309235 19880 309240
rect 19840 309205 19845 309235
rect 19875 309205 19880 309235
rect 19840 309200 19880 309205
rect 19680 309155 19720 309160
rect 19680 309125 19685 309155
rect 19715 309125 19720 309155
rect 19680 309120 19720 309125
rect 19840 309155 19880 309160
rect 19840 309125 19845 309155
rect 19875 309125 19880 309155
rect 19840 309120 19880 309125
rect 19680 309075 19720 309080
rect 19680 309045 19685 309075
rect 19715 309045 19720 309075
rect 19680 309040 19720 309045
rect 19840 309075 19880 309080
rect 19840 309045 19845 309075
rect 19875 309045 19880 309075
rect 19840 309040 19880 309045
rect 19680 308995 19720 309000
rect 19680 308965 19685 308995
rect 19715 308965 19720 308995
rect 19680 308960 19720 308965
rect 19840 308995 19880 309000
rect 19840 308965 19845 308995
rect 19875 308965 19880 308995
rect 19840 308960 19880 308965
rect 19680 308915 19720 308920
rect 19680 308885 19685 308915
rect 19715 308885 19720 308915
rect 19680 308880 19720 308885
rect 19840 308915 19880 308920
rect 19840 308885 19845 308915
rect 19875 308885 19880 308915
rect 19840 308880 19880 308885
rect 19680 308835 19720 308840
rect 19680 308805 19685 308835
rect 19715 308805 19720 308835
rect 19680 308800 19720 308805
rect 19840 308835 19880 308840
rect 19840 308805 19845 308835
rect 19875 308805 19880 308835
rect 19840 308800 19880 308805
rect 19680 308755 19720 308760
rect 19680 308725 19685 308755
rect 19715 308725 19720 308755
rect 19680 308720 19720 308725
rect 19840 308755 19880 308760
rect 19840 308725 19845 308755
rect 19875 308725 19880 308755
rect 19840 308720 19880 308725
rect 19680 308675 19720 308680
rect 19680 308645 19685 308675
rect 19715 308645 19720 308675
rect 19680 308640 19720 308645
rect 19840 308675 19880 308680
rect 19840 308645 19845 308675
rect 19875 308645 19880 308675
rect 19840 308640 19880 308645
rect 19680 308595 19720 308600
rect 19680 308565 19685 308595
rect 19715 308565 19720 308595
rect 19680 308560 19720 308565
rect 19840 308595 19880 308600
rect 19840 308565 19845 308595
rect 19875 308565 19880 308595
rect 19840 308560 19880 308565
rect 19680 308515 19720 308520
rect 19680 308485 19685 308515
rect 19715 308485 19720 308515
rect 19680 308480 19720 308485
rect 19840 308515 19880 308520
rect 19840 308485 19845 308515
rect 19875 308485 19880 308515
rect 19840 308480 19880 308485
rect 19680 308435 19720 308440
rect 19680 308405 19685 308435
rect 19715 308405 19720 308435
rect 19680 308400 19720 308405
rect 19840 308435 19880 308440
rect 19840 308405 19845 308435
rect 19875 308405 19880 308435
rect 19840 308400 19880 308405
rect 19680 308355 19720 308360
rect 19680 308325 19685 308355
rect 19715 308325 19720 308355
rect 19680 308320 19720 308325
rect 19840 308355 19880 308360
rect 19840 308325 19845 308355
rect 19875 308325 19880 308355
rect 19840 308320 19880 308325
rect 19680 308275 19720 308280
rect 19680 308245 19685 308275
rect 19715 308245 19720 308275
rect 19680 308240 19720 308245
rect 19840 308275 19880 308280
rect 19840 308245 19845 308275
rect 19875 308245 19880 308275
rect 19840 308240 19880 308245
rect 19680 308195 19720 308200
rect 19680 308165 19685 308195
rect 19715 308165 19720 308195
rect 19680 308160 19720 308165
rect 19840 308195 19880 308200
rect 19840 308165 19845 308195
rect 19875 308165 19880 308195
rect 19840 308160 19880 308165
rect 19680 308115 19720 308120
rect 19680 308085 19685 308115
rect 19715 308085 19720 308115
rect 19680 308080 19720 308085
rect 19840 308115 19880 308120
rect 19840 308085 19845 308115
rect 19875 308085 19880 308115
rect 19840 308080 19880 308085
rect 19680 308035 19720 308040
rect 19680 308005 19685 308035
rect 19715 308005 19720 308035
rect 19680 308000 19720 308005
rect 19840 308035 19880 308040
rect 19840 308005 19845 308035
rect 19875 308005 19880 308035
rect 19840 308000 19880 308005
rect 19680 307955 19720 307960
rect 19680 307925 19685 307955
rect 19715 307925 19720 307955
rect 19680 307920 19720 307925
rect 19840 307955 19880 307960
rect 19840 307925 19845 307955
rect 19875 307925 19880 307955
rect 19840 307920 19880 307925
rect 19680 307875 19720 307880
rect 19680 307845 19685 307875
rect 19715 307845 19720 307875
rect 19680 307840 19720 307845
rect 19840 307875 19880 307880
rect 19840 307845 19845 307875
rect 19875 307845 19880 307875
rect 19840 307840 19880 307845
rect 19680 307795 19720 307800
rect 19680 307765 19685 307795
rect 19715 307765 19720 307795
rect 19680 307760 19720 307765
rect 19840 307795 19880 307800
rect 19840 307765 19845 307795
rect 19875 307765 19880 307795
rect 19840 307760 19880 307765
rect 19680 307715 19720 307720
rect 19680 307685 19685 307715
rect 19715 307685 19720 307715
rect 19680 307680 19720 307685
rect 19840 307715 19880 307720
rect 19840 307685 19845 307715
rect 19875 307685 19880 307715
rect 19840 307680 19880 307685
rect 19680 307635 19720 307640
rect 19680 307605 19685 307635
rect 19715 307605 19720 307635
rect 19680 307600 19720 307605
rect 19840 307635 19880 307640
rect 19840 307605 19845 307635
rect 19875 307605 19880 307635
rect 19840 307600 19880 307605
rect 19680 307555 19720 307560
rect 19680 307525 19685 307555
rect 19715 307525 19720 307555
rect 19680 307520 19720 307525
rect 19840 307555 19880 307560
rect 19840 307525 19845 307555
rect 19875 307525 19880 307555
rect 19840 307520 19880 307525
rect 19680 307475 19720 307480
rect 19680 307445 19685 307475
rect 19715 307445 19720 307475
rect 19680 307440 19720 307445
rect 19840 307475 19880 307480
rect 19840 307445 19845 307475
rect 19875 307445 19880 307475
rect 19840 307440 19880 307445
rect 19680 307395 19720 307400
rect 19680 307365 19685 307395
rect 19715 307365 19720 307395
rect 19680 307360 19720 307365
rect 19840 307395 19880 307400
rect 19840 307365 19845 307395
rect 19875 307365 19880 307395
rect 19840 307360 19880 307365
rect 19680 307315 19720 307320
rect 19680 307285 19685 307315
rect 19715 307285 19720 307315
rect 19680 307280 19720 307285
rect 19840 307315 19880 307320
rect 19840 307285 19845 307315
rect 19875 307285 19880 307315
rect 19840 307280 19880 307285
rect 19680 307235 19720 307240
rect 19680 307205 19685 307235
rect 19715 307205 19720 307235
rect 19680 307200 19720 307205
rect 19840 307235 19880 307240
rect 19840 307205 19845 307235
rect 19875 307205 19880 307235
rect 19840 307200 19880 307205
rect 19680 307155 19720 307160
rect 19680 307125 19685 307155
rect 19715 307125 19720 307155
rect 19680 307120 19720 307125
rect 19840 307155 19880 307160
rect 19840 307125 19845 307155
rect 19875 307125 19880 307155
rect 19840 307120 19880 307125
rect 19680 307075 19720 307080
rect 19680 307045 19685 307075
rect 19715 307045 19720 307075
rect 19680 307040 19720 307045
rect 19840 307075 19880 307080
rect 19840 307045 19845 307075
rect 19875 307045 19880 307075
rect 19840 307040 19880 307045
rect 19680 306995 19720 307000
rect 19680 306965 19685 306995
rect 19715 306965 19720 306995
rect 19680 306960 19720 306965
rect 19840 306995 19880 307000
rect 19840 306965 19845 306995
rect 19875 306965 19880 306995
rect 19840 306960 19880 306965
rect 19680 306915 19720 306920
rect 19680 306885 19685 306915
rect 19715 306885 19720 306915
rect 19680 306880 19720 306885
rect 19840 306915 19880 306920
rect 19840 306885 19845 306915
rect 19875 306885 19880 306915
rect 19840 306880 19880 306885
rect 19680 306835 19720 306840
rect 19680 306805 19685 306835
rect 19715 306805 19720 306835
rect 19680 306800 19720 306805
rect 19840 306835 19880 306840
rect 19840 306805 19845 306835
rect 19875 306805 19880 306835
rect 19840 306800 19880 306805
rect 19680 306755 19720 306760
rect 19680 306725 19685 306755
rect 19715 306725 19720 306755
rect 19680 306720 19720 306725
rect 19840 306755 19880 306760
rect 19840 306725 19845 306755
rect 19875 306725 19880 306755
rect 19840 306720 19880 306725
rect 19680 306675 19720 306680
rect 19680 306645 19685 306675
rect 19715 306645 19720 306675
rect 19680 306640 19720 306645
rect 19840 306675 19880 306680
rect 19840 306645 19845 306675
rect 19875 306645 19880 306675
rect 19840 306640 19880 306645
rect 19680 306595 19720 306600
rect 19680 306565 19685 306595
rect 19715 306565 19720 306595
rect 19680 306560 19720 306565
rect 19840 306595 19880 306600
rect 19840 306565 19845 306595
rect 19875 306565 19880 306595
rect 19840 306560 19880 306565
rect 19680 306515 19720 306520
rect 19680 306485 19685 306515
rect 19715 306485 19720 306515
rect 19680 306480 19720 306485
rect 19840 306515 19880 306520
rect 19840 306485 19845 306515
rect 19875 306485 19880 306515
rect 19840 306480 19880 306485
rect 19680 306435 19720 306440
rect 19680 306405 19685 306435
rect 19715 306405 19720 306435
rect 19680 306400 19720 306405
rect 19840 306435 19880 306440
rect 19840 306405 19845 306435
rect 19875 306405 19880 306435
rect 19840 306400 19880 306405
rect 19680 306355 19720 306360
rect 19680 306325 19685 306355
rect 19715 306325 19720 306355
rect 19680 306320 19720 306325
rect 19840 306355 19880 306360
rect 19840 306325 19845 306355
rect 19875 306325 19880 306355
rect 19840 306320 19880 306325
rect 19680 306275 19720 306280
rect 19680 306245 19685 306275
rect 19715 306245 19720 306275
rect 19680 306240 19720 306245
rect 19840 306275 19880 306280
rect 19840 306245 19845 306275
rect 19875 306245 19880 306275
rect 19840 306240 19880 306245
rect 19680 306195 19720 306200
rect 19680 306165 19685 306195
rect 19715 306165 19720 306195
rect 19680 306160 19720 306165
rect 19840 306195 19880 306200
rect 19840 306165 19845 306195
rect 19875 306165 19880 306195
rect 19840 306160 19880 306165
rect 19680 306115 19720 306120
rect 19680 306085 19685 306115
rect 19715 306085 19720 306115
rect 19680 306080 19720 306085
rect 19840 306115 19880 306120
rect 19840 306085 19845 306115
rect 19875 306085 19880 306115
rect 19840 306080 19880 306085
rect 19680 306035 19720 306040
rect 19680 306005 19685 306035
rect 19715 306005 19720 306035
rect 19680 306000 19720 306005
rect 19840 306035 19880 306040
rect 19840 306005 19845 306035
rect 19875 306005 19880 306035
rect 19840 306000 19880 306005
rect 19680 305955 19720 305960
rect 19680 305925 19685 305955
rect 19715 305925 19720 305955
rect 19680 305920 19720 305925
rect 19840 305955 19880 305960
rect 19840 305925 19845 305955
rect 19875 305925 19880 305955
rect 19840 305920 19880 305925
rect 19680 305875 19720 305880
rect 19680 305845 19685 305875
rect 19715 305845 19720 305875
rect 19680 305840 19720 305845
rect 19840 305875 19880 305880
rect 19840 305845 19845 305875
rect 19875 305845 19880 305875
rect 19840 305840 19880 305845
rect 19680 305795 19720 305800
rect 19680 305765 19685 305795
rect 19715 305765 19720 305795
rect 19680 305760 19720 305765
rect 19840 305795 19880 305800
rect 19840 305765 19845 305795
rect 19875 305765 19880 305795
rect 19840 305760 19880 305765
rect 19680 305715 19720 305720
rect 19680 305685 19685 305715
rect 19715 305685 19720 305715
rect 19680 305680 19720 305685
rect 19840 305715 19880 305720
rect 19840 305685 19845 305715
rect 19875 305685 19880 305715
rect 19840 305680 19880 305685
rect 19680 305635 19720 305640
rect 19680 305605 19685 305635
rect 19715 305605 19720 305635
rect 19680 305600 19720 305605
rect 19840 305635 19880 305640
rect 19840 305605 19845 305635
rect 19875 305605 19880 305635
rect 19840 305600 19880 305605
rect 19680 305555 19720 305560
rect 19680 305525 19685 305555
rect 19715 305525 19720 305555
rect 19680 305520 19720 305525
rect 19840 305555 19880 305560
rect 19840 305525 19845 305555
rect 19875 305525 19880 305555
rect 19840 305520 19880 305525
rect 19680 305475 19720 305480
rect 19680 305445 19685 305475
rect 19715 305445 19720 305475
rect 19680 305440 19720 305445
rect 19840 305475 19880 305480
rect 19840 305445 19845 305475
rect 19875 305445 19880 305475
rect 19840 305440 19880 305445
rect 19680 305395 19720 305400
rect 19680 305365 19685 305395
rect 19715 305365 19720 305395
rect 19680 305360 19720 305365
rect 19840 305395 19880 305400
rect 19840 305365 19845 305395
rect 19875 305365 19880 305395
rect 19840 305360 19880 305365
rect 19680 305315 19720 305320
rect 19680 305285 19685 305315
rect 19715 305285 19720 305315
rect 19680 305280 19720 305285
rect 19840 305315 19880 305320
rect 19840 305285 19845 305315
rect 19875 305285 19880 305315
rect 19840 305280 19880 305285
rect 19680 305235 19720 305240
rect 19680 305205 19685 305235
rect 19715 305205 19720 305235
rect 19680 305200 19720 305205
rect 19840 305235 19880 305240
rect 19840 305205 19845 305235
rect 19875 305205 19880 305235
rect 19840 305200 19880 305205
rect 19680 305155 19720 305160
rect 19680 305125 19685 305155
rect 19715 305125 19720 305155
rect 19680 305120 19720 305125
rect 19840 305155 19880 305160
rect 19840 305125 19845 305155
rect 19875 305125 19880 305155
rect 19840 305120 19880 305125
rect 19680 305075 19720 305080
rect 19680 305045 19685 305075
rect 19715 305045 19720 305075
rect 19680 305040 19720 305045
rect 19840 305075 19880 305080
rect 19840 305045 19845 305075
rect 19875 305045 19880 305075
rect 19840 305040 19880 305045
rect 19680 304995 19720 305000
rect 19680 304965 19685 304995
rect 19715 304965 19720 304995
rect 19680 304960 19720 304965
rect 19840 304995 19880 305000
rect 19840 304965 19845 304995
rect 19875 304965 19880 304995
rect 19840 304960 19880 304965
rect 19680 304915 19720 304920
rect 19680 304885 19685 304915
rect 19715 304885 19720 304915
rect 19680 304880 19720 304885
rect 19840 304915 19880 304920
rect 19840 304885 19845 304915
rect 19875 304885 19880 304915
rect 19840 304880 19880 304885
rect 19680 304835 19720 304840
rect 19680 304805 19685 304835
rect 19715 304805 19720 304835
rect 19680 304800 19720 304805
rect 19840 304835 19880 304840
rect 19840 304805 19845 304835
rect 19875 304805 19880 304835
rect 19840 304800 19880 304805
rect 19680 304755 19720 304760
rect 19680 304725 19685 304755
rect 19715 304725 19720 304755
rect 19680 304720 19720 304725
rect 19840 304755 19880 304760
rect 19840 304725 19845 304755
rect 19875 304725 19880 304755
rect 19840 304720 19880 304725
rect 19680 304675 19720 304680
rect 19680 304645 19685 304675
rect 19715 304645 19720 304675
rect 19680 304640 19720 304645
rect 19840 304675 19880 304680
rect 19840 304645 19845 304675
rect 19875 304645 19880 304675
rect 19840 304640 19880 304645
rect 19680 304595 19720 304600
rect 19680 304565 19685 304595
rect 19715 304565 19720 304595
rect 19680 304560 19720 304565
rect 19840 304595 19880 304600
rect 19840 304565 19845 304595
rect 19875 304565 19880 304595
rect 19840 304560 19880 304565
rect 19680 304515 19720 304520
rect 19680 304485 19685 304515
rect 19715 304485 19720 304515
rect 19680 304480 19720 304485
rect 19840 304515 19880 304520
rect 19840 304485 19845 304515
rect 19875 304485 19880 304515
rect 19840 304480 19880 304485
rect 19680 304435 19720 304440
rect 19680 304405 19685 304435
rect 19715 304405 19720 304435
rect 19680 304400 19720 304405
rect 19840 304435 19880 304440
rect 19840 304405 19845 304435
rect 19875 304405 19880 304435
rect 19840 304400 19880 304405
rect 19680 304355 19720 304360
rect 19680 304325 19685 304355
rect 19715 304325 19720 304355
rect 19680 304320 19720 304325
rect 19840 304355 19880 304360
rect 19840 304325 19845 304355
rect 19875 304325 19880 304355
rect 19840 304320 19880 304325
rect 19680 304275 19720 304280
rect 19680 304245 19685 304275
rect 19715 304245 19720 304275
rect 19680 304240 19720 304245
rect 19840 304275 19880 304280
rect 19840 304245 19845 304275
rect 19875 304245 19880 304275
rect 19840 304240 19880 304245
rect 19680 304195 19720 304200
rect 19680 304165 19685 304195
rect 19715 304165 19720 304195
rect 19680 304160 19720 304165
rect 19840 304195 19880 304200
rect 19840 304165 19845 304195
rect 19875 304165 19880 304195
rect 19840 304160 19880 304165
rect 19680 304115 19720 304120
rect 19680 304085 19685 304115
rect 19715 304085 19720 304115
rect 19680 304080 19720 304085
rect 19840 304115 19880 304120
rect 19840 304085 19845 304115
rect 19875 304085 19880 304115
rect 19840 304080 19880 304085
rect 19680 304035 19720 304040
rect 19680 304005 19685 304035
rect 19715 304005 19720 304035
rect 19680 304000 19720 304005
rect 19840 304035 19880 304040
rect 19840 304005 19845 304035
rect 19875 304005 19880 304035
rect 19840 304000 19880 304005
rect 19680 303955 19720 303960
rect 19680 303925 19685 303955
rect 19715 303925 19720 303955
rect 19680 303920 19720 303925
rect 19840 303955 19880 303960
rect 19840 303925 19845 303955
rect 19875 303925 19880 303955
rect 19840 303920 19880 303925
rect 19680 303875 19720 303880
rect 19680 303845 19685 303875
rect 19715 303845 19720 303875
rect 19680 303840 19720 303845
rect 19840 303875 19880 303880
rect 19840 303845 19845 303875
rect 19875 303845 19880 303875
rect 19840 303840 19880 303845
rect 19680 303795 19720 303800
rect 19680 303765 19685 303795
rect 19715 303765 19720 303795
rect 19680 303760 19720 303765
rect 19840 303795 19880 303800
rect 19840 303765 19845 303795
rect 19875 303765 19880 303795
rect 19840 303760 19880 303765
rect 19680 303715 19720 303720
rect 19680 303685 19685 303715
rect 19715 303685 19720 303715
rect 19680 303680 19720 303685
rect 19840 303715 19880 303720
rect 19840 303685 19845 303715
rect 19875 303685 19880 303715
rect 19840 303680 19880 303685
rect 19680 303635 19720 303640
rect 19680 303605 19685 303635
rect 19715 303605 19720 303635
rect 19680 303600 19720 303605
rect 19840 303635 19880 303640
rect 19840 303605 19845 303635
rect 19875 303605 19880 303635
rect 19840 303600 19880 303605
rect 19680 303555 19720 303560
rect 19680 303525 19685 303555
rect 19715 303525 19720 303555
rect 19680 303520 19720 303525
rect 19840 303555 19880 303560
rect 19840 303525 19845 303555
rect 19875 303525 19880 303555
rect 19840 303520 19880 303525
rect 19680 303475 19720 303480
rect 19680 303445 19685 303475
rect 19715 303445 19720 303475
rect 19680 303440 19720 303445
rect 19840 303475 19880 303480
rect 19840 303445 19845 303475
rect 19875 303445 19880 303475
rect 19840 303440 19880 303445
rect 19680 303395 19720 303400
rect 19680 303365 19685 303395
rect 19715 303365 19720 303395
rect 19680 303360 19720 303365
rect 19840 303395 19880 303400
rect 19840 303365 19845 303395
rect 19875 303365 19880 303395
rect 19840 303360 19880 303365
rect 19680 303315 19720 303320
rect 19680 303285 19685 303315
rect 19715 303285 19720 303315
rect 19680 303280 19720 303285
rect 19840 303315 19880 303320
rect 19840 303285 19845 303315
rect 19875 303285 19880 303315
rect 19840 303280 19880 303285
rect 19680 303235 19720 303240
rect 19680 303205 19685 303235
rect 19715 303205 19720 303235
rect 19680 303200 19720 303205
rect 19840 303235 19880 303240
rect 19840 303205 19845 303235
rect 19875 303205 19880 303235
rect 19840 303200 19880 303205
rect 19680 303155 19720 303160
rect 19680 303125 19685 303155
rect 19715 303125 19720 303155
rect 19680 303120 19720 303125
rect 19840 303155 19880 303160
rect 19840 303125 19845 303155
rect 19875 303125 19880 303155
rect 19840 303120 19880 303125
rect 19680 303075 19720 303080
rect 19680 303045 19685 303075
rect 19715 303045 19720 303075
rect 19680 303040 19720 303045
rect 19840 303075 19880 303080
rect 19840 303045 19845 303075
rect 19875 303045 19880 303075
rect 19840 303040 19880 303045
rect 19680 302995 19720 303000
rect 19680 302965 19685 302995
rect 19715 302965 19720 302995
rect 19680 302960 19720 302965
rect 19840 302995 19880 303000
rect 19840 302965 19845 302995
rect 19875 302965 19880 302995
rect 19840 302960 19880 302965
rect 19680 302915 19720 302920
rect 19680 302885 19685 302915
rect 19715 302885 19720 302915
rect 19680 302880 19720 302885
rect 19840 302915 19880 302920
rect 19840 302885 19845 302915
rect 19875 302885 19880 302915
rect 19840 302880 19880 302885
rect 19680 302835 19720 302840
rect 19680 302805 19685 302835
rect 19715 302805 19720 302835
rect 19680 302800 19720 302805
rect 19840 302835 19880 302840
rect 19840 302805 19845 302835
rect 19875 302805 19880 302835
rect 19840 302800 19880 302805
rect 19680 302755 19720 302760
rect 19680 302725 19685 302755
rect 19715 302725 19720 302755
rect 19680 302720 19720 302725
rect 19840 302755 19880 302760
rect 19840 302725 19845 302755
rect 19875 302725 19880 302755
rect 19840 302720 19880 302725
rect 19680 302675 19720 302680
rect 19680 302645 19685 302675
rect 19715 302645 19720 302675
rect 19680 302640 19720 302645
rect 19840 302675 19880 302680
rect 19840 302645 19845 302675
rect 19875 302645 19880 302675
rect 19840 302640 19880 302645
rect 19680 302595 19720 302600
rect 19680 302565 19685 302595
rect 19715 302565 19720 302595
rect 19680 302560 19720 302565
rect 19840 302595 19880 302600
rect 19840 302565 19845 302595
rect 19875 302565 19880 302595
rect 19840 302560 19880 302565
rect 19680 302515 19720 302520
rect 19680 302485 19685 302515
rect 19715 302485 19720 302515
rect 19680 302480 19720 302485
rect 19840 302515 19880 302520
rect 19840 302485 19845 302515
rect 19875 302485 19880 302515
rect 19840 302480 19880 302485
rect 19680 302435 19720 302440
rect 19680 302405 19685 302435
rect 19715 302405 19720 302435
rect 19680 302400 19720 302405
rect 19840 302435 19880 302440
rect 19840 302405 19845 302435
rect 19875 302405 19880 302435
rect 19840 302400 19880 302405
rect 19680 302355 19720 302360
rect 19680 302325 19685 302355
rect 19715 302325 19720 302355
rect 19680 302320 19720 302325
rect 19840 302355 19880 302360
rect 19840 302325 19845 302355
rect 19875 302325 19880 302355
rect 19840 302320 19880 302325
rect 19680 302275 19720 302280
rect 19680 302245 19685 302275
rect 19715 302245 19720 302275
rect 19680 302240 19720 302245
rect 19840 302275 19880 302280
rect 19840 302245 19845 302275
rect 19875 302245 19880 302275
rect 19840 302240 19880 302245
rect 19680 302195 19720 302200
rect 19680 302165 19685 302195
rect 19715 302165 19720 302195
rect 19680 302160 19720 302165
rect 19840 302195 19880 302200
rect 19840 302165 19845 302195
rect 19875 302165 19880 302195
rect 19840 302160 19880 302165
rect 19680 302115 19720 302120
rect 19680 302085 19685 302115
rect 19715 302085 19720 302115
rect 19680 302080 19720 302085
rect 19840 302115 19880 302120
rect 19840 302085 19845 302115
rect 19875 302085 19880 302115
rect 19840 302080 19880 302085
rect 19680 302035 19720 302040
rect 19680 302005 19685 302035
rect 19715 302005 19720 302035
rect 19680 302000 19720 302005
rect 19840 302035 19880 302040
rect 19840 302005 19845 302035
rect 19875 302005 19880 302035
rect 19840 302000 19880 302005
rect 19680 301955 19720 301960
rect 19680 301925 19685 301955
rect 19715 301925 19720 301955
rect 19680 301920 19720 301925
rect 19840 301955 19880 301960
rect 19840 301925 19845 301955
rect 19875 301925 19880 301955
rect 19840 301920 19880 301925
rect 19680 301875 19720 301880
rect 19680 301845 19685 301875
rect 19715 301845 19720 301875
rect 19680 301840 19720 301845
rect 19840 301875 19880 301880
rect 19840 301845 19845 301875
rect 19875 301845 19880 301875
rect 19840 301840 19880 301845
rect 19680 301795 19720 301800
rect 19680 301765 19685 301795
rect 19715 301765 19720 301795
rect 19680 301760 19720 301765
rect 19840 301795 19880 301800
rect 19840 301765 19845 301795
rect 19875 301765 19880 301795
rect 19840 301760 19880 301765
rect 19680 301715 19720 301720
rect 19680 301685 19685 301715
rect 19715 301685 19720 301715
rect 19680 301680 19720 301685
rect 19840 301715 19880 301720
rect 19840 301685 19845 301715
rect 19875 301685 19880 301715
rect 19840 301680 19880 301685
rect 19680 301635 19720 301640
rect 19680 301605 19685 301635
rect 19715 301605 19720 301635
rect 19680 301600 19720 301605
rect 19840 301635 19880 301640
rect 19840 301605 19845 301635
rect 19875 301605 19880 301635
rect 19840 301600 19880 301605
rect 19680 301555 19720 301560
rect 19680 301525 19685 301555
rect 19715 301525 19720 301555
rect 19680 301520 19720 301525
rect 19840 301555 19880 301560
rect 19840 301525 19845 301555
rect 19875 301525 19880 301555
rect 19840 301520 19880 301525
rect 19680 301475 19720 301480
rect 19680 301445 19685 301475
rect 19715 301445 19720 301475
rect 19680 301440 19720 301445
rect 19840 301475 19880 301480
rect 19840 301445 19845 301475
rect 19875 301445 19880 301475
rect 19840 301440 19880 301445
rect 19680 301395 19720 301400
rect 19680 301365 19685 301395
rect 19715 301365 19720 301395
rect 19680 301360 19720 301365
rect 19840 301395 19880 301400
rect 19840 301365 19845 301395
rect 19875 301365 19880 301395
rect 19840 301360 19880 301365
rect 19680 301315 19720 301320
rect 19680 301285 19685 301315
rect 19715 301285 19720 301315
rect 19680 301280 19720 301285
rect 19840 301315 19880 301320
rect 19840 301285 19845 301315
rect 19875 301285 19880 301315
rect 19840 301280 19880 301285
rect 19680 301235 19720 301240
rect 19680 301205 19685 301235
rect 19715 301205 19720 301235
rect 19680 301200 19720 301205
rect 19840 301235 19880 301240
rect 19840 301205 19845 301235
rect 19875 301205 19880 301235
rect 19840 301200 19880 301205
rect 19680 301155 19720 301160
rect 19680 301125 19685 301155
rect 19715 301125 19720 301155
rect 19680 301120 19720 301125
rect 19840 301155 19880 301160
rect 19840 301125 19845 301155
rect 19875 301125 19880 301155
rect 19840 301120 19880 301125
rect 19680 301075 19720 301080
rect 19680 301045 19685 301075
rect 19715 301045 19720 301075
rect 19680 301040 19720 301045
rect 19840 301075 19880 301080
rect 19840 301045 19845 301075
rect 19875 301045 19880 301075
rect 19840 301040 19880 301045
rect 19680 300995 19720 301000
rect 19680 300965 19685 300995
rect 19715 300965 19720 300995
rect 19680 300960 19720 300965
rect 19840 300995 19880 301000
rect 19840 300965 19845 300995
rect 19875 300965 19880 300995
rect 19840 300960 19880 300965
rect 19680 300915 19720 300920
rect 19680 300885 19685 300915
rect 19715 300885 19720 300915
rect 19680 300880 19720 300885
rect 19840 300915 19880 300920
rect 19840 300885 19845 300915
rect 19875 300885 19880 300915
rect 19840 300880 19880 300885
rect 19680 300835 19720 300840
rect 19680 300805 19685 300835
rect 19715 300805 19720 300835
rect 19680 300800 19720 300805
rect 19840 300835 19880 300840
rect 19840 300805 19845 300835
rect 19875 300805 19880 300835
rect 19840 300800 19880 300805
rect 19680 300755 19720 300760
rect 19680 300725 19685 300755
rect 19715 300725 19720 300755
rect 19680 300720 19720 300725
rect 19840 300755 19880 300760
rect 19840 300725 19845 300755
rect 19875 300725 19880 300755
rect 19840 300720 19880 300725
rect 19680 300675 19720 300680
rect 19680 300645 19685 300675
rect 19715 300645 19720 300675
rect 19680 300640 19720 300645
rect 19840 300675 19880 300680
rect 19840 300645 19845 300675
rect 19875 300645 19880 300675
rect 19840 300640 19880 300645
rect 19680 300595 19720 300600
rect 19680 300565 19685 300595
rect 19715 300565 19720 300595
rect 19680 300560 19720 300565
rect 19840 300595 19880 300600
rect 19840 300565 19845 300595
rect 19875 300565 19880 300595
rect 19840 300560 19880 300565
rect 19680 300515 19720 300520
rect 19680 300485 19685 300515
rect 19715 300485 19720 300515
rect 19680 300480 19720 300485
rect 19840 300515 19880 300520
rect 19840 300485 19845 300515
rect 19875 300485 19880 300515
rect 19840 300480 19880 300485
rect 19680 300435 19720 300440
rect 19680 300405 19685 300435
rect 19715 300405 19720 300435
rect 19680 300400 19720 300405
rect 19840 300435 19880 300440
rect 19840 300405 19845 300435
rect 19875 300405 19880 300435
rect 19840 300400 19880 300405
rect 19680 300355 19720 300360
rect 19680 300325 19685 300355
rect 19715 300325 19720 300355
rect 19680 300320 19720 300325
rect 19840 300355 19880 300360
rect 19840 300325 19845 300355
rect 19875 300325 19880 300355
rect 19840 300320 19880 300325
rect 19680 300275 19720 300280
rect 19680 300245 19685 300275
rect 19715 300245 19720 300275
rect 19680 300240 19720 300245
rect 19840 300275 19880 300280
rect 19840 300245 19845 300275
rect 19875 300245 19880 300275
rect 19840 300240 19880 300245
rect 19680 300195 19720 300200
rect 19680 300165 19685 300195
rect 19715 300165 19720 300195
rect 19680 300160 19720 300165
rect 19840 300195 19880 300200
rect 19840 300165 19845 300195
rect 19875 300165 19880 300195
rect 19840 300160 19880 300165
rect 19680 300115 19720 300120
rect 19680 300085 19685 300115
rect 19715 300085 19720 300115
rect 19680 300080 19720 300085
rect 19840 300115 19880 300120
rect 19840 300085 19845 300115
rect 19875 300085 19880 300115
rect 19840 300080 19880 300085
rect 19680 300035 19720 300040
rect 19680 300005 19685 300035
rect 19715 300005 19720 300035
rect 19680 300000 19720 300005
rect 19840 300035 19880 300040
rect 19840 300005 19845 300035
rect 19875 300005 19880 300035
rect 19840 300000 19880 300005
rect 19680 299955 19720 299960
rect 19680 299925 19685 299955
rect 19715 299925 19720 299955
rect 19680 299920 19720 299925
rect 19840 299955 19880 299960
rect 19840 299925 19845 299955
rect 19875 299925 19880 299955
rect 19840 299920 19880 299925
rect 19680 299875 19720 299880
rect 19680 299845 19685 299875
rect 19715 299845 19720 299875
rect 19680 299840 19720 299845
rect 19840 299875 19880 299880
rect 19840 299845 19845 299875
rect 19875 299845 19880 299875
rect 19840 299840 19880 299845
rect 19680 299795 19720 299800
rect 19680 299765 19685 299795
rect 19715 299765 19720 299795
rect 19680 299760 19720 299765
rect 19840 299795 19880 299800
rect 19840 299765 19845 299795
rect 19875 299765 19880 299795
rect 19840 299760 19880 299765
rect 19680 299715 19720 299720
rect 19680 299685 19685 299715
rect 19715 299685 19720 299715
rect 19680 299680 19720 299685
rect 19840 299715 19880 299720
rect 19840 299685 19845 299715
rect 19875 299685 19880 299715
rect 19840 299680 19880 299685
rect 19680 299635 19720 299640
rect 19680 299605 19685 299635
rect 19715 299605 19720 299635
rect 19680 299600 19720 299605
rect 19840 299635 19880 299640
rect 19840 299605 19845 299635
rect 19875 299605 19880 299635
rect 19840 299600 19880 299605
rect 19680 299555 19720 299560
rect 19680 299525 19685 299555
rect 19715 299525 19720 299555
rect 19680 299520 19720 299525
rect 19840 299555 19880 299560
rect 19840 299525 19845 299555
rect 19875 299525 19880 299555
rect 19840 299520 19880 299525
rect 19680 299475 19720 299480
rect 19680 299445 19685 299475
rect 19715 299445 19720 299475
rect 19680 299440 19720 299445
rect 19840 299475 19880 299480
rect 19840 299445 19845 299475
rect 19875 299445 19880 299475
rect 19840 299440 19880 299445
rect 19680 299395 19720 299400
rect 19680 299365 19685 299395
rect 19715 299365 19720 299395
rect 19680 299360 19720 299365
rect 19840 299395 19880 299400
rect 19840 299365 19845 299395
rect 19875 299365 19880 299395
rect 19840 299360 19880 299365
rect 19680 299315 19720 299320
rect 19680 299285 19685 299315
rect 19715 299285 19720 299315
rect 19680 299280 19720 299285
rect 19840 299315 19880 299320
rect 19840 299285 19845 299315
rect 19875 299285 19880 299315
rect 19840 299280 19880 299285
rect 19680 299235 19720 299240
rect 19680 299205 19685 299235
rect 19715 299205 19720 299235
rect 19680 299200 19720 299205
rect 19840 299235 19880 299240
rect 19840 299205 19845 299235
rect 19875 299205 19880 299235
rect 19840 299200 19880 299205
rect 19680 299155 19720 299160
rect 19680 299125 19685 299155
rect 19715 299125 19720 299155
rect 19680 299120 19720 299125
rect 19840 299155 19880 299160
rect 19840 299125 19845 299155
rect 19875 299125 19880 299155
rect 19840 299120 19880 299125
rect 19680 299075 19720 299080
rect 19680 299045 19685 299075
rect 19715 299045 19720 299075
rect 19680 299040 19720 299045
rect 19840 299075 19880 299080
rect 19840 299045 19845 299075
rect 19875 299045 19880 299075
rect 19840 299040 19880 299045
rect 19680 298995 19720 299000
rect 19680 298965 19685 298995
rect 19715 298965 19720 298995
rect 19680 298960 19720 298965
rect 19840 298995 19880 299000
rect 19840 298965 19845 298995
rect 19875 298965 19880 298995
rect 19840 298960 19880 298965
rect 19680 298915 19720 298920
rect 19680 298885 19685 298915
rect 19715 298885 19720 298915
rect 19680 298880 19720 298885
rect 19840 298915 19880 298920
rect 19840 298885 19845 298915
rect 19875 298885 19880 298915
rect 19840 298880 19880 298885
rect 19680 298835 19720 298840
rect 19680 298805 19685 298835
rect 19715 298805 19720 298835
rect 19680 298800 19720 298805
rect 19840 298835 19880 298840
rect 19840 298805 19845 298835
rect 19875 298805 19880 298835
rect 19840 298800 19880 298805
rect 19680 298755 19720 298760
rect 19680 298725 19685 298755
rect 19715 298725 19720 298755
rect 19680 298720 19720 298725
rect 19840 298755 19880 298760
rect 19840 298725 19845 298755
rect 19875 298725 19880 298755
rect 19840 298720 19880 298725
rect 19680 298675 19720 298680
rect 19680 298645 19685 298675
rect 19715 298645 19720 298675
rect 19680 298640 19720 298645
rect 19840 298675 19880 298680
rect 19840 298645 19845 298675
rect 19875 298645 19880 298675
rect 19840 298640 19880 298645
rect 19680 298595 19720 298600
rect 19680 298565 19685 298595
rect 19715 298565 19720 298595
rect 19680 298560 19720 298565
rect 19840 298595 19880 298600
rect 19840 298565 19845 298595
rect 19875 298565 19880 298595
rect 19840 298560 19880 298565
rect 19680 298515 19720 298520
rect 19680 298485 19685 298515
rect 19715 298485 19720 298515
rect 19680 298480 19720 298485
rect 19840 298515 19880 298520
rect 19840 298485 19845 298515
rect 19875 298485 19880 298515
rect 19840 298480 19880 298485
rect 19680 298435 19720 298440
rect 19680 298405 19685 298435
rect 19715 298405 19720 298435
rect 19680 298400 19720 298405
rect 19840 298435 19880 298440
rect 19840 298405 19845 298435
rect 19875 298405 19880 298435
rect 19840 298400 19880 298405
rect 19680 298355 19720 298360
rect 19680 298325 19685 298355
rect 19715 298325 19720 298355
rect 19680 298320 19720 298325
rect 19840 298355 19880 298360
rect 19840 298325 19845 298355
rect 19875 298325 19880 298355
rect 19840 298320 19880 298325
rect 19680 298275 19720 298280
rect 19680 298245 19685 298275
rect 19715 298245 19720 298275
rect 19680 298240 19720 298245
rect 19840 298275 19880 298280
rect 19840 298245 19845 298275
rect 19875 298245 19880 298275
rect 19840 298240 19880 298245
rect 19680 298195 19720 298200
rect 19680 298165 19685 298195
rect 19715 298165 19720 298195
rect 19680 298160 19720 298165
rect 19840 298195 19880 298200
rect 19840 298165 19845 298195
rect 19875 298165 19880 298195
rect 19840 298160 19880 298165
rect 19680 298115 19720 298120
rect 19680 298085 19685 298115
rect 19715 298085 19720 298115
rect 19680 298080 19720 298085
rect 19840 298115 19880 298120
rect 19840 298085 19845 298115
rect 19875 298085 19880 298115
rect 19840 298080 19880 298085
rect 19680 298035 19720 298040
rect 19680 298005 19685 298035
rect 19715 298005 19720 298035
rect 19680 298000 19720 298005
rect 19840 298035 19880 298040
rect 19840 298005 19845 298035
rect 19875 298005 19880 298035
rect 19840 298000 19880 298005
rect 19680 297955 19720 297960
rect 19680 297925 19685 297955
rect 19715 297925 19720 297955
rect 19680 297920 19720 297925
rect 19840 297955 19880 297960
rect 19840 297925 19845 297955
rect 19875 297925 19880 297955
rect 19840 297920 19880 297925
rect 19680 297875 19720 297880
rect 19680 297845 19685 297875
rect 19715 297845 19720 297875
rect 19680 297840 19720 297845
rect 19840 297875 19880 297880
rect 19840 297845 19845 297875
rect 19875 297845 19880 297875
rect 19840 297840 19880 297845
rect 19680 297795 19720 297800
rect 19680 297765 19685 297795
rect 19715 297765 19720 297795
rect 19680 297760 19720 297765
rect 19840 297795 19880 297800
rect 19840 297765 19845 297795
rect 19875 297765 19880 297795
rect 19840 297760 19880 297765
rect 19680 297715 19720 297720
rect 19680 297685 19685 297715
rect 19715 297685 19720 297715
rect 19680 297680 19720 297685
rect 19840 297715 19880 297720
rect 19840 297685 19845 297715
rect 19875 297685 19880 297715
rect 19840 297680 19880 297685
rect 19680 297635 19720 297640
rect 19680 297605 19685 297635
rect 19715 297605 19720 297635
rect 19680 297600 19720 297605
rect 19840 297635 19880 297640
rect 19840 297605 19845 297635
rect 19875 297605 19880 297635
rect 19840 297600 19880 297605
rect 19680 297555 19720 297560
rect 19680 297525 19685 297555
rect 19715 297525 19720 297555
rect 19680 297520 19720 297525
rect 19840 297555 19880 297560
rect 19840 297525 19845 297555
rect 19875 297525 19880 297555
rect 19840 297520 19880 297525
rect 19680 297475 19720 297480
rect 19680 297445 19685 297475
rect 19715 297445 19720 297475
rect 19680 297440 19720 297445
rect 19840 297475 19880 297480
rect 19840 297445 19845 297475
rect 19875 297445 19880 297475
rect 19840 297440 19880 297445
rect 19680 297395 19720 297400
rect 19680 297365 19685 297395
rect 19715 297365 19720 297395
rect 19680 297360 19720 297365
rect 19840 297395 19880 297400
rect 19840 297365 19845 297395
rect 19875 297365 19880 297395
rect 19840 297360 19880 297365
rect 19680 297315 19720 297320
rect 19680 297285 19685 297315
rect 19715 297285 19720 297315
rect 19680 297280 19720 297285
rect 19840 297315 19880 297320
rect 19840 297285 19845 297315
rect 19875 297285 19880 297315
rect 19840 297280 19880 297285
rect 19680 297235 19720 297240
rect 19680 297205 19685 297235
rect 19715 297205 19720 297235
rect 19680 297200 19720 297205
rect 19840 297235 19880 297240
rect 19840 297205 19845 297235
rect 19875 297205 19880 297235
rect 19840 297200 19880 297205
rect 19680 297155 19720 297160
rect 19680 297125 19685 297155
rect 19715 297125 19720 297155
rect 19680 297120 19720 297125
rect 19840 297155 19880 297160
rect 19840 297125 19845 297155
rect 19875 297125 19880 297155
rect 19840 297120 19880 297125
rect 19680 297075 19720 297080
rect 19680 297045 19685 297075
rect 19715 297045 19720 297075
rect 19680 297040 19720 297045
rect 19840 297075 19880 297080
rect 19840 297045 19845 297075
rect 19875 297045 19880 297075
rect 19840 297040 19880 297045
rect 19680 296995 19720 297000
rect 19680 296965 19685 296995
rect 19715 296965 19720 296995
rect 19680 296960 19720 296965
rect 19840 296995 19880 297000
rect 19840 296965 19845 296995
rect 19875 296965 19880 296995
rect 19840 296960 19880 296965
rect 19680 296915 19720 296920
rect 19680 296885 19685 296915
rect 19715 296885 19720 296915
rect 19680 296880 19720 296885
rect 19840 296915 19880 296920
rect 19840 296885 19845 296915
rect 19875 296885 19880 296915
rect 19840 296880 19880 296885
rect 19680 296835 19720 296840
rect 19680 296805 19685 296835
rect 19715 296805 19720 296835
rect 19680 296800 19720 296805
rect 19840 296835 19880 296840
rect 19840 296805 19845 296835
rect 19875 296805 19880 296835
rect 19840 296800 19880 296805
rect 19680 296755 19720 296760
rect 19680 296725 19685 296755
rect 19715 296725 19720 296755
rect 19680 296720 19720 296725
rect 19840 296755 19880 296760
rect 19840 296725 19845 296755
rect 19875 296725 19880 296755
rect 19840 296720 19880 296725
rect 19680 296675 19720 296680
rect 19680 296645 19685 296675
rect 19715 296645 19720 296675
rect 19680 296640 19720 296645
rect 19840 296675 19880 296680
rect 19840 296645 19845 296675
rect 19875 296645 19880 296675
rect 19840 296640 19880 296645
rect 19680 296595 19720 296600
rect 19680 296565 19685 296595
rect 19715 296565 19720 296595
rect 19680 296560 19720 296565
rect 19840 296595 19880 296600
rect 19840 296565 19845 296595
rect 19875 296565 19880 296595
rect 19840 296560 19880 296565
rect 19680 296515 19720 296520
rect 19680 296485 19685 296515
rect 19715 296485 19720 296515
rect 19680 296480 19720 296485
rect 19840 296515 19880 296520
rect 19840 296485 19845 296515
rect 19875 296485 19880 296515
rect 19840 296480 19880 296485
rect 19680 296435 19720 296440
rect 19680 296405 19685 296435
rect 19715 296405 19720 296435
rect 19680 296400 19720 296405
rect 19840 296435 19880 296440
rect 19840 296405 19845 296435
rect 19875 296405 19880 296435
rect 19840 296400 19880 296405
rect 19680 296355 19720 296360
rect 19680 296325 19685 296355
rect 19715 296325 19720 296355
rect 19680 296320 19720 296325
rect 19840 296355 19880 296360
rect 19840 296325 19845 296355
rect 19875 296325 19880 296355
rect 19840 296320 19880 296325
rect 19680 296275 19720 296280
rect 19680 296245 19685 296275
rect 19715 296245 19720 296275
rect 19680 296240 19720 296245
rect 19840 296275 19880 296280
rect 19840 296245 19845 296275
rect 19875 296245 19880 296275
rect 19840 296240 19880 296245
rect 19680 296195 19720 296200
rect 19680 296165 19685 296195
rect 19715 296165 19720 296195
rect 19680 296160 19720 296165
rect 19840 296195 19880 296200
rect 19840 296165 19845 296195
rect 19875 296165 19880 296195
rect 19840 296160 19880 296165
rect 19680 296115 19720 296120
rect 19680 296085 19685 296115
rect 19715 296085 19720 296115
rect 19680 296080 19720 296085
rect 19840 296115 19880 296120
rect 19840 296085 19845 296115
rect 19875 296085 19880 296115
rect 19840 296080 19880 296085
rect 19680 296035 19720 296040
rect 19680 296005 19685 296035
rect 19715 296005 19720 296035
rect 19680 296000 19720 296005
rect 19840 296035 19880 296040
rect 19840 296005 19845 296035
rect 19875 296005 19880 296035
rect 19840 296000 19880 296005
rect 19680 295955 19720 295960
rect 19680 295925 19685 295955
rect 19715 295925 19720 295955
rect 19680 295920 19720 295925
rect 19840 295955 19880 295960
rect 19840 295925 19845 295955
rect 19875 295925 19880 295955
rect 19840 295920 19880 295925
rect 19680 295875 19720 295880
rect 19680 295845 19685 295875
rect 19715 295845 19720 295875
rect 19680 295840 19720 295845
rect 19840 295875 19880 295880
rect 19840 295845 19845 295875
rect 19875 295845 19880 295875
rect 19840 295840 19880 295845
rect 19680 295795 19720 295800
rect 19680 295765 19685 295795
rect 19715 295765 19720 295795
rect 19680 295760 19720 295765
rect 19840 295795 19880 295800
rect 19840 295765 19845 295795
rect 19875 295765 19880 295795
rect 19840 295760 19880 295765
rect 19680 295715 19720 295720
rect 19680 295685 19685 295715
rect 19715 295685 19720 295715
rect 19680 295680 19720 295685
rect 19840 295715 19880 295720
rect 19840 295685 19845 295715
rect 19875 295685 19880 295715
rect 19840 295680 19880 295685
rect 19680 295635 19720 295640
rect 19680 295605 19685 295635
rect 19715 295605 19720 295635
rect 19680 295600 19720 295605
rect 19840 295635 19880 295640
rect 19840 295605 19845 295635
rect 19875 295605 19880 295635
rect 19840 295600 19880 295605
rect 19680 295555 19720 295560
rect 19680 295525 19685 295555
rect 19715 295525 19720 295555
rect 19680 295520 19720 295525
rect 19840 295555 19880 295560
rect 19840 295525 19845 295555
rect 19875 295525 19880 295555
rect 19840 295520 19880 295525
rect 19680 295475 19720 295480
rect 19680 295445 19685 295475
rect 19715 295445 19720 295475
rect 19680 295440 19720 295445
rect 19840 295475 19880 295480
rect 19840 295445 19845 295475
rect 19875 295445 19880 295475
rect 19840 295440 19880 295445
rect 19680 295395 19720 295400
rect 19680 295365 19685 295395
rect 19715 295365 19720 295395
rect 19680 295360 19720 295365
rect 19840 295395 19880 295400
rect 19840 295365 19845 295395
rect 19875 295365 19880 295395
rect 19840 295360 19880 295365
rect 19680 295315 19720 295320
rect 19680 295285 19685 295315
rect 19715 295285 19720 295315
rect 19680 295280 19720 295285
rect 19840 295315 19880 295320
rect 19840 295285 19845 295315
rect 19875 295285 19880 295315
rect 19840 295280 19880 295285
rect 19680 295235 19720 295240
rect 19680 295205 19685 295235
rect 19715 295205 19720 295235
rect 19680 295200 19720 295205
rect 19840 295235 19880 295240
rect 19840 295205 19845 295235
rect 19875 295205 19880 295235
rect 19840 295200 19880 295205
rect 19680 295155 19720 295160
rect 19680 295125 19685 295155
rect 19715 295125 19720 295155
rect 19680 295120 19720 295125
rect 19840 295155 19880 295160
rect 19840 295125 19845 295155
rect 19875 295125 19880 295155
rect 19840 295120 19880 295125
rect 19680 295075 19720 295080
rect 19680 295045 19685 295075
rect 19715 295045 19720 295075
rect 19680 295040 19720 295045
rect 19840 295075 19880 295080
rect 19840 295045 19845 295075
rect 19875 295045 19880 295075
rect 19840 295040 19880 295045
rect 19680 294995 19720 295000
rect 19680 294965 19685 294995
rect 19715 294965 19720 294995
rect 19680 294960 19720 294965
rect 19840 294995 19880 295000
rect 19840 294965 19845 294995
rect 19875 294965 19880 294995
rect 19840 294960 19880 294965
rect 19680 294915 19720 294920
rect 19680 294885 19685 294915
rect 19715 294885 19720 294915
rect 19680 294880 19720 294885
rect 19840 294915 19880 294920
rect 19840 294885 19845 294915
rect 19875 294885 19880 294915
rect 19840 294880 19880 294885
rect 19680 294835 19720 294840
rect 19680 294805 19685 294835
rect 19715 294805 19720 294835
rect 19680 294800 19720 294805
rect 19840 294835 19880 294840
rect 19840 294805 19845 294835
rect 19875 294805 19880 294835
rect 19840 294800 19880 294805
rect 19680 294755 19720 294760
rect 19680 294725 19685 294755
rect 19715 294725 19720 294755
rect 19680 294720 19720 294725
rect 19840 294755 19880 294760
rect 19840 294725 19845 294755
rect 19875 294725 19880 294755
rect 19840 294720 19880 294725
rect 19680 294675 19720 294680
rect 19680 294645 19685 294675
rect 19715 294645 19720 294675
rect 19680 294640 19720 294645
rect 19840 294675 19880 294680
rect 19840 294645 19845 294675
rect 19875 294645 19880 294675
rect 19840 294640 19880 294645
rect 19680 294595 19720 294600
rect 19680 294565 19685 294595
rect 19715 294565 19720 294595
rect 19680 294560 19720 294565
rect 19840 294595 19880 294600
rect 19840 294565 19845 294595
rect 19875 294565 19880 294595
rect 19840 294560 19880 294565
rect 19680 294515 19720 294520
rect 19680 294485 19685 294515
rect 19715 294485 19720 294515
rect 19680 294480 19720 294485
rect 19840 294515 19880 294520
rect 19840 294485 19845 294515
rect 19875 294485 19880 294515
rect 19840 294480 19880 294485
rect 19680 294435 19720 294440
rect 19680 294405 19685 294435
rect 19715 294405 19720 294435
rect 19680 294400 19720 294405
rect 19840 294435 19880 294440
rect 19840 294405 19845 294435
rect 19875 294405 19880 294435
rect 19840 294400 19880 294405
rect 19680 294355 19720 294360
rect 19680 294325 19685 294355
rect 19715 294325 19720 294355
rect 19680 294320 19720 294325
rect 19840 294355 19880 294360
rect 19840 294325 19845 294355
rect 19875 294325 19880 294355
rect 19840 294320 19880 294325
rect 19680 294275 19720 294280
rect 19680 294245 19685 294275
rect 19715 294245 19720 294275
rect 19680 294240 19720 294245
rect 19840 294275 19880 294280
rect 19840 294245 19845 294275
rect 19875 294245 19880 294275
rect 19840 294240 19880 294245
rect 19680 294195 19720 294200
rect 19680 294165 19685 294195
rect 19715 294165 19720 294195
rect 19680 294160 19720 294165
rect 19840 294195 19880 294200
rect 19840 294165 19845 294195
rect 19875 294165 19880 294195
rect 19840 294160 19880 294165
rect 19680 294115 19720 294120
rect 19680 294085 19685 294115
rect 19715 294085 19720 294115
rect 19680 294080 19720 294085
rect 19840 294115 19880 294120
rect 19840 294085 19845 294115
rect 19875 294085 19880 294115
rect 19840 294080 19880 294085
rect 19680 294035 19720 294040
rect 19680 294005 19685 294035
rect 19715 294005 19720 294035
rect 19680 294000 19720 294005
rect 19840 294035 19880 294040
rect 19840 294005 19845 294035
rect 19875 294005 19880 294035
rect 19840 294000 19880 294005
rect 19680 293955 19720 293960
rect 19680 293925 19685 293955
rect 19715 293925 19720 293955
rect 19680 293920 19720 293925
rect 19840 293955 19880 293960
rect 19840 293925 19845 293955
rect 19875 293925 19880 293955
rect 19840 293920 19880 293925
rect 19680 293875 19720 293880
rect 19680 293845 19685 293875
rect 19715 293845 19720 293875
rect 19680 293840 19720 293845
rect 19840 293875 19880 293880
rect 19840 293845 19845 293875
rect 19875 293845 19880 293875
rect 19840 293840 19880 293845
rect 19680 293795 19720 293800
rect 19680 293765 19685 293795
rect 19715 293765 19720 293795
rect 19680 293760 19720 293765
rect 19840 293795 19880 293800
rect 19840 293765 19845 293795
rect 19875 293765 19880 293795
rect 19840 293760 19880 293765
rect 19680 293715 19720 293720
rect 19680 293685 19685 293715
rect 19715 293685 19720 293715
rect 19680 293680 19720 293685
rect 19840 293715 19880 293720
rect 19840 293685 19845 293715
rect 19875 293685 19880 293715
rect 19840 293680 19880 293685
rect 19680 293635 19720 293640
rect 19680 293605 19685 293635
rect 19715 293605 19720 293635
rect 19680 293600 19720 293605
rect 19840 293635 19880 293640
rect 19840 293605 19845 293635
rect 19875 293605 19880 293635
rect 19840 293600 19880 293605
rect 19680 293555 19720 293560
rect 19680 293525 19685 293555
rect 19715 293525 19720 293555
rect 19680 293520 19720 293525
rect 19840 293555 19880 293560
rect 19840 293525 19845 293555
rect 19875 293525 19880 293555
rect 19840 293520 19880 293525
rect 19680 293475 19720 293480
rect 19680 293445 19685 293475
rect 19715 293445 19720 293475
rect 19680 293440 19720 293445
rect 19840 293475 19880 293480
rect 19840 293445 19845 293475
rect 19875 293445 19880 293475
rect 19840 293440 19880 293445
rect 19680 293395 19720 293400
rect 19680 293365 19685 293395
rect 19715 293365 19720 293395
rect 19680 293360 19720 293365
rect 19840 293395 19880 293400
rect 19840 293365 19845 293395
rect 19875 293365 19880 293395
rect 19840 293360 19880 293365
rect 19680 293315 19720 293320
rect 19680 293285 19685 293315
rect 19715 293285 19720 293315
rect 19680 293280 19720 293285
rect 19840 293315 19880 293320
rect 19840 293285 19845 293315
rect 19875 293285 19880 293315
rect 19840 293280 19880 293285
rect 19680 293235 19720 293240
rect 19680 293205 19685 293235
rect 19715 293205 19720 293235
rect 19680 293200 19720 293205
rect 19840 293235 19880 293240
rect 19840 293205 19845 293235
rect 19875 293205 19880 293235
rect 19840 293200 19880 293205
rect 19680 293155 19720 293160
rect 19680 293125 19685 293155
rect 19715 293125 19720 293155
rect 19680 293120 19720 293125
rect 19840 293155 19880 293160
rect 19840 293125 19845 293155
rect 19875 293125 19880 293155
rect 19840 293120 19880 293125
rect 19680 293075 19720 293080
rect 19680 293045 19685 293075
rect 19715 293045 19720 293075
rect 19680 293040 19720 293045
rect 19840 293075 19880 293080
rect 19840 293045 19845 293075
rect 19875 293045 19880 293075
rect 19840 293040 19880 293045
rect 19680 292995 19720 293000
rect 19680 292965 19685 292995
rect 19715 292965 19720 292995
rect 19680 292960 19720 292965
rect 19840 292995 19880 293000
rect 19840 292965 19845 292995
rect 19875 292965 19880 292995
rect 19840 292960 19880 292965
rect 19680 292915 19720 292920
rect 19680 292885 19685 292915
rect 19715 292885 19720 292915
rect 19680 292880 19720 292885
rect 19840 292915 19880 292920
rect 19840 292885 19845 292915
rect 19875 292885 19880 292915
rect 19840 292880 19880 292885
rect 19680 292835 19720 292840
rect 19680 292805 19685 292835
rect 19715 292805 19720 292835
rect 19680 292800 19720 292805
rect 19840 292835 19880 292840
rect 19840 292805 19845 292835
rect 19875 292805 19880 292835
rect 19840 292800 19880 292805
rect 19680 292755 19720 292760
rect 19680 292725 19685 292755
rect 19715 292725 19720 292755
rect 19680 292720 19720 292725
rect 19840 292755 19880 292760
rect 19840 292725 19845 292755
rect 19875 292725 19880 292755
rect 19840 292720 19880 292725
rect 19680 292675 19720 292680
rect 19680 292645 19685 292675
rect 19715 292645 19720 292675
rect 19680 292640 19720 292645
rect 19840 292675 19880 292680
rect 19840 292645 19845 292675
rect 19875 292645 19880 292675
rect 19840 292640 19880 292645
rect 19680 292595 19720 292600
rect 19680 292565 19685 292595
rect 19715 292565 19720 292595
rect 19680 292560 19720 292565
rect 19840 292595 19880 292600
rect 19840 292565 19845 292595
rect 19875 292565 19880 292595
rect 19840 292560 19880 292565
rect 19680 292515 19720 292520
rect 19680 292485 19685 292515
rect 19715 292485 19720 292515
rect 19680 292480 19720 292485
rect 19840 292515 19880 292520
rect 19840 292485 19845 292515
rect 19875 292485 19880 292515
rect 19840 292480 19880 292485
rect 19680 292435 19720 292440
rect 19680 292405 19685 292435
rect 19715 292405 19720 292435
rect 19680 292400 19720 292405
rect 19840 292435 19880 292440
rect 19840 292405 19845 292435
rect 19875 292405 19880 292435
rect 19840 292400 19880 292405
rect 19680 292355 19720 292360
rect 19680 292325 19685 292355
rect 19715 292325 19720 292355
rect 19680 292320 19720 292325
rect 19840 292355 19880 292360
rect 19840 292325 19845 292355
rect 19875 292325 19880 292355
rect 19840 292320 19880 292325
rect 19680 292275 19720 292280
rect 19680 292245 19685 292275
rect 19715 292245 19720 292275
rect 19680 292240 19720 292245
rect 19840 292275 19880 292280
rect 19840 292245 19845 292275
rect 19875 292245 19880 292275
rect 19840 292240 19880 292245
rect 19680 292195 19720 292200
rect 19680 292165 19685 292195
rect 19715 292165 19720 292195
rect 19680 292160 19720 292165
rect 19840 292195 19880 292200
rect 19840 292165 19845 292195
rect 19875 292165 19880 292195
rect 19840 292160 19880 292165
rect 19680 292115 19720 292120
rect 19680 292085 19685 292115
rect 19715 292085 19720 292115
rect 19680 292080 19720 292085
rect 19840 292115 19880 292120
rect 19840 292085 19845 292115
rect 19875 292085 19880 292115
rect 19840 292080 19880 292085
rect 19680 292035 19720 292040
rect 19680 292005 19685 292035
rect 19715 292005 19720 292035
rect 19680 292000 19720 292005
rect 19840 292035 19880 292040
rect 19840 292005 19845 292035
rect 19875 292005 19880 292035
rect 19840 292000 19880 292005
rect 19680 291955 19720 291960
rect 19680 291925 19685 291955
rect 19715 291925 19720 291955
rect 19680 291920 19720 291925
rect 19840 291955 19880 291960
rect 19840 291925 19845 291955
rect 19875 291925 19880 291955
rect 19840 291920 19880 291925
rect 19680 291875 19720 291880
rect 19680 291845 19685 291875
rect 19715 291845 19720 291875
rect 19680 291840 19720 291845
rect 19840 291875 19880 291880
rect 19840 291845 19845 291875
rect 19875 291845 19880 291875
rect 19840 291840 19880 291845
rect 19680 291795 19720 291800
rect 19680 291765 19685 291795
rect 19715 291765 19720 291795
rect 19680 291760 19720 291765
rect 19840 291795 19880 291800
rect 19840 291765 19845 291795
rect 19875 291765 19880 291795
rect 19840 291760 19880 291765
rect 19680 291715 19720 291720
rect 19680 291685 19685 291715
rect 19715 291685 19720 291715
rect 19680 291680 19720 291685
rect 19840 291715 19880 291720
rect 19840 291685 19845 291715
rect 19875 291685 19880 291715
rect 19840 291680 19880 291685
rect 19680 291635 19720 291640
rect 19680 291605 19685 291635
rect 19715 291605 19720 291635
rect 19680 291600 19720 291605
rect 19840 291635 19880 291640
rect 19840 291605 19845 291635
rect 19875 291605 19880 291635
rect 19840 291600 19880 291605
rect 19680 291555 19720 291560
rect 19680 291525 19685 291555
rect 19715 291525 19720 291555
rect 19680 291520 19720 291525
rect 19840 291555 19880 291560
rect 19840 291525 19845 291555
rect 19875 291525 19880 291555
rect 19840 291520 19880 291525
rect 19680 291475 19720 291480
rect 19680 291445 19685 291475
rect 19715 291445 19720 291475
rect 19680 291440 19720 291445
rect 19840 291475 19880 291480
rect 19840 291445 19845 291475
rect 19875 291445 19880 291475
rect 19840 291440 19880 291445
rect 19680 291395 19720 291400
rect 19680 291365 19685 291395
rect 19715 291365 19720 291395
rect 19680 291360 19720 291365
rect 19840 291395 19880 291400
rect 19840 291365 19845 291395
rect 19875 291365 19880 291395
rect 19840 291360 19880 291365
rect 19680 291315 19720 291320
rect 19680 291285 19685 291315
rect 19715 291285 19720 291315
rect 19680 291280 19720 291285
rect 19840 291315 19880 291320
rect 19840 291285 19845 291315
rect 19875 291285 19880 291315
rect 19840 291280 19880 291285
rect 19680 291235 19720 291240
rect 19680 291205 19685 291235
rect 19715 291205 19720 291235
rect 19680 291200 19720 291205
rect 19840 291235 19880 291240
rect 19840 291205 19845 291235
rect 19875 291205 19880 291235
rect 19840 291200 19880 291205
rect 19680 291155 19720 291160
rect 19680 291125 19685 291155
rect 19715 291125 19720 291155
rect 19680 291120 19720 291125
rect 19840 291155 19880 291160
rect 19840 291125 19845 291155
rect 19875 291125 19880 291155
rect 19840 291120 19880 291125
rect 19680 291075 19720 291080
rect 19680 291045 19685 291075
rect 19715 291045 19720 291075
rect 19680 291040 19720 291045
rect 19840 291075 19880 291080
rect 19840 291045 19845 291075
rect 19875 291045 19880 291075
rect 19840 291040 19880 291045
rect 19680 290995 19720 291000
rect 19680 290965 19685 290995
rect 19715 290965 19720 290995
rect 19680 290960 19720 290965
rect 19840 290995 19880 291000
rect 19840 290965 19845 290995
rect 19875 290965 19880 290995
rect 19840 290960 19880 290965
rect 19680 290915 19720 290920
rect 19680 290885 19685 290915
rect 19715 290885 19720 290915
rect 19680 290880 19720 290885
rect 19840 290915 19880 290920
rect 19840 290885 19845 290915
rect 19875 290885 19880 290915
rect 19840 290880 19880 290885
rect 19680 290835 19720 290840
rect 19680 290805 19685 290835
rect 19715 290805 19720 290835
rect 19680 290800 19720 290805
rect 19840 290835 19880 290840
rect 19840 290805 19845 290835
rect 19875 290805 19880 290835
rect 19840 290800 19880 290805
rect 19680 290755 19720 290760
rect 19680 290725 19685 290755
rect 19715 290725 19720 290755
rect 19680 290720 19720 290725
rect 19840 290755 19880 290760
rect 19840 290725 19845 290755
rect 19875 290725 19880 290755
rect 19840 290720 19880 290725
rect 19680 290675 19720 290680
rect 19680 290645 19685 290675
rect 19715 290645 19720 290675
rect 19680 290640 19720 290645
rect 19840 290675 19880 290680
rect 19840 290645 19845 290675
rect 19875 290645 19880 290675
rect 19840 290640 19880 290645
rect 19680 290595 19720 290600
rect 19680 290565 19685 290595
rect 19715 290565 19720 290595
rect 19680 290560 19720 290565
rect 19840 290595 19880 290600
rect 19840 290565 19845 290595
rect 19875 290565 19880 290595
rect 19840 290560 19880 290565
rect 19680 290515 19720 290520
rect 19680 290485 19685 290515
rect 19715 290485 19720 290515
rect 19680 290480 19720 290485
rect 19840 290515 19880 290520
rect 19840 290485 19845 290515
rect 19875 290485 19880 290515
rect 19840 290480 19880 290485
rect 19680 290435 19720 290440
rect 19680 290405 19685 290435
rect 19715 290405 19720 290435
rect 19680 290400 19720 290405
rect 19840 290435 19880 290440
rect 19840 290405 19845 290435
rect 19875 290405 19880 290435
rect 19840 290400 19880 290405
rect 19680 290355 19720 290360
rect 19680 290325 19685 290355
rect 19715 290325 19720 290355
rect 19680 290320 19720 290325
rect 19840 290355 19880 290360
rect 19840 290325 19845 290355
rect 19875 290325 19880 290355
rect 19840 290320 19880 290325
rect 19680 290275 19720 290280
rect 19680 290245 19685 290275
rect 19715 290245 19720 290275
rect 19680 290240 19720 290245
rect 19840 290275 19880 290280
rect 19840 290245 19845 290275
rect 19875 290245 19880 290275
rect 19840 290240 19880 290245
rect 19680 290195 19720 290200
rect 19680 290165 19685 290195
rect 19715 290165 19720 290195
rect 19680 290160 19720 290165
rect 19840 290195 19880 290200
rect 19840 290165 19845 290195
rect 19875 290165 19880 290195
rect 19840 290160 19880 290165
rect 19680 290115 19720 290120
rect 19680 290085 19685 290115
rect 19715 290085 19720 290115
rect 19680 290080 19720 290085
rect 19840 290115 19880 290120
rect 19840 290085 19845 290115
rect 19875 290085 19880 290115
rect 19840 290080 19880 290085
rect 19680 290035 19720 290040
rect 19680 290005 19685 290035
rect 19715 290005 19720 290035
rect 19680 290000 19720 290005
rect 19840 290035 19880 290040
rect 19840 290005 19845 290035
rect 19875 290005 19880 290035
rect 19840 290000 19880 290005
rect 19680 289955 19720 289960
rect 19680 289925 19685 289955
rect 19715 289925 19720 289955
rect 19680 289920 19720 289925
rect 19840 289955 19880 289960
rect 19840 289925 19845 289955
rect 19875 289925 19880 289955
rect 19840 289920 19880 289925
rect 19680 289875 19720 289880
rect 19680 289845 19685 289875
rect 19715 289845 19720 289875
rect 19680 289840 19720 289845
rect 19840 289875 19880 289880
rect 19840 289845 19845 289875
rect 19875 289845 19880 289875
rect 19840 289840 19880 289845
rect 19680 289795 19720 289800
rect 19680 289765 19685 289795
rect 19715 289765 19720 289795
rect 19680 289760 19720 289765
rect 19840 289795 19880 289800
rect 19840 289765 19845 289795
rect 19875 289765 19880 289795
rect 19840 289760 19880 289765
rect 19680 289715 19720 289720
rect 19680 289685 19685 289715
rect 19715 289685 19720 289715
rect 19680 289680 19720 289685
rect 19840 289715 19880 289720
rect 19840 289685 19845 289715
rect 19875 289685 19880 289715
rect 19840 289680 19880 289685
rect 19680 289635 19720 289640
rect 19680 289605 19685 289635
rect 19715 289605 19720 289635
rect 19680 289600 19720 289605
rect 19840 289635 19880 289640
rect 19840 289605 19845 289635
rect 19875 289605 19880 289635
rect 19840 289600 19880 289605
rect 19680 289555 19720 289560
rect 19680 289525 19685 289555
rect 19715 289525 19720 289555
rect 19680 289520 19720 289525
rect 19840 289555 19880 289560
rect 19840 289525 19845 289555
rect 19875 289525 19880 289555
rect 19840 289520 19880 289525
rect 19680 289475 19720 289480
rect 19680 289445 19685 289475
rect 19715 289445 19720 289475
rect 19680 289440 19720 289445
rect 19840 289475 19880 289480
rect 19840 289445 19845 289475
rect 19875 289445 19880 289475
rect 19840 289440 19880 289445
rect 19680 289395 19720 289400
rect 19680 289365 19685 289395
rect 19715 289365 19720 289395
rect 19680 289360 19720 289365
rect 19840 289395 19880 289400
rect 19840 289365 19845 289395
rect 19875 289365 19880 289395
rect 19840 289360 19880 289365
rect 19680 289315 19720 289320
rect 19680 289285 19685 289315
rect 19715 289285 19720 289315
rect 19680 289280 19720 289285
rect 19840 289315 19880 289320
rect 19840 289285 19845 289315
rect 19875 289285 19880 289315
rect 19840 289280 19880 289285
rect 19680 289235 19720 289240
rect 19680 289205 19685 289235
rect 19715 289205 19720 289235
rect 19680 289200 19720 289205
rect 19840 289235 19880 289240
rect 19840 289205 19845 289235
rect 19875 289205 19880 289235
rect 19840 289200 19880 289205
rect 19680 289155 19720 289160
rect 19680 289125 19685 289155
rect 19715 289125 19720 289155
rect 19680 289120 19720 289125
rect 19840 289155 19880 289160
rect 19840 289125 19845 289155
rect 19875 289125 19880 289155
rect 19840 289120 19880 289125
rect 19680 289075 19720 289080
rect 19680 289045 19685 289075
rect 19715 289045 19720 289075
rect 19680 289040 19720 289045
rect 19840 289075 19880 289080
rect 19840 289045 19845 289075
rect 19875 289045 19880 289075
rect 19840 289040 19880 289045
rect 19680 288995 19720 289000
rect 19680 288965 19685 288995
rect 19715 288965 19720 288995
rect 19680 288960 19720 288965
rect 19840 288995 19880 289000
rect 19840 288965 19845 288995
rect 19875 288965 19880 288995
rect 19840 288960 19880 288965
rect 19680 288915 19720 288920
rect 19680 288885 19685 288915
rect 19715 288885 19720 288915
rect 19680 288880 19720 288885
rect 19840 288915 19880 288920
rect 19840 288885 19845 288915
rect 19875 288885 19880 288915
rect 19840 288880 19880 288885
rect 19680 288835 19720 288840
rect 19680 288805 19685 288835
rect 19715 288805 19720 288835
rect 19680 288800 19720 288805
rect 19840 288835 19880 288840
rect 19840 288805 19845 288835
rect 19875 288805 19880 288835
rect 19840 288800 19880 288805
rect 19680 288755 19720 288760
rect 19680 288725 19685 288755
rect 19715 288725 19720 288755
rect 19680 288720 19720 288725
rect 19840 288755 19880 288760
rect 19840 288725 19845 288755
rect 19875 288725 19880 288755
rect 19840 288720 19880 288725
rect 19680 288675 19720 288680
rect 19680 288645 19685 288675
rect 19715 288645 19720 288675
rect 19680 288640 19720 288645
rect 19840 288675 19880 288680
rect 19840 288645 19845 288675
rect 19875 288645 19880 288675
rect 19840 288640 19880 288645
rect 19680 288595 19720 288600
rect 19680 288565 19685 288595
rect 19715 288565 19720 288595
rect 19680 288560 19720 288565
rect 19840 288595 19880 288600
rect 19840 288565 19845 288595
rect 19875 288565 19880 288595
rect 19840 288560 19880 288565
rect 19680 288515 19720 288520
rect 19680 288485 19685 288515
rect 19715 288485 19720 288515
rect 19680 288480 19720 288485
rect 19840 288515 19880 288520
rect 19840 288485 19845 288515
rect 19875 288485 19880 288515
rect 19840 288480 19880 288485
rect 19680 288435 19720 288440
rect 19680 288405 19685 288435
rect 19715 288405 19720 288435
rect 19680 288400 19720 288405
rect 19840 288435 19880 288440
rect 19840 288405 19845 288435
rect 19875 288405 19880 288435
rect 19840 288400 19880 288405
rect 19680 288355 19720 288360
rect 19680 288325 19685 288355
rect 19715 288325 19720 288355
rect 19680 288320 19720 288325
rect 19840 288355 19880 288360
rect 19840 288325 19845 288355
rect 19875 288325 19880 288355
rect 19840 288320 19880 288325
rect 19680 288275 19720 288280
rect 19680 288245 19685 288275
rect 19715 288245 19720 288275
rect 19680 288240 19720 288245
rect 19840 288275 19880 288280
rect 19840 288245 19845 288275
rect 19875 288245 19880 288275
rect 19840 288240 19880 288245
rect 19680 288195 19720 288200
rect 19680 288165 19685 288195
rect 19715 288165 19720 288195
rect 19680 288160 19720 288165
rect 19840 288195 19880 288200
rect 19840 288165 19845 288195
rect 19875 288165 19880 288195
rect 19840 288160 19880 288165
rect 19680 288115 19720 288120
rect 19680 288085 19685 288115
rect 19715 288085 19720 288115
rect 19680 288080 19720 288085
rect 19840 288115 19880 288120
rect 19840 288085 19845 288115
rect 19875 288085 19880 288115
rect 19840 288080 19880 288085
rect 19680 288035 19720 288040
rect 19680 288005 19685 288035
rect 19715 288005 19720 288035
rect 19680 288000 19720 288005
rect 19840 288035 19880 288040
rect 19840 288005 19845 288035
rect 19875 288005 19880 288035
rect 19840 288000 19880 288005
rect 19680 287955 19720 287960
rect 19680 287925 19685 287955
rect 19715 287925 19720 287955
rect 19680 287920 19720 287925
rect 19840 287955 19880 287960
rect 19840 287925 19845 287955
rect 19875 287925 19880 287955
rect 19840 287920 19880 287925
rect 19680 287875 19720 287880
rect 19680 287845 19685 287875
rect 19715 287845 19720 287875
rect 19680 287840 19720 287845
rect 19840 287875 19880 287880
rect 19840 287845 19845 287875
rect 19875 287845 19880 287875
rect 19840 287840 19880 287845
rect 19680 287795 19720 287800
rect 19680 287765 19685 287795
rect 19715 287765 19720 287795
rect 19680 287760 19720 287765
rect 19840 287795 19880 287800
rect 19840 287765 19845 287795
rect 19875 287765 19880 287795
rect 19840 287760 19880 287765
rect 19680 287715 19720 287720
rect 19680 287685 19685 287715
rect 19715 287685 19720 287715
rect 19680 287680 19720 287685
rect 19840 287715 19880 287720
rect 19840 287685 19845 287715
rect 19875 287685 19880 287715
rect 19840 287680 19880 287685
rect 19680 287635 19720 287640
rect 19680 287605 19685 287635
rect 19715 287605 19720 287635
rect 19680 287600 19720 287605
rect 19840 287635 19880 287640
rect 19840 287605 19845 287635
rect 19875 287605 19880 287635
rect 19840 287600 19880 287605
rect 19680 287555 19720 287560
rect 19680 287525 19685 287555
rect 19715 287525 19720 287555
rect 19680 287520 19720 287525
rect 19840 287555 19880 287560
rect 19840 287525 19845 287555
rect 19875 287525 19880 287555
rect 19840 287520 19880 287525
rect 19680 287475 19720 287480
rect 19680 287445 19685 287475
rect 19715 287445 19720 287475
rect 19680 287440 19720 287445
rect 19840 287475 19880 287480
rect 19840 287445 19845 287475
rect 19875 287445 19880 287475
rect 19840 287440 19880 287445
rect 19680 287395 19720 287400
rect 19680 287365 19685 287395
rect 19715 287365 19720 287395
rect 19680 287360 19720 287365
rect 19840 287395 19880 287400
rect 19840 287365 19845 287395
rect 19875 287365 19880 287395
rect 19840 287360 19880 287365
rect 19680 287315 19720 287320
rect 19680 287285 19685 287315
rect 19715 287285 19720 287315
rect 19680 287280 19720 287285
rect 19840 287315 19880 287320
rect 19840 287285 19845 287315
rect 19875 287285 19880 287315
rect 19840 287280 19880 287285
rect 19680 287235 19720 287240
rect 19680 287205 19685 287235
rect 19715 287205 19720 287235
rect 19680 287200 19720 287205
rect 19840 287235 19880 287240
rect 19840 287205 19845 287235
rect 19875 287205 19880 287235
rect 19840 287200 19880 287205
rect 19680 287155 19720 287160
rect 19680 287125 19685 287155
rect 19715 287125 19720 287155
rect 19680 287120 19720 287125
rect 19840 287155 19880 287160
rect 19840 287125 19845 287155
rect 19875 287125 19880 287155
rect 19840 287120 19880 287125
rect 19680 287075 19720 287080
rect 19680 287045 19685 287075
rect 19715 287045 19720 287075
rect 19680 287040 19720 287045
rect 19840 287075 19880 287080
rect 19840 287045 19845 287075
rect 19875 287045 19880 287075
rect 19840 287040 19880 287045
rect 19680 286995 19720 287000
rect 19680 286965 19685 286995
rect 19715 286965 19720 286995
rect 19680 286960 19720 286965
rect 19840 286995 19880 287000
rect 19840 286965 19845 286995
rect 19875 286965 19880 286995
rect 19840 286960 19880 286965
rect 19680 286915 19720 286920
rect 19680 286885 19685 286915
rect 19715 286885 19720 286915
rect 19680 286880 19720 286885
rect 19840 286915 19880 286920
rect 19840 286885 19845 286915
rect 19875 286885 19880 286915
rect 19840 286880 19880 286885
rect 19680 286835 19720 286840
rect 19680 286805 19685 286835
rect 19715 286805 19720 286835
rect 19680 286800 19720 286805
rect 19840 286835 19880 286840
rect 19840 286805 19845 286835
rect 19875 286805 19880 286835
rect 19840 286800 19880 286805
rect 19680 286755 19720 286760
rect 19680 286725 19685 286755
rect 19715 286725 19720 286755
rect 19680 286720 19720 286725
rect 19840 286755 19880 286760
rect 19840 286725 19845 286755
rect 19875 286725 19880 286755
rect 19840 286720 19880 286725
rect 19680 286675 19720 286680
rect 19680 286645 19685 286675
rect 19715 286645 19720 286675
rect 19680 286640 19720 286645
rect 19840 286675 19880 286680
rect 19840 286645 19845 286675
rect 19875 286645 19880 286675
rect 19840 286640 19880 286645
rect 19680 286595 19720 286600
rect 19680 286565 19685 286595
rect 19715 286565 19720 286595
rect 19680 286560 19720 286565
rect 19840 286595 19880 286600
rect 19840 286565 19845 286595
rect 19875 286565 19880 286595
rect 19840 286560 19880 286565
rect 19680 286515 19720 286520
rect 19680 286485 19685 286515
rect 19715 286485 19720 286515
rect 19680 286480 19720 286485
rect 19840 286515 19880 286520
rect 19840 286485 19845 286515
rect 19875 286485 19880 286515
rect 19840 286480 19880 286485
rect 19680 286435 19720 286440
rect 19680 286405 19685 286435
rect 19715 286405 19720 286435
rect 19680 286400 19720 286405
rect 19840 286435 19880 286440
rect 19840 286405 19845 286435
rect 19875 286405 19880 286435
rect 19840 286400 19880 286405
rect 19680 286355 19720 286360
rect 19680 286325 19685 286355
rect 19715 286325 19720 286355
rect 19680 286320 19720 286325
rect 19840 286355 19880 286360
rect 19840 286325 19845 286355
rect 19875 286325 19880 286355
rect 19840 286320 19880 286325
rect 19680 286275 19720 286280
rect 19680 286245 19685 286275
rect 19715 286245 19720 286275
rect 19680 286240 19720 286245
rect 19840 286275 19880 286280
rect 19840 286245 19845 286275
rect 19875 286245 19880 286275
rect 19840 286240 19880 286245
rect 19680 286195 19720 286200
rect 19680 286165 19685 286195
rect 19715 286165 19720 286195
rect 19680 286160 19720 286165
rect 19840 286195 19880 286200
rect 19840 286165 19845 286195
rect 19875 286165 19880 286195
rect 19840 286160 19880 286165
rect 19680 286115 19720 286120
rect 19680 286085 19685 286115
rect 19715 286085 19720 286115
rect 19680 286080 19720 286085
rect 19840 286115 19880 286120
rect 19840 286085 19845 286115
rect 19875 286085 19880 286115
rect 19840 286080 19880 286085
rect 19680 286035 19720 286040
rect 19680 286005 19685 286035
rect 19715 286005 19720 286035
rect 19680 286000 19720 286005
rect 19840 286035 19880 286040
rect 19840 286005 19845 286035
rect 19875 286005 19880 286035
rect 19840 286000 19880 286005
rect 19680 285955 19720 285960
rect 19680 285925 19685 285955
rect 19715 285925 19720 285955
rect 19680 285920 19720 285925
rect 19840 285955 19880 285960
rect 19840 285925 19845 285955
rect 19875 285925 19880 285955
rect 19840 285920 19880 285925
rect 19680 285875 19720 285880
rect 19680 285845 19685 285875
rect 19715 285845 19720 285875
rect 19680 285840 19720 285845
rect 19840 285875 19880 285880
rect 19840 285845 19845 285875
rect 19875 285845 19880 285875
rect 19840 285840 19880 285845
rect 19680 285795 19720 285800
rect 19680 285765 19685 285795
rect 19715 285765 19720 285795
rect 19680 285760 19720 285765
rect 19840 285795 19880 285800
rect 19840 285765 19845 285795
rect 19875 285765 19880 285795
rect 19840 285760 19880 285765
rect 19680 285715 19720 285720
rect 19680 285685 19685 285715
rect 19715 285685 19720 285715
rect 19680 285680 19720 285685
rect 19840 285715 19880 285720
rect 19840 285685 19845 285715
rect 19875 285685 19880 285715
rect 19840 285680 19880 285685
rect 19680 285635 19720 285640
rect 19680 285605 19685 285635
rect 19715 285605 19720 285635
rect 19680 285600 19720 285605
rect 19840 285635 19880 285640
rect 19840 285605 19845 285635
rect 19875 285605 19880 285635
rect 19840 285600 19880 285605
rect 19680 285555 19720 285560
rect 19680 285525 19685 285555
rect 19715 285525 19720 285555
rect 19680 285520 19720 285525
rect 19840 285555 19880 285560
rect 19840 285525 19845 285555
rect 19875 285525 19880 285555
rect 19840 285520 19880 285525
rect 19680 285475 19720 285480
rect 19680 285445 19685 285475
rect 19715 285445 19720 285475
rect 19680 285440 19720 285445
rect 19840 285475 19880 285480
rect 19840 285445 19845 285475
rect 19875 285445 19880 285475
rect 19840 285440 19880 285445
rect 19680 285395 19720 285400
rect 19680 285365 19685 285395
rect 19715 285365 19720 285395
rect 19680 285360 19720 285365
rect 19840 285395 19880 285400
rect 19840 285365 19845 285395
rect 19875 285365 19880 285395
rect 19840 285360 19880 285365
rect 19680 285315 19720 285320
rect 19680 285285 19685 285315
rect 19715 285285 19720 285315
rect 19680 285280 19720 285285
rect 19840 285315 19880 285320
rect 19840 285285 19845 285315
rect 19875 285285 19880 285315
rect 19840 285280 19880 285285
rect 19680 285235 19720 285240
rect 19680 285205 19685 285235
rect 19715 285205 19720 285235
rect 19680 285200 19720 285205
rect 19840 285235 19880 285240
rect 19840 285205 19845 285235
rect 19875 285205 19880 285235
rect 19840 285200 19880 285205
rect 19680 285155 19720 285160
rect 19680 285125 19685 285155
rect 19715 285125 19720 285155
rect 19680 285120 19720 285125
rect 19840 285155 19880 285160
rect 19840 285125 19845 285155
rect 19875 285125 19880 285155
rect 19840 285120 19880 285125
rect 19680 285075 19720 285080
rect 19680 285045 19685 285075
rect 19715 285045 19720 285075
rect 19680 285040 19720 285045
rect 19840 285075 19880 285080
rect 19840 285045 19845 285075
rect 19875 285045 19880 285075
rect 19840 285040 19880 285045
rect 19680 284995 19720 285000
rect 19680 284965 19685 284995
rect 19715 284965 19720 284995
rect 19680 284960 19720 284965
rect 19840 284995 19880 285000
rect 19840 284965 19845 284995
rect 19875 284965 19880 284995
rect 19840 284960 19880 284965
rect 19680 284915 19720 284920
rect 19680 284885 19685 284915
rect 19715 284885 19720 284915
rect 19680 284880 19720 284885
rect 19840 284915 19880 284920
rect 19840 284885 19845 284915
rect 19875 284885 19880 284915
rect 19840 284880 19880 284885
rect 19680 284835 19720 284840
rect 19680 284805 19685 284835
rect 19715 284805 19720 284835
rect 19680 284800 19720 284805
rect 19840 284835 19880 284840
rect 19840 284805 19845 284835
rect 19875 284805 19880 284835
rect 19840 284800 19880 284805
rect 19680 284755 19720 284760
rect 19680 284725 19685 284755
rect 19715 284725 19720 284755
rect 19680 284720 19720 284725
rect 19840 284755 19880 284760
rect 19840 284725 19845 284755
rect 19875 284725 19880 284755
rect 19840 284720 19880 284725
rect 19680 284675 19720 284680
rect 19680 284645 19685 284675
rect 19715 284645 19720 284675
rect 19680 284640 19720 284645
rect 19840 284675 19880 284680
rect 19840 284645 19845 284675
rect 19875 284645 19880 284675
rect 19840 284640 19880 284645
rect 19680 284595 19720 284600
rect 19680 284565 19685 284595
rect 19715 284565 19720 284595
rect 19680 284560 19720 284565
rect 19840 284595 19880 284600
rect 19840 284565 19845 284595
rect 19875 284565 19880 284595
rect 19840 284560 19880 284565
rect 19680 284515 19720 284520
rect 19680 284485 19685 284515
rect 19715 284485 19720 284515
rect 19680 284480 19720 284485
rect 19840 284515 19880 284520
rect 19840 284485 19845 284515
rect 19875 284485 19880 284515
rect 19840 284480 19880 284485
rect 19680 284435 19720 284440
rect 19680 284405 19685 284435
rect 19715 284405 19720 284435
rect 19680 284400 19720 284405
rect 19840 284435 19880 284440
rect 19840 284405 19845 284435
rect 19875 284405 19880 284435
rect 19840 284400 19880 284405
rect 19680 284355 19720 284360
rect 19680 284325 19685 284355
rect 19715 284325 19720 284355
rect 19680 284320 19720 284325
rect 19840 284355 19880 284360
rect 19840 284325 19845 284355
rect 19875 284325 19880 284355
rect 19840 284320 19880 284325
rect 19680 284275 19720 284280
rect 19680 284245 19685 284275
rect 19715 284245 19720 284275
rect 19680 284240 19720 284245
rect 19840 284275 19880 284280
rect 19840 284245 19845 284275
rect 19875 284245 19880 284275
rect 19840 284240 19880 284245
rect 19680 284195 19720 284200
rect 19680 284165 19685 284195
rect 19715 284165 19720 284195
rect 19680 284160 19720 284165
rect 19840 284195 19880 284200
rect 19840 284165 19845 284195
rect 19875 284165 19880 284195
rect 19840 284160 19880 284165
rect 19680 284115 19720 284120
rect 19680 284085 19685 284115
rect 19715 284085 19720 284115
rect 19680 284080 19720 284085
rect 19840 284115 19880 284120
rect 19840 284085 19845 284115
rect 19875 284085 19880 284115
rect 19840 284080 19880 284085
rect 19680 284035 19720 284040
rect 19680 284005 19685 284035
rect 19715 284005 19720 284035
rect 19680 284000 19720 284005
rect 19840 284035 19880 284040
rect 19840 284005 19845 284035
rect 19875 284005 19880 284035
rect 19840 284000 19880 284005
rect 19680 283955 19720 283960
rect 19680 283925 19685 283955
rect 19715 283925 19720 283955
rect 19680 283920 19720 283925
rect 19840 283955 19880 283960
rect 19840 283925 19845 283955
rect 19875 283925 19880 283955
rect 19840 283920 19880 283925
rect 19680 283875 19720 283880
rect 19680 283845 19685 283875
rect 19715 283845 19720 283875
rect 19680 283840 19720 283845
rect 19840 283875 19880 283880
rect 19840 283845 19845 283875
rect 19875 283845 19880 283875
rect 19840 283840 19880 283845
rect 19680 283795 19720 283800
rect 19680 283765 19685 283795
rect 19715 283765 19720 283795
rect 19680 283760 19720 283765
rect 19840 283795 19880 283800
rect 19840 283765 19845 283795
rect 19875 283765 19880 283795
rect 19840 283760 19880 283765
rect 19680 283715 19720 283720
rect 19680 283685 19685 283715
rect 19715 283685 19720 283715
rect 19680 283680 19720 283685
rect 19840 283715 19880 283720
rect 19840 283685 19845 283715
rect 19875 283685 19880 283715
rect 19840 283680 19880 283685
rect 19680 283635 19720 283640
rect 19680 283605 19685 283635
rect 19715 283605 19720 283635
rect 19680 283600 19720 283605
rect 19840 283635 19880 283640
rect 19840 283605 19845 283635
rect 19875 283605 19880 283635
rect 19840 283600 19880 283605
rect 19680 283555 19720 283560
rect 19680 283525 19685 283555
rect 19715 283525 19720 283555
rect 19680 283520 19720 283525
rect 19840 283555 19880 283560
rect 19840 283525 19845 283555
rect 19875 283525 19880 283555
rect 19840 283520 19880 283525
rect 19680 283475 19720 283480
rect 19680 283445 19685 283475
rect 19715 283445 19720 283475
rect 19680 283440 19720 283445
rect 19840 283475 19880 283480
rect 19840 283445 19845 283475
rect 19875 283445 19880 283475
rect 19840 283440 19880 283445
rect 19680 283395 19720 283400
rect 19680 283365 19685 283395
rect 19715 283365 19720 283395
rect 19680 283360 19720 283365
rect 19840 283395 19880 283400
rect 19840 283365 19845 283395
rect 19875 283365 19880 283395
rect 19840 283360 19880 283365
rect 19680 283315 19720 283320
rect 19680 283285 19685 283315
rect 19715 283285 19720 283315
rect 19680 283280 19720 283285
rect 19840 283315 19880 283320
rect 19840 283285 19845 283315
rect 19875 283285 19880 283315
rect 19840 283280 19880 283285
rect 19680 283235 19720 283240
rect 19680 283205 19685 283235
rect 19715 283205 19720 283235
rect 19680 283200 19720 283205
rect 19840 283235 19880 283240
rect 19840 283205 19845 283235
rect 19875 283205 19880 283235
rect 19840 283200 19880 283205
rect 19680 283155 19720 283160
rect 19680 283125 19685 283155
rect 19715 283125 19720 283155
rect 19680 283120 19720 283125
rect 19840 283155 19880 283160
rect 19840 283125 19845 283155
rect 19875 283125 19880 283155
rect 19840 283120 19880 283125
rect 19680 283075 19720 283080
rect 19680 283045 19685 283075
rect 19715 283045 19720 283075
rect 19680 283040 19720 283045
rect 19840 283075 19880 283080
rect 19840 283045 19845 283075
rect 19875 283045 19880 283075
rect 19840 283040 19880 283045
rect 19680 282995 19720 283000
rect 19680 282965 19685 282995
rect 19715 282965 19720 282995
rect 19680 282960 19720 282965
rect 19840 282995 19880 283000
rect 19840 282965 19845 282995
rect 19875 282965 19880 282995
rect 19840 282960 19880 282965
rect 19680 282915 19720 282920
rect 19680 282885 19685 282915
rect 19715 282885 19720 282915
rect 19680 282880 19720 282885
rect 19840 282915 19880 282920
rect 19840 282885 19845 282915
rect 19875 282885 19880 282915
rect 19840 282880 19880 282885
rect 19680 282835 19720 282840
rect 19680 282805 19685 282835
rect 19715 282805 19720 282835
rect 19680 282800 19720 282805
rect 19840 282835 19880 282840
rect 19840 282805 19845 282835
rect 19875 282805 19880 282835
rect 19840 282800 19880 282805
rect 19680 282755 19720 282760
rect 19680 282725 19685 282755
rect 19715 282725 19720 282755
rect 19680 282720 19720 282725
rect 19840 282755 19880 282760
rect 19840 282725 19845 282755
rect 19875 282725 19880 282755
rect 19840 282720 19880 282725
rect 19680 282675 19720 282680
rect 19680 282645 19685 282675
rect 19715 282645 19720 282675
rect 19680 282640 19720 282645
rect 19840 282675 19880 282680
rect 19840 282645 19845 282675
rect 19875 282645 19880 282675
rect 19840 282640 19880 282645
rect 19680 282595 19720 282600
rect 19680 282565 19685 282595
rect 19715 282565 19720 282595
rect 19680 282560 19720 282565
rect 19840 282595 19880 282600
rect 19840 282565 19845 282595
rect 19875 282565 19880 282595
rect 19840 282560 19880 282565
rect 19680 282515 19720 282520
rect 19680 282485 19685 282515
rect 19715 282485 19720 282515
rect 19680 282480 19720 282485
rect 19840 282515 19880 282520
rect 19840 282485 19845 282515
rect 19875 282485 19880 282515
rect 19840 282480 19880 282485
rect 19680 282435 19720 282440
rect 19680 282405 19685 282435
rect 19715 282405 19720 282435
rect 19680 282400 19720 282405
rect 19840 282435 19880 282440
rect 19840 282405 19845 282435
rect 19875 282405 19880 282435
rect 19840 282400 19880 282405
rect 19680 282355 19720 282360
rect 19680 282325 19685 282355
rect 19715 282325 19720 282355
rect 19680 282320 19720 282325
rect 19840 282355 19880 282360
rect 19840 282325 19845 282355
rect 19875 282325 19880 282355
rect 19840 282320 19880 282325
rect 19680 282275 19720 282280
rect 19680 282245 19685 282275
rect 19715 282245 19720 282275
rect 19680 282240 19720 282245
rect 19840 282275 19880 282280
rect 19840 282245 19845 282275
rect 19875 282245 19880 282275
rect 19840 282240 19880 282245
rect 19680 282195 19720 282200
rect 19680 282165 19685 282195
rect 19715 282165 19720 282195
rect 19680 282160 19720 282165
rect 19840 282195 19880 282200
rect 19840 282165 19845 282195
rect 19875 282165 19880 282195
rect 19840 282160 19880 282165
rect 19680 282115 19720 282120
rect 19680 282085 19685 282115
rect 19715 282085 19720 282115
rect 19680 282080 19720 282085
rect 19840 282115 19880 282120
rect 19840 282085 19845 282115
rect 19875 282085 19880 282115
rect 19840 282080 19880 282085
rect 19680 282035 19720 282040
rect 19680 282005 19685 282035
rect 19715 282005 19720 282035
rect 19680 282000 19720 282005
rect 19840 282035 19880 282040
rect 19840 282005 19845 282035
rect 19875 282005 19880 282035
rect 19840 282000 19880 282005
rect 19680 281955 19720 281960
rect 19680 281925 19685 281955
rect 19715 281925 19720 281955
rect 19680 281920 19720 281925
rect 19840 281955 19880 281960
rect 19840 281925 19845 281955
rect 19875 281925 19880 281955
rect 19840 281920 19880 281925
rect 19680 281875 19720 281880
rect 19680 281845 19685 281875
rect 19715 281845 19720 281875
rect 19680 281840 19720 281845
rect 19840 281875 19880 281880
rect 19840 281845 19845 281875
rect 19875 281845 19880 281875
rect 19840 281840 19880 281845
rect 19680 281795 19720 281800
rect 19680 281765 19685 281795
rect 19715 281765 19720 281795
rect 19680 281760 19720 281765
rect 19840 281795 19880 281800
rect 19840 281765 19845 281795
rect 19875 281765 19880 281795
rect 19840 281760 19880 281765
rect 19680 281715 19720 281720
rect 19680 281685 19685 281715
rect 19715 281685 19720 281715
rect 19680 281680 19720 281685
rect 19840 281715 19880 281720
rect 19840 281685 19845 281715
rect 19875 281685 19880 281715
rect 19840 281680 19880 281685
rect 19680 281635 19720 281640
rect 19680 281605 19685 281635
rect 19715 281605 19720 281635
rect 19680 281600 19720 281605
rect 19840 281635 19880 281640
rect 19840 281605 19845 281635
rect 19875 281605 19880 281635
rect 19840 281600 19880 281605
rect 19680 281555 19720 281560
rect 19680 281525 19685 281555
rect 19715 281525 19720 281555
rect 19680 281520 19720 281525
rect 19840 281555 19880 281560
rect 19840 281525 19845 281555
rect 19875 281525 19880 281555
rect 19840 281520 19880 281525
rect 19680 281475 19720 281480
rect 19680 281445 19685 281475
rect 19715 281445 19720 281475
rect 19680 281440 19720 281445
rect 19840 281475 19880 281480
rect 19840 281445 19845 281475
rect 19875 281445 19880 281475
rect 19840 281440 19880 281445
rect 19680 281395 19720 281400
rect 19680 281365 19685 281395
rect 19715 281365 19720 281395
rect 19680 281360 19720 281365
rect 19840 281395 19880 281400
rect 19840 281365 19845 281395
rect 19875 281365 19880 281395
rect 19840 281360 19880 281365
rect 19680 281315 19720 281320
rect 19680 281285 19685 281315
rect 19715 281285 19720 281315
rect 19680 281280 19720 281285
rect 19840 281315 19880 281320
rect 19840 281285 19845 281315
rect 19875 281285 19880 281315
rect 19840 281280 19880 281285
rect 19680 281235 19720 281240
rect 19680 281205 19685 281235
rect 19715 281205 19720 281235
rect 19680 281200 19720 281205
rect 19840 281235 19880 281240
rect 19840 281205 19845 281235
rect 19875 281205 19880 281235
rect 19840 281200 19880 281205
rect 19680 281155 19720 281160
rect 19680 281125 19685 281155
rect 19715 281125 19720 281155
rect 19680 281120 19720 281125
rect 19840 281155 19880 281160
rect 19840 281125 19845 281155
rect 19875 281125 19880 281155
rect 19840 281120 19880 281125
rect 19680 281075 19720 281080
rect 19680 281045 19685 281075
rect 19715 281045 19720 281075
rect 19680 281040 19720 281045
rect 19840 281075 19880 281080
rect 19840 281045 19845 281075
rect 19875 281045 19880 281075
rect 19840 281040 19880 281045
rect 19680 280995 19720 281000
rect 19680 280965 19685 280995
rect 19715 280965 19720 280995
rect 19680 280960 19720 280965
rect 19840 280995 19880 281000
rect 19840 280965 19845 280995
rect 19875 280965 19880 280995
rect 19840 280960 19880 280965
rect 19680 280915 19720 280920
rect 19680 280885 19685 280915
rect 19715 280885 19720 280915
rect 19680 280880 19720 280885
rect 19840 280915 19880 280920
rect 19840 280885 19845 280915
rect 19875 280885 19880 280915
rect 19840 280880 19880 280885
rect 19680 280835 19720 280840
rect 19680 280805 19685 280835
rect 19715 280805 19720 280835
rect 19680 280800 19720 280805
rect 19840 280835 19880 280840
rect 19840 280805 19845 280835
rect 19875 280805 19880 280835
rect 19840 280800 19880 280805
rect 19680 280755 19720 280760
rect 19680 280725 19685 280755
rect 19715 280725 19720 280755
rect 19680 280720 19720 280725
rect 19840 280755 19880 280760
rect 19840 280725 19845 280755
rect 19875 280725 19880 280755
rect 19840 280720 19880 280725
rect 19680 280675 19720 280680
rect 19680 280645 19685 280675
rect 19715 280645 19720 280675
rect 19680 280640 19720 280645
rect 19840 280675 19880 280680
rect 19840 280645 19845 280675
rect 19875 280645 19880 280675
rect 19840 280640 19880 280645
rect 19680 280595 19720 280600
rect 19680 280565 19685 280595
rect 19715 280565 19720 280595
rect 19680 280560 19720 280565
rect 19840 280595 19880 280600
rect 19840 280565 19845 280595
rect 19875 280565 19880 280595
rect 19840 280560 19880 280565
rect 19680 280515 19720 280520
rect 19680 280485 19685 280515
rect 19715 280485 19720 280515
rect 19680 280480 19720 280485
rect 19840 280515 19880 280520
rect 19840 280485 19845 280515
rect 19875 280485 19880 280515
rect 19840 280480 19880 280485
rect 19680 280435 19720 280440
rect 19680 280405 19685 280435
rect 19715 280405 19720 280435
rect 19680 280400 19720 280405
rect 19840 280435 19880 280440
rect 19840 280405 19845 280435
rect 19875 280405 19880 280435
rect 19840 280400 19880 280405
rect 19680 280355 19720 280360
rect 19680 280325 19685 280355
rect 19715 280325 19720 280355
rect 19680 280320 19720 280325
rect 19840 280355 19880 280360
rect 19840 280325 19845 280355
rect 19875 280325 19880 280355
rect 19840 280320 19880 280325
rect 19680 280275 19720 280280
rect 19680 280245 19685 280275
rect 19715 280245 19720 280275
rect 19680 280240 19720 280245
rect 19840 280275 19880 280280
rect 19840 280245 19845 280275
rect 19875 280245 19880 280275
rect 19840 280240 19880 280245
rect 19680 280195 19720 280200
rect 19680 280165 19685 280195
rect 19715 280165 19720 280195
rect 19680 280160 19720 280165
rect 19840 280195 19880 280200
rect 19840 280165 19845 280195
rect 19875 280165 19880 280195
rect 19840 280160 19880 280165
rect 19680 280115 19720 280120
rect 19680 280085 19685 280115
rect 19715 280085 19720 280115
rect 19680 280080 19720 280085
rect 19840 280115 19880 280120
rect 19840 280085 19845 280115
rect 19875 280085 19880 280115
rect 19840 280080 19880 280085
rect 19680 280035 19720 280040
rect 19680 280005 19685 280035
rect 19715 280005 19720 280035
rect 19680 280000 19720 280005
rect 19840 280035 19880 280040
rect 19840 280005 19845 280035
rect 19875 280005 19880 280035
rect 19840 280000 19880 280005
rect 19680 279955 19720 279960
rect 19680 279925 19685 279955
rect 19715 279925 19720 279955
rect 19680 279920 19720 279925
rect 19840 279955 19880 279960
rect 19840 279925 19845 279955
rect 19875 279925 19880 279955
rect 19840 279920 19880 279925
rect 19680 279875 19720 279880
rect 19680 279845 19685 279875
rect 19715 279845 19720 279875
rect 19680 279840 19720 279845
rect 19840 279875 19880 279880
rect 19840 279845 19845 279875
rect 19875 279845 19880 279875
rect 19840 279840 19880 279845
rect 19680 279795 19720 279800
rect 19680 279765 19685 279795
rect 19715 279765 19720 279795
rect 19680 279760 19720 279765
rect 19840 279795 19880 279800
rect 19840 279765 19845 279795
rect 19875 279765 19880 279795
rect 19840 279760 19880 279765
rect 19680 279715 19720 279720
rect 19680 279685 19685 279715
rect 19715 279685 19720 279715
rect 19680 279680 19720 279685
rect 19840 279715 19880 279720
rect 19840 279685 19845 279715
rect 19875 279685 19880 279715
rect 19840 279680 19880 279685
rect 19680 279635 19720 279640
rect 19680 279605 19685 279635
rect 19715 279605 19720 279635
rect 19680 279600 19720 279605
rect 19840 279635 19880 279640
rect 19840 279605 19845 279635
rect 19875 279605 19880 279635
rect 19840 279600 19880 279605
rect 19680 279555 19720 279560
rect 19680 279525 19685 279555
rect 19715 279525 19720 279555
rect 19680 279520 19720 279525
rect 19840 279555 19880 279560
rect 19840 279525 19845 279555
rect 19875 279525 19880 279555
rect 19840 279520 19880 279525
rect 19680 279475 19720 279480
rect 19680 279445 19685 279475
rect 19715 279445 19720 279475
rect 19680 279440 19720 279445
rect 19840 279475 19880 279480
rect 19840 279445 19845 279475
rect 19875 279445 19880 279475
rect 19840 279440 19880 279445
rect 19680 279395 19720 279400
rect 19680 279365 19685 279395
rect 19715 279365 19720 279395
rect 19680 279360 19720 279365
rect 19840 279395 19880 279400
rect 19840 279365 19845 279395
rect 19875 279365 19880 279395
rect 19840 279360 19880 279365
rect 19680 279315 19720 279320
rect 19680 279285 19685 279315
rect 19715 279285 19720 279315
rect 19680 279280 19720 279285
rect 19840 279315 19880 279320
rect 19840 279285 19845 279315
rect 19875 279285 19880 279315
rect 19840 279280 19880 279285
rect 19680 279235 19720 279240
rect 19680 279205 19685 279235
rect 19715 279205 19720 279235
rect 19680 279200 19720 279205
rect 19840 279235 19880 279240
rect 19840 279205 19845 279235
rect 19875 279205 19880 279235
rect 19840 279200 19880 279205
rect 19680 279155 19720 279160
rect 19680 279125 19685 279155
rect 19715 279125 19720 279155
rect 19680 279120 19720 279125
rect 19840 279155 19880 279160
rect 19840 279125 19845 279155
rect 19875 279125 19880 279155
rect 19840 279120 19880 279125
rect 19680 279075 19720 279080
rect 19680 279045 19685 279075
rect 19715 279045 19720 279075
rect 19680 279040 19720 279045
rect 19840 279075 19880 279080
rect 19840 279045 19845 279075
rect 19875 279045 19880 279075
rect 19840 279040 19880 279045
rect 19680 278995 19720 279000
rect 19680 278965 19685 278995
rect 19715 278965 19720 278995
rect 19680 278960 19720 278965
rect 19840 278995 19880 279000
rect 19840 278965 19845 278995
rect 19875 278965 19880 278995
rect 19840 278960 19880 278965
rect 19680 278915 19720 278920
rect 19680 278885 19685 278915
rect 19715 278885 19720 278915
rect 19680 278880 19720 278885
rect 19840 278915 19880 278920
rect 19840 278885 19845 278915
rect 19875 278885 19880 278915
rect 19840 278880 19880 278885
rect 19680 278835 19720 278840
rect 19680 278805 19685 278835
rect 19715 278805 19720 278835
rect 19680 278800 19720 278805
rect 19840 278835 19880 278840
rect 19840 278805 19845 278835
rect 19875 278805 19880 278835
rect 19840 278800 19880 278805
rect 19680 278755 19720 278760
rect 19680 278725 19685 278755
rect 19715 278725 19720 278755
rect 19680 278720 19720 278725
rect 19840 278755 19880 278760
rect 19840 278725 19845 278755
rect 19875 278725 19880 278755
rect 19840 278720 19880 278725
rect 17040 278675 17080 278680
rect 17040 278645 17045 278675
rect 17075 278645 17080 278675
rect 17040 278640 17080 278645
rect 17200 278675 17240 278680
rect 17200 278645 17205 278675
rect 17235 278645 17240 278675
rect 17200 278640 17240 278645
rect 17280 278675 17320 278680
rect 17280 278645 17285 278675
rect 17315 278645 17320 278675
rect 17280 278640 17320 278645
rect 17360 278675 17400 278680
rect 17360 278645 17365 278675
rect 17395 278645 17400 278675
rect 17360 278640 17400 278645
rect 17440 278675 17480 278680
rect 17440 278645 17445 278675
rect 17475 278645 17480 278675
rect 17440 278640 17480 278645
rect 17520 278675 17560 278680
rect 17520 278645 17525 278675
rect 17555 278645 17560 278675
rect 17520 278640 17560 278645
rect 17600 278675 17640 278680
rect 17600 278645 17605 278675
rect 17635 278645 17640 278675
rect 17600 278640 17640 278645
rect 17680 278675 17720 278680
rect 17680 278645 17685 278675
rect 17715 278645 17720 278675
rect 17680 278640 17720 278645
rect 17760 278675 17800 278680
rect 17760 278645 17765 278675
rect 17795 278645 17800 278675
rect 17760 278640 17800 278645
rect 19520 278675 19560 278680
rect 19520 278645 19525 278675
rect 19555 278645 19560 278675
rect 19520 278640 19560 278645
rect 19600 278675 19640 278680
rect 19600 278645 19605 278675
rect 19635 278645 19640 278675
rect 19600 278640 19640 278645
rect 19680 278675 19720 278680
rect 19680 278645 19685 278675
rect 19715 278645 19720 278675
rect 19680 278640 19720 278645
rect 19840 278675 19880 278680
rect 19840 278645 19845 278675
rect 19875 278645 19880 278675
rect 19840 278640 19880 278645
rect 17040 278515 17080 278520
rect 17040 278485 17045 278515
rect 17075 278485 17080 278515
rect 17040 278480 17080 278485
rect 17200 278515 17240 278520
rect 17200 278485 17205 278515
rect 17235 278485 17240 278515
rect 17200 278480 17240 278485
rect 17280 278515 17320 278520
rect 17280 278485 17285 278515
rect 17315 278485 17320 278515
rect 17280 278480 17320 278485
rect 17360 278515 17400 278520
rect 17360 278485 17365 278515
rect 17395 278485 17400 278515
rect 17360 278480 17400 278485
rect 17440 278515 17480 278520
rect 17440 278485 17445 278515
rect 17475 278485 17480 278515
rect 17440 278480 17480 278485
rect 17520 278515 17560 278520
rect 17520 278485 17525 278515
rect 17555 278485 17560 278515
rect 17520 278480 17560 278485
rect 17600 278515 17640 278520
rect 17600 278485 17605 278515
rect 17635 278485 17640 278515
rect 17600 278480 17640 278485
rect 17680 278515 17720 278520
rect 17680 278485 17685 278515
rect 17715 278485 17720 278515
rect 17680 278480 17720 278485
rect 17760 278515 17800 278520
rect 17760 278485 17765 278515
rect 17795 278485 17800 278515
rect 17760 278480 17800 278485
rect 19520 278515 19560 278520
rect 19520 278485 19525 278515
rect 19555 278485 19560 278515
rect 19520 278480 19560 278485
rect 19600 278515 19640 278520
rect 19600 278485 19605 278515
rect 19635 278485 19640 278515
rect 19600 278480 19640 278485
rect 19680 278515 19720 278520
rect 19680 278485 19685 278515
rect 19715 278485 19720 278515
rect 19680 278480 19720 278485
rect 19840 278515 19880 278520
rect 19840 278485 19845 278515
rect 19875 278485 19880 278515
rect 19840 278480 19880 278485
rect 17040 278435 17080 278440
rect 17040 278405 17045 278435
rect 17075 278405 17080 278435
rect 17040 278400 17080 278405
rect 17200 278435 17240 278440
rect 17200 278405 17205 278435
rect 17235 278405 17240 278435
rect 17200 278400 17240 278405
rect 17040 278355 17080 278360
rect 17040 278325 17045 278355
rect 17075 278325 17080 278355
rect 17040 278320 17080 278325
rect 17200 278355 17240 278360
rect 17200 278325 17205 278355
rect 17235 278325 17240 278355
rect 17200 278320 17240 278325
rect 17040 278275 17080 278280
rect 17040 278245 17045 278275
rect 17075 278245 17080 278275
rect 17040 278240 17080 278245
rect 17200 278275 17240 278280
rect 17200 278245 17205 278275
rect 17235 278245 17240 278275
rect 17200 278240 17240 278245
rect 17040 278195 17080 278200
rect 17040 278165 17045 278195
rect 17075 278165 17080 278195
rect 17040 278160 17080 278165
rect 17200 278195 17240 278200
rect 17200 278165 17205 278195
rect 17235 278165 17240 278195
rect 17200 278160 17240 278165
rect 17040 278115 17080 278120
rect 17040 278085 17045 278115
rect 17075 278085 17080 278115
rect 17040 278080 17080 278085
rect 17200 278115 17240 278120
rect 17200 278085 17205 278115
rect 17235 278085 17240 278115
rect 17200 278080 17240 278085
rect 17040 278035 17080 278040
rect 17040 278005 17045 278035
rect 17075 278005 17080 278035
rect 17040 278000 17080 278005
rect 17200 278035 17240 278040
rect 17200 278005 17205 278035
rect 17235 278005 17240 278035
rect 17200 278000 17240 278005
rect 17040 277955 17080 277960
rect 17040 277925 17045 277955
rect 17075 277925 17080 277955
rect 17040 277920 17080 277925
rect 17200 277955 17240 277960
rect 17200 277925 17205 277955
rect 17235 277925 17240 277955
rect 17200 277920 17240 277925
rect 17040 277875 17080 277880
rect 17040 277845 17045 277875
rect 17075 277845 17080 277875
rect 17040 277840 17080 277845
rect 17200 277875 17240 277880
rect 17200 277845 17205 277875
rect 17235 277845 17240 277875
rect 17200 277840 17240 277845
<< via1 >>
rect 10725 351365 10755 351395
rect 10805 351365 10835 351395
rect 10885 351365 10915 351395
rect 10965 351365 10995 351395
rect 11045 351365 11075 351395
rect 11125 351365 11155 351395
rect 11205 351365 11235 351395
rect 11285 351365 11315 351395
rect 11365 351365 11395 351395
rect 11445 351365 11475 351395
rect 11525 351365 11555 351395
rect 11605 351365 11635 351395
rect 11685 351365 11715 351395
rect 11765 351365 11795 351395
rect 11845 351365 11875 351395
rect 11925 351365 11955 351395
rect 12005 351365 12035 351395
rect 12085 351365 12115 351395
rect 12165 351365 12195 351395
rect 12245 351365 12275 351395
rect 12325 351365 12355 351395
rect 12405 351365 12435 351395
rect 12485 351365 12515 351395
rect 12565 351365 12595 351395
rect 12645 351365 12675 351395
rect 12725 351365 12755 351395
rect 12805 351365 12835 351395
rect 12885 351365 12915 351395
rect 12965 351365 12995 351395
rect 13045 351365 13075 351395
rect 13125 351365 13155 351395
rect 13205 351365 13235 351395
rect 13285 351365 13315 351395
rect 13365 351365 13395 351395
rect 13445 351365 13475 351395
rect 13525 351365 13555 351395
rect 13605 351365 13635 351395
rect 13685 351365 13715 351395
rect 13765 351365 13795 351395
rect 13845 351365 13875 351395
rect 13925 351365 13955 351395
rect 14005 351365 14035 351395
rect 14085 351365 14115 351395
rect 14165 351365 14195 351395
rect 14245 351365 14275 351395
rect 14325 351365 14355 351395
rect 14405 351365 14435 351395
rect 14485 351365 14515 351395
rect 14565 351365 14595 351395
rect 14645 351365 14675 351395
rect 14725 351365 14755 351395
rect 14805 351365 14835 351395
rect 14885 351365 14915 351395
rect 14965 351365 14995 351395
rect 15045 351365 15075 351395
rect 15125 351365 15155 351395
rect 15205 351365 15235 351395
rect 15285 351365 15315 351395
rect 15365 351365 15395 351395
rect 15445 351365 15475 351395
rect 15525 351365 15555 351395
rect 15605 351365 15635 351395
rect 15685 351365 15715 351395
rect 15765 351365 15795 351395
rect 15845 351365 15875 351395
rect 15925 351365 15955 351395
rect 16005 351365 16035 351395
rect 16085 351365 16115 351395
rect 16165 351365 16195 351395
rect 16245 351365 16275 351395
rect 16325 351365 16355 351395
rect 16405 351365 16435 351395
rect 16485 351365 16515 351395
rect 16565 351365 16595 351395
rect 16645 351365 16675 351395
rect 16725 351365 16755 351395
rect 16805 351365 16835 351395
rect 16885 351365 16915 351395
rect 16965 351365 16995 351395
rect 17045 351365 17075 351395
rect 17125 351365 17155 351395
rect 17205 351365 17235 351395
rect 17285 351365 17315 351395
rect 17365 351365 17395 351395
rect 17445 351365 17475 351395
rect 17525 351365 17555 351395
rect 17605 351365 17635 351395
rect 17685 351365 17715 351395
rect 17765 351365 17795 351395
rect 17845 351365 17875 351395
rect 17925 351365 17955 351395
rect 18005 351365 18035 351395
rect 18085 351365 18115 351395
rect 18165 351365 18195 351395
rect 18245 351365 18275 351395
rect 18325 351365 18355 351395
rect 18405 351365 18435 351395
rect 18485 351365 18515 351395
rect 18565 351365 18595 351395
rect 18645 351365 18675 351395
rect 18725 351365 18755 351395
rect 18805 351365 18835 351395
rect 18885 351365 18915 351395
rect 18965 351365 18995 351395
rect 19045 351365 19075 351395
rect 19125 351365 19155 351395
rect 19205 351365 19235 351395
rect 19285 351365 19315 351395
rect 19365 351365 19395 351395
rect 19445 351365 19475 351395
rect 19525 351365 19555 351395
rect 19605 351365 19635 351395
rect 19685 351365 19715 351395
rect 19845 351365 19875 351395
rect 10725 351205 10755 351235
rect 10805 351205 10835 351235
rect 10885 351205 10915 351235
rect 10965 351205 10995 351235
rect 11045 351205 11075 351235
rect 11125 351205 11155 351235
rect 11205 351205 11235 351235
rect 11285 351205 11315 351235
rect 11365 351205 11395 351235
rect 11445 351205 11475 351235
rect 11525 351205 11555 351235
rect 11605 351205 11635 351235
rect 11685 351205 11715 351235
rect 11765 351205 11795 351235
rect 11845 351205 11875 351235
rect 11925 351205 11955 351235
rect 12005 351205 12035 351235
rect 12085 351205 12115 351235
rect 12165 351205 12195 351235
rect 12245 351205 12275 351235
rect 12325 351205 12355 351235
rect 12405 351205 12435 351235
rect 12485 351205 12515 351235
rect 12565 351205 12595 351235
rect 12645 351205 12675 351235
rect 12725 351205 12755 351235
rect 12805 351205 12835 351235
rect 12885 351205 12915 351235
rect 12965 351205 12995 351235
rect 13045 351205 13075 351235
rect 13125 351205 13155 351235
rect 13205 351205 13235 351235
rect 13285 351205 13315 351235
rect 13365 351205 13395 351235
rect 13445 351205 13475 351235
rect 13525 351205 13555 351235
rect 13605 351205 13635 351235
rect 13685 351205 13715 351235
rect 13765 351205 13795 351235
rect 13845 351205 13875 351235
rect 13925 351205 13955 351235
rect 14005 351205 14035 351235
rect 14085 351205 14115 351235
rect 14165 351205 14195 351235
rect 14245 351205 14275 351235
rect 14325 351205 14355 351235
rect 14405 351205 14435 351235
rect 14485 351205 14515 351235
rect 14565 351205 14595 351235
rect 14645 351205 14675 351235
rect 14725 351205 14755 351235
rect 14805 351205 14835 351235
rect 14885 351205 14915 351235
rect 14965 351205 14995 351235
rect 15045 351205 15075 351235
rect 15125 351205 15155 351235
rect 15205 351205 15235 351235
rect 15285 351205 15315 351235
rect 15365 351205 15395 351235
rect 15445 351205 15475 351235
rect 15525 351205 15555 351235
rect 15605 351205 15635 351235
rect 15685 351205 15715 351235
rect 15765 351205 15795 351235
rect 15845 351205 15875 351235
rect 15925 351205 15955 351235
rect 16005 351205 16035 351235
rect 16085 351205 16115 351235
rect 16165 351205 16195 351235
rect 16245 351205 16275 351235
rect 16325 351205 16355 351235
rect 16405 351205 16435 351235
rect 16485 351205 16515 351235
rect 16565 351205 16595 351235
rect 16645 351205 16675 351235
rect 16725 351205 16755 351235
rect 16805 351205 16835 351235
rect 16885 351205 16915 351235
rect 16965 351205 16995 351235
rect 17045 351205 17075 351235
rect 17125 351205 17155 351235
rect 17205 351205 17235 351235
rect 17285 351205 17315 351235
rect 17365 351205 17395 351235
rect 17445 351205 17475 351235
rect 17525 351205 17555 351235
rect 17605 351205 17635 351235
rect 17685 351205 17715 351235
rect 17765 351205 17795 351235
rect 17845 351205 17875 351235
rect 17925 351205 17955 351235
rect 18005 351205 18035 351235
rect 18085 351205 18115 351235
rect 18165 351205 18195 351235
rect 18245 351205 18275 351235
rect 18325 351205 18355 351235
rect 18405 351205 18435 351235
rect 18485 351205 18515 351235
rect 18565 351205 18595 351235
rect 18645 351205 18675 351235
rect 18725 351205 18755 351235
rect 18805 351205 18835 351235
rect 18885 351205 18915 351235
rect 18965 351205 18995 351235
rect 19045 351205 19075 351235
rect 19125 351205 19155 351235
rect 19205 351205 19235 351235
rect 19285 351205 19315 351235
rect 19365 351205 19395 351235
rect 19445 351205 19475 351235
rect 19525 351205 19555 351235
rect 19605 351205 19635 351235
rect 19685 351205 19715 351235
rect 19845 351205 19875 351235
rect 19685 351125 19715 351155
rect 19845 351125 19875 351155
rect 19685 351045 19715 351075
rect 19845 351045 19875 351075
rect 19685 350965 19715 350995
rect 19845 350965 19875 350995
rect 19685 350885 19715 350915
rect 19845 350885 19875 350915
rect 19685 350805 19715 350835
rect 19845 350805 19875 350835
rect 19685 350725 19715 350755
rect 19845 350725 19875 350755
rect 19685 350645 19715 350675
rect 19845 350645 19875 350675
rect 19685 350565 19715 350595
rect 19845 350565 19875 350595
rect 19685 350485 19715 350515
rect 19845 350485 19875 350515
rect 19685 350405 19715 350435
rect 19845 350405 19875 350435
rect 19685 350325 19715 350355
rect 19845 350325 19875 350355
rect 19685 350245 19715 350275
rect 19845 350245 19875 350275
rect 19685 350165 19715 350195
rect 19845 350165 19875 350195
rect 19685 350085 19715 350115
rect 19845 350085 19875 350115
rect 19685 350005 19715 350035
rect 19845 350005 19875 350035
rect 19685 349925 19715 349955
rect 19845 349925 19875 349955
rect 19685 349845 19715 349875
rect 19845 349845 19875 349875
rect 19685 349765 19715 349795
rect 19845 349765 19875 349795
rect 19685 349685 19715 349715
rect 19845 349685 19875 349715
rect 19685 349605 19715 349635
rect 19845 349605 19875 349635
rect 19685 349525 19715 349555
rect 19845 349525 19875 349555
rect 19685 349445 19715 349475
rect 19845 349445 19875 349475
rect 19685 349365 19715 349395
rect 19845 349365 19875 349395
rect 19685 349285 19715 349315
rect 19845 349285 19875 349315
rect 19685 349205 19715 349235
rect 19845 349205 19875 349235
rect 19685 349125 19715 349155
rect 19845 349125 19875 349155
rect 19685 349045 19715 349075
rect 19845 349045 19875 349075
rect 19685 348965 19715 348995
rect 19845 348965 19875 348995
rect 19685 348885 19715 348915
rect 19845 348885 19875 348915
rect 19685 348805 19715 348835
rect 19845 348805 19875 348835
rect 19685 348725 19715 348755
rect 19845 348725 19875 348755
rect 19685 348645 19715 348675
rect 19845 348645 19875 348675
rect 19685 348565 19715 348595
rect 19845 348565 19875 348595
rect 19685 348485 19715 348515
rect 19845 348485 19875 348515
rect 19685 348405 19715 348435
rect 19845 348405 19875 348435
rect 19685 348325 19715 348355
rect 19845 348325 19875 348355
rect 19685 348245 19715 348275
rect 19845 348245 19875 348275
rect 19685 348165 19715 348195
rect 19845 348165 19875 348195
rect 19685 348085 19715 348115
rect 19845 348085 19875 348115
rect 19685 348005 19715 348035
rect 19845 348005 19875 348035
rect 19685 347925 19715 347955
rect 19845 347925 19875 347955
rect 19685 347845 19715 347875
rect 19845 347845 19875 347875
rect 19685 347765 19715 347795
rect 19845 347765 19875 347795
rect 19685 347685 19715 347715
rect 19845 347685 19875 347715
rect 19685 347605 19715 347635
rect 19845 347605 19875 347635
rect 19685 347525 19715 347555
rect 19845 347525 19875 347555
rect 19685 347445 19715 347475
rect 19845 347445 19875 347475
rect 19685 347365 19715 347395
rect 19845 347365 19875 347395
rect 19685 347285 19715 347315
rect 19845 347285 19875 347315
rect 19685 347205 19715 347235
rect 19845 347205 19875 347235
rect 19685 347125 19715 347155
rect 19845 347125 19875 347155
rect 19685 347045 19715 347075
rect 19845 347045 19875 347075
rect 19685 346965 19715 346995
rect 19845 346965 19875 346995
rect 19685 346885 19715 346915
rect 19845 346885 19875 346915
rect 19685 346805 19715 346835
rect 19845 346805 19875 346835
rect 19685 346725 19715 346755
rect 19845 346725 19875 346755
rect 19685 346645 19715 346675
rect 19845 346645 19875 346675
rect 19685 346565 19715 346595
rect 19845 346565 19875 346595
rect 19685 346485 19715 346515
rect 19845 346485 19875 346515
rect 19685 346405 19715 346435
rect 19845 346405 19875 346435
rect 19685 346325 19715 346355
rect 19845 346325 19875 346355
rect 19685 346245 19715 346275
rect 19845 346245 19875 346275
rect 19685 346165 19715 346195
rect 19845 346165 19875 346195
rect 19685 346085 19715 346115
rect 19845 346085 19875 346115
rect 19685 346005 19715 346035
rect 19845 346005 19875 346035
rect 19685 345925 19715 345955
rect 19845 345925 19875 345955
rect 19685 345845 19715 345875
rect 19845 345845 19875 345875
rect 19685 345765 19715 345795
rect 19845 345765 19875 345795
rect 19685 345685 19715 345715
rect 19845 345685 19875 345715
rect 19685 345605 19715 345635
rect 19845 345605 19875 345635
rect 19685 345525 19715 345555
rect 19845 345525 19875 345555
rect 19685 345445 19715 345475
rect 19845 345445 19875 345475
rect 19685 345365 19715 345395
rect 19845 345365 19875 345395
rect 19685 345285 19715 345315
rect 19845 345285 19875 345315
rect 19685 345205 19715 345235
rect 19845 345205 19875 345235
rect 19685 345125 19715 345155
rect 19845 345125 19875 345155
rect 19685 345045 19715 345075
rect 19845 345045 19875 345075
rect 19685 344965 19715 344995
rect 19845 344965 19875 344995
rect 19685 344885 19715 344915
rect 19845 344885 19875 344915
rect 19685 344805 19715 344835
rect 19845 344805 19875 344835
rect 19685 344725 19715 344755
rect 19845 344725 19875 344755
rect 19685 344645 19715 344675
rect 19845 344645 19875 344675
rect 19685 344565 19715 344595
rect 19845 344565 19875 344595
rect 19685 344485 19715 344515
rect 19845 344485 19875 344515
rect 19685 344405 19715 344435
rect 19845 344405 19875 344435
rect 19685 344325 19715 344355
rect 19845 344325 19875 344355
rect 19685 344245 19715 344275
rect 19845 344245 19875 344275
rect 19685 344165 19715 344195
rect 19845 344165 19875 344195
rect 19685 344085 19715 344115
rect 19845 344085 19875 344115
rect 19685 344005 19715 344035
rect 19845 344005 19875 344035
rect 19685 343925 19715 343955
rect 19845 343925 19875 343955
rect 19685 343845 19715 343875
rect 19845 343845 19875 343875
rect 19685 343765 19715 343795
rect 19845 343765 19875 343795
rect 19685 343685 19715 343715
rect 19845 343685 19875 343715
rect 19685 343605 19715 343635
rect 19845 343605 19875 343635
rect 19685 343525 19715 343555
rect 19845 343525 19875 343555
rect 19685 343445 19715 343475
rect 19845 343445 19875 343475
rect 19685 343365 19715 343395
rect 19845 343365 19875 343395
rect 19685 343285 19715 343315
rect 19845 343285 19875 343315
rect 19685 343205 19715 343235
rect 19845 343205 19875 343235
rect 19685 343125 19715 343155
rect 19845 343125 19875 343155
rect 19685 343045 19715 343075
rect 19845 343045 19875 343075
rect 19685 342965 19715 342995
rect 19845 342965 19875 342995
rect 19685 342885 19715 342915
rect 19845 342885 19875 342915
rect 19685 342805 19715 342835
rect 19845 342805 19875 342835
rect 19685 342725 19715 342755
rect 19845 342725 19875 342755
rect 19685 342645 19715 342675
rect 19845 342645 19875 342675
rect 19685 342565 19715 342595
rect 19845 342565 19875 342595
rect 19685 342485 19715 342515
rect 19845 342485 19875 342515
rect 19685 342405 19715 342435
rect 19845 342405 19875 342435
rect 19685 342325 19715 342355
rect 19845 342325 19875 342355
rect 19685 342245 19715 342275
rect 19845 342245 19875 342275
rect 19685 342165 19715 342195
rect 19845 342165 19875 342195
rect 19685 342085 19715 342115
rect 19845 342085 19875 342115
rect 19685 342005 19715 342035
rect 19845 342005 19875 342035
rect 19685 341925 19715 341955
rect 19845 341925 19875 341955
rect 19685 341845 19715 341875
rect 19845 341845 19875 341875
rect 19685 341765 19715 341795
rect 19845 341765 19875 341795
rect 19685 341685 19715 341715
rect 19845 341685 19875 341715
rect 19685 341605 19715 341635
rect 19845 341605 19875 341635
rect 19685 341525 19715 341555
rect 19845 341525 19875 341555
rect 19685 341445 19715 341475
rect 19845 341445 19875 341475
rect 19685 341365 19715 341395
rect 19845 341365 19875 341395
rect 19685 341285 19715 341315
rect 19845 341285 19875 341315
rect 19685 341205 19715 341235
rect 19845 341205 19875 341235
rect 19685 341125 19715 341155
rect 19845 341125 19875 341155
rect 19685 341045 19715 341075
rect 19845 341045 19875 341075
rect 19685 340965 19715 340995
rect 19845 340965 19875 340995
rect 19685 340885 19715 340915
rect 19845 340885 19875 340915
rect 19685 340805 19715 340835
rect 19845 340805 19875 340835
rect 19685 340725 19715 340755
rect 19845 340725 19875 340755
rect 19685 340645 19715 340675
rect 19845 340645 19875 340675
rect 19685 340565 19715 340595
rect 19845 340565 19875 340595
rect 19685 340485 19715 340515
rect 19845 340485 19875 340515
rect 19685 340405 19715 340435
rect 19845 340405 19875 340435
rect 19685 340325 19715 340355
rect 19845 340325 19875 340355
rect 19685 340245 19715 340275
rect 19845 340245 19875 340275
rect 19685 340165 19715 340195
rect 19845 340165 19875 340195
rect 19685 340085 19715 340115
rect 19845 340085 19875 340115
rect 19685 340005 19715 340035
rect 19845 340005 19875 340035
rect 19685 339925 19715 339955
rect 19845 339925 19875 339955
rect 19685 339845 19715 339875
rect 19845 339845 19875 339875
rect 19685 339765 19715 339795
rect 19845 339765 19875 339795
rect 19685 339685 19715 339715
rect 19845 339685 19875 339715
rect 19685 339605 19715 339635
rect 19845 339605 19875 339635
rect 19685 339525 19715 339555
rect 19845 339525 19875 339555
rect 19685 339445 19715 339475
rect 19845 339445 19875 339475
rect 19685 339365 19715 339395
rect 19845 339365 19875 339395
rect 19685 339285 19715 339315
rect 19845 339285 19875 339315
rect 19685 339205 19715 339235
rect 19845 339205 19875 339235
rect 19685 339125 19715 339155
rect 19845 339125 19875 339155
rect 19685 339045 19715 339075
rect 19845 339045 19875 339075
rect 19685 338965 19715 338995
rect 19845 338965 19875 338995
rect 19685 338885 19715 338915
rect 19845 338885 19875 338915
rect 19685 338805 19715 338835
rect 19845 338805 19875 338835
rect 19685 338725 19715 338755
rect 19845 338725 19875 338755
rect 19685 338645 19715 338675
rect 19845 338645 19875 338675
rect 19685 338565 19715 338595
rect 19845 338565 19875 338595
rect 19685 338485 19715 338515
rect 19845 338485 19875 338515
rect 19685 338405 19715 338435
rect 19845 338405 19875 338435
rect 19685 338325 19715 338355
rect 19845 338325 19875 338355
rect 19685 338245 19715 338275
rect 19845 338245 19875 338275
rect 19685 338165 19715 338195
rect 19845 338165 19875 338195
rect 19685 338085 19715 338115
rect 19845 338085 19875 338115
rect 19685 338005 19715 338035
rect 19845 338005 19875 338035
rect 19685 337925 19715 337955
rect 19845 337925 19875 337955
rect 19685 337845 19715 337875
rect 19845 337845 19875 337875
rect 19685 337765 19715 337795
rect 19845 337765 19875 337795
rect 19685 337685 19715 337715
rect 19845 337685 19875 337715
rect 19685 337605 19715 337635
rect 19845 337605 19875 337635
rect 19685 337525 19715 337555
rect 19845 337525 19875 337555
rect 19685 337445 19715 337475
rect 19845 337445 19875 337475
rect 19685 337365 19715 337395
rect 19845 337365 19875 337395
rect 19685 337285 19715 337315
rect 19845 337285 19875 337315
rect 19685 337205 19715 337235
rect 19845 337205 19875 337235
rect 19685 337125 19715 337155
rect 19845 337125 19875 337155
rect 19685 337045 19715 337075
rect 19845 337045 19875 337075
rect 19685 336965 19715 336995
rect 19845 336965 19875 336995
rect 19685 336885 19715 336915
rect 19845 336885 19875 336915
rect 19685 336805 19715 336835
rect 19845 336805 19875 336835
rect 19685 336725 19715 336755
rect 19845 336725 19875 336755
rect 19685 336645 19715 336675
rect 19845 336645 19875 336675
rect 19685 336565 19715 336595
rect 19845 336565 19875 336595
rect 19685 336485 19715 336515
rect 19845 336485 19875 336515
rect 19685 336405 19715 336435
rect 19845 336405 19875 336435
rect 19685 336325 19715 336355
rect 19845 336325 19875 336355
rect 19685 336245 19715 336275
rect 19845 336245 19875 336275
rect 19685 336165 19715 336195
rect 19845 336165 19875 336195
rect 19685 336085 19715 336115
rect 19845 336085 19875 336115
rect 19685 336005 19715 336035
rect 19845 336005 19875 336035
rect 19685 335925 19715 335955
rect 19845 335925 19875 335955
rect 19685 335845 19715 335875
rect 19845 335845 19875 335875
rect 19685 335765 19715 335795
rect 19845 335765 19875 335795
rect 19685 335685 19715 335715
rect 19845 335685 19875 335715
rect 19685 335605 19715 335635
rect 19845 335605 19875 335635
rect 19685 335525 19715 335555
rect 19845 335525 19875 335555
rect 19685 335445 19715 335475
rect 19845 335445 19875 335475
rect 19685 335365 19715 335395
rect 19845 335365 19875 335395
rect 19685 335285 19715 335315
rect 19845 335285 19875 335315
rect 19685 335205 19715 335235
rect 19845 335205 19875 335235
rect 19685 335125 19715 335155
rect 19845 335125 19875 335155
rect 19685 335045 19715 335075
rect 19845 335045 19875 335075
rect 19685 334965 19715 334995
rect 19845 334965 19875 334995
rect 19685 334885 19715 334915
rect 19845 334885 19875 334915
rect 19685 334805 19715 334835
rect 19845 334805 19875 334835
rect 19685 334725 19715 334755
rect 19845 334725 19875 334755
rect 19685 334645 19715 334675
rect 19845 334645 19875 334675
rect 19685 334565 19715 334595
rect 19845 334565 19875 334595
rect 19685 334485 19715 334515
rect 19845 334485 19875 334515
rect 19685 334405 19715 334435
rect 19845 334405 19875 334435
rect 19685 334325 19715 334355
rect 19845 334325 19875 334355
rect 19685 334245 19715 334275
rect 19845 334245 19875 334275
rect 19685 334165 19715 334195
rect 19845 334165 19875 334195
rect 19685 334085 19715 334115
rect 19845 334085 19875 334115
rect 19685 334005 19715 334035
rect 19845 334005 19875 334035
rect 19685 333925 19715 333955
rect 19845 333925 19875 333955
rect 19685 333845 19715 333875
rect 19845 333845 19875 333875
rect 19685 333765 19715 333795
rect 19845 333765 19875 333795
rect 19685 333685 19715 333715
rect 19845 333685 19875 333715
rect 19685 333605 19715 333635
rect 19845 333605 19875 333635
rect 19685 333525 19715 333555
rect 19845 333525 19875 333555
rect 19685 333445 19715 333475
rect 19845 333445 19875 333475
rect 19685 333365 19715 333395
rect 19845 333365 19875 333395
rect 19685 333285 19715 333315
rect 19845 333285 19875 333315
rect 19685 333205 19715 333235
rect 19845 333205 19875 333235
rect 19685 333125 19715 333155
rect 19845 333125 19875 333155
rect 19685 333045 19715 333075
rect 19845 333045 19875 333075
rect 19685 332965 19715 332995
rect 19845 332965 19875 332995
rect 19685 332885 19715 332915
rect 19845 332885 19875 332915
rect 19685 332805 19715 332835
rect 19845 332805 19875 332835
rect 19685 332725 19715 332755
rect 19845 332725 19875 332755
rect 19685 332645 19715 332675
rect 19845 332645 19875 332675
rect 19685 332565 19715 332595
rect 19845 332565 19875 332595
rect 19685 332485 19715 332515
rect 19845 332485 19875 332515
rect 19685 332405 19715 332435
rect 19845 332405 19875 332435
rect 19685 332325 19715 332355
rect 19845 332325 19875 332355
rect 19685 332245 19715 332275
rect 19845 332245 19875 332275
rect 19685 332165 19715 332195
rect 19845 332165 19875 332195
rect 19685 332085 19715 332115
rect 19845 332085 19875 332115
rect 19685 332005 19715 332035
rect 19845 332005 19875 332035
rect 19685 331925 19715 331955
rect 19845 331925 19875 331955
rect 19685 331845 19715 331875
rect 19845 331845 19875 331875
rect 19685 331765 19715 331795
rect 19845 331765 19875 331795
rect 19685 331685 19715 331715
rect 19845 331685 19875 331715
rect 19685 331605 19715 331635
rect 19845 331605 19875 331635
rect 19685 331525 19715 331555
rect 19845 331525 19875 331555
rect 19685 331445 19715 331475
rect 19845 331445 19875 331475
rect 19685 331365 19715 331395
rect 19845 331365 19875 331395
rect 19685 331285 19715 331315
rect 19845 331285 19875 331315
rect 19685 331205 19715 331235
rect 19845 331205 19875 331235
rect 19685 331125 19715 331155
rect 19845 331125 19875 331155
rect 19685 331045 19715 331075
rect 19845 331045 19875 331075
rect 19685 330965 19715 330995
rect 19845 330965 19875 330995
rect 19685 330885 19715 330915
rect 19845 330885 19875 330915
rect 19685 330805 19715 330835
rect 19845 330805 19875 330835
rect 19685 330725 19715 330755
rect 19845 330725 19875 330755
rect 19685 330645 19715 330675
rect 19845 330645 19875 330675
rect 19685 330565 19715 330595
rect 19845 330565 19875 330595
rect 19685 330485 19715 330515
rect 19845 330485 19875 330515
rect 19685 330405 19715 330435
rect 19845 330405 19875 330435
rect 19685 330325 19715 330355
rect 19845 330325 19875 330355
rect 19685 330245 19715 330275
rect 19845 330245 19875 330275
rect 19685 330165 19715 330195
rect 19845 330165 19875 330195
rect 19685 330085 19715 330115
rect 19845 330085 19875 330115
rect 19685 330005 19715 330035
rect 19845 330005 19875 330035
rect 19685 329925 19715 329955
rect 19845 329925 19875 329955
rect 19685 329845 19715 329875
rect 19845 329845 19875 329875
rect 19685 329765 19715 329795
rect 19845 329765 19875 329795
rect 19685 329685 19715 329715
rect 19845 329685 19875 329715
rect 19685 329605 19715 329635
rect 19845 329605 19875 329635
rect 19685 329525 19715 329555
rect 19845 329525 19875 329555
rect 19685 329445 19715 329475
rect 19845 329445 19875 329475
rect 19685 329365 19715 329395
rect 19845 329365 19875 329395
rect 19685 329285 19715 329315
rect 19845 329285 19875 329315
rect 19685 329205 19715 329235
rect 19845 329205 19875 329235
rect 19685 329125 19715 329155
rect 19845 329125 19875 329155
rect 19685 329045 19715 329075
rect 19845 329045 19875 329075
rect 19685 328965 19715 328995
rect 19845 328965 19875 328995
rect 19685 328885 19715 328915
rect 19845 328885 19875 328915
rect 19685 328805 19715 328835
rect 19845 328805 19875 328835
rect 19685 328725 19715 328755
rect 19845 328725 19875 328755
rect 19685 328645 19715 328675
rect 19845 328645 19875 328675
rect 19685 328565 19715 328595
rect 19845 328565 19875 328595
rect 19685 328485 19715 328515
rect 19845 328485 19875 328515
rect 19685 328405 19715 328435
rect 19845 328405 19875 328435
rect 19685 328325 19715 328355
rect 19845 328325 19875 328355
rect 19685 328245 19715 328275
rect 19845 328245 19875 328275
rect 19685 328165 19715 328195
rect 19845 328165 19875 328195
rect 19685 328085 19715 328115
rect 19845 328085 19875 328115
rect 19685 328005 19715 328035
rect 19845 328005 19875 328035
rect 19685 327925 19715 327955
rect 19845 327925 19875 327955
rect 19685 327845 19715 327875
rect 19845 327845 19875 327875
rect 19685 327765 19715 327795
rect 19845 327765 19875 327795
rect 19685 327685 19715 327715
rect 19845 327685 19875 327715
rect 19685 327605 19715 327635
rect 19845 327605 19875 327635
rect 19685 327525 19715 327555
rect 19845 327525 19875 327555
rect 19685 327445 19715 327475
rect 19845 327445 19875 327475
rect 19685 327365 19715 327395
rect 19845 327365 19875 327395
rect 19685 327285 19715 327315
rect 19845 327285 19875 327315
rect 19685 327205 19715 327235
rect 19845 327205 19875 327235
rect 19685 327125 19715 327155
rect 19845 327125 19875 327155
rect 19685 327045 19715 327075
rect 19845 327045 19875 327075
rect 19685 326965 19715 326995
rect 19845 326965 19875 326995
rect 19685 326885 19715 326915
rect 19845 326885 19875 326915
rect 19685 326805 19715 326835
rect 19845 326805 19875 326835
rect 19685 326725 19715 326755
rect 19845 326725 19875 326755
rect 19685 326645 19715 326675
rect 19845 326645 19875 326675
rect 19685 326565 19715 326595
rect 19845 326565 19875 326595
rect 19685 326485 19715 326515
rect 19845 326485 19875 326515
rect 19685 326405 19715 326435
rect 19845 326405 19875 326435
rect 19685 326325 19715 326355
rect 19845 326325 19875 326355
rect 19685 326245 19715 326275
rect 19845 326245 19875 326275
rect 19685 326165 19715 326195
rect 19845 326165 19875 326195
rect 19685 326085 19715 326115
rect 19845 326085 19875 326115
rect 19685 326005 19715 326035
rect 19845 326005 19875 326035
rect 19685 325925 19715 325955
rect 19845 325925 19875 325955
rect 19685 325845 19715 325875
rect 19845 325845 19875 325875
rect 19685 325765 19715 325795
rect 19845 325765 19875 325795
rect 19685 325685 19715 325715
rect 19845 325685 19875 325715
rect 19685 325605 19715 325635
rect 19845 325605 19875 325635
rect 19685 325525 19715 325555
rect 19845 325525 19875 325555
rect 19685 325445 19715 325475
rect 19845 325445 19875 325475
rect 19685 325365 19715 325395
rect 19845 325365 19875 325395
rect 19685 325285 19715 325315
rect 19845 325285 19875 325315
rect 19685 325205 19715 325235
rect 19845 325205 19875 325235
rect 19685 325125 19715 325155
rect 19845 325125 19875 325155
rect 19685 325045 19715 325075
rect 19845 325045 19875 325075
rect 19685 324965 19715 324995
rect 19845 324965 19875 324995
rect 19685 324885 19715 324915
rect 19845 324885 19875 324915
rect 19685 324805 19715 324835
rect 19845 324805 19875 324835
rect 19685 324725 19715 324755
rect 19845 324725 19875 324755
rect 19685 324645 19715 324675
rect 19845 324645 19875 324675
rect 19685 324565 19715 324595
rect 19845 324565 19875 324595
rect 19685 324485 19715 324515
rect 19845 324485 19875 324515
rect 19685 324405 19715 324435
rect 19845 324405 19875 324435
rect 19685 324325 19715 324355
rect 19845 324325 19875 324355
rect 19685 324245 19715 324275
rect 19845 324245 19875 324275
rect 19685 324165 19715 324195
rect 19845 324165 19875 324195
rect 19685 324085 19715 324115
rect 19845 324085 19875 324115
rect 19685 324005 19715 324035
rect 19845 324005 19875 324035
rect 19685 323925 19715 323955
rect 19845 323925 19875 323955
rect 19685 323845 19715 323875
rect 19845 323845 19875 323875
rect 19685 323765 19715 323795
rect 19845 323765 19875 323795
rect 19685 323685 19715 323715
rect 19845 323685 19875 323715
rect 19685 323605 19715 323635
rect 19845 323605 19875 323635
rect 19685 323525 19715 323555
rect 19845 323525 19875 323555
rect 19685 323445 19715 323475
rect 19845 323445 19875 323475
rect 19685 323365 19715 323395
rect 19845 323365 19875 323395
rect 19685 323285 19715 323315
rect 19845 323285 19875 323315
rect 19685 323205 19715 323235
rect 19845 323205 19875 323235
rect 19685 323125 19715 323155
rect 19845 323125 19875 323155
rect 19685 323045 19715 323075
rect 19845 323045 19875 323075
rect 19685 322965 19715 322995
rect 19845 322965 19875 322995
rect 19685 322885 19715 322915
rect 19845 322885 19875 322915
rect 19685 322805 19715 322835
rect 19845 322805 19875 322835
rect 19685 322725 19715 322755
rect 19845 322725 19875 322755
rect 19685 322645 19715 322675
rect 19845 322645 19875 322675
rect 19685 322565 19715 322595
rect 19845 322565 19875 322595
rect 19685 322485 19715 322515
rect 19845 322485 19875 322515
rect 19685 322405 19715 322435
rect 19845 322405 19875 322435
rect 19685 322325 19715 322355
rect 19845 322325 19875 322355
rect 19685 322245 19715 322275
rect 19845 322245 19875 322275
rect 19685 322165 19715 322195
rect 19845 322165 19875 322195
rect 19685 322085 19715 322115
rect 19845 322085 19875 322115
rect 19685 322005 19715 322035
rect 19845 322005 19875 322035
rect 19685 321925 19715 321955
rect 19845 321925 19875 321955
rect 19685 321845 19715 321875
rect 19845 321845 19875 321875
rect 19685 321765 19715 321795
rect 19845 321765 19875 321795
rect 19685 321685 19715 321715
rect 19845 321685 19875 321715
rect 19685 321605 19715 321635
rect 19845 321605 19875 321635
rect 19685 321525 19715 321555
rect 19845 321525 19875 321555
rect 19685 321445 19715 321475
rect 19845 321445 19875 321475
rect 19685 321365 19715 321395
rect 19845 321365 19875 321395
rect 19685 321285 19715 321315
rect 19845 321285 19875 321315
rect 19685 321205 19715 321235
rect 19845 321205 19875 321235
rect 19685 321125 19715 321155
rect 19845 321125 19875 321155
rect 19685 321045 19715 321075
rect 19845 321045 19875 321075
rect 19685 320965 19715 320995
rect 19845 320965 19875 320995
rect 19685 320885 19715 320915
rect 19845 320885 19875 320915
rect 19685 320805 19715 320835
rect 19845 320805 19875 320835
rect 19685 320725 19715 320755
rect 19845 320725 19875 320755
rect 19685 320645 19715 320675
rect 19845 320645 19875 320675
rect 19685 320565 19715 320595
rect 19845 320565 19875 320595
rect 19685 320485 19715 320515
rect 19845 320485 19875 320515
rect 19685 320405 19715 320435
rect 19845 320405 19875 320435
rect 19685 320325 19715 320355
rect 19845 320325 19875 320355
rect 19685 320245 19715 320275
rect 19845 320245 19875 320275
rect 19685 320165 19715 320195
rect 19845 320165 19875 320195
rect 19685 320085 19715 320115
rect 19845 320085 19875 320115
rect 19685 320005 19715 320035
rect 19845 320005 19875 320035
rect 19685 319925 19715 319955
rect 19845 319925 19875 319955
rect 19685 319845 19715 319875
rect 19845 319845 19875 319875
rect 19685 319765 19715 319795
rect 19845 319765 19875 319795
rect 19685 319685 19715 319715
rect 19845 319685 19875 319715
rect 19685 319605 19715 319635
rect 19845 319605 19875 319635
rect 19685 319525 19715 319555
rect 19845 319525 19875 319555
rect 19685 319445 19715 319475
rect 19845 319445 19875 319475
rect 19685 319365 19715 319395
rect 19845 319365 19875 319395
rect 19685 319285 19715 319315
rect 19845 319285 19875 319315
rect 19685 319205 19715 319235
rect 19845 319205 19875 319235
rect 19685 319125 19715 319155
rect 19845 319125 19875 319155
rect 19685 319045 19715 319075
rect 19845 319045 19875 319075
rect 19685 318965 19715 318995
rect 19845 318965 19875 318995
rect 19685 318885 19715 318915
rect 19845 318885 19875 318915
rect 19685 318805 19715 318835
rect 19845 318805 19875 318835
rect 19685 318725 19715 318755
rect 19845 318725 19875 318755
rect 19685 318645 19715 318675
rect 19845 318645 19875 318675
rect 19685 318565 19715 318595
rect 19845 318565 19875 318595
rect 19685 318485 19715 318515
rect 19845 318485 19875 318515
rect 19685 318405 19715 318435
rect 19845 318405 19875 318435
rect 19685 318325 19715 318355
rect 19845 318325 19875 318355
rect 19685 318245 19715 318275
rect 19845 318245 19875 318275
rect 19685 318165 19715 318195
rect 19845 318165 19875 318195
rect 19685 318085 19715 318115
rect 19845 318085 19875 318115
rect 19685 318005 19715 318035
rect 19845 318005 19875 318035
rect 19685 317925 19715 317955
rect 19845 317925 19875 317955
rect 19685 317845 19715 317875
rect 19845 317845 19875 317875
rect 19685 317765 19715 317795
rect 19845 317765 19875 317795
rect 19685 317685 19715 317715
rect 19845 317685 19875 317715
rect 19685 317605 19715 317635
rect 19845 317605 19875 317635
rect 19685 317525 19715 317555
rect 19845 317525 19875 317555
rect 19685 317445 19715 317475
rect 19845 317445 19875 317475
rect 19685 317365 19715 317395
rect 19845 317365 19875 317395
rect 19685 317285 19715 317315
rect 19845 317285 19875 317315
rect 19685 317205 19715 317235
rect 19845 317205 19875 317235
rect 19685 317125 19715 317155
rect 19845 317125 19875 317155
rect 19685 317045 19715 317075
rect 19845 317045 19875 317075
rect 19685 316965 19715 316995
rect 19845 316965 19875 316995
rect 19685 316885 19715 316915
rect 19845 316885 19875 316915
rect 19685 316805 19715 316835
rect 19845 316805 19875 316835
rect 19685 316725 19715 316755
rect 19845 316725 19875 316755
rect 19685 316645 19715 316675
rect 19845 316645 19875 316675
rect 19685 316565 19715 316595
rect 19845 316565 19875 316595
rect 19685 316485 19715 316515
rect 19845 316485 19875 316515
rect 19685 316405 19715 316435
rect 19845 316405 19875 316435
rect 19685 316325 19715 316355
rect 19845 316325 19875 316355
rect 19685 316245 19715 316275
rect 19845 316245 19875 316275
rect 19685 316165 19715 316195
rect 19845 316165 19875 316195
rect 19685 316085 19715 316115
rect 19845 316085 19875 316115
rect 19685 316005 19715 316035
rect 19845 316005 19875 316035
rect 19685 315925 19715 315955
rect 19845 315925 19875 315955
rect 19685 315845 19715 315875
rect 19845 315845 19875 315875
rect 19685 315765 19715 315795
rect 19845 315765 19875 315795
rect 19685 315685 19715 315715
rect 19845 315685 19875 315715
rect 19685 315605 19715 315635
rect 19845 315605 19875 315635
rect 19685 315525 19715 315555
rect 19845 315525 19875 315555
rect 19685 315445 19715 315475
rect 19845 315445 19875 315475
rect 19685 315365 19715 315395
rect 19845 315365 19875 315395
rect 19685 315285 19715 315315
rect 19845 315285 19875 315315
rect 19685 315205 19715 315235
rect 19845 315205 19875 315235
rect 19685 315125 19715 315155
rect 19845 315125 19875 315155
rect 19685 315045 19715 315075
rect 19845 315045 19875 315075
rect 19685 314965 19715 314995
rect 19845 314965 19875 314995
rect 19685 314885 19715 314915
rect 19845 314885 19875 314915
rect 19685 314805 19715 314835
rect 19845 314805 19875 314835
rect 19685 314725 19715 314755
rect 19845 314725 19875 314755
rect 19685 314645 19715 314675
rect 19845 314645 19875 314675
rect 19685 314565 19715 314595
rect 19845 314565 19875 314595
rect 19685 314485 19715 314515
rect 19845 314485 19875 314515
rect 19685 314405 19715 314435
rect 19845 314405 19875 314435
rect 19685 314325 19715 314355
rect 19845 314325 19875 314355
rect 19685 314245 19715 314275
rect 19845 314245 19875 314275
rect 19685 314165 19715 314195
rect 19845 314165 19875 314195
rect 19685 314085 19715 314115
rect 19845 314085 19875 314115
rect 19685 314005 19715 314035
rect 19845 314005 19875 314035
rect 19685 313925 19715 313955
rect 19845 313925 19875 313955
rect 19685 313845 19715 313875
rect 19845 313845 19875 313875
rect 19685 313765 19715 313795
rect 19845 313765 19875 313795
rect 19685 313685 19715 313715
rect 19845 313685 19875 313715
rect 19685 313605 19715 313635
rect 19845 313605 19875 313635
rect 19685 313525 19715 313555
rect 19845 313525 19875 313555
rect 19685 313445 19715 313475
rect 19845 313445 19875 313475
rect 19685 313365 19715 313395
rect 19845 313365 19875 313395
rect 19685 313285 19715 313315
rect 19845 313285 19875 313315
rect 19685 313205 19715 313235
rect 19845 313205 19875 313235
rect 19685 313125 19715 313155
rect 19845 313125 19875 313155
rect 19685 313045 19715 313075
rect 19845 313045 19875 313075
rect 19685 312965 19715 312995
rect 19845 312965 19875 312995
rect 19685 312885 19715 312915
rect 19845 312885 19875 312915
rect 19685 312805 19715 312835
rect 19845 312805 19875 312835
rect 19685 312725 19715 312755
rect 19845 312725 19875 312755
rect 19685 312645 19715 312675
rect 19845 312645 19875 312675
rect 19685 312565 19715 312595
rect 19845 312565 19875 312595
rect 19685 312485 19715 312515
rect 19845 312485 19875 312515
rect 19685 312405 19715 312435
rect 19845 312405 19875 312435
rect 19685 312325 19715 312355
rect 19845 312325 19875 312355
rect 19685 312245 19715 312275
rect 19845 312245 19875 312275
rect 19685 312165 19715 312195
rect 19845 312165 19875 312195
rect 19685 312085 19715 312115
rect 19845 312085 19875 312115
rect 19685 312005 19715 312035
rect 19845 312005 19875 312035
rect 19685 311925 19715 311955
rect 19845 311925 19875 311955
rect 19685 311845 19715 311875
rect 19845 311845 19875 311875
rect 19685 311765 19715 311795
rect 19845 311765 19875 311795
rect 19685 311685 19715 311715
rect 19845 311685 19875 311715
rect 19685 311605 19715 311635
rect 19845 311605 19875 311635
rect 19685 311525 19715 311555
rect 19845 311525 19875 311555
rect 19685 311445 19715 311475
rect 19845 311445 19875 311475
rect 19685 311365 19715 311395
rect 19845 311365 19875 311395
rect 19685 311285 19715 311315
rect 19845 311285 19875 311315
rect 19685 311205 19715 311235
rect 19845 311205 19875 311235
rect 19685 311125 19715 311155
rect 19845 311125 19875 311155
rect 19685 311045 19715 311075
rect 19845 311045 19875 311075
rect 19685 310965 19715 310995
rect 19845 310965 19875 310995
rect 19685 310885 19715 310915
rect 19845 310885 19875 310915
rect 19685 310805 19715 310835
rect 19845 310805 19875 310835
rect 19685 310725 19715 310755
rect 19845 310725 19875 310755
rect 19685 310645 19715 310675
rect 19845 310645 19875 310675
rect 19685 310565 19715 310595
rect 19845 310565 19875 310595
rect 19685 310485 19715 310515
rect 19845 310485 19875 310515
rect 19685 310405 19715 310435
rect 19845 310405 19875 310435
rect 19685 310325 19715 310355
rect 19845 310325 19875 310355
rect 19685 310245 19715 310275
rect 19845 310245 19875 310275
rect 19685 310165 19715 310195
rect 19845 310165 19875 310195
rect 19685 310085 19715 310115
rect 19845 310085 19875 310115
rect 19685 310005 19715 310035
rect 19845 310005 19875 310035
rect 19685 309925 19715 309955
rect 19845 309925 19875 309955
rect 19685 309845 19715 309875
rect 19845 309845 19875 309875
rect 19685 309765 19715 309795
rect 19845 309765 19875 309795
rect 19685 309685 19715 309715
rect 19845 309685 19875 309715
rect 19685 309605 19715 309635
rect 19845 309605 19875 309635
rect 19685 309525 19715 309555
rect 19845 309525 19875 309555
rect 19685 309445 19715 309475
rect 19845 309445 19875 309475
rect 19685 309365 19715 309395
rect 19845 309365 19875 309395
rect 19685 309285 19715 309315
rect 19845 309285 19875 309315
rect 19685 309205 19715 309235
rect 19845 309205 19875 309235
rect 19685 309125 19715 309155
rect 19845 309125 19875 309155
rect 19685 309045 19715 309075
rect 19845 309045 19875 309075
rect 19685 308965 19715 308995
rect 19845 308965 19875 308995
rect 19685 308885 19715 308915
rect 19845 308885 19875 308915
rect 19685 308805 19715 308835
rect 19845 308805 19875 308835
rect 19685 308725 19715 308755
rect 19845 308725 19875 308755
rect 19685 308645 19715 308675
rect 19845 308645 19875 308675
rect 19685 308565 19715 308595
rect 19845 308565 19875 308595
rect 19685 308485 19715 308515
rect 19845 308485 19875 308515
rect 19685 308405 19715 308435
rect 19845 308405 19875 308435
rect 19685 308325 19715 308355
rect 19845 308325 19875 308355
rect 19685 308245 19715 308275
rect 19845 308245 19875 308275
rect 19685 308165 19715 308195
rect 19845 308165 19875 308195
rect 19685 308085 19715 308115
rect 19845 308085 19875 308115
rect 19685 308005 19715 308035
rect 19845 308005 19875 308035
rect 19685 307925 19715 307955
rect 19845 307925 19875 307955
rect 19685 307845 19715 307875
rect 19845 307845 19875 307875
rect 19685 307765 19715 307795
rect 19845 307765 19875 307795
rect 19685 307685 19715 307715
rect 19845 307685 19875 307715
rect 19685 307605 19715 307635
rect 19845 307605 19875 307635
rect 19685 307525 19715 307555
rect 19845 307525 19875 307555
rect 19685 307445 19715 307475
rect 19845 307445 19875 307475
rect 19685 307365 19715 307395
rect 19845 307365 19875 307395
rect 19685 307285 19715 307315
rect 19845 307285 19875 307315
rect 19685 307205 19715 307235
rect 19845 307205 19875 307235
rect 19685 307125 19715 307155
rect 19845 307125 19875 307155
rect 19685 307045 19715 307075
rect 19845 307045 19875 307075
rect 19685 306965 19715 306995
rect 19845 306965 19875 306995
rect 19685 306885 19715 306915
rect 19845 306885 19875 306915
rect 19685 306805 19715 306835
rect 19845 306805 19875 306835
rect 19685 306725 19715 306755
rect 19845 306725 19875 306755
rect 19685 306645 19715 306675
rect 19845 306645 19875 306675
rect 19685 306565 19715 306595
rect 19845 306565 19875 306595
rect 19685 306485 19715 306515
rect 19845 306485 19875 306515
rect 19685 306405 19715 306435
rect 19845 306405 19875 306435
rect 19685 306325 19715 306355
rect 19845 306325 19875 306355
rect 19685 306245 19715 306275
rect 19845 306245 19875 306275
rect 19685 306165 19715 306195
rect 19845 306165 19875 306195
rect 19685 306085 19715 306115
rect 19845 306085 19875 306115
rect 19685 306005 19715 306035
rect 19845 306005 19875 306035
rect 19685 305925 19715 305955
rect 19845 305925 19875 305955
rect 19685 305845 19715 305875
rect 19845 305845 19875 305875
rect 19685 305765 19715 305795
rect 19845 305765 19875 305795
rect 19685 305685 19715 305715
rect 19845 305685 19875 305715
rect 19685 305605 19715 305635
rect 19845 305605 19875 305635
rect 19685 305525 19715 305555
rect 19845 305525 19875 305555
rect 19685 305445 19715 305475
rect 19845 305445 19875 305475
rect 19685 305365 19715 305395
rect 19845 305365 19875 305395
rect 19685 305285 19715 305315
rect 19845 305285 19875 305315
rect 19685 305205 19715 305235
rect 19845 305205 19875 305235
rect 19685 305125 19715 305155
rect 19845 305125 19875 305155
rect 19685 305045 19715 305075
rect 19845 305045 19875 305075
rect 19685 304965 19715 304995
rect 19845 304965 19875 304995
rect 19685 304885 19715 304915
rect 19845 304885 19875 304915
rect 19685 304805 19715 304835
rect 19845 304805 19875 304835
rect 19685 304725 19715 304755
rect 19845 304725 19875 304755
rect 19685 304645 19715 304675
rect 19845 304645 19875 304675
rect 19685 304565 19715 304595
rect 19845 304565 19875 304595
rect 19685 304485 19715 304515
rect 19845 304485 19875 304515
rect 19685 304405 19715 304435
rect 19845 304405 19875 304435
rect 19685 304325 19715 304355
rect 19845 304325 19875 304355
rect 19685 304245 19715 304275
rect 19845 304245 19875 304275
rect 19685 304165 19715 304195
rect 19845 304165 19875 304195
rect 19685 304085 19715 304115
rect 19845 304085 19875 304115
rect 19685 304005 19715 304035
rect 19845 304005 19875 304035
rect 19685 303925 19715 303955
rect 19845 303925 19875 303955
rect 19685 303845 19715 303875
rect 19845 303845 19875 303875
rect 19685 303765 19715 303795
rect 19845 303765 19875 303795
rect 19685 303685 19715 303715
rect 19845 303685 19875 303715
rect 19685 303605 19715 303635
rect 19845 303605 19875 303635
rect 19685 303525 19715 303555
rect 19845 303525 19875 303555
rect 19685 303445 19715 303475
rect 19845 303445 19875 303475
rect 19685 303365 19715 303395
rect 19845 303365 19875 303395
rect 19685 303285 19715 303315
rect 19845 303285 19875 303315
rect 19685 303205 19715 303235
rect 19845 303205 19875 303235
rect 19685 303125 19715 303155
rect 19845 303125 19875 303155
rect 19685 303045 19715 303075
rect 19845 303045 19875 303075
rect 19685 302965 19715 302995
rect 19845 302965 19875 302995
rect 19685 302885 19715 302915
rect 19845 302885 19875 302915
rect 19685 302805 19715 302835
rect 19845 302805 19875 302835
rect 19685 302725 19715 302755
rect 19845 302725 19875 302755
rect 19685 302645 19715 302675
rect 19845 302645 19875 302675
rect 19685 302565 19715 302595
rect 19845 302565 19875 302595
rect 19685 302485 19715 302515
rect 19845 302485 19875 302515
rect 19685 302405 19715 302435
rect 19845 302405 19875 302435
rect 19685 302325 19715 302355
rect 19845 302325 19875 302355
rect 19685 302245 19715 302275
rect 19845 302245 19875 302275
rect 19685 302165 19715 302195
rect 19845 302165 19875 302195
rect 19685 302085 19715 302115
rect 19845 302085 19875 302115
rect 19685 302005 19715 302035
rect 19845 302005 19875 302035
rect 19685 301925 19715 301955
rect 19845 301925 19875 301955
rect 19685 301845 19715 301875
rect 19845 301845 19875 301875
rect 19685 301765 19715 301795
rect 19845 301765 19875 301795
rect 19685 301685 19715 301715
rect 19845 301685 19875 301715
rect 19685 301605 19715 301635
rect 19845 301605 19875 301635
rect 19685 301525 19715 301555
rect 19845 301525 19875 301555
rect 19685 301445 19715 301475
rect 19845 301445 19875 301475
rect 19685 301365 19715 301395
rect 19845 301365 19875 301395
rect 19685 301285 19715 301315
rect 19845 301285 19875 301315
rect 19685 301205 19715 301235
rect 19845 301205 19875 301235
rect 19685 301125 19715 301155
rect 19845 301125 19875 301155
rect 19685 301045 19715 301075
rect 19845 301045 19875 301075
rect 19685 300965 19715 300995
rect 19845 300965 19875 300995
rect 19685 300885 19715 300915
rect 19845 300885 19875 300915
rect 19685 300805 19715 300835
rect 19845 300805 19875 300835
rect 19685 300725 19715 300755
rect 19845 300725 19875 300755
rect 19685 300645 19715 300675
rect 19845 300645 19875 300675
rect 19685 300565 19715 300595
rect 19845 300565 19875 300595
rect 19685 300485 19715 300515
rect 19845 300485 19875 300515
rect 19685 300405 19715 300435
rect 19845 300405 19875 300435
rect 19685 300325 19715 300355
rect 19845 300325 19875 300355
rect 19685 300245 19715 300275
rect 19845 300245 19875 300275
rect 19685 300165 19715 300195
rect 19845 300165 19875 300195
rect 19685 300085 19715 300115
rect 19845 300085 19875 300115
rect 19685 300005 19715 300035
rect 19845 300005 19875 300035
rect 19685 299925 19715 299955
rect 19845 299925 19875 299955
rect 19685 299845 19715 299875
rect 19845 299845 19875 299875
rect 19685 299765 19715 299795
rect 19845 299765 19875 299795
rect 19685 299685 19715 299715
rect 19845 299685 19875 299715
rect 19685 299605 19715 299635
rect 19845 299605 19875 299635
rect 19685 299525 19715 299555
rect 19845 299525 19875 299555
rect 19685 299445 19715 299475
rect 19845 299445 19875 299475
rect 19685 299365 19715 299395
rect 19845 299365 19875 299395
rect 19685 299285 19715 299315
rect 19845 299285 19875 299315
rect 19685 299205 19715 299235
rect 19845 299205 19875 299235
rect 19685 299125 19715 299155
rect 19845 299125 19875 299155
rect 19685 299045 19715 299075
rect 19845 299045 19875 299075
rect 19685 298965 19715 298995
rect 19845 298965 19875 298995
rect 19685 298885 19715 298915
rect 19845 298885 19875 298915
rect 19685 298805 19715 298835
rect 19845 298805 19875 298835
rect 19685 298725 19715 298755
rect 19845 298725 19875 298755
rect 19685 298645 19715 298675
rect 19845 298645 19875 298675
rect 19685 298565 19715 298595
rect 19845 298565 19875 298595
rect 19685 298485 19715 298515
rect 19845 298485 19875 298515
rect 19685 298405 19715 298435
rect 19845 298405 19875 298435
rect 19685 298325 19715 298355
rect 19845 298325 19875 298355
rect 19685 298245 19715 298275
rect 19845 298245 19875 298275
rect 19685 298165 19715 298195
rect 19845 298165 19875 298195
rect 19685 298085 19715 298115
rect 19845 298085 19875 298115
rect 19685 298005 19715 298035
rect 19845 298005 19875 298035
rect 19685 297925 19715 297955
rect 19845 297925 19875 297955
rect 19685 297845 19715 297875
rect 19845 297845 19875 297875
rect 19685 297765 19715 297795
rect 19845 297765 19875 297795
rect 19685 297685 19715 297715
rect 19845 297685 19875 297715
rect 19685 297605 19715 297635
rect 19845 297605 19875 297635
rect 19685 297525 19715 297555
rect 19845 297525 19875 297555
rect 19685 297445 19715 297475
rect 19845 297445 19875 297475
rect 19685 297365 19715 297395
rect 19845 297365 19875 297395
rect 19685 297285 19715 297315
rect 19845 297285 19875 297315
rect 19685 297205 19715 297235
rect 19845 297205 19875 297235
rect 19685 297125 19715 297155
rect 19845 297125 19875 297155
rect 19685 297045 19715 297075
rect 19845 297045 19875 297075
rect 19685 296965 19715 296995
rect 19845 296965 19875 296995
rect 19685 296885 19715 296915
rect 19845 296885 19875 296915
rect 19685 296805 19715 296835
rect 19845 296805 19875 296835
rect 19685 296725 19715 296755
rect 19845 296725 19875 296755
rect 19685 296645 19715 296675
rect 19845 296645 19875 296675
rect 19685 296565 19715 296595
rect 19845 296565 19875 296595
rect 19685 296485 19715 296515
rect 19845 296485 19875 296515
rect 19685 296405 19715 296435
rect 19845 296405 19875 296435
rect 19685 296325 19715 296355
rect 19845 296325 19875 296355
rect 19685 296245 19715 296275
rect 19845 296245 19875 296275
rect 19685 296165 19715 296195
rect 19845 296165 19875 296195
rect 19685 296085 19715 296115
rect 19845 296085 19875 296115
rect 19685 296005 19715 296035
rect 19845 296005 19875 296035
rect 19685 295925 19715 295955
rect 19845 295925 19875 295955
rect 19685 295845 19715 295875
rect 19845 295845 19875 295875
rect 19685 295765 19715 295795
rect 19845 295765 19875 295795
rect 19685 295685 19715 295715
rect 19845 295685 19875 295715
rect 19685 295605 19715 295635
rect 19845 295605 19875 295635
rect 19685 295525 19715 295555
rect 19845 295525 19875 295555
rect 19685 295445 19715 295475
rect 19845 295445 19875 295475
rect 19685 295365 19715 295395
rect 19845 295365 19875 295395
rect 19685 295285 19715 295315
rect 19845 295285 19875 295315
rect 19685 295205 19715 295235
rect 19845 295205 19875 295235
rect 19685 295125 19715 295155
rect 19845 295125 19875 295155
rect 19685 295045 19715 295075
rect 19845 295045 19875 295075
rect 19685 294965 19715 294995
rect 19845 294965 19875 294995
rect 19685 294885 19715 294915
rect 19845 294885 19875 294915
rect 19685 294805 19715 294835
rect 19845 294805 19875 294835
rect 19685 294725 19715 294755
rect 19845 294725 19875 294755
rect 19685 294645 19715 294675
rect 19845 294645 19875 294675
rect 19685 294565 19715 294595
rect 19845 294565 19875 294595
rect 19685 294485 19715 294515
rect 19845 294485 19875 294515
rect 19685 294405 19715 294435
rect 19845 294405 19875 294435
rect 19685 294325 19715 294355
rect 19845 294325 19875 294355
rect 19685 294245 19715 294275
rect 19845 294245 19875 294275
rect 19685 294165 19715 294195
rect 19845 294165 19875 294195
rect 19685 294085 19715 294115
rect 19845 294085 19875 294115
rect 19685 294005 19715 294035
rect 19845 294005 19875 294035
rect 19685 293925 19715 293955
rect 19845 293925 19875 293955
rect 19685 293845 19715 293875
rect 19845 293845 19875 293875
rect 19685 293765 19715 293795
rect 19845 293765 19875 293795
rect 19685 293685 19715 293715
rect 19845 293685 19875 293715
rect 19685 293605 19715 293635
rect 19845 293605 19875 293635
rect 19685 293525 19715 293555
rect 19845 293525 19875 293555
rect 19685 293445 19715 293475
rect 19845 293445 19875 293475
rect 19685 293365 19715 293395
rect 19845 293365 19875 293395
rect 19685 293285 19715 293315
rect 19845 293285 19875 293315
rect 19685 293205 19715 293235
rect 19845 293205 19875 293235
rect 19685 293125 19715 293155
rect 19845 293125 19875 293155
rect 19685 293045 19715 293075
rect 19845 293045 19875 293075
rect 19685 292965 19715 292995
rect 19845 292965 19875 292995
rect 19685 292885 19715 292915
rect 19845 292885 19875 292915
rect 19685 292805 19715 292835
rect 19845 292805 19875 292835
rect 19685 292725 19715 292755
rect 19845 292725 19875 292755
rect 19685 292645 19715 292675
rect 19845 292645 19875 292675
rect 19685 292565 19715 292595
rect 19845 292565 19875 292595
rect 19685 292485 19715 292515
rect 19845 292485 19875 292515
rect 19685 292405 19715 292435
rect 19845 292405 19875 292435
rect 19685 292325 19715 292355
rect 19845 292325 19875 292355
rect 19685 292245 19715 292275
rect 19845 292245 19875 292275
rect 19685 292165 19715 292195
rect 19845 292165 19875 292195
rect 19685 292085 19715 292115
rect 19845 292085 19875 292115
rect 19685 292005 19715 292035
rect 19845 292005 19875 292035
rect 19685 291925 19715 291955
rect 19845 291925 19875 291955
rect 19685 291845 19715 291875
rect 19845 291845 19875 291875
rect 19685 291765 19715 291795
rect 19845 291765 19875 291795
rect 19685 291685 19715 291715
rect 19845 291685 19875 291715
rect 19685 291605 19715 291635
rect 19845 291605 19875 291635
rect 19685 291525 19715 291555
rect 19845 291525 19875 291555
rect 19685 291445 19715 291475
rect 19845 291445 19875 291475
rect 19685 291365 19715 291395
rect 19845 291365 19875 291395
rect 19685 291285 19715 291315
rect 19845 291285 19875 291315
rect 19685 291205 19715 291235
rect 19845 291205 19875 291235
rect 19685 291125 19715 291155
rect 19845 291125 19875 291155
rect 19685 291045 19715 291075
rect 19845 291045 19875 291075
rect 19685 290965 19715 290995
rect 19845 290965 19875 290995
rect 19685 290885 19715 290915
rect 19845 290885 19875 290915
rect 19685 290805 19715 290835
rect 19845 290805 19875 290835
rect 19685 290725 19715 290755
rect 19845 290725 19875 290755
rect 19685 290645 19715 290675
rect 19845 290645 19875 290675
rect 19685 290565 19715 290595
rect 19845 290565 19875 290595
rect 19685 290485 19715 290515
rect 19845 290485 19875 290515
rect 19685 290405 19715 290435
rect 19845 290405 19875 290435
rect 19685 290325 19715 290355
rect 19845 290325 19875 290355
rect 19685 290245 19715 290275
rect 19845 290245 19875 290275
rect 19685 290165 19715 290195
rect 19845 290165 19875 290195
rect 19685 290085 19715 290115
rect 19845 290085 19875 290115
rect 19685 290005 19715 290035
rect 19845 290005 19875 290035
rect 19685 289925 19715 289955
rect 19845 289925 19875 289955
rect 19685 289845 19715 289875
rect 19845 289845 19875 289875
rect 19685 289765 19715 289795
rect 19845 289765 19875 289795
rect 19685 289685 19715 289715
rect 19845 289685 19875 289715
rect 19685 289605 19715 289635
rect 19845 289605 19875 289635
rect 19685 289525 19715 289555
rect 19845 289525 19875 289555
rect 19685 289445 19715 289475
rect 19845 289445 19875 289475
rect 19685 289365 19715 289395
rect 19845 289365 19875 289395
rect 19685 289285 19715 289315
rect 19845 289285 19875 289315
rect 19685 289205 19715 289235
rect 19845 289205 19875 289235
rect 19685 289125 19715 289155
rect 19845 289125 19875 289155
rect 19685 289045 19715 289075
rect 19845 289045 19875 289075
rect 19685 288965 19715 288995
rect 19845 288965 19875 288995
rect 19685 288885 19715 288915
rect 19845 288885 19875 288915
rect 19685 288805 19715 288835
rect 19845 288805 19875 288835
rect 19685 288725 19715 288755
rect 19845 288725 19875 288755
rect 19685 288645 19715 288675
rect 19845 288645 19875 288675
rect 19685 288565 19715 288595
rect 19845 288565 19875 288595
rect 19685 288485 19715 288515
rect 19845 288485 19875 288515
rect 19685 288405 19715 288435
rect 19845 288405 19875 288435
rect 19685 288325 19715 288355
rect 19845 288325 19875 288355
rect 19685 288245 19715 288275
rect 19845 288245 19875 288275
rect 19685 288165 19715 288195
rect 19845 288165 19875 288195
rect 19685 288085 19715 288115
rect 19845 288085 19875 288115
rect 19685 288005 19715 288035
rect 19845 288005 19875 288035
rect 19685 287925 19715 287955
rect 19845 287925 19875 287955
rect 19685 287845 19715 287875
rect 19845 287845 19875 287875
rect 19685 287765 19715 287795
rect 19845 287765 19875 287795
rect 19685 287685 19715 287715
rect 19845 287685 19875 287715
rect 19685 287605 19715 287635
rect 19845 287605 19875 287635
rect 19685 287525 19715 287555
rect 19845 287525 19875 287555
rect 19685 287445 19715 287475
rect 19845 287445 19875 287475
rect 19685 287365 19715 287395
rect 19845 287365 19875 287395
rect 19685 287285 19715 287315
rect 19845 287285 19875 287315
rect 19685 287205 19715 287235
rect 19845 287205 19875 287235
rect 19685 287125 19715 287155
rect 19845 287125 19875 287155
rect 19685 287045 19715 287075
rect 19845 287045 19875 287075
rect 19685 286965 19715 286995
rect 19845 286965 19875 286995
rect 19685 286885 19715 286915
rect 19845 286885 19875 286915
rect 19685 286805 19715 286835
rect 19845 286805 19875 286835
rect 19685 286725 19715 286755
rect 19845 286725 19875 286755
rect 19685 286645 19715 286675
rect 19845 286645 19875 286675
rect 19685 286565 19715 286595
rect 19845 286565 19875 286595
rect 19685 286485 19715 286515
rect 19845 286485 19875 286515
rect 19685 286405 19715 286435
rect 19845 286405 19875 286435
rect 19685 286325 19715 286355
rect 19845 286325 19875 286355
rect 19685 286245 19715 286275
rect 19845 286245 19875 286275
rect 19685 286165 19715 286195
rect 19845 286165 19875 286195
rect 19685 286085 19715 286115
rect 19845 286085 19875 286115
rect 19685 286005 19715 286035
rect 19845 286005 19875 286035
rect 19685 285925 19715 285955
rect 19845 285925 19875 285955
rect 19685 285845 19715 285875
rect 19845 285845 19875 285875
rect 19685 285765 19715 285795
rect 19845 285765 19875 285795
rect 19685 285685 19715 285715
rect 19845 285685 19875 285715
rect 19685 285605 19715 285635
rect 19845 285605 19875 285635
rect 19685 285525 19715 285555
rect 19845 285525 19875 285555
rect 19685 285445 19715 285475
rect 19845 285445 19875 285475
rect 19685 285365 19715 285395
rect 19845 285365 19875 285395
rect 19685 285285 19715 285315
rect 19845 285285 19875 285315
rect 19685 285205 19715 285235
rect 19845 285205 19875 285235
rect 19685 285125 19715 285155
rect 19845 285125 19875 285155
rect 19685 285045 19715 285075
rect 19845 285045 19875 285075
rect 19685 284965 19715 284995
rect 19845 284965 19875 284995
rect 19685 284885 19715 284915
rect 19845 284885 19875 284915
rect 19685 284805 19715 284835
rect 19845 284805 19875 284835
rect 19685 284725 19715 284755
rect 19845 284725 19875 284755
rect 19685 284645 19715 284675
rect 19845 284645 19875 284675
rect 19685 284565 19715 284595
rect 19845 284565 19875 284595
rect 19685 284485 19715 284515
rect 19845 284485 19875 284515
rect 19685 284405 19715 284435
rect 19845 284405 19875 284435
rect 19685 284325 19715 284355
rect 19845 284325 19875 284355
rect 19685 284245 19715 284275
rect 19845 284245 19875 284275
rect 19685 284165 19715 284195
rect 19845 284165 19875 284195
rect 19685 284085 19715 284115
rect 19845 284085 19875 284115
rect 19685 284005 19715 284035
rect 19845 284005 19875 284035
rect 19685 283925 19715 283955
rect 19845 283925 19875 283955
rect 19685 283845 19715 283875
rect 19845 283845 19875 283875
rect 19685 283765 19715 283795
rect 19845 283765 19875 283795
rect 19685 283685 19715 283715
rect 19845 283685 19875 283715
rect 19685 283605 19715 283635
rect 19845 283605 19875 283635
rect 19685 283525 19715 283555
rect 19845 283525 19875 283555
rect 19685 283445 19715 283475
rect 19845 283445 19875 283475
rect 19685 283365 19715 283395
rect 19845 283365 19875 283395
rect 19685 283285 19715 283315
rect 19845 283285 19875 283315
rect 19685 283205 19715 283235
rect 19845 283205 19875 283235
rect 19685 283125 19715 283155
rect 19845 283125 19875 283155
rect 19685 283045 19715 283075
rect 19845 283045 19875 283075
rect 19685 282965 19715 282995
rect 19845 282965 19875 282995
rect 19685 282885 19715 282915
rect 19845 282885 19875 282915
rect 19685 282805 19715 282835
rect 19845 282805 19875 282835
rect 19685 282725 19715 282755
rect 19845 282725 19875 282755
rect 19685 282645 19715 282675
rect 19845 282645 19875 282675
rect 19685 282565 19715 282595
rect 19845 282565 19875 282595
rect 19685 282485 19715 282515
rect 19845 282485 19875 282515
rect 19685 282405 19715 282435
rect 19845 282405 19875 282435
rect 19685 282325 19715 282355
rect 19845 282325 19875 282355
rect 19685 282245 19715 282275
rect 19845 282245 19875 282275
rect 19685 282165 19715 282195
rect 19845 282165 19875 282195
rect 19685 282085 19715 282115
rect 19845 282085 19875 282115
rect 19685 282005 19715 282035
rect 19845 282005 19875 282035
rect 19685 281925 19715 281955
rect 19845 281925 19875 281955
rect 19685 281845 19715 281875
rect 19845 281845 19875 281875
rect 19685 281765 19715 281795
rect 19845 281765 19875 281795
rect 19685 281685 19715 281715
rect 19845 281685 19875 281715
rect 19685 281605 19715 281635
rect 19845 281605 19875 281635
rect 19685 281525 19715 281555
rect 19845 281525 19875 281555
rect 19685 281445 19715 281475
rect 19845 281445 19875 281475
rect 19685 281365 19715 281395
rect 19845 281365 19875 281395
rect 19685 281285 19715 281315
rect 19845 281285 19875 281315
rect 19685 281205 19715 281235
rect 19845 281205 19875 281235
rect 19685 281125 19715 281155
rect 19845 281125 19875 281155
rect 19685 281045 19715 281075
rect 19845 281045 19875 281075
rect 19685 280965 19715 280995
rect 19845 280965 19875 280995
rect 19685 280885 19715 280915
rect 19845 280885 19875 280915
rect 19685 280805 19715 280835
rect 19845 280805 19875 280835
rect 19685 280725 19715 280755
rect 19845 280725 19875 280755
rect 19685 280645 19715 280675
rect 19845 280645 19875 280675
rect 19685 280565 19715 280595
rect 19845 280565 19875 280595
rect 19685 280485 19715 280515
rect 19845 280485 19875 280515
rect 19685 280405 19715 280435
rect 19845 280405 19875 280435
rect 19685 280325 19715 280355
rect 19845 280325 19875 280355
rect 19685 280245 19715 280275
rect 19845 280245 19875 280275
rect 19685 280165 19715 280195
rect 19845 280165 19875 280195
rect 19685 280085 19715 280115
rect 19845 280085 19875 280115
rect 19685 280005 19715 280035
rect 19845 280005 19875 280035
rect 19685 279925 19715 279955
rect 19845 279925 19875 279955
rect 19685 279845 19715 279875
rect 19845 279845 19875 279875
rect 19685 279765 19715 279795
rect 19845 279765 19875 279795
rect 19685 279685 19715 279715
rect 19845 279685 19875 279715
rect 19685 279605 19715 279635
rect 19845 279605 19875 279635
rect 19685 279525 19715 279555
rect 19845 279525 19875 279555
rect 19685 279445 19715 279475
rect 19845 279445 19875 279475
rect 19685 279365 19715 279395
rect 19845 279365 19875 279395
rect 19685 279285 19715 279315
rect 19845 279285 19875 279315
rect 19685 279205 19715 279235
rect 19845 279205 19875 279235
rect 19685 279125 19715 279155
rect 19845 279125 19875 279155
rect 19685 279045 19715 279075
rect 19845 279045 19875 279075
rect 19685 278965 19715 278995
rect 19845 278965 19875 278995
rect 19685 278885 19715 278915
rect 19845 278885 19875 278915
rect 19685 278805 19715 278835
rect 19845 278805 19875 278835
rect 19685 278725 19715 278755
rect 19845 278725 19875 278755
rect 17045 278645 17075 278675
rect 17205 278645 17235 278675
rect 17285 278645 17315 278675
rect 17365 278645 17395 278675
rect 17445 278645 17475 278675
rect 17525 278645 17555 278675
rect 17605 278645 17635 278675
rect 17685 278645 17715 278675
rect 17765 278645 17795 278675
rect 19525 278645 19555 278675
rect 19605 278645 19635 278675
rect 19685 278645 19715 278675
rect 19845 278645 19875 278675
rect 17045 278485 17075 278515
rect 17205 278485 17235 278515
rect 17285 278485 17315 278515
rect 17365 278485 17395 278515
rect 17445 278485 17475 278515
rect 17525 278485 17555 278515
rect 17605 278485 17635 278515
rect 17685 278485 17715 278515
rect 17765 278485 17795 278515
rect 19525 278485 19555 278515
rect 19605 278485 19635 278515
rect 19685 278485 19715 278515
rect 19845 278485 19875 278515
rect 17045 278405 17075 278435
rect 17205 278405 17235 278435
rect 17045 278325 17075 278355
rect 17205 278325 17235 278355
rect 17045 278245 17075 278275
rect 17205 278245 17235 278275
rect 17045 278165 17075 278195
rect 17205 278165 17235 278195
rect 17045 278085 17075 278115
rect 17205 278085 17235 278115
rect 17045 278005 17075 278035
rect 17205 278005 17235 278035
rect 17045 277925 17075 277955
rect 17205 277925 17235 277955
rect 17045 277845 17075 277875
rect 17205 277845 17235 277875
<< metal2 >>
rect 10720 351395 19880 351400
rect 10720 351365 10725 351395
rect 10755 351365 10805 351395
rect 10835 351365 10885 351395
rect 10915 351365 10965 351395
rect 10995 351365 11045 351395
rect 11075 351365 11125 351395
rect 11155 351365 11205 351395
rect 11235 351365 11285 351395
rect 11315 351365 11365 351395
rect 11395 351365 11445 351395
rect 11475 351365 11525 351395
rect 11555 351365 11605 351395
rect 11635 351365 11685 351395
rect 11715 351365 11765 351395
rect 11795 351365 11845 351395
rect 11875 351365 11925 351395
rect 11955 351365 12005 351395
rect 12035 351365 12085 351395
rect 12115 351365 12165 351395
rect 12195 351365 12245 351395
rect 12275 351365 12325 351395
rect 12355 351365 12405 351395
rect 12435 351365 12485 351395
rect 12515 351365 12565 351395
rect 12595 351365 12645 351395
rect 12675 351365 12725 351395
rect 12755 351365 12805 351395
rect 12835 351365 12885 351395
rect 12915 351365 12965 351395
rect 12995 351365 13045 351395
rect 13075 351365 13125 351395
rect 13155 351365 13205 351395
rect 13235 351365 13285 351395
rect 13315 351365 13365 351395
rect 13395 351365 13445 351395
rect 13475 351365 13525 351395
rect 13555 351365 13605 351395
rect 13635 351365 13685 351395
rect 13715 351365 13765 351395
rect 13795 351365 13845 351395
rect 13875 351365 13925 351395
rect 13955 351365 14005 351395
rect 14035 351365 14085 351395
rect 14115 351365 14165 351395
rect 14195 351365 14245 351395
rect 14275 351365 14325 351395
rect 14355 351365 14405 351395
rect 14435 351365 14485 351395
rect 14515 351365 14565 351395
rect 14595 351365 14645 351395
rect 14675 351365 14725 351395
rect 14755 351365 14805 351395
rect 14835 351365 14885 351395
rect 14915 351365 14965 351395
rect 14995 351365 15045 351395
rect 15075 351365 15125 351395
rect 15155 351365 15205 351395
rect 15235 351365 15285 351395
rect 15315 351365 15365 351395
rect 15395 351365 15445 351395
rect 15475 351365 15525 351395
rect 15555 351365 15605 351395
rect 15635 351365 15685 351395
rect 15715 351365 15765 351395
rect 15795 351365 15845 351395
rect 15875 351365 15925 351395
rect 15955 351365 16005 351395
rect 16035 351365 16085 351395
rect 16115 351365 16165 351395
rect 16195 351365 16245 351395
rect 16275 351365 16325 351395
rect 16355 351365 16405 351395
rect 16435 351365 16485 351395
rect 16515 351365 16565 351395
rect 16595 351365 16645 351395
rect 16675 351365 16725 351395
rect 16755 351365 16805 351395
rect 16835 351365 16885 351395
rect 16915 351365 16965 351395
rect 16995 351365 17045 351395
rect 17075 351365 17125 351395
rect 17155 351365 17205 351395
rect 17235 351365 17285 351395
rect 17315 351365 17365 351395
rect 17395 351365 17445 351395
rect 17475 351365 17525 351395
rect 17555 351365 17605 351395
rect 17635 351365 17685 351395
rect 17715 351365 17765 351395
rect 17795 351365 17845 351395
rect 17875 351365 17925 351395
rect 17955 351365 18005 351395
rect 18035 351365 18085 351395
rect 18115 351365 18165 351395
rect 18195 351365 18245 351395
rect 18275 351365 18325 351395
rect 18355 351365 18405 351395
rect 18435 351365 18485 351395
rect 18515 351365 18565 351395
rect 18595 351365 18645 351395
rect 18675 351365 18725 351395
rect 18755 351365 18805 351395
rect 18835 351365 18885 351395
rect 18915 351365 18965 351395
rect 18995 351365 19045 351395
rect 19075 351365 19125 351395
rect 19155 351365 19205 351395
rect 19235 351365 19285 351395
rect 19315 351365 19365 351395
rect 19395 351365 19445 351395
rect 19475 351365 19525 351395
rect 19555 351365 19605 351395
rect 19635 351365 19685 351395
rect 19715 351365 19845 351395
rect 19875 351365 19880 351395
rect 10720 351360 19880 351365
rect 10640 351315 19800 351320
rect 10640 351285 10645 351315
rect 10675 351285 19765 351315
rect 19795 351285 19800 351315
rect 10640 351280 19800 351285
rect 10720 351235 19880 351240
rect 10720 351205 10725 351235
rect 10755 351205 10805 351235
rect 10835 351205 10885 351235
rect 10915 351205 10965 351235
rect 10995 351205 11045 351235
rect 11075 351205 11125 351235
rect 11155 351205 11205 351235
rect 11235 351205 11285 351235
rect 11315 351205 11365 351235
rect 11395 351205 11445 351235
rect 11475 351205 11525 351235
rect 11555 351205 11605 351235
rect 11635 351205 11685 351235
rect 11715 351205 11765 351235
rect 11795 351205 11845 351235
rect 11875 351205 11925 351235
rect 11955 351205 12005 351235
rect 12035 351205 12085 351235
rect 12115 351205 12165 351235
rect 12195 351205 12245 351235
rect 12275 351205 12325 351235
rect 12355 351205 12405 351235
rect 12435 351205 12485 351235
rect 12515 351205 12565 351235
rect 12595 351205 12645 351235
rect 12675 351205 12725 351235
rect 12755 351205 12805 351235
rect 12835 351205 12885 351235
rect 12915 351205 12965 351235
rect 12995 351205 13045 351235
rect 13075 351205 13125 351235
rect 13155 351205 13205 351235
rect 13235 351205 13285 351235
rect 13315 351205 13365 351235
rect 13395 351205 13445 351235
rect 13475 351205 13525 351235
rect 13555 351205 13605 351235
rect 13635 351205 13685 351235
rect 13715 351205 13765 351235
rect 13795 351205 13845 351235
rect 13875 351205 13925 351235
rect 13955 351205 14005 351235
rect 14035 351205 14085 351235
rect 14115 351205 14165 351235
rect 14195 351205 14245 351235
rect 14275 351205 14325 351235
rect 14355 351205 14405 351235
rect 14435 351205 14485 351235
rect 14515 351205 14565 351235
rect 14595 351205 14645 351235
rect 14675 351205 14725 351235
rect 14755 351205 14805 351235
rect 14835 351205 14885 351235
rect 14915 351205 14965 351235
rect 14995 351205 15045 351235
rect 15075 351205 15125 351235
rect 15155 351205 15205 351235
rect 15235 351205 15285 351235
rect 15315 351205 15365 351235
rect 15395 351205 15445 351235
rect 15475 351205 15525 351235
rect 15555 351205 15605 351235
rect 15635 351205 15685 351235
rect 15715 351205 15765 351235
rect 15795 351205 15845 351235
rect 15875 351205 15925 351235
rect 15955 351205 16005 351235
rect 16035 351205 16085 351235
rect 16115 351205 16165 351235
rect 16195 351205 16245 351235
rect 16275 351205 16325 351235
rect 16355 351205 16405 351235
rect 16435 351205 16485 351235
rect 16515 351205 16565 351235
rect 16595 351205 16645 351235
rect 16675 351205 16725 351235
rect 16755 351205 16805 351235
rect 16835 351205 16885 351235
rect 16915 351205 16965 351235
rect 16995 351205 17045 351235
rect 17075 351205 17125 351235
rect 17155 351205 17205 351235
rect 17235 351205 17285 351235
rect 17315 351205 17365 351235
rect 17395 351205 17445 351235
rect 17475 351205 17525 351235
rect 17555 351205 17605 351235
rect 17635 351205 17685 351235
rect 17715 351205 17765 351235
rect 17795 351205 17845 351235
rect 17875 351205 17925 351235
rect 17955 351205 18005 351235
rect 18035 351205 18085 351235
rect 18115 351205 18165 351235
rect 18195 351205 18245 351235
rect 18275 351205 18325 351235
rect 18355 351205 18405 351235
rect 18435 351205 18485 351235
rect 18515 351205 18565 351235
rect 18595 351205 18645 351235
rect 18675 351205 18725 351235
rect 18755 351205 18805 351235
rect 18835 351205 18885 351235
rect 18915 351205 18965 351235
rect 18995 351205 19045 351235
rect 19075 351205 19125 351235
rect 19155 351205 19205 351235
rect 19235 351205 19285 351235
rect 19315 351205 19365 351235
rect 19395 351205 19445 351235
rect 19475 351205 19525 351235
rect 19555 351205 19605 351235
rect 19635 351205 19685 351235
rect 19715 351205 19845 351235
rect 19875 351205 19880 351235
rect 10720 351200 19880 351205
rect 19680 351155 19880 351160
rect 19680 351125 19685 351155
rect 19715 351125 19845 351155
rect 19875 351125 19880 351155
rect 19680 351120 19880 351125
rect 19680 351075 19880 351080
rect 19680 351045 19685 351075
rect 19715 351045 19845 351075
rect 19875 351045 19880 351075
rect 19680 351040 19880 351045
rect 19680 350995 19880 351000
rect 19680 350965 19685 350995
rect 19715 350965 19845 350995
rect 19875 350965 19880 350995
rect 19680 350960 19880 350965
rect 19680 350915 19880 350920
rect 19680 350885 19685 350915
rect 19715 350885 19845 350915
rect 19875 350885 19880 350915
rect 19680 350880 19880 350885
rect 19680 350835 19880 350840
rect 19680 350805 19685 350835
rect 19715 350805 19845 350835
rect 19875 350805 19880 350835
rect 19680 350800 19880 350805
rect 19680 350755 19880 350760
rect 19680 350725 19685 350755
rect 19715 350725 19845 350755
rect 19875 350725 19880 350755
rect 19680 350720 19880 350725
rect 19680 350675 19880 350680
rect 19680 350645 19685 350675
rect 19715 350645 19845 350675
rect 19875 350645 19880 350675
rect 19680 350640 19880 350645
rect 19680 350595 19880 350600
rect 19680 350565 19685 350595
rect 19715 350565 19845 350595
rect 19875 350565 19880 350595
rect 19680 350560 19880 350565
rect 19680 350515 19880 350520
rect 19680 350485 19685 350515
rect 19715 350485 19845 350515
rect 19875 350485 19880 350515
rect 19680 350480 19880 350485
rect 19680 350435 19880 350440
rect 19680 350405 19685 350435
rect 19715 350405 19845 350435
rect 19875 350405 19880 350435
rect 19680 350400 19880 350405
rect 19680 350355 19880 350360
rect 19680 350325 19685 350355
rect 19715 350325 19845 350355
rect 19875 350325 19880 350355
rect 19680 350320 19880 350325
rect 19680 350275 19880 350280
rect 19680 350245 19685 350275
rect 19715 350245 19845 350275
rect 19875 350245 19880 350275
rect 19680 350240 19880 350245
rect 19680 350195 19880 350200
rect 19680 350165 19685 350195
rect 19715 350165 19845 350195
rect 19875 350165 19880 350195
rect 19680 350160 19880 350165
rect 19680 350115 19880 350120
rect 19680 350085 19685 350115
rect 19715 350085 19845 350115
rect 19875 350085 19880 350115
rect 19680 350080 19880 350085
rect 19680 350035 19880 350040
rect 19680 350005 19685 350035
rect 19715 350005 19845 350035
rect 19875 350005 19880 350035
rect 19680 350000 19880 350005
rect 19680 349955 19880 349960
rect 19680 349925 19685 349955
rect 19715 349925 19845 349955
rect 19875 349925 19880 349955
rect 19680 349920 19880 349925
rect 19680 349875 19880 349880
rect 19680 349845 19685 349875
rect 19715 349845 19845 349875
rect 19875 349845 19880 349875
rect 19680 349840 19880 349845
rect 19680 349795 19880 349800
rect 19680 349765 19685 349795
rect 19715 349765 19845 349795
rect 19875 349765 19880 349795
rect 19680 349760 19880 349765
rect 19680 349715 19880 349720
rect 19680 349685 19685 349715
rect 19715 349685 19845 349715
rect 19875 349685 19880 349715
rect 19680 349680 19880 349685
rect 19680 349635 19880 349640
rect 19680 349605 19685 349635
rect 19715 349605 19845 349635
rect 19875 349605 19880 349635
rect 19680 349600 19880 349605
rect 19680 349555 19880 349560
rect 19680 349525 19685 349555
rect 19715 349525 19845 349555
rect 19875 349525 19880 349555
rect 19680 349520 19880 349525
rect 19680 349475 19880 349480
rect 19680 349445 19685 349475
rect 19715 349445 19845 349475
rect 19875 349445 19880 349475
rect 19680 349440 19880 349445
rect 19680 349395 19880 349400
rect 19680 349365 19685 349395
rect 19715 349365 19845 349395
rect 19875 349365 19880 349395
rect 19680 349360 19880 349365
rect 19680 349315 19880 349320
rect 19680 349285 19685 349315
rect 19715 349285 19845 349315
rect 19875 349285 19880 349315
rect 19680 349280 19880 349285
rect 19680 349235 19880 349240
rect 19680 349205 19685 349235
rect 19715 349205 19845 349235
rect 19875 349205 19880 349235
rect 19680 349200 19880 349205
rect 19680 349155 19880 349160
rect 19680 349125 19685 349155
rect 19715 349125 19845 349155
rect 19875 349125 19880 349155
rect 19680 349120 19880 349125
rect 19680 349075 19880 349080
rect 19680 349045 19685 349075
rect 19715 349045 19845 349075
rect 19875 349045 19880 349075
rect 19680 349040 19880 349045
rect 19680 348995 19880 349000
rect 19680 348965 19685 348995
rect 19715 348965 19845 348995
rect 19875 348965 19880 348995
rect 19680 348960 19880 348965
rect 19680 348915 19880 348920
rect 19680 348885 19685 348915
rect 19715 348885 19845 348915
rect 19875 348885 19880 348915
rect 19680 348880 19880 348885
rect 19680 348835 19880 348840
rect 19680 348805 19685 348835
rect 19715 348805 19845 348835
rect 19875 348805 19880 348835
rect 19680 348800 19880 348805
rect 19680 348755 19880 348760
rect 19680 348725 19685 348755
rect 19715 348725 19845 348755
rect 19875 348725 19880 348755
rect 19680 348720 19880 348725
rect 19680 348675 19880 348680
rect 19680 348645 19685 348675
rect 19715 348645 19845 348675
rect 19875 348645 19880 348675
rect 19680 348640 19880 348645
rect 19680 348595 19880 348600
rect 19680 348565 19685 348595
rect 19715 348565 19845 348595
rect 19875 348565 19880 348595
rect 19680 348560 19880 348565
rect 19680 348515 19880 348520
rect 19680 348485 19685 348515
rect 19715 348485 19845 348515
rect 19875 348485 19880 348515
rect 19680 348480 19880 348485
rect 19680 348435 19880 348440
rect 19680 348405 19685 348435
rect 19715 348405 19845 348435
rect 19875 348405 19880 348435
rect 19680 348400 19880 348405
rect 19680 348355 19880 348360
rect 19680 348325 19685 348355
rect 19715 348325 19845 348355
rect 19875 348325 19880 348355
rect 19680 348320 19880 348325
rect 19680 348275 19880 348280
rect 19680 348245 19685 348275
rect 19715 348245 19845 348275
rect 19875 348245 19880 348275
rect 19680 348240 19880 348245
rect 19680 348195 19880 348200
rect 19680 348165 19685 348195
rect 19715 348165 19845 348195
rect 19875 348165 19880 348195
rect 19680 348160 19880 348165
rect 19680 348115 19880 348120
rect 19680 348085 19685 348115
rect 19715 348085 19845 348115
rect 19875 348085 19880 348115
rect 19680 348080 19880 348085
rect 19680 348035 19880 348040
rect 19680 348005 19685 348035
rect 19715 348005 19845 348035
rect 19875 348005 19880 348035
rect 19680 348000 19880 348005
rect 19680 347955 19880 347960
rect 19680 347925 19685 347955
rect 19715 347925 19845 347955
rect 19875 347925 19880 347955
rect 19680 347920 19880 347925
rect 19680 347875 19880 347880
rect 19680 347845 19685 347875
rect 19715 347845 19845 347875
rect 19875 347845 19880 347875
rect 19680 347840 19880 347845
rect 19680 347795 19880 347800
rect 19680 347765 19685 347795
rect 19715 347765 19845 347795
rect 19875 347765 19880 347795
rect 19680 347760 19880 347765
rect 19680 347715 19880 347720
rect 19680 347685 19685 347715
rect 19715 347685 19845 347715
rect 19875 347685 19880 347715
rect 19680 347680 19880 347685
rect 19680 347635 19880 347640
rect 19680 347605 19685 347635
rect 19715 347605 19845 347635
rect 19875 347605 19880 347635
rect 19680 347600 19880 347605
rect 19680 347555 19880 347560
rect 19680 347525 19685 347555
rect 19715 347525 19845 347555
rect 19875 347525 19880 347555
rect 19680 347520 19880 347525
rect 19680 347475 19880 347480
rect 19680 347445 19685 347475
rect 19715 347445 19845 347475
rect 19875 347445 19880 347475
rect 19680 347440 19880 347445
rect 19680 347395 19880 347400
rect 19680 347365 19685 347395
rect 19715 347365 19845 347395
rect 19875 347365 19880 347395
rect 19680 347360 19880 347365
rect 19680 347315 19880 347320
rect 19680 347285 19685 347315
rect 19715 347285 19845 347315
rect 19875 347285 19880 347315
rect 19680 347280 19880 347285
rect 19680 347235 19880 347240
rect 19680 347205 19685 347235
rect 19715 347205 19845 347235
rect 19875 347205 19880 347235
rect 19680 347200 19880 347205
rect 19680 347155 19880 347160
rect 19680 347125 19685 347155
rect 19715 347125 19845 347155
rect 19875 347125 19880 347155
rect 19680 347120 19880 347125
rect 19680 347075 19880 347080
rect 19680 347045 19685 347075
rect 19715 347045 19845 347075
rect 19875 347045 19880 347075
rect 19680 347040 19880 347045
rect 19680 346995 19880 347000
rect 19680 346965 19685 346995
rect 19715 346965 19845 346995
rect 19875 346965 19880 346995
rect 19680 346960 19880 346965
rect 19680 346915 19880 346920
rect 19680 346885 19685 346915
rect 19715 346885 19845 346915
rect 19875 346885 19880 346915
rect 19680 346880 19880 346885
rect 19680 346835 19880 346840
rect 19680 346805 19685 346835
rect 19715 346805 19845 346835
rect 19875 346805 19880 346835
rect 19680 346800 19880 346805
rect 19680 346755 19880 346760
rect 19680 346725 19685 346755
rect 19715 346725 19845 346755
rect 19875 346725 19880 346755
rect 19680 346720 19880 346725
rect 19680 346675 19880 346680
rect 19680 346645 19685 346675
rect 19715 346645 19845 346675
rect 19875 346645 19880 346675
rect 19680 346640 19880 346645
rect 19680 346595 19880 346600
rect 19680 346565 19685 346595
rect 19715 346565 19845 346595
rect 19875 346565 19880 346595
rect 19680 346560 19880 346565
rect 19680 346515 19880 346520
rect 19680 346485 19685 346515
rect 19715 346485 19845 346515
rect 19875 346485 19880 346515
rect 19680 346480 19880 346485
rect 19680 346435 19880 346440
rect 19680 346405 19685 346435
rect 19715 346405 19845 346435
rect 19875 346405 19880 346435
rect 19680 346400 19880 346405
rect 19680 346355 19880 346360
rect 19680 346325 19685 346355
rect 19715 346325 19845 346355
rect 19875 346325 19880 346355
rect 19680 346320 19880 346325
rect 19680 346275 19880 346280
rect 19680 346245 19685 346275
rect 19715 346245 19845 346275
rect 19875 346245 19880 346275
rect 19680 346240 19880 346245
rect 19680 346195 19880 346200
rect 19680 346165 19685 346195
rect 19715 346165 19845 346195
rect 19875 346165 19880 346195
rect 19680 346160 19880 346165
rect 19680 346115 19880 346120
rect 19680 346085 19685 346115
rect 19715 346085 19845 346115
rect 19875 346085 19880 346115
rect 19680 346080 19880 346085
rect 19680 346035 19880 346040
rect 19680 346005 19685 346035
rect 19715 346005 19845 346035
rect 19875 346005 19880 346035
rect 19680 346000 19880 346005
rect 19680 345955 19880 345960
rect 19680 345925 19685 345955
rect 19715 345925 19845 345955
rect 19875 345925 19880 345955
rect 19680 345920 19880 345925
rect 19680 345875 19880 345880
rect 19680 345845 19685 345875
rect 19715 345845 19845 345875
rect 19875 345845 19880 345875
rect 19680 345840 19880 345845
rect 19680 345795 19880 345800
rect 19680 345765 19685 345795
rect 19715 345765 19845 345795
rect 19875 345765 19880 345795
rect 19680 345760 19880 345765
rect 19680 345715 19880 345720
rect 19680 345685 19685 345715
rect 19715 345685 19845 345715
rect 19875 345685 19880 345715
rect 19680 345680 19880 345685
rect 19680 345635 19880 345640
rect 19680 345605 19685 345635
rect 19715 345605 19845 345635
rect 19875 345605 19880 345635
rect 19680 345600 19880 345605
rect 19680 345555 19880 345560
rect 19680 345525 19685 345555
rect 19715 345525 19845 345555
rect 19875 345525 19880 345555
rect 19680 345520 19880 345525
rect 19680 345475 19880 345480
rect 19680 345445 19685 345475
rect 19715 345445 19845 345475
rect 19875 345445 19880 345475
rect 19680 345440 19880 345445
rect 19680 345395 19880 345400
rect 19680 345365 19685 345395
rect 19715 345365 19845 345395
rect 19875 345365 19880 345395
rect 19680 345360 19880 345365
rect 19680 345315 19880 345320
rect 19680 345285 19685 345315
rect 19715 345285 19845 345315
rect 19875 345285 19880 345315
rect 19680 345280 19880 345285
rect 19680 345235 19880 345240
rect 19680 345205 19685 345235
rect 19715 345205 19845 345235
rect 19875 345205 19880 345235
rect 19680 345200 19880 345205
rect 19680 345155 19880 345160
rect 19680 345125 19685 345155
rect 19715 345125 19845 345155
rect 19875 345125 19880 345155
rect 19680 345120 19880 345125
rect 19680 345075 19880 345080
rect 19680 345045 19685 345075
rect 19715 345045 19845 345075
rect 19875 345045 19880 345075
rect 19680 345040 19880 345045
rect 19680 344995 19880 345000
rect 19680 344965 19685 344995
rect 19715 344965 19845 344995
rect 19875 344965 19880 344995
rect 19680 344960 19880 344965
rect 19680 344915 19880 344920
rect 19680 344885 19685 344915
rect 19715 344885 19845 344915
rect 19875 344885 19880 344915
rect 19680 344880 19880 344885
rect 19680 344835 19880 344840
rect 19680 344805 19685 344835
rect 19715 344805 19845 344835
rect 19875 344805 19880 344835
rect 19680 344800 19880 344805
rect 19680 344755 19880 344760
rect 19680 344725 19685 344755
rect 19715 344725 19845 344755
rect 19875 344725 19880 344755
rect 19680 344720 19880 344725
rect 19680 344675 19880 344680
rect 19680 344645 19685 344675
rect 19715 344645 19845 344675
rect 19875 344645 19880 344675
rect 19680 344640 19880 344645
rect 19680 344595 19880 344600
rect 19680 344565 19685 344595
rect 19715 344565 19845 344595
rect 19875 344565 19880 344595
rect 19680 344560 19880 344565
rect 19680 344515 19880 344520
rect 19680 344485 19685 344515
rect 19715 344485 19845 344515
rect 19875 344485 19880 344515
rect 19680 344480 19880 344485
rect 19680 344435 19880 344440
rect 19680 344405 19685 344435
rect 19715 344405 19845 344435
rect 19875 344405 19880 344435
rect 19680 344400 19880 344405
rect 19680 344355 19880 344360
rect 19680 344325 19685 344355
rect 19715 344325 19845 344355
rect 19875 344325 19880 344355
rect 19680 344320 19880 344325
rect 19680 344275 19880 344280
rect 19680 344245 19685 344275
rect 19715 344245 19845 344275
rect 19875 344245 19880 344275
rect 19680 344240 19880 344245
rect 19680 344195 19880 344200
rect 19680 344165 19685 344195
rect 19715 344165 19845 344195
rect 19875 344165 19880 344195
rect 19680 344160 19880 344165
rect 19680 344115 19880 344120
rect 19680 344085 19685 344115
rect 19715 344085 19845 344115
rect 19875 344085 19880 344115
rect 19680 344080 19880 344085
rect 19680 344035 19880 344040
rect 19680 344005 19685 344035
rect 19715 344005 19845 344035
rect 19875 344005 19880 344035
rect 19680 344000 19880 344005
rect 19680 343955 19880 343960
rect 19680 343925 19685 343955
rect 19715 343925 19845 343955
rect 19875 343925 19880 343955
rect 19680 343920 19880 343925
rect 19680 343875 19880 343880
rect 19680 343845 19685 343875
rect 19715 343845 19845 343875
rect 19875 343845 19880 343875
rect 19680 343840 19880 343845
rect 19680 343795 19880 343800
rect 19680 343765 19685 343795
rect 19715 343765 19845 343795
rect 19875 343765 19880 343795
rect 19680 343760 19880 343765
rect 19680 343715 19880 343720
rect 19680 343685 19685 343715
rect 19715 343685 19845 343715
rect 19875 343685 19880 343715
rect 19680 343680 19880 343685
rect 19680 343635 19880 343640
rect 19680 343605 19685 343635
rect 19715 343605 19845 343635
rect 19875 343605 19880 343635
rect 19680 343600 19880 343605
rect 19680 343555 19880 343560
rect 19680 343525 19685 343555
rect 19715 343525 19845 343555
rect 19875 343525 19880 343555
rect 19680 343520 19880 343525
rect 19680 343475 19880 343480
rect 19680 343445 19685 343475
rect 19715 343445 19845 343475
rect 19875 343445 19880 343475
rect 19680 343440 19880 343445
rect 19680 343395 19880 343400
rect 19680 343365 19685 343395
rect 19715 343365 19845 343395
rect 19875 343365 19880 343395
rect 19680 343360 19880 343365
rect 19680 343315 19880 343320
rect 19680 343285 19685 343315
rect 19715 343285 19845 343315
rect 19875 343285 19880 343315
rect 19680 343280 19880 343285
rect 19680 343235 19880 343240
rect 19680 343205 19685 343235
rect 19715 343205 19845 343235
rect 19875 343205 19880 343235
rect 19680 343200 19880 343205
rect 19680 343155 19880 343160
rect 19680 343125 19685 343155
rect 19715 343125 19845 343155
rect 19875 343125 19880 343155
rect 19680 343120 19880 343125
rect 19680 343075 19880 343080
rect 19680 343045 19685 343075
rect 19715 343045 19845 343075
rect 19875 343045 19880 343075
rect 19680 343040 19880 343045
rect 19680 342995 19880 343000
rect 19680 342965 19685 342995
rect 19715 342965 19845 342995
rect 19875 342965 19880 342995
rect 19680 342960 19880 342965
rect 19680 342915 19880 342920
rect 19680 342885 19685 342915
rect 19715 342885 19845 342915
rect 19875 342885 19880 342915
rect 19680 342880 19880 342885
rect 19680 342835 19880 342840
rect 19680 342805 19685 342835
rect 19715 342805 19845 342835
rect 19875 342805 19880 342835
rect 19680 342800 19880 342805
rect 19680 342755 19880 342760
rect 19680 342725 19685 342755
rect 19715 342725 19845 342755
rect 19875 342725 19880 342755
rect 19680 342720 19880 342725
rect 19680 342675 19880 342680
rect 19680 342645 19685 342675
rect 19715 342645 19845 342675
rect 19875 342645 19880 342675
rect 19680 342640 19880 342645
rect 19680 342595 19880 342600
rect 19680 342565 19685 342595
rect 19715 342565 19845 342595
rect 19875 342565 19880 342595
rect 19680 342560 19880 342565
rect 19680 342515 19880 342520
rect 19680 342485 19685 342515
rect 19715 342485 19845 342515
rect 19875 342485 19880 342515
rect 19680 342480 19880 342485
rect 19680 342435 19880 342440
rect 19680 342405 19685 342435
rect 19715 342405 19845 342435
rect 19875 342405 19880 342435
rect 19680 342400 19880 342405
rect 19680 342355 19880 342360
rect 19680 342325 19685 342355
rect 19715 342325 19845 342355
rect 19875 342325 19880 342355
rect 19680 342320 19880 342325
rect 19680 342275 19880 342280
rect 19680 342245 19685 342275
rect 19715 342245 19845 342275
rect 19875 342245 19880 342275
rect 19680 342240 19880 342245
rect 19680 342195 19880 342200
rect 19680 342165 19685 342195
rect 19715 342165 19845 342195
rect 19875 342165 19880 342195
rect 19680 342160 19880 342165
rect 19680 342115 19880 342120
rect 19680 342085 19685 342115
rect 19715 342085 19845 342115
rect 19875 342085 19880 342115
rect 19680 342080 19880 342085
rect 19680 342035 19880 342040
rect 19680 342005 19685 342035
rect 19715 342005 19845 342035
rect 19875 342005 19880 342035
rect 19680 342000 19880 342005
rect 19680 341955 19880 341960
rect 19680 341925 19685 341955
rect 19715 341925 19845 341955
rect 19875 341925 19880 341955
rect 19680 341920 19880 341925
rect 19680 341875 19880 341880
rect 19680 341845 19685 341875
rect 19715 341845 19845 341875
rect 19875 341845 19880 341875
rect 19680 341840 19880 341845
rect 19680 341795 19880 341800
rect 19680 341765 19685 341795
rect 19715 341765 19845 341795
rect 19875 341765 19880 341795
rect 19680 341760 19880 341765
rect 19680 341715 19880 341720
rect 19680 341685 19685 341715
rect 19715 341685 19845 341715
rect 19875 341685 19880 341715
rect 19680 341680 19880 341685
rect 19680 341635 19880 341640
rect 19680 341605 19685 341635
rect 19715 341605 19845 341635
rect 19875 341605 19880 341635
rect 19680 341600 19880 341605
rect 19680 341555 19880 341560
rect 19680 341525 19685 341555
rect 19715 341525 19845 341555
rect 19875 341525 19880 341555
rect 19680 341520 19880 341525
rect 19680 341475 19880 341480
rect 19680 341445 19685 341475
rect 19715 341445 19845 341475
rect 19875 341445 19880 341475
rect 19680 341440 19880 341445
rect 19680 341395 19880 341400
rect 19680 341365 19685 341395
rect 19715 341365 19845 341395
rect 19875 341365 19880 341395
rect 19680 341360 19880 341365
rect 19680 341315 19880 341320
rect 19680 341285 19685 341315
rect 19715 341285 19845 341315
rect 19875 341285 19880 341315
rect 19680 341280 19880 341285
rect 19680 341235 19880 341240
rect 19680 341205 19685 341235
rect 19715 341205 19845 341235
rect 19875 341205 19880 341235
rect 19680 341200 19880 341205
rect 19680 341155 19880 341160
rect 19680 341125 19685 341155
rect 19715 341125 19845 341155
rect 19875 341125 19880 341155
rect 19680 341120 19880 341125
rect 19680 341075 19880 341080
rect 19680 341045 19685 341075
rect 19715 341045 19845 341075
rect 19875 341045 19880 341075
rect 19680 341040 19880 341045
rect 19680 340995 19880 341000
rect 19680 340965 19685 340995
rect 19715 340965 19845 340995
rect 19875 340965 19880 340995
rect 19680 340960 19880 340965
rect 19680 340915 19880 340920
rect 19680 340885 19685 340915
rect 19715 340885 19845 340915
rect 19875 340885 19880 340915
rect 19680 340880 19880 340885
rect 19680 340835 19880 340840
rect 19680 340805 19685 340835
rect 19715 340805 19845 340835
rect 19875 340805 19880 340835
rect 19680 340800 19880 340805
rect 19680 340755 19880 340760
rect 19680 340725 19685 340755
rect 19715 340725 19845 340755
rect 19875 340725 19880 340755
rect 19680 340720 19880 340725
rect 19680 340675 19880 340680
rect 19680 340645 19685 340675
rect 19715 340645 19845 340675
rect 19875 340645 19880 340675
rect 19680 340640 19880 340645
rect 19680 340595 19880 340600
rect 19680 340565 19685 340595
rect 19715 340565 19845 340595
rect 19875 340565 19880 340595
rect 19680 340560 19880 340565
rect 19680 340515 19880 340520
rect 19680 340485 19685 340515
rect 19715 340485 19845 340515
rect 19875 340485 19880 340515
rect 19680 340480 19880 340485
rect 19680 340435 19880 340440
rect 19680 340405 19685 340435
rect 19715 340405 19845 340435
rect 19875 340405 19880 340435
rect 19680 340400 19880 340405
rect 19680 340355 19880 340360
rect 19680 340325 19685 340355
rect 19715 340325 19845 340355
rect 19875 340325 19880 340355
rect 19680 340320 19880 340325
rect 19680 340275 19880 340280
rect 19680 340245 19685 340275
rect 19715 340245 19845 340275
rect 19875 340245 19880 340275
rect 19680 340240 19880 340245
rect 19680 340195 19880 340200
rect 19680 340165 19685 340195
rect 19715 340165 19845 340195
rect 19875 340165 19880 340195
rect 19680 340160 19880 340165
rect 19680 340115 19880 340120
rect 19680 340085 19685 340115
rect 19715 340085 19845 340115
rect 19875 340085 19880 340115
rect 19680 340080 19880 340085
rect 19680 340035 19880 340040
rect 19680 340005 19685 340035
rect 19715 340005 19845 340035
rect 19875 340005 19880 340035
rect 19680 340000 19880 340005
rect 19680 339955 19880 339960
rect 19680 339925 19685 339955
rect 19715 339925 19845 339955
rect 19875 339925 19880 339955
rect 19680 339920 19880 339925
rect 19680 339875 19880 339880
rect 19680 339845 19685 339875
rect 19715 339845 19845 339875
rect 19875 339845 19880 339875
rect 19680 339840 19880 339845
rect 19680 339795 19880 339800
rect 19680 339765 19685 339795
rect 19715 339765 19845 339795
rect 19875 339765 19880 339795
rect 19680 339760 19880 339765
rect 19680 339715 19880 339720
rect 19680 339685 19685 339715
rect 19715 339685 19845 339715
rect 19875 339685 19880 339715
rect 19680 339680 19880 339685
rect 19680 339635 19880 339640
rect 19680 339605 19685 339635
rect 19715 339605 19845 339635
rect 19875 339605 19880 339635
rect 19680 339600 19880 339605
rect 19680 339555 19880 339560
rect 19680 339525 19685 339555
rect 19715 339525 19845 339555
rect 19875 339525 19880 339555
rect 19680 339520 19880 339525
rect 19680 339475 19880 339480
rect 19680 339445 19685 339475
rect 19715 339445 19845 339475
rect 19875 339445 19880 339475
rect 19680 339440 19880 339445
rect 19680 339395 19880 339400
rect 19680 339365 19685 339395
rect 19715 339365 19845 339395
rect 19875 339365 19880 339395
rect 19680 339360 19880 339365
rect 19680 339315 19880 339320
rect 19680 339285 19685 339315
rect 19715 339285 19845 339315
rect 19875 339285 19880 339315
rect 19680 339280 19880 339285
rect 19680 339235 19880 339240
rect 19680 339205 19685 339235
rect 19715 339205 19845 339235
rect 19875 339205 19880 339235
rect 19680 339200 19880 339205
rect 19680 339155 19880 339160
rect 19680 339125 19685 339155
rect 19715 339125 19845 339155
rect 19875 339125 19880 339155
rect 19680 339120 19880 339125
rect 19680 339075 19880 339080
rect 19680 339045 19685 339075
rect 19715 339045 19845 339075
rect 19875 339045 19880 339075
rect 19680 339040 19880 339045
rect 19680 338995 19880 339000
rect 19680 338965 19685 338995
rect 19715 338965 19845 338995
rect 19875 338965 19880 338995
rect 19680 338960 19880 338965
rect 19680 338915 19880 338920
rect 19680 338885 19685 338915
rect 19715 338885 19845 338915
rect 19875 338885 19880 338915
rect 19680 338880 19880 338885
rect 19680 338835 19880 338840
rect 19680 338805 19685 338835
rect 19715 338805 19845 338835
rect 19875 338805 19880 338835
rect 19680 338800 19880 338805
rect 19680 338755 19880 338760
rect 19680 338725 19685 338755
rect 19715 338725 19845 338755
rect 19875 338725 19880 338755
rect 19680 338720 19880 338725
rect 19680 338675 19880 338680
rect 19680 338645 19685 338675
rect 19715 338645 19845 338675
rect 19875 338645 19880 338675
rect 19680 338640 19880 338645
rect 19680 338595 19880 338600
rect 19680 338565 19685 338595
rect 19715 338565 19845 338595
rect 19875 338565 19880 338595
rect 19680 338560 19880 338565
rect 19680 338515 19880 338520
rect 19680 338485 19685 338515
rect 19715 338485 19845 338515
rect 19875 338485 19880 338515
rect 19680 338480 19880 338485
rect 19680 338435 19880 338440
rect 19680 338405 19685 338435
rect 19715 338405 19845 338435
rect 19875 338405 19880 338435
rect 19680 338400 19880 338405
rect 19680 338355 19880 338360
rect 19680 338325 19685 338355
rect 19715 338325 19845 338355
rect 19875 338325 19880 338355
rect 19680 338320 19880 338325
rect 19680 338275 19880 338280
rect 19680 338245 19685 338275
rect 19715 338245 19845 338275
rect 19875 338245 19880 338275
rect 19680 338240 19880 338245
rect 19680 338195 19880 338200
rect 19680 338165 19685 338195
rect 19715 338165 19845 338195
rect 19875 338165 19880 338195
rect 19680 338160 19880 338165
rect 19680 338115 19880 338120
rect 19680 338085 19685 338115
rect 19715 338085 19845 338115
rect 19875 338085 19880 338115
rect 19680 338080 19880 338085
rect 19680 338035 19880 338040
rect 19680 338005 19685 338035
rect 19715 338005 19845 338035
rect 19875 338005 19880 338035
rect 19680 338000 19880 338005
rect 19680 337955 19880 337960
rect 19680 337925 19685 337955
rect 19715 337925 19845 337955
rect 19875 337925 19880 337955
rect 19680 337920 19880 337925
rect 19680 337875 19880 337880
rect 19680 337845 19685 337875
rect 19715 337845 19845 337875
rect 19875 337845 19880 337875
rect 19680 337840 19880 337845
rect 19680 337795 19880 337800
rect 19680 337765 19685 337795
rect 19715 337765 19845 337795
rect 19875 337765 19880 337795
rect 19680 337760 19880 337765
rect 19680 337715 19880 337720
rect 19680 337685 19685 337715
rect 19715 337685 19845 337715
rect 19875 337685 19880 337715
rect 19680 337680 19880 337685
rect 19680 337635 19880 337640
rect 19680 337605 19685 337635
rect 19715 337605 19845 337635
rect 19875 337605 19880 337635
rect 19680 337600 19880 337605
rect 19680 337555 19880 337560
rect 19680 337525 19685 337555
rect 19715 337525 19845 337555
rect 19875 337525 19880 337555
rect 19680 337520 19880 337525
rect 19680 337475 19880 337480
rect 19680 337445 19685 337475
rect 19715 337445 19845 337475
rect 19875 337445 19880 337475
rect 19680 337440 19880 337445
rect 19680 337395 19880 337400
rect 19680 337365 19685 337395
rect 19715 337365 19845 337395
rect 19875 337365 19880 337395
rect 19680 337360 19880 337365
rect 19680 337315 19880 337320
rect 19680 337285 19685 337315
rect 19715 337285 19845 337315
rect 19875 337285 19880 337315
rect 19680 337280 19880 337285
rect 19680 337235 19880 337240
rect 19680 337205 19685 337235
rect 19715 337205 19845 337235
rect 19875 337205 19880 337235
rect 19680 337200 19880 337205
rect 19680 337155 19880 337160
rect 19680 337125 19685 337155
rect 19715 337125 19845 337155
rect 19875 337125 19880 337155
rect 19680 337120 19880 337125
rect 19680 337075 19880 337080
rect 19680 337045 19685 337075
rect 19715 337045 19845 337075
rect 19875 337045 19880 337075
rect 19680 337040 19880 337045
rect 19680 336995 19880 337000
rect 19680 336965 19685 336995
rect 19715 336965 19845 336995
rect 19875 336965 19880 336995
rect 19680 336960 19880 336965
rect 19680 336915 19880 336920
rect 19680 336885 19685 336915
rect 19715 336885 19845 336915
rect 19875 336885 19880 336915
rect 19680 336880 19880 336885
rect 19680 336835 19880 336840
rect 19680 336805 19685 336835
rect 19715 336805 19845 336835
rect 19875 336805 19880 336835
rect 19680 336800 19880 336805
rect 19680 336755 19880 336760
rect 19680 336725 19685 336755
rect 19715 336725 19845 336755
rect 19875 336725 19880 336755
rect 19680 336720 19880 336725
rect 19680 336675 19880 336680
rect 19680 336645 19685 336675
rect 19715 336645 19845 336675
rect 19875 336645 19880 336675
rect 19680 336640 19880 336645
rect 19680 336595 19880 336600
rect 19680 336565 19685 336595
rect 19715 336565 19845 336595
rect 19875 336565 19880 336595
rect 19680 336560 19880 336565
rect 19680 336515 19880 336520
rect 19680 336485 19685 336515
rect 19715 336485 19845 336515
rect 19875 336485 19880 336515
rect 19680 336480 19880 336485
rect 19680 336435 19880 336440
rect 19680 336405 19685 336435
rect 19715 336405 19845 336435
rect 19875 336405 19880 336435
rect 19680 336400 19880 336405
rect 19680 336355 19880 336360
rect 19680 336325 19685 336355
rect 19715 336325 19845 336355
rect 19875 336325 19880 336355
rect 19680 336320 19880 336325
rect 19680 336275 19880 336280
rect 19680 336245 19685 336275
rect 19715 336245 19845 336275
rect 19875 336245 19880 336275
rect 19680 336240 19880 336245
rect 19680 336195 19880 336200
rect 19680 336165 19685 336195
rect 19715 336165 19845 336195
rect 19875 336165 19880 336195
rect 19680 336160 19880 336165
rect 19680 336115 19880 336120
rect 19680 336085 19685 336115
rect 19715 336085 19845 336115
rect 19875 336085 19880 336115
rect 19680 336080 19880 336085
rect 19680 336035 19880 336040
rect 19680 336005 19685 336035
rect 19715 336005 19845 336035
rect 19875 336005 19880 336035
rect 19680 336000 19880 336005
rect 19680 335955 19880 335960
rect 19680 335925 19685 335955
rect 19715 335925 19845 335955
rect 19875 335925 19880 335955
rect 19680 335920 19880 335925
rect 19680 335875 19880 335880
rect 19680 335845 19685 335875
rect 19715 335845 19845 335875
rect 19875 335845 19880 335875
rect 19680 335840 19880 335845
rect 19680 335795 19880 335800
rect 19680 335765 19685 335795
rect 19715 335765 19845 335795
rect 19875 335765 19880 335795
rect 19680 335760 19880 335765
rect 19680 335715 19880 335720
rect 19680 335685 19685 335715
rect 19715 335685 19845 335715
rect 19875 335685 19880 335715
rect 19680 335680 19880 335685
rect 19680 335635 19880 335640
rect 19680 335605 19685 335635
rect 19715 335605 19845 335635
rect 19875 335605 19880 335635
rect 19680 335600 19880 335605
rect 19680 335555 19880 335560
rect 19680 335525 19685 335555
rect 19715 335525 19845 335555
rect 19875 335525 19880 335555
rect 19680 335520 19880 335525
rect 19680 335475 19880 335480
rect 19680 335445 19685 335475
rect 19715 335445 19845 335475
rect 19875 335445 19880 335475
rect 19680 335440 19880 335445
rect 19680 335395 19880 335400
rect 19680 335365 19685 335395
rect 19715 335365 19845 335395
rect 19875 335365 19880 335395
rect 19680 335360 19880 335365
rect 19680 335315 19880 335320
rect 19680 335285 19685 335315
rect 19715 335285 19845 335315
rect 19875 335285 19880 335315
rect 19680 335280 19880 335285
rect 19680 335235 19880 335240
rect 19680 335205 19685 335235
rect 19715 335205 19845 335235
rect 19875 335205 19880 335235
rect 19680 335200 19880 335205
rect 19680 335155 19880 335160
rect 19680 335125 19685 335155
rect 19715 335125 19845 335155
rect 19875 335125 19880 335155
rect 19680 335120 19880 335125
rect 19680 335075 19880 335080
rect 19680 335045 19685 335075
rect 19715 335045 19845 335075
rect 19875 335045 19880 335075
rect 19680 335040 19880 335045
rect 19680 334995 19880 335000
rect 19680 334965 19685 334995
rect 19715 334965 19845 334995
rect 19875 334965 19880 334995
rect 19680 334960 19880 334965
rect 19680 334915 19880 334920
rect 19680 334885 19685 334915
rect 19715 334885 19845 334915
rect 19875 334885 19880 334915
rect 19680 334880 19880 334885
rect 19680 334835 19880 334840
rect 19680 334805 19685 334835
rect 19715 334805 19845 334835
rect 19875 334805 19880 334835
rect 19680 334800 19880 334805
rect 19680 334755 19880 334760
rect 19680 334725 19685 334755
rect 19715 334725 19845 334755
rect 19875 334725 19880 334755
rect 19680 334720 19880 334725
rect 19680 334675 19880 334680
rect 19680 334645 19685 334675
rect 19715 334645 19845 334675
rect 19875 334645 19880 334675
rect 19680 334640 19880 334645
rect 19680 334595 19880 334600
rect 19680 334565 19685 334595
rect 19715 334565 19845 334595
rect 19875 334565 19880 334595
rect 19680 334560 19880 334565
rect 19680 334515 19880 334520
rect 19680 334485 19685 334515
rect 19715 334485 19845 334515
rect 19875 334485 19880 334515
rect 19680 334480 19880 334485
rect 19680 334435 19880 334440
rect 19680 334405 19685 334435
rect 19715 334405 19845 334435
rect 19875 334405 19880 334435
rect 19680 334400 19880 334405
rect 19680 334355 19880 334360
rect 19680 334325 19685 334355
rect 19715 334325 19845 334355
rect 19875 334325 19880 334355
rect 19680 334320 19880 334325
rect 19680 334275 19880 334280
rect 19680 334245 19685 334275
rect 19715 334245 19845 334275
rect 19875 334245 19880 334275
rect 19680 334240 19880 334245
rect 19680 334195 19880 334200
rect 19680 334165 19685 334195
rect 19715 334165 19845 334195
rect 19875 334165 19880 334195
rect 19680 334160 19880 334165
rect 19680 334115 19880 334120
rect 19680 334085 19685 334115
rect 19715 334085 19845 334115
rect 19875 334085 19880 334115
rect 19680 334080 19880 334085
rect 19680 334035 19880 334040
rect 19680 334005 19685 334035
rect 19715 334005 19845 334035
rect 19875 334005 19880 334035
rect 19680 334000 19880 334005
rect 19680 333955 19880 333960
rect 19680 333925 19685 333955
rect 19715 333925 19845 333955
rect 19875 333925 19880 333955
rect 19680 333920 19880 333925
rect 19680 333875 19880 333880
rect 19680 333845 19685 333875
rect 19715 333845 19845 333875
rect 19875 333845 19880 333875
rect 19680 333840 19880 333845
rect 19680 333795 19880 333800
rect 19680 333765 19685 333795
rect 19715 333765 19845 333795
rect 19875 333765 19880 333795
rect 19680 333760 19880 333765
rect 19680 333715 19880 333720
rect 19680 333685 19685 333715
rect 19715 333685 19845 333715
rect 19875 333685 19880 333715
rect 19680 333680 19880 333685
rect 19680 333635 19880 333640
rect 19680 333605 19685 333635
rect 19715 333605 19845 333635
rect 19875 333605 19880 333635
rect 19680 333600 19880 333605
rect 19680 333555 19880 333560
rect 19680 333525 19685 333555
rect 19715 333525 19845 333555
rect 19875 333525 19880 333555
rect 19680 333520 19880 333525
rect 19680 333475 19880 333480
rect 19680 333445 19685 333475
rect 19715 333445 19845 333475
rect 19875 333445 19880 333475
rect 19680 333440 19880 333445
rect 19680 333395 19880 333400
rect 19680 333365 19685 333395
rect 19715 333365 19845 333395
rect 19875 333365 19880 333395
rect 19680 333360 19880 333365
rect 19680 333315 19880 333320
rect 19680 333285 19685 333315
rect 19715 333285 19845 333315
rect 19875 333285 19880 333315
rect 19680 333280 19880 333285
rect 19680 333235 19880 333240
rect 19680 333205 19685 333235
rect 19715 333205 19845 333235
rect 19875 333205 19880 333235
rect 19680 333200 19880 333205
rect 19680 333155 19880 333160
rect 19680 333125 19685 333155
rect 19715 333125 19845 333155
rect 19875 333125 19880 333155
rect 19680 333120 19880 333125
rect 19680 333075 19880 333080
rect 19680 333045 19685 333075
rect 19715 333045 19845 333075
rect 19875 333045 19880 333075
rect 19680 333040 19880 333045
rect 19680 332995 19880 333000
rect 19680 332965 19685 332995
rect 19715 332965 19845 332995
rect 19875 332965 19880 332995
rect 19680 332960 19880 332965
rect 19680 332915 19880 332920
rect 19680 332885 19685 332915
rect 19715 332885 19845 332915
rect 19875 332885 19880 332915
rect 19680 332880 19880 332885
rect 19680 332835 19880 332840
rect 19680 332805 19685 332835
rect 19715 332805 19845 332835
rect 19875 332805 19880 332835
rect 19680 332800 19880 332805
rect 19680 332755 19880 332760
rect 19680 332725 19685 332755
rect 19715 332725 19845 332755
rect 19875 332725 19880 332755
rect 19680 332720 19880 332725
rect 19680 332675 19880 332680
rect 19680 332645 19685 332675
rect 19715 332645 19845 332675
rect 19875 332645 19880 332675
rect 19680 332640 19880 332645
rect 19680 332595 19880 332600
rect 19680 332565 19685 332595
rect 19715 332565 19845 332595
rect 19875 332565 19880 332595
rect 19680 332560 19880 332565
rect 19680 332515 19880 332520
rect 19680 332485 19685 332515
rect 19715 332485 19845 332515
rect 19875 332485 19880 332515
rect 19680 332480 19880 332485
rect 19680 332435 19880 332440
rect 19680 332405 19685 332435
rect 19715 332405 19845 332435
rect 19875 332405 19880 332435
rect 19680 332400 19880 332405
rect 19680 332355 19880 332360
rect 19680 332325 19685 332355
rect 19715 332325 19845 332355
rect 19875 332325 19880 332355
rect 19680 332320 19880 332325
rect 19680 332275 19880 332280
rect 19680 332245 19685 332275
rect 19715 332245 19845 332275
rect 19875 332245 19880 332275
rect 19680 332240 19880 332245
rect 19680 332195 19880 332200
rect 19680 332165 19685 332195
rect 19715 332165 19845 332195
rect 19875 332165 19880 332195
rect 19680 332160 19880 332165
rect 19680 332115 19880 332120
rect 19680 332085 19685 332115
rect 19715 332085 19845 332115
rect 19875 332085 19880 332115
rect 19680 332080 19880 332085
rect 19680 332035 19880 332040
rect 19680 332005 19685 332035
rect 19715 332005 19845 332035
rect 19875 332005 19880 332035
rect 19680 332000 19880 332005
rect 19680 331955 19880 331960
rect 19680 331925 19685 331955
rect 19715 331925 19845 331955
rect 19875 331925 19880 331955
rect 19680 331920 19880 331925
rect 19680 331875 19880 331880
rect 19680 331845 19685 331875
rect 19715 331845 19845 331875
rect 19875 331845 19880 331875
rect 19680 331840 19880 331845
rect 19680 331795 19880 331800
rect 19680 331765 19685 331795
rect 19715 331765 19845 331795
rect 19875 331765 19880 331795
rect 19680 331760 19880 331765
rect 19680 331715 19880 331720
rect 19680 331685 19685 331715
rect 19715 331685 19845 331715
rect 19875 331685 19880 331715
rect 19680 331680 19880 331685
rect 19680 331635 19880 331640
rect 19680 331605 19685 331635
rect 19715 331605 19845 331635
rect 19875 331605 19880 331635
rect 19680 331600 19880 331605
rect 19680 331555 19880 331560
rect 19680 331525 19685 331555
rect 19715 331525 19845 331555
rect 19875 331525 19880 331555
rect 19680 331520 19880 331525
rect 19680 331475 19880 331480
rect 19680 331445 19685 331475
rect 19715 331445 19845 331475
rect 19875 331445 19880 331475
rect 19680 331440 19880 331445
rect 19680 331395 19880 331400
rect 19680 331365 19685 331395
rect 19715 331365 19845 331395
rect 19875 331365 19880 331395
rect 19680 331360 19880 331365
rect 19680 331315 19880 331320
rect 19680 331285 19685 331315
rect 19715 331285 19845 331315
rect 19875 331285 19880 331315
rect 19680 331280 19880 331285
rect 19680 331235 19880 331240
rect 19680 331205 19685 331235
rect 19715 331205 19845 331235
rect 19875 331205 19880 331235
rect 19680 331200 19880 331205
rect 19680 331155 19880 331160
rect 19680 331125 19685 331155
rect 19715 331125 19845 331155
rect 19875 331125 19880 331155
rect 19680 331120 19880 331125
rect 19680 331075 19880 331080
rect 19680 331045 19685 331075
rect 19715 331045 19845 331075
rect 19875 331045 19880 331075
rect 19680 331040 19880 331045
rect 19680 330995 19880 331000
rect 19680 330965 19685 330995
rect 19715 330965 19845 330995
rect 19875 330965 19880 330995
rect 19680 330960 19880 330965
rect 19680 330915 19880 330920
rect 19680 330885 19685 330915
rect 19715 330885 19845 330915
rect 19875 330885 19880 330915
rect 19680 330880 19880 330885
rect 19680 330835 19880 330840
rect 19680 330805 19685 330835
rect 19715 330805 19845 330835
rect 19875 330805 19880 330835
rect 19680 330800 19880 330805
rect 19680 330755 19880 330760
rect 19680 330725 19685 330755
rect 19715 330725 19845 330755
rect 19875 330725 19880 330755
rect 19680 330720 19880 330725
rect 19680 330675 19880 330680
rect 19680 330645 19685 330675
rect 19715 330645 19845 330675
rect 19875 330645 19880 330675
rect 19680 330640 19880 330645
rect 19680 330595 19880 330600
rect 19680 330565 19685 330595
rect 19715 330565 19845 330595
rect 19875 330565 19880 330595
rect 19680 330560 19880 330565
rect 19680 330515 19880 330520
rect 19680 330485 19685 330515
rect 19715 330485 19845 330515
rect 19875 330485 19880 330515
rect 19680 330480 19880 330485
rect 19680 330435 19880 330440
rect 19680 330405 19685 330435
rect 19715 330405 19845 330435
rect 19875 330405 19880 330435
rect 19680 330400 19880 330405
rect 19680 330355 19880 330360
rect 19680 330325 19685 330355
rect 19715 330325 19845 330355
rect 19875 330325 19880 330355
rect 19680 330320 19880 330325
rect 19680 330275 19880 330280
rect 19680 330245 19685 330275
rect 19715 330245 19845 330275
rect 19875 330245 19880 330275
rect 19680 330240 19880 330245
rect 19680 330195 19880 330200
rect 19680 330165 19685 330195
rect 19715 330165 19845 330195
rect 19875 330165 19880 330195
rect 19680 330160 19880 330165
rect 19680 330115 19880 330120
rect 19680 330085 19685 330115
rect 19715 330085 19845 330115
rect 19875 330085 19880 330115
rect 19680 330080 19880 330085
rect 19680 330035 19880 330040
rect 19680 330005 19685 330035
rect 19715 330005 19845 330035
rect 19875 330005 19880 330035
rect 19680 330000 19880 330005
rect 19680 329955 19880 329960
rect 19680 329925 19685 329955
rect 19715 329925 19845 329955
rect 19875 329925 19880 329955
rect 19680 329920 19880 329925
rect 19680 329875 19880 329880
rect 19680 329845 19685 329875
rect 19715 329845 19845 329875
rect 19875 329845 19880 329875
rect 19680 329840 19880 329845
rect 19680 329795 19880 329800
rect 19680 329765 19685 329795
rect 19715 329765 19845 329795
rect 19875 329765 19880 329795
rect 19680 329760 19880 329765
rect 19680 329715 19880 329720
rect 19680 329685 19685 329715
rect 19715 329685 19845 329715
rect 19875 329685 19880 329715
rect 19680 329680 19880 329685
rect 19680 329635 19880 329640
rect 19680 329605 19685 329635
rect 19715 329605 19845 329635
rect 19875 329605 19880 329635
rect 19680 329600 19880 329605
rect 19680 329555 19880 329560
rect 19680 329525 19685 329555
rect 19715 329525 19845 329555
rect 19875 329525 19880 329555
rect 19680 329520 19880 329525
rect 19680 329475 19880 329480
rect 19680 329445 19685 329475
rect 19715 329445 19845 329475
rect 19875 329445 19880 329475
rect 19680 329440 19880 329445
rect 19680 329395 19880 329400
rect 19680 329365 19685 329395
rect 19715 329365 19845 329395
rect 19875 329365 19880 329395
rect 19680 329360 19880 329365
rect 19680 329315 19880 329320
rect 19680 329285 19685 329315
rect 19715 329285 19845 329315
rect 19875 329285 19880 329315
rect 19680 329280 19880 329285
rect 19680 329235 19880 329240
rect 19680 329205 19685 329235
rect 19715 329205 19845 329235
rect 19875 329205 19880 329235
rect 19680 329200 19880 329205
rect 19680 329155 19880 329160
rect 19680 329125 19685 329155
rect 19715 329125 19845 329155
rect 19875 329125 19880 329155
rect 19680 329120 19880 329125
rect 19680 329075 19880 329080
rect 19680 329045 19685 329075
rect 19715 329045 19845 329075
rect 19875 329045 19880 329075
rect 19680 329040 19880 329045
rect 19680 328995 19880 329000
rect 19680 328965 19685 328995
rect 19715 328965 19845 328995
rect 19875 328965 19880 328995
rect 19680 328960 19880 328965
rect 19680 328915 19880 328920
rect 19680 328885 19685 328915
rect 19715 328885 19845 328915
rect 19875 328885 19880 328915
rect 19680 328880 19880 328885
rect 19680 328835 19880 328840
rect 19680 328805 19685 328835
rect 19715 328805 19845 328835
rect 19875 328805 19880 328835
rect 19680 328800 19880 328805
rect 19680 328755 19880 328760
rect 19680 328725 19685 328755
rect 19715 328725 19845 328755
rect 19875 328725 19880 328755
rect 19680 328720 19880 328725
rect 19680 328675 19880 328680
rect 19680 328645 19685 328675
rect 19715 328645 19845 328675
rect 19875 328645 19880 328675
rect 19680 328640 19880 328645
rect 19680 328595 19880 328600
rect 19680 328565 19685 328595
rect 19715 328565 19845 328595
rect 19875 328565 19880 328595
rect 19680 328560 19880 328565
rect 19680 328515 19880 328520
rect 19680 328485 19685 328515
rect 19715 328485 19845 328515
rect 19875 328485 19880 328515
rect 19680 328480 19880 328485
rect 19680 328435 19880 328440
rect 19680 328405 19685 328435
rect 19715 328405 19845 328435
rect 19875 328405 19880 328435
rect 19680 328400 19880 328405
rect 19680 328355 19880 328360
rect 19680 328325 19685 328355
rect 19715 328325 19845 328355
rect 19875 328325 19880 328355
rect 19680 328320 19880 328325
rect 19680 328275 19880 328280
rect 19680 328245 19685 328275
rect 19715 328245 19845 328275
rect 19875 328245 19880 328275
rect 19680 328240 19880 328245
rect 19680 328195 19880 328200
rect 19680 328165 19685 328195
rect 19715 328165 19845 328195
rect 19875 328165 19880 328195
rect 19680 328160 19880 328165
rect 19680 328115 19880 328120
rect 19680 328085 19685 328115
rect 19715 328085 19845 328115
rect 19875 328085 19880 328115
rect 19680 328080 19880 328085
rect 19680 328035 19880 328040
rect 19680 328005 19685 328035
rect 19715 328005 19845 328035
rect 19875 328005 19880 328035
rect 19680 328000 19880 328005
rect 19680 327955 19880 327960
rect 19680 327925 19685 327955
rect 19715 327925 19845 327955
rect 19875 327925 19880 327955
rect 19680 327920 19880 327925
rect 19680 327875 19880 327880
rect 19680 327845 19685 327875
rect 19715 327845 19845 327875
rect 19875 327845 19880 327875
rect 19680 327840 19880 327845
rect 19680 327795 19880 327800
rect 19680 327765 19685 327795
rect 19715 327765 19845 327795
rect 19875 327765 19880 327795
rect 19680 327760 19880 327765
rect 19680 327715 19880 327720
rect 19680 327685 19685 327715
rect 19715 327685 19845 327715
rect 19875 327685 19880 327715
rect 19680 327680 19880 327685
rect 19680 327635 19880 327640
rect 19680 327605 19685 327635
rect 19715 327605 19845 327635
rect 19875 327605 19880 327635
rect 19680 327600 19880 327605
rect 19680 327555 19880 327560
rect 19680 327525 19685 327555
rect 19715 327525 19845 327555
rect 19875 327525 19880 327555
rect 19680 327520 19880 327525
rect 19680 327475 19880 327480
rect 19680 327445 19685 327475
rect 19715 327445 19845 327475
rect 19875 327445 19880 327475
rect 19680 327440 19880 327445
rect 19680 327395 19880 327400
rect 19680 327365 19685 327395
rect 19715 327365 19845 327395
rect 19875 327365 19880 327395
rect 19680 327360 19880 327365
rect 19680 327315 19880 327320
rect 19680 327285 19685 327315
rect 19715 327285 19845 327315
rect 19875 327285 19880 327315
rect 19680 327280 19880 327285
rect 19680 327235 19880 327240
rect 19680 327205 19685 327235
rect 19715 327205 19845 327235
rect 19875 327205 19880 327235
rect 19680 327200 19880 327205
rect 19680 327155 19880 327160
rect 19680 327125 19685 327155
rect 19715 327125 19845 327155
rect 19875 327125 19880 327155
rect 19680 327120 19880 327125
rect 19680 327075 19880 327080
rect 19680 327045 19685 327075
rect 19715 327045 19845 327075
rect 19875 327045 19880 327075
rect 19680 327040 19880 327045
rect 19680 326995 19880 327000
rect 19680 326965 19685 326995
rect 19715 326965 19845 326995
rect 19875 326965 19880 326995
rect 19680 326960 19880 326965
rect 19680 326915 19880 326920
rect 19680 326885 19685 326915
rect 19715 326885 19845 326915
rect 19875 326885 19880 326915
rect 19680 326880 19880 326885
rect 19680 326835 19880 326840
rect 19680 326805 19685 326835
rect 19715 326805 19845 326835
rect 19875 326805 19880 326835
rect 19680 326800 19880 326805
rect 19680 326755 19880 326760
rect 19680 326725 19685 326755
rect 19715 326725 19845 326755
rect 19875 326725 19880 326755
rect 19680 326720 19880 326725
rect 19680 326675 19880 326680
rect 19680 326645 19685 326675
rect 19715 326645 19845 326675
rect 19875 326645 19880 326675
rect 19680 326640 19880 326645
rect 19680 326595 19880 326600
rect 19680 326565 19685 326595
rect 19715 326565 19845 326595
rect 19875 326565 19880 326595
rect 19680 326560 19880 326565
rect 19680 326515 19880 326520
rect 19680 326485 19685 326515
rect 19715 326485 19845 326515
rect 19875 326485 19880 326515
rect 19680 326480 19880 326485
rect 19680 326435 19880 326440
rect 19680 326405 19685 326435
rect 19715 326405 19845 326435
rect 19875 326405 19880 326435
rect 19680 326400 19880 326405
rect 19680 326355 19880 326360
rect 19680 326325 19685 326355
rect 19715 326325 19845 326355
rect 19875 326325 19880 326355
rect 19680 326320 19880 326325
rect 19680 326275 19880 326280
rect 19680 326245 19685 326275
rect 19715 326245 19845 326275
rect 19875 326245 19880 326275
rect 19680 326240 19880 326245
rect 19680 326195 19880 326200
rect 19680 326165 19685 326195
rect 19715 326165 19845 326195
rect 19875 326165 19880 326195
rect 19680 326160 19880 326165
rect 19680 326115 19880 326120
rect 19680 326085 19685 326115
rect 19715 326085 19845 326115
rect 19875 326085 19880 326115
rect 19680 326080 19880 326085
rect 19680 326035 19880 326040
rect 19680 326005 19685 326035
rect 19715 326005 19845 326035
rect 19875 326005 19880 326035
rect 19680 326000 19880 326005
rect 19680 325955 19880 325960
rect 19680 325925 19685 325955
rect 19715 325925 19845 325955
rect 19875 325925 19880 325955
rect 19680 325920 19880 325925
rect 19680 325875 19880 325880
rect 19680 325845 19685 325875
rect 19715 325845 19845 325875
rect 19875 325845 19880 325875
rect 19680 325840 19880 325845
rect 19680 325795 19880 325800
rect 19680 325765 19685 325795
rect 19715 325765 19845 325795
rect 19875 325765 19880 325795
rect 19680 325760 19880 325765
rect 19680 325715 19880 325720
rect 19680 325685 19685 325715
rect 19715 325685 19845 325715
rect 19875 325685 19880 325715
rect 19680 325680 19880 325685
rect 19680 325635 19880 325640
rect 19680 325605 19685 325635
rect 19715 325605 19845 325635
rect 19875 325605 19880 325635
rect 19680 325600 19880 325605
rect 19680 325555 19880 325560
rect 19680 325525 19685 325555
rect 19715 325525 19845 325555
rect 19875 325525 19880 325555
rect 19680 325520 19880 325525
rect 19680 325475 19880 325480
rect 19680 325445 19685 325475
rect 19715 325445 19845 325475
rect 19875 325445 19880 325475
rect 19680 325440 19880 325445
rect 19680 325395 19880 325400
rect 19680 325365 19685 325395
rect 19715 325365 19845 325395
rect 19875 325365 19880 325395
rect 19680 325360 19880 325365
rect 19680 325315 19880 325320
rect 19680 325285 19685 325315
rect 19715 325285 19845 325315
rect 19875 325285 19880 325315
rect 19680 325280 19880 325285
rect 19680 325235 19880 325240
rect 19680 325205 19685 325235
rect 19715 325205 19845 325235
rect 19875 325205 19880 325235
rect 19680 325200 19880 325205
rect 19680 325155 19880 325160
rect 19680 325125 19685 325155
rect 19715 325125 19845 325155
rect 19875 325125 19880 325155
rect 19680 325120 19880 325125
rect 19680 325075 19880 325080
rect 19680 325045 19685 325075
rect 19715 325045 19845 325075
rect 19875 325045 19880 325075
rect 19680 325040 19880 325045
rect 19680 324995 19880 325000
rect 19680 324965 19685 324995
rect 19715 324965 19845 324995
rect 19875 324965 19880 324995
rect 19680 324960 19880 324965
rect 19680 324915 19880 324920
rect 19680 324885 19685 324915
rect 19715 324885 19845 324915
rect 19875 324885 19880 324915
rect 19680 324880 19880 324885
rect 19680 324835 19880 324840
rect 19680 324805 19685 324835
rect 19715 324805 19845 324835
rect 19875 324805 19880 324835
rect 19680 324800 19880 324805
rect 19680 324755 19880 324760
rect 19680 324725 19685 324755
rect 19715 324725 19845 324755
rect 19875 324725 19880 324755
rect 19680 324720 19880 324725
rect 19680 324675 19880 324680
rect 19680 324645 19685 324675
rect 19715 324645 19845 324675
rect 19875 324645 19880 324675
rect 19680 324640 19880 324645
rect 19680 324595 19880 324600
rect 19680 324565 19685 324595
rect 19715 324565 19845 324595
rect 19875 324565 19880 324595
rect 19680 324560 19880 324565
rect 19680 324515 19880 324520
rect 19680 324485 19685 324515
rect 19715 324485 19845 324515
rect 19875 324485 19880 324515
rect 19680 324480 19880 324485
rect 19680 324435 19880 324440
rect 19680 324405 19685 324435
rect 19715 324405 19845 324435
rect 19875 324405 19880 324435
rect 19680 324400 19880 324405
rect 19680 324355 19880 324360
rect 19680 324325 19685 324355
rect 19715 324325 19845 324355
rect 19875 324325 19880 324355
rect 19680 324320 19880 324325
rect 19680 324275 19880 324280
rect 19680 324245 19685 324275
rect 19715 324245 19845 324275
rect 19875 324245 19880 324275
rect 19680 324240 19880 324245
rect 19680 324195 19880 324200
rect 19680 324165 19685 324195
rect 19715 324165 19845 324195
rect 19875 324165 19880 324195
rect 19680 324160 19880 324165
rect 19680 324115 19880 324120
rect 19680 324085 19685 324115
rect 19715 324085 19845 324115
rect 19875 324085 19880 324115
rect 19680 324080 19880 324085
rect 19680 324035 19880 324040
rect 19680 324005 19685 324035
rect 19715 324005 19845 324035
rect 19875 324005 19880 324035
rect 19680 324000 19880 324005
rect 19680 323955 19880 323960
rect 19680 323925 19685 323955
rect 19715 323925 19845 323955
rect 19875 323925 19880 323955
rect 19680 323920 19880 323925
rect 19680 323875 19880 323880
rect 19680 323845 19685 323875
rect 19715 323845 19845 323875
rect 19875 323845 19880 323875
rect 19680 323840 19880 323845
rect 19680 323795 19880 323800
rect 19680 323765 19685 323795
rect 19715 323765 19845 323795
rect 19875 323765 19880 323795
rect 19680 323760 19880 323765
rect 19680 323715 19880 323720
rect 19680 323685 19685 323715
rect 19715 323685 19845 323715
rect 19875 323685 19880 323715
rect 19680 323680 19880 323685
rect 19680 323635 19880 323640
rect 19680 323605 19685 323635
rect 19715 323605 19845 323635
rect 19875 323605 19880 323635
rect 19680 323600 19880 323605
rect 19680 323555 19880 323560
rect 19680 323525 19685 323555
rect 19715 323525 19845 323555
rect 19875 323525 19880 323555
rect 19680 323520 19880 323525
rect 19680 323475 19880 323480
rect 19680 323445 19685 323475
rect 19715 323445 19845 323475
rect 19875 323445 19880 323475
rect 19680 323440 19880 323445
rect 19680 323395 19880 323400
rect 19680 323365 19685 323395
rect 19715 323365 19845 323395
rect 19875 323365 19880 323395
rect 19680 323360 19880 323365
rect 19680 323315 19880 323320
rect 19680 323285 19685 323315
rect 19715 323285 19845 323315
rect 19875 323285 19880 323315
rect 19680 323280 19880 323285
rect 19680 323235 19880 323240
rect 19680 323205 19685 323235
rect 19715 323205 19845 323235
rect 19875 323205 19880 323235
rect 19680 323200 19880 323205
rect 19680 323155 19880 323160
rect 19680 323125 19685 323155
rect 19715 323125 19845 323155
rect 19875 323125 19880 323155
rect 19680 323120 19880 323125
rect 19680 323075 19880 323080
rect 19680 323045 19685 323075
rect 19715 323045 19845 323075
rect 19875 323045 19880 323075
rect 19680 323040 19880 323045
rect 19680 322995 19880 323000
rect 19680 322965 19685 322995
rect 19715 322965 19845 322995
rect 19875 322965 19880 322995
rect 19680 322960 19880 322965
rect 19680 322915 19880 322920
rect 19680 322885 19685 322915
rect 19715 322885 19845 322915
rect 19875 322885 19880 322915
rect 19680 322880 19880 322885
rect 19680 322835 19880 322840
rect 19680 322805 19685 322835
rect 19715 322805 19845 322835
rect 19875 322805 19880 322835
rect 19680 322800 19880 322805
rect 19680 322755 19880 322760
rect 19680 322725 19685 322755
rect 19715 322725 19845 322755
rect 19875 322725 19880 322755
rect 19680 322720 19880 322725
rect 19680 322675 19880 322680
rect 19680 322645 19685 322675
rect 19715 322645 19845 322675
rect 19875 322645 19880 322675
rect 19680 322640 19880 322645
rect 19680 322595 19880 322600
rect 19680 322565 19685 322595
rect 19715 322565 19845 322595
rect 19875 322565 19880 322595
rect 19680 322560 19880 322565
rect 19680 322515 19880 322520
rect 19680 322485 19685 322515
rect 19715 322485 19845 322515
rect 19875 322485 19880 322515
rect 19680 322480 19880 322485
rect 19680 322435 19880 322440
rect 19680 322405 19685 322435
rect 19715 322405 19845 322435
rect 19875 322405 19880 322435
rect 19680 322400 19880 322405
rect 19680 322355 19880 322360
rect 19680 322325 19685 322355
rect 19715 322325 19845 322355
rect 19875 322325 19880 322355
rect 19680 322320 19880 322325
rect 19680 322275 19880 322280
rect 19680 322245 19685 322275
rect 19715 322245 19845 322275
rect 19875 322245 19880 322275
rect 19680 322240 19880 322245
rect 19680 322195 19880 322200
rect 19680 322165 19685 322195
rect 19715 322165 19845 322195
rect 19875 322165 19880 322195
rect 19680 322160 19880 322165
rect 19680 322115 19880 322120
rect 19680 322085 19685 322115
rect 19715 322085 19845 322115
rect 19875 322085 19880 322115
rect 19680 322080 19880 322085
rect 19680 322035 19880 322040
rect 19680 322005 19685 322035
rect 19715 322005 19845 322035
rect 19875 322005 19880 322035
rect 19680 322000 19880 322005
rect 19680 321955 19880 321960
rect 19680 321925 19685 321955
rect 19715 321925 19845 321955
rect 19875 321925 19880 321955
rect 19680 321920 19880 321925
rect 19680 321875 19880 321880
rect 19680 321845 19685 321875
rect 19715 321845 19845 321875
rect 19875 321845 19880 321875
rect 19680 321840 19880 321845
rect 19680 321795 19880 321800
rect 19680 321765 19685 321795
rect 19715 321765 19845 321795
rect 19875 321765 19880 321795
rect 19680 321760 19880 321765
rect 19680 321715 19880 321720
rect 19680 321685 19685 321715
rect 19715 321685 19845 321715
rect 19875 321685 19880 321715
rect 19680 321680 19880 321685
rect 19680 321635 19880 321640
rect 19680 321605 19685 321635
rect 19715 321605 19845 321635
rect 19875 321605 19880 321635
rect 19680 321600 19880 321605
rect 19680 321555 19880 321560
rect 19680 321525 19685 321555
rect 19715 321525 19845 321555
rect 19875 321525 19880 321555
rect 19680 321520 19880 321525
rect 19680 321475 19880 321480
rect 19680 321445 19685 321475
rect 19715 321445 19845 321475
rect 19875 321445 19880 321475
rect 19680 321440 19880 321445
rect 19680 321395 19880 321400
rect 19680 321365 19685 321395
rect 19715 321365 19845 321395
rect 19875 321365 19880 321395
rect 19680 321360 19880 321365
rect 19680 321315 19880 321320
rect 19680 321285 19685 321315
rect 19715 321285 19845 321315
rect 19875 321285 19880 321315
rect 19680 321280 19880 321285
rect 19680 321235 19880 321240
rect 19680 321205 19685 321235
rect 19715 321205 19845 321235
rect 19875 321205 19880 321235
rect 19680 321200 19880 321205
rect 19680 321155 19880 321160
rect 19680 321125 19685 321155
rect 19715 321125 19845 321155
rect 19875 321125 19880 321155
rect 19680 321120 19880 321125
rect 19680 321075 19880 321080
rect 19680 321045 19685 321075
rect 19715 321045 19845 321075
rect 19875 321045 19880 321075
rect 19680 321040 19880 321045
rect 19680 320995 19880 321000
rect 19680 320965 19685 320995
rect 19715 320965 19845 320995
rect 19875 320965 19880 320995
rect 19680 320960 19880 320965
rect 19680 320915 19880 320920
rect 19680 320885 19685 320915
rect 19715 320885 19845 320915
rect 19875 320885 19880 320915
rect 19680 320880 19880 320885
rect 19680 320835 19880 320840
rect 19680 320805 19685 320835
rect 19715 320805 19845 320835
rect 19875 320805 19880 320835
rect 19680 320800 19880 320805
rect 19680 320755 19880 320760
rect 19680 320725 19685 320755
rect 19715 320725 19845 320755
rect 19875 320725 19880 320755
rect 19680 320720 19880 320725
rect 19680 320675 19880 320680
rect 19680 320645 19685 320675
rect 19715 320645 19845 320675
rect 19875 320645 19880 320675
rect 19680 320640 19880 320645
rect 19680 320595 19880 320600
rect 19680 320565 19685 320595
rect 19715 320565 19845 320595
rect 19875 320565 19880 320595
rect 19680 320560 19880 320565
rect 19680 320515 19880 320520
rect 19680 320485 19685 320515
rect 19715 320485 19845 320515
rect 19875 320485 19880 320515
rect 19680 320480 19880 320485
rect 19680 320435 19880 320440
rect 19680 320405 19685 320435
rect 19715 320405 19845 320435
rect 19875 320405 19880 320435
rect 19680 320400 19880 320405
rect 19680 320355 19880 320360
rect 19680 320325 19685 320355
rect 19715 320325 19845 320355
rect 19875 320325 19880 320355
rect 19680 320320 19880 320325
rect 19680 320275 19880 320280
rect 19680 320245 19685 320275
rect 19715 320245 19845 320275
rect 19875 320245 19880 320275
rect 19680 320240 19880 320245
rect 19680 320195 19880 320200
rect 19680 320165 19685 320195
rect 19715 320165 19845 320195
rect 19875 320165 19880 320195
rect 19680 320160 19880 320165
rect 19680 320115 19880 320120
rect 19680 320085 19685 320115
rect 19715 320085 19845 320115
rect 19875 320085 19880 320115
rect 19680 320080 19880 320085
rect 19680 320035 19880 320040
rect 19680 320005 19685 320035
rect 19715 320005 19845 320035
rect 19875 320005 19880 320035
rect 19680 320000 19880 320005
rect 19680 319955 19880 319960
rect 19680 319925 19685 319955
rect 19715 319925 19845 319955
rect 19875 319925 19880 319955
rect 19680 319920 19880 319925
rect 19680 319875 19880 319880
rect 19680 319845 19685 319875
rect 19715 319845 19845 319875
rect 19875 319845 19880 319875
rect 19680 319840 19880 319845
rect 19680 319795 19880 319800
rect 19680 319765 19685 319795
rect 19715 319765 19845 319795
rect 19875 319765 19880 319795
rect 19680 319760 19880 319765
rect 19680 319715 19880 319720
rect 19680 319685 19685 319715
rect 19715 319685 19845 319715
rect 19875 319685 19880 319715
rect 19680 319680 19880 319685
rect 19680 319635 19880 319640
rect 19680 319605 19685 319635
rect 19715 319605 19845 319635
rect 19875 319605 19880 319635
rect 19680 319600 19880 319605
rect 19680 319555 19880 319560
rect 19680 319525 19685 319555
rect 19715 319525 19845 319555
rect 19875 319525 19880 319555
rect 19680 319520 19880 319525
rect 19680 319475 19880 319480
rect 19680 319445 19685 319475
rect 19715 319445 19845 319475
rect 19875 319445 19880 319475
rect 19680 319440 19880 319445
rect 19680 319395 19880 319400
rect 19680 319365 19685 319395
rect 19715 319365 19845 319395
rect 19875 319365 19880 319395
rect 19680 319360 19880 319365
rect 19680 319315 19880 319320
rect 19680 319285 19685 319315
rect 19715 319285 19845 319315
rect 19875 319285 19880 319315
rect 19680 319280 19880 319285
rect 19680 319235 19880 319240
rect 19680 319205 19685 319235
rect 19715 319205 19845 319235
rect 19875 319205 19880 319235
rect 19680 319200 19880 319205
rect 19680 319155 19880 319160
rect 19680 319125 19685 319155
rect 19715 319125 19845 319155
rect 19875 319125 19880 319155
rect 19680 319120 19880 319125
rect 19680 319075 19880 319080
rect 19680 319045 19685 319075
rect 19715 319045 19845 319075
rect 19875 319045 19880 319075
rect 19680 319040 19880 319045
rect 19680 318995 19880 319000
rect 19680 318965 19685 318995
rect 19715 318965 19845 318995
rect 19875 318965 19880 318995
rect 19680 318960 19880 318965
rect 19680 318915 19880 318920
rect 19680 318885 19685 318915
rect 19715 318885 19845 318915
rect 19875 318885 19880 318915
rect 19680 318880 19880 318885
rect 19680 318835 19880 318840
rect 19680 318805 19685 318835
rect 19715 318805 19845 318835
rect 19875 318805 19880 318835
rect 19680 318800 19880 318805
rect 19680 318755 19880 318760
rect 19680 318725 19685 318755
rect 19715 318725 19845 318755
rect 19875 318725 19880 318755
rect 19680 318720 19880 318725
rect 19680 318675 19880 318680
rect 19680 318645 19685 318675
rect 19715 318645 19845 318675
rect 19875 318645 19880 318675
rect 19680 318640 19880 318645
rect 19680 318595 19880 318600
rect 19680 318565 19685 318595
rect 19715 318565 19845 318595
rect 19875 318565 19880 318595
rect 19680 318560 19880 318565
rect 19680 318515 19880 318520
rect 19680 318485 19685 318515
rect 19715 318485 19845 318515
rect 19875 318485 19880 318515
rect 19680 318480 19880 318485
rect 19680 318435 19880 318440
rect 19680 318405 19685 318435
rect 19715 318405 19845 318435
rect 19875 318405 19880 318435
rect 19680 318400 19880 318405
rect 19680 318355 19880 318360
rect 19680 318325 19685 318355
rect 19715 318325 19845 318355
rect 19875 318325 19880 318355
rect 19680 318320 19880 318325
rect 19680 318275 19880 318280
rect 19680 318245 19685 318275
rect 19715 318245 19845 318275
rect 19875 318245 19880 318275
rect 19680 318240 19880 318245
rect 19680 318195 19880 318200
rect 19680 318165 19685 318195
rect 19715 318165 19845 318195
rect 19875 318165 19880 318195
rect 19680 318160 19880 318165
rect 19680 318115 19880 318120
rect 19680 318085 19685 318115
rect 19715 318085 19845 318115
rect 19875 318085 19880 318115
rect 19680 318080 19880 318085
rect 19680 318035 19880 318040
rect 19680 318005 19685 318035
rect 19715 318005 19845 318035
rect 19875 318005 19880 318035
rect 19680 318000 19880 318005
rect 19680 317955 19880 317960
rect 19680 317925 19685 317955
rect 19715 317925 19845 317955
rect 19875 317925 19880 317955
rect 19680 317920 19880 317925
rect 19680 317875 19880 317880
rect 19680 317845 19685 317875
rect 19715 317845 19845 317875
rect 19875 317845 19880 317875
rect 19680 317840 19880 317845
rect 19680 317795 19880 317800
rect 19680 317765 19685 317795
rect 19715 317765 19845 317795
rect 19875 317765 19880 317795
rect 19680 317760 19880 317765
rect 19680 317715 19880 317720
rect 19680 317685 19685 317715
rect 19715 317685 19845 317715
rect 19875 317685 19880 317715
rect 19680 317680 19880 317685
rect 19680 317635 19880 317640
rect 19680 317605 19685 317635
rect 19715 317605 19845 317635
rect 19875 317605 19880 317635
rect 19680 317600 19880 317605
rect 19680 317555 19880 317560
rect 19680 317525 19685 317555
rect 19715 317525 19845 317555
rect 19875 317525 19880 317555
rect 19680 317520 19880 317525
rect 19680 317475 19880 317480
rect 19680 317445 19685 317475
rect 19715 317445 19845 317475
rect 19875 317445 19880 317475
rect 19680 317440 19880 317445
rect 19680 317395 19880 317400
rect 19680 317365 19685 317395
rect 19715 317365 19845 317395
rect 19875 317365 19880 317395
rect 19680 317360 19880 317365
rect 19680 317315 19880 317320
rect 19680 317285 19685 317315
rect 19715 317285 19845 317315
rect 19875 317285 19880 317315
rect 19680 317280 19880 317285
rect 19680 317235 19880 317240
rect 19680 317205 19685 317235
rect 19715 317205 19845 317235
rect 19875 317205 19880 317235
rect 19680 317200 19880 317205
rect 19680 317155 19880 317160
rect 19680 317125 19685 317155
rect 19715 317125 19845 317155
rect 19875 317125 19880 317155
rect 19680 317120 19880 317125
rect 19680 317075 19880 317080
rect 19680 317045 19685 317075
rect 19715 317045 19845 317075
rect 19875 317045 19880 317075
rect 19680 317040 19880 317045
rect 19680 316995 19880 317000
rect 19680 316965 19685 316995
rect 19715 316965 19845 316995
rect 19875 316965 19880 316995
rect 19680 316960 19880 316965
rect 19680 316915 19880 316920
rect 19680 316885 19685 316915
rect 19715 316885 19845 316915
rect 19875 316885 19880 316915
rect 19680 316880 19880 316885
rect 19680 316835 19880 316840
rect 19680 316805 19685 316835
rect 19715 316805 19845 316835
rect 19875 316805 19880 316835
rect 19680 316800 19880 316805
rect 19680 316755 19880 316760
rect 19680 316725 19685 316755
rect 19715 316725 19845 316755
rect 19875 316725 19880 316755
rect 19680 316720 19880 316725
rect 19680 316675 19880 316680
rect 19680 316645 19685 316675
rect 19715 316645 19845 316675
rect 19875 316645 19880 316675
rect 19680 316640 19880 316645
rect 19680 316595 19880 316600
rect 19680 316565 19685 316595
rect 19715 316565 19845 316595
rect 19875 316565 19880 316595
rect 19680 316560 19880 316565
rect 19680 316515 19880 316520
rect 19680 316485 19685 316515
rect 19715 316485 19845 316515
rect 19875 316485 19880 316515
rect 19680 316480 19880 316485
rect 19680 316435 19880 316440
rect 19680 316405 19685 316435
rect 19715 316405 19845 316435
rect 19875 316405 19880 316435
rect 19680 316400 19880 316405
rect 19680 316355 19880 316360
rect 19680 316325 19685 316355
rect 19715 316325 19845 316355
rect 19875 316325 19880 316355
rect 19680 316320 19880 316325
rect 19680 316275 19880 316280
rect 19680 316245 19685 316275
rect 19715 316245 19845 316275
rect 19875 316245 19880 316275
rect 19680 316240 19880 316245
rect 19680 316195 19880 316200
rect 19680 316165 19685 316195
rect 19715 316165 19845 316195
rect 19875 316165 19880 316195
rect 19680 316160 19880 316165
rect 19680 316115 19880 316120
rect 19680 316085 19685 316115
rect 19715 316085 19845 316115
rect 19875 316085 19880 316115
rect 19680 316080 19880 316085
rect 19680 316035 19880 316040
rect 19680 316005 19685 316035
rect 19715 316005 19845 316035
rect 19875 316005 19880 316035
rect 19680 316000 19880 316005
rect 19680 315955 19880 315960
rect 19680 315925 19685 315955
rect 19715 315925 19845 315955
rect 19875 315925 19880 315955
rect 19680 315920 19880 315925
rect 19680 315875 19880 315880
rect 19680 315845 19685 315875
rect 19715 315845 19845 315875
rect 19875 315845 19880 315875
rect 19680 315840 19880 315845
rect 19680 315795 19880 315800
rect 19680 315765 19685 315795
rect 19715 315765 19845 315795
rect 19875 315765 19880 315795
rect 19680 315760 19880 315765
rect 19680 315715 19880 315720
rect 19680 315685 19685 315715
rect 19715 315685 19845 315715
rect 19875 315685 19880 315715
rect 19680 315680 19880 315685
rect 19680 315635 19880 315640
rect 19680 315605 19685 315635
rect 19715 315605 19845 315635
rect 19875 315605 19880 315635
rect 19680 315600 19880 315605
rect 19680 315555 19880 315560
rect 19680 315525 19685 315555
rect 19715 315525 19845 315555
rect 19875 315525 19880 315555
rect 19680 315520 19880 315525
rect 19680 315475 19880 315480
rect 19680 315445 19685 315475
rect 19715 315445 19845 315475
rect 19875 315445 19880 315475
rect 19680 315440 19880 315445
rect 19680 315395 19880 315400
rect 19680 315365 19685 315395
rect 19715 315365 19845 315395
rect 19875 315365 19880 315395
rect 19680 315360 19880 315365
rect 19680 315315 19880 315320
rect 19680 315285 19685 315315
rect 19715 315285 19845 315315
rect 19875 315285 19880 315315
rect 19680 315280 19880 315285
rect 19680 315235 19880 315240
rect 19680 315205 19685 315235
rect 19715 315205 19845 315235
rect 19875 315205 19880 315235
rect 19680 315200 19880 315205
rect 19680 315155 19880 315160
rect 19680 315125 19685 315155
rect 19715 315125 19845 315155
rect 19875 315125 19880 315155
rect 19680 315120 19880 315125
rect 19680 315075 19880 315080
rect 19680 315045 19685 315075
rect 19715 315045 19845 315075
rect 19875 315045 19880 315075
rect 19680 315040 19880 315045
rect 19680 314995 19880 315000
rect 19680 314965 19685 314995
rect 19715 314965 19845 314995
rect 19875 314965 19880 314995
rect 19680 314960 19880 314965
rect 19680 314915 19880 314920
rect 19680 314885 19685 314915
rect 19715 314885 19845 314915
rect 19875 314885 19880 314915
rect 19680 314880 19880 314885
rect 19680 314835 19880 314840
rect 19680 314805 19685 314835
rect 19715 314805 19845 314835
rect 19875 314805 19880 314835
rect 19680 314800 19880 314805
rect 19680 314755 19880 314760
rect 19680 314725 19685 314755
rect 19715 314725 19845 314755
rect 19875 314725 19880 314755
rect 19680 314720 19880 314725
rect 19680 314675 19880 314680
rect 19680 314645 19685 314675
rect 19715 314645 19845 314675
rect 19875 314645 19880 314675
rect 19680 314640 19880 314645
rect 19680 314595 19880 314600
rect 19680 314565 19685 314595
rect 19715 314565 19845 314595
rect 19875 314565 19880 314595
rect 19680 314560 19880 314565
rect 19680 314515 19880 314520
rect 19680 314485 19685 314515
rect 19715 314485 19845 314515
rect 19875 314485 19880 314515
rect 19680 314480 19880 314485
rect 19680 314435 19880 314440
rect 19680 314405 19685 314435
rect 19715 314405 19845 314435
rect 19875 314405 19880 314435
rect 19680 314400 19880 314405
rect 19680 314355 19880 314360
rect 19680 314325 19685 314355
rect 19715 314325 19845 314355
rect 19875 314325 19880 314355
rect 19680 314320 19880 314325
rect 19680 314275 19880 314280
rect 19680 314245 19685 314275
rect 19715 314245 19845 314275
rect 19875 314245 19880 314275
rect 19680 314240 19880 314245
rect 19680 314195 19880 314200
rect 19680 314165 19685 314195
rect 19715 314165 19845 314195
rect 19875 314165 19880 314195
rect 19680 314160 19880 314165
rect 19680 314115 19880 314120
rect 19680 314085 19685 314115
rect 19715 314085 19845 314115
rect 19875 314085 19880 314115
rect 19680 314080 19880 314085
rect 19680 314035 19880 314040
rect 19680 314005 19685 314035
rect 19715 314005 19845 314035
rect 19875 314005 19880 314035
rect 19680 314000 19880 314005
rect 19680 313955 19880 313960
rect 19680 313925 19685 313955
rect 19715 313925 19845 313955
rect 19875 313925 19880 313955
rect 19680 313920 19880 313925
rect 19680 313875 19880 313880
rect 19680 313845 19685 313875
rect 19715 313845 19845 313875
rect 19875 313845 19880 313875
rect 19680 313840 19880 313845
rect 19680 313795 19880 313800
rect 19680 313765 19685 313795
rect 19715 313765 19845 313795
rect 19875 313765 19880 313795
rect 19680 313760 19880 313765
rect 19680 313715 19880 313720
rect 19680 313685 19685 313715
rect 19715 313685 19845 313715
rect 19875 313685 19880 313715
rect 19680 313680 19880 313685
rect 19680 313635 19880 313640
rect 19680 313605 19685 313635
rect 19715 313605 19845 313635
rect 19875 313605 19880 313635
rect 19680 313600 19880 313605
rect 19680 313555 19880 313560
rect 19680 313525 19685 313555
rect 19715 313525 19845 313555
rect 19875 313525 19880 313555
rect 19680 313520 19880 313525
rect 19680 313475 19880 313480
rect 19680 313445 19685 313475
rect 19715 313445 19845 313475
rect 19875 313445 19880 313475
rect 19680 313440 19880 313445
rect 19680 313395 19880 313400
rect 19680 313365 19685 313395
rect 19715 313365 19845 313395
rect 19875 313365 19880 313395
rect 19680 313360 19880 313365
rect 19680 313315 19880 313320
rect 19680 313285 19685 313315
rect 19715 313285 19845 313315
rect 19875 313285 19880 313315
rect 19680 313280 19880 313285
rect 19680 313235 19880 313240
rect 19680 313205 19685 313235
rect 19715 313205 19845 313235
rect 19875 313205 19880 313235
rect 19680 313200 19880 313205
rect 19680 313155 19880 313160
rect 19680 313125 19685 313155
rect 19715 313125 19845 313155
rect 19875 313125 19880 313155
rect 19680 313120 19880 313125
rect 19680 313075 19880 313080
rect 19680 313045 19685 313075
rect 19715 313045 19845 313075
rect 19875 313045 19880 313075
rect 19680 313040 19880 313045
rect 19680 312995 19880 313000
rect 19680 312965 19685 312995
rect 19715 312965 19845 312995
rect 19875 312965 19880 312995
rect 19680 312960 19880 312965
rect 19680 312915 19880 312920
rect 19680 312885 19685 312915
rect 19715 312885 19845 312915
rect 19875 312885 19880 312915
rect 19680 312880 19880 312885
rect 19680 312835 19880 312840
rect 19680 312805 19685 312835
rect 19715 312805 19845 312835
rect 19875 312805 19880 312835
rect 19680 312800 19880 312805
rect 19680 312755 19880 312760
rect 19680 312725 19685 312755
rect 19715 312725 19845 312755
rect 19875 312725 19880 312755
rect 19680 312720 19880 312725
rect 19680 312675 19880 312680
rect 19680 312645 19685 312675
rect 19715 312645 19845 312675
rect 19875 312645 19880 312675
rect 19680 312640 19880 312645
rect 19680 312595 19880 312600
rect 19680 312565 19685 312595
rect 19715 312565 19845 312595
rect 19875 312565 19880 312595
rect 19680 312560 19880 312565
rect 19680 312515 19880 312520
rect 19680 312485 19685 312515
rect 19715 312485 19845 312515
rect 19875 312485 19880 312515
rect 19680 312480 19880 312485
rect 19680 312435 19880 312440
rect 19680 312405 19685 312435
rect 19715 312405 19845 312435
rect 19875 312405 19880 312435
rect 19680 312400 19880 312405
rect 19680 312355 19880 312360
rect 19680 312325 19685 312355
rect 19715 312325 19845 312355
rect 19875 312325 19880 312355
rect 19680 312320 19880 312325
rect 19680 312275 19880 312280
rect 19680 312245 19685 312275
rect 19715 312245 19845 312275
rect 19875 312245 19880 312275
rect 19680 312240 19880 312245
rect 19680 312195 19880 312200
rect 19680 312165 19685 312195
rect 19715 312165 19845 312195
rect 19875 312165 19880 312195
rect 19680 312160 19880 312165
rect 19680 312115 19880 312120
rect 19680 312085 19685 312115
rect 19715 312085 19845 312115
rect 19875 312085 19880 312115
rect 19680 312080 19880 312085
rect 19680 312035 19880 312040
rect 19680 312005 19685 312035
rect 19715 312005 19845 312035
rect 19875 312005 19880 312035
rect 19680 312000 19880 312005
rect 19680 311955 19880 311960
rect 19680 311925 19685 311955
rect 19715 311925 19845 311955
rect 19875 311925 19880 311955
rect 19680 311920 19880 311925
rect 19680 311875 19880 311880
rect 19680 311845 19685 311875
rect 19715 311845 19845 311875
rect 19875 311845 19880 311875
rect 19680 311840 19880 311845
rect 19680 311795 19880 311800
rect 19680 311765 19685 311795
rect 19715 311765 19845 311795
rect 19875 311765 19880 311795
rect 19680 311760 19880 311765
rect 19680 311715 19880 311720
rect 19680 311685 19685 311715
rect 19715 311685 19845 311715
rect 19875 311685 19880 311715
rect 19680 311680 19880 311685
rect 19680 311635 19880 311640
rect 19680 311605 19685 311635
rect 19715 311605 19845 311635
rect 19875 311605 19880 311635
rect 19680 311600 19880 311605
rect 19680 311555 19880 311560
rect 19680 311525 19685 311555
rect 19715 311525 19845 311555
rect 19875 311525 19880 311555
rect 19680 311520 19880 311525
rect 19680 311475 19880 311480
rect 19680 311445 19685 311475
rect 19715 311445 19845 311475
rect 19875 311445 19880 311475
rect 19680 311440 19880 311445
rect 19680 311395 19880 311400
rect 19680 311365 19685 311395
rect 19715 311365 19845 311395
rect 19875 311365 19880 311395
rect 19680 311360 19880 311365
rect 19680 311315 19880 311320
rect 19680 311285 19685 311315
rect 19715 311285 19845 311315
rect 19875 311285 19880 311315
rect 19680 311280 19880 311285
rect 19680 311235 19880 311240
rect 19680 311205 19685 311235
rect 19715 311205 19845 311235
rect 19875 311205 19880 311235
rect 19680 311200 19880 311205
rect 19680 311155 19880 311160
rect 19680 311125 19685 311155
rect 19715 311125 19845 311155
rect 19875 311125 19880 311155
rect 19680 311120 19880 311125
rect 19680 311075 19880 311080
rect 19680 311045 19685 311075
rect 19715 311045 19845 311075
rect 19875 311045 19880 311075
rect 19680 311040 19880 311045
rect 19680 310995 19880 311000
rect 19680 310965 19685 310995
rect 19715 310965 19845 310995
rect 19875 310965 19880 310995
rect 19680 310960 19880 310965
rect 19680 310915 19880 310920
rect 19680 310885 19685 310915
rect 19715 310885 19845 310915
rect 19875 310885 19880 310915
rect 19680 310880 19880 310885
rect 19680 310835 19880 310840
rect 19680 310805 19685 310835
rect 19715 310805 19845 310835
rect 19875 310805 19880 310835
rect 19680 310800 19880 310805
rect 19680 310755 19880 310760
rect 19680 310725 19685 310755
rect 19715 310725 19845 310755
rect 19875 310725 19880 310755
rect 19680 310720 19880 310725
rect 19680 310675 19880 310680
rect 19680 310645 19685 310675
rect 19715 310645 19845 310675
rect 19875 310645 19880 310675
rect 19680 310640 19880 310645
rect 19680 310595 19880 310600
rect 19680 310565 19685 310595
rect 19715 310565 19845 310595
rect 19875 310565 19880 310595
rect 19680 310560 19880 310565
rect 19680 310515 19880 310520
rect 19680 310485 19685 310515
rect 19715 310485 19845 310515
rect 19875 310485 19880 310515
rect 19680 310480 19880 310485
rect 19680 310435 19880 310440
rect 19680 310405 19685 310435
rect 19715 310405 19845 310435
rect 19875 310405 19880 310435
rect 19680 310400 19880 310405
rect 19680 310355 19880 310360
rect 19680 310325 19685 310355
rect 19715 310325 19845 310355
rect 19875 310325 19880 310355
rect 19680 310320 19880 310325
rect 19680 310275 19880 310280
rect 19680 310245 19685 310275
rect 19715 310245 19845 310275
rect 19875 310245 19880 310275
rect 19680 310240 19880 310245
rect 19680 310195 19880 310200
rect 19680 310165 19685 310195
rect 19715 310165 19845 310195
rect 19875 310165 19880 310195
rect 19680 310160 19880 310165
rect 19680 310115 19880 310120
rect 19680 310085 19685 310115
rect 19715 310085 19845 310115
rect 19875 310085 19880 310115
rect 19680 310080 19880 310085
rect 19680 310035 19880 310040
rect 19680 310005 19685 310035
rect 19715 310005 19845 310035
rect 19875 310005 19880 310035
rect 19680 310000 19880 310005
rect 19680 309955 19880 309960
rect 19680 309925 19685 309955
rect 19715 309925 19845 309955
rect 19875 309925 19880 309955
rect 19680 309920 19880 309925
rect 19680 309875 19880 309880
rect 19680 309845 19685 309875
rect 19715 309845 19845 309875
rect 19875 309845 19880 309875
rect 19680 309840 19880 309845
rect 19680 309795 19880 309800
rect 19680 309765 19685 309795
rect 19715 309765 19845 309795
rect 19875 309765 19880 309795
rect 19680 309760 19880 309765
rect 19680 309715 19880 309720
rect 19680 309685 19685 309715
rect 19715 309685 19845 309715
rect 19875 309685 19880 309715
rect 19680 309680 19880 309685
rect 19680 309635 19880 309640
rect 19680 309605 19685 309635
rect 19715 309605 19845 309635
rect 19875 309605 19880 309635
rect 19680 309600 19880 309605
rect 19680 309555 19880 309560
rect 19680 309525 19685 309555
rect 19715 309525 19845 309555
rect 19875 309525 19880 309555
rect 19680 309520 19880 309525
rect 19680 309475 19880 309480
rect 19680 309445 19685 309475
rect 19715 309445 19845 309475
rect 19875 309445 19880 309475
rect 19680 309440 19880 309445
rect 19680 309395 19880 309400
rect 19680 309365 19685 309395
rect 19715 309365 19845 309395
rect 19875 309365 19880 309395
rect 19680 309360 19880 309365
rect 19680 309315 19880 309320
rect 19680 309285 19685 309315
rect 19715 309285 19845 309315
rect 19875 309285 19880 309315
rect 19680 309280 19880 309285
rect 19680 309235 19880 309240
rect 19680 309205 19685 309235
rect 19715 309205 19845 309235
rect 19875 309205 19880 309235
rect 19680 309200 19880 309205
rect 19680 309155 19880 309160
rect 19680 309125 19685 309155
rect 19715 309125 19845 309155
rect 19875 309125 19880 309155
rect 19680 309120 19880 309125
rect 19680 309075 19880 309080
rect 19680 309045 19685 309075
rect 19715 309045 19845 309075
rect 19875 309045 19880 309075
rect 19680 309040 19880 309045
rect 19680 308995 19880 309000
rect 19680 308965 19685 308995
rect 19715 308965 19845 308995
rect 19875 308965 19880 308995
rect 19680 308960 19880 308965
rect 19680 308915 19880 308920
rect 19680 308885 19685 308915
rect 19715 308885 19845 308915
rect 19875 308885 19880 308915
rect 19680 308880 19880 308885
rect 19680 308835 19880 308840
rect 19680 308805 19685 308835
rect 19715 308805 19845 308835
rect 19875 308805 19880 308835
rect 19680 308800 19880 308805
rect 19680 308755 19880 308760
rect 19680 308725 19685 308755
rect 19715 308725 19845 308755
rect 19875 308725 19880 308755
rect 19680 308720 19880 308725
rect 19680 308675 19880 308680
rect 19680 308645 19685 308675
rect 19715 308645 19845 308675
rect 19875 308645 19880 308675
rect 19680 308640 19880 308645
rect 19680 308595 19880 308600
rect 19680 308565 19685 308595
rect 19715 308565 19845 308595
rect 19875 308565 19880 308595
rect 19680 308560 19880 308565
rect 19680 308515 19880 308520
rect 19680 308485 19685 308515
rect 19715 308485 19845 308515
rect 19875 308485 19880 308515
rect 19680 308480 19880 308485
rect 19680 308435 19880 308440
rect 19680 308405 19685 308435
rect 19715 308405 19845 308435
rect 19875 308405 19880 308435
rect 19680 308400 19880 308405
rect 19680 308355 19880 308360
rect 19680 308325 19685 308355
rect 19715 308325 19845 308355
rect 19875 308325 19880 308355
rect 19680 308320 19880 308325
rect 19680 308275 19880 308280
rect 19680 308245 19685 308275
rect 19715 308245 19845 308275
rect 19875 308245 19880 308275
rect 19680 308240 19880 308245
rect 19680 308195 19880 308200
rect 19680 308165 19685 308195
rect 19715 308165 19845 308195
rect 19875 308165 19880 308195
rect 19680 308160 19880 308165
rect 19680 308115 19880 308120
rect 19680 308085 19685 308115
rect 19715 308085 19845 308115
rect 19875 308085 19880 308115
rect 19680 308080 19880 308085
rect 19680 308035 19880 308040
rect 19680 308005 19685 308035
rect 19715 308005 19845 308035
rect 19875 308005 19880 308035
rect 19680 308000 19880 308005
rect 19680 307955 19880 307960
rect 19680 307925 19685 307955
rect 19715 307925 19845 307955
rect 19875 307925 19880 307955
rect 19680 307920 19880 307925
rect 19680 307875 19880 307880
rect 19680 307845 19685 307875
rect 19715 307845 19845 307875
rect 19875 307845 19880 307875
rect 19680 307840 19880 307845
rect 19680 307795 19880 307800
rect 19680 307765 19685 307795
rect 19715 307765 19845 307795
rect 19875 307765 19880 307795
rect 19680 307760 19880 307765
rect 19680 307715 19880 307720
rect 19680 307685 19685 307715
rect 19715 307685 19845 307715
rect 19875 307685 19880 307715
rect 19680 307680 19880 307685
rect 19680 307635 19880 307640
rect 19680 307605 19685 307635
rect 19715 307605 19845 307635
rect 19875 307605 19880 307635
rect 19680 307600 19880 307605
rect 19680 307555 19880 307560
rect 19680 307525 19685 307555
rect 19715 307525 19845 307555
rect 19875 307525 19880 307555
rect 19680 307520 19880 307525
rect 19680 307475 19880 307480
rect 19680 307445 19685 307475
rect 19715 307445 19845 307475
rect 19875 307445 19880 307475
rect 19680 307440 19880 307445
rect 19680 307395 19880 307400
rect 19680 307365 19685 307395
rect 19715 307365 19845 307395
rect 19875 307365 19880 307395
rect 19680 307360 19880 307365
rect 19680 307315 19880 307320
rect 19680 307285 19685 307315
rect 19715 307285 19845 307315
rect 19875 307285 19880 307315
rect 19680 307280 19880 307285
rect 19680 307235 19880 307240
rect 19680 307205 19685 307235
rect 19715 307205 19845 307235
rect 19875 307205 19880 307235
rect 19680 307200 19880 307205
rect 19680 307155 19880 307160
rect 19680 307125 19685 307155
rect 19715 307125 19845 307155
rect 19875 307125 19880 307155
rect 19680 307120 19880 307125
rect 19680 307075 19880 307080
rect 19680 307045 19685 307075
rect 19715 307045 19845 307075
rect 19875 307045 19880 307075
rect 19680 307040 19880 307045
rect 19680 306995 19880 307000
rect 19680 306965 19685 306995
rect 19715 306965 19845 306995
rect 19875 306965 19880 306995
rect 19680 306960 19880 306965
rect 19680 306915 19880 306920
rect 19680 306885 19685 306915
rect 19715 306885 19845 306915
rect 19875 306885 19880 306915
rect 19680 306880 19880 306885
rect 19680 306835 19880 306840
rect 19680 306805 19685 306835
rect 19715 306805 19845 306835
rect 19875 306805 19880 306835
rect 19680 306800 19880 306805
rect 19680 306755 19880 306760
rect 19680 306725 19685 306755
rect 19715 306725 19845 306755
rect 19875 306725 19880 306755
rect 19680 306720 19880 306725
rect 19680 306675 19880 306680
rect 19680 306645 19685 306675
rect 19715 306645 19845 306675
rect 19875 306645 19880 306675
rect 19680 306640 19880 306645
rect 19680 306595 19880 306600
rect 19680 306565 19685 306595
rect 19715 306565 19845 306595
rect 19875 306565 19880 306595
rect 19680 306560 19880 306565
rect 19680 306515 19880 306520
rect 19680 306485 19685 306515
rect 19715 306485 19845 306515
rect 19875 306485 19880 306515
rect 19680 306480 19880 306485
rect 19680 306435 19880 306440
rect 19680 306405 19685 306435
rect 19715 306405 19845 306435
rect 19875 306405 19880 306435
rect 19680 306400 19880 306405
rect 19680 306355 19880 306360
rect 19680 306325 19685 306355
rect 19715 306325 19845 306355
rect 19875 306325 19880 306355
rect 19680 306320 19880 306325
rect 19680 306275 19880 306280
rect 19680 306245 19685 306275
rect 19715 306245 19845 306275
rect 19875 306245 19880 306275
rect 19680 306240 19880 306245
rect 19680 306195 19880 306200
rect 19680 306165 19685 306195
rect 19715 306165 19845 306195
rect 19875 306165 19880 306195
rect 19680 306160 19880 306165
rect 19680 306115 19880 306120
rect 19680 306085 19685 306115
rect 19715 306085 19845 306115
rect 19875 306085 19880 306115
rect 19680 306080 19880 306085
rect 19680 306035 19880 306040
rect 19680 306005 19685 306035
rect 19715 306005 19845 306035
rect 19875 306005 19880 306035
rect 19680 306000 19880 306005
rect 19680 305955 19880 305960
rect 19680 305925 19685 305955
rect 19715 305925 19845 305955
rect 19875 305925 19880 305955
rect 19680 305920 19880 305925
rect 19680 305875 19880 305880
rect 19680 305845 19685 305875
rect 19715 305845 19845 305875
rect 19875 305845 19880 305875
rect 19680 305840 19880 305845
rect 19680 305795 19880 305800
rect 19680 305765 19685 305795
rect 19715 305765 19845 305795
rect 19875 305765 19880 305795
rect 19680 305760 19880 305765
rect 19680 305715 19880 305720
rect 19680 305685 19685 305715
rect 19715 305685 19845 305715
rect 19875 305685 19880 305715
rect 19680 305680 19880 305685
rect 19680 305635 19880 305640
rect 19680 305605 19685 305635
rect 19715 305605 19845 305635
rect 19875 305605 19880 305635
rect 19680 305600 19880 305605
rect 19680 305555 19880 305560
rect 19680 305525 19685 305555
rect 19715 305525 19845 305555
rect 19875 305525 19880 305555
rect 19680 305520 19880 305525
rect 19680 305475 19880 305480
rect 19680 305445 19685 305475
rect 19715 305445 19845 305475
rect 19875 305445 19880 305475
rect 19680 305440 19880 305445
rect 19680 305395 19880 305400
rect 19680 305365 19685 305395
rect 19715 305365 19845 305395
rect 19875 305365 19880 305395
rect 19680 305360 19880 305365
rect 19680 305315 19880 305320
rect 19680 305285 19685 305315
rect 19715 305285 19845 305315
rect 19875 305285 19880 305315
rect 19680 305280 19880 305285
rect 19680 305235 19880 305240
rect 19680 305205 19685 305235
rect 19715 305205 19845 305235
rect 19875 305205 19880 305235
rect 19680 305200 19880 305205
rect 19680 305155 19880 305160
rect 19680 305125 19685 305155
rect 19715 305125 19845 305155
rect 19875 305125 19880 305155
rect 19680 305120 19880 305125
rect 19680 305075 19880 305080
rect 19680 305045 19685 305075
rect 19715 305045 19845 305075
rect 19875 305045 19880 305075
rect 19680 305040 19880 305045
rect 19680 304995 19880 305000
rect 19680 304965 19685 304995
rect 19715 304965 19845 304995
rect 19875 304965 19880 304995
rect 19680 304960 19880 304965
rect 19680 304915 19880 304920
rect 19680 304885 19685 304915
rect 19715 304885 19845 304915
rect 19875 304885 19880 304915
rect 19680 304880 19880 304885
rect 19680 304835 19880 304840
rect 19680 304805 19685 304835
rect 19715 304805 19845 304835
rect 19875 304805 19880 304835
rect 19680 304800 19880 304805
rect 19680 304755 19880 304760
rect 19680 304725 19685 304755
rect 19715 304725 19845 304755
rect 19875 304725 19880 304755
rect 19680 304720 19880 304725
rect 19680 304675 19880 304680
rect 19680 304645 19685 304675
rect 19715 304645 19845 304675
rect 19875 304645 19880 304675
rect 19680 304640 19880 304645
rect 19680 304595 19880 304600
rect 19680 304565 19685 304595
rect 19715 304565 19845 304595
rect 19875 304565 19880 304595
rect 19680 304560 19880 304565
rect 19680 304515 19880 304520
rect 19680 304485 19685 304515
rect 19715 304485 19845 304515
rect 19875 304485 19880 304515
rect 19680 304480 19880 304485
rect 19680 304435 19880 304440
rect 19680 304405 19685 304435
rect 19715 304405 19845 304435
rect 19875 304405 19880 304435
rect 19680 304400 19880 304405
rect 19680 304355 19880 304360
rect 19680 304325 19685 304355
rect 19715 304325 19845 304355
rect 19875 304325 19880 304355
rect 19680 304320 19880 304325
rect 19680 304275 19880 304280
rect 19680 304245 19685 304275
rect 19715 304245 19845 304275
rect 19875 304245 19880 304275
rect 19680 304240 19880 304245
rect 19680 304195 19880 304200
rect 19680 304165 19685 304195
rect 19715 304165 19845 304195
rect 19875 304165 19880 304195
rect 19680 304160 19880 304165
rect 19680 304115 19880 304120
rect 19680 304085 19685 304115
rect 19715 304085 19845 304115
rect 19875 304085 19880 304115
rect 19680 304080 19880 304085
rect 19680 304035 19880 304040
rect 19680 304005 19685 304035
rect 19715 304005 19845 304035
rect 19875 304005 19880 304035
rect 19680 304000 19880 304005
rect 19680 303955 19880 303960
rect 19680 303925 19685 303955
rect 19715 303925 19845 303955
rect 19875 303925 19880 303955
rect 19680 303920 19880 303925
rect 19680 303875 19880 303880
rect 19680 303845 19685 303875
rect 19715 303845 19845 303875
rect 19875 303845 19880 303875
rect 19680 303840 19880 303845
rect 19680 303795 19880 303800
rect 19680 303765 19685 303795
rect 19715 303765 19845 303795
rect 19875 303765 19880 303795
rect 19680 303760 19880 303765
rect 19680 303715 19880 303720
rect 19680 303685 19685 303715
rect 19715 303685 19845 303715
rect 19875 303685 19880 303715
rect 19680 303680 19880 303685
rect 19680 303635 19880 303640
rect 19680 303605 19685 303635
rect 19715 303605 19845 303635
rect 19875 303605 19880 303635
rect 19680 303600 19880 303605
rect 19680 303555 19880 303560
rect 19680 303525 19685 303555
rect 19715 303525 19845 303555
rect 19875 303525 19880 303555
rect 19680 303520 19880 303525
rect 19680 303475 19880 303480
rect 19680 303445 19685 303475
rect 19715 303445 19845 303475
rect 19875 303445 19880 303475
rect 19680 303440 19880 303445
rect 19680 303395 19880 303400
rect 19680 303365 19685 303395
rect 19715 303365 19845 303395
rect 19875 303365 19880 303395
rect 19680 303360 19880 303365
rect 19680 303315 19880 303320
rect 19680 303285 19685 303315
rect 19715 303285 19845 303315
rect 19875 303285 19880 303315
rect 19680 303280 19880 303285
rect 19680 303235 19880 303240
rect 19680 303205 19685 303235
rect 19715 303205 19845 303235
rect 19875 303205 19880 303235
rect 19680 303200 19880 303205
rect 19680 303155 19880 303160
rect 19680 303125 19685 303155
rect 19715 303125 19845 303155
rect 19875 303125 19880 303155
rect 19680 303120 19880 303125
rect 19680 303075 19880 303080
rect 19680 303045 19685 303075
rect 19715 303045 19845 303075
rect 19875 303045 19880 303075
rect 19680 303040 19880 303045
rect 19680 302995 19880 303000
rect 19680 302965 19685 302995
rect 19715 302965 19845 302995
rect 19875 302965 19880 302995
rect 19680 302960 19880 302965
rect 19680 302915 19880 302920
rect 19680 302885 19685 302915
rect 19715 302885 19845 302915
rect 19875 302885 19880 302915
rect 19680 302880 19880 302885
rect 19680 302835 19880 302840
rect 19680 302805 19685 302835
rect 19715 302805 19845 302835
rect 19875 302805 19880 302835
rect 19680 302800 19880 302805
rect 19680 302755 19880 302760
rect 19680 302725 19685 302755
rect 19715 302725 19845 302755
rect 19875 302725 19880 302755
rect 19680 302720 19880 302725
rect 19680 302675 19880 302680
rect 19680 302645 19685 302675
rect 19715 302645 19845 302675
rect 19875 302645 19880 302675
rect 19680 302640 19880 302645
rect 19680 302595 19880 302600
rect 19680 302565 19685 302595
rect 19715 302565 19845 302595
rect 19875 302565 19880 302595
rect 19680 302560 19880 302565
rect 19680 302515 19880 302520
rect 19680 302485 19685 302515
rect 19715 302485 19845 302515
rect 19875 302485 19880 302515
rect 19680 302480 19880 302485
rect 19680 302435 19880 302440
rect 19680 302405 19685 302435
rect 19715 302405 19845 302435
rect 19875 302405 19880 302435
rect 19680 302400 19880 302405
rect 19680 302355 19880 302360
rect 19680 302325 19685 302355
rect 19715 302325 19845 302355
rect 19875 302325 19880 302355
rect 19680 302320 19880 302325
rect 19680 302275 19880 302280
rect 19680 302245 19685 302275
rect 19715 302245 19845 302275
rect 19875 302245 19880 302275
rect 19680 302240 19880 302245
rect 19680 302195 19880 302200
rect 19680 302165 19685 302195
rect 19715 302165 19845 302195
rect 19875 302165 19880 302195
rect 19680 302160 19880 302165
rect 19680 302115 19880 302120
rect 19680 302085 19685 302115
rect 19715 302085 19845 302115
rect 19875 302085 19880 302115
rect 19680 302080 19880 302085
rect 19680 302035 19880 302040
rect 19680 302005 19685 302035
rect 19715 302005 19845 302035
rect 19875 302005 19880 302035
rect 19680 302000 19880 302005
rect 19680 301955 19880 301960
rect 19680 301925 19685 301955
rect 19715 301925 19845 301955
rect 19875 301925 19880 301955
rect 19680 301920 19880 301925
rect 19680 301875 19880 301880
rect 19680 301845 19685 301875
rect 19715 301845 19845 301875
rect 19875 301845 19880 301875
rect 19680 301840 19880 301845
rect 19680 301795 19880 301800
rect 19680 301765 19685 301795
rect 19715 301765 19845 301795
rect 19875 301765 19880 301795
rect 19680 301760 19880 301765
rect 19680 301715 19880 301720
rect 19680 301685 19685 301715
rect 19715 301685 19845 301715
rect 19875 301685 19880 301715
rect 19680 301680 19880 301685
rect 19680 301635 19880 301640
rect 19680 301605 19685 301635
rect 19715 301605 19845 301635
rect 19875 301605 19880 301635
rect 19680 301600 19880 301605
rect 19680 301555 19880 301560
rect 19680 301525 19685 301555
rect 19715 301525 19845 301555
rect 19875 301525 19880 301555
rect 19680 301520 19880 301525
rect 19680 301475 19880 301480
rect 19680 301445 19685 301475
rect 19715 301445 19845 301475
rect 19875 301445 19880 301475
rect 19680 301440 19880 301445
rect 19680 301395 19880 301400
rect 19680 301365 19685 301395
rect 19715 301365 19845 301395
rect 19875 301365 19880 301395
rect 19680 301360 19880 301365
rect 19680 301315 19880 301320
rect 19680 301285 19685 301315
rect 19715 301285 19845 301315
rect 19875 301285 19880 301315
rect 19680 301280 19880 301285
rect 19680 301235 19880 301240
rect 19680 301205 19685 301235
rect 19715 301205 19845 301235
rect 19875 301205 19880 301235
rect 19680 301200 19880 301205
rect 19680 301155 19880 301160
rect 19680 301125 19685 301155
rect 19715 301125 19845 301155
rect 19875 301125 19880 301155
rect 19680 301120 19880 301125
rect 19680 301075 19880 301080
rect 19680 301045 19685 301075
rect 19715 301045 19845 301075
rect 19875 301045 19880 301075
rect 19680 301040 19880 301045
rect 19680 300995 19880 301000
rect 19680 300965 19685 300995
rect 19715 300965 19845 300995
rect 19875 300965 19880 300995
rect 19680 300960 19880 300965
rect 19680 300915 19880 300920
rect 19680 300885 19685 300915
rect 19715 300885 19845 300915
rect 19875 300885 19880 300915
rect 19680 300880 19880 300885
rect 19680 300835 19880 300840
rect 19680 300805 19685 300835
rect 19715 300805 19845 300835
rect 19875 300805 19880 300835
rect 19680 300800 19880 300805
rect 19680 300755 19880 300760
rect 19680 300725 19685 300755
rect 19715 300725 19845 300755
rect 19875 300725 19880 300755
rect 19680 300720 19880 300725
rect 19680 300675 19880 300680
rect 19680 300645 19685 300675
rect 19715 300645 19845 300675
rect 19875 300645 19880 300675
rect 19680 300640 19880 300645
rect 19680 300595 19880 300600
rect 19680 300565 19685 300595
rect 19715 300565 19845 300595
rect 19875 300565 19880 300595
rect 19680 300560 19880 300565
rect 19680 300515 19880 300520
rect 19680 300485 19685 300515
rect 19715 300485 19845 300515
rect 19875 300485 19880 300515
rect 19680 300480 19880 300485
rect 19680 300435 19880 300440
rect 19680 300405 19685 300435
rect 19715 300405 19845 300435
rect 19875 300405 19880 300435
rect 19680 300400 19880 300405
rect 19680 300355 19880 300360
rect 19680 300325 19685 300355
rect 19715 300325 19845 300355
rect 19875 300325 19880 300355
rect 19680 300320 19880 300325
rect 19680 300275 19880 300280
rect 19680 300245 19685 300275
rect 19715 300245 19845 300275
rect 19875 300245 19880 300275
rect 19680 300240 19880 300245
rect 19680 300195 19880 300200
rect 19680 300165 19685 300195
rect 19715 300165 19845 300195
rect 19875 300165 19880 300195
rect 19680 300160 19880 300165
rect 19680 300115 19880 300120
rect 19680 300085 19685 300115
rect 19715 300085 19845 300115
rect 19875 300085 19880 300115
rect 19680 300080 19880 300085
rect 19680 300035 19880 300040
rect 19680 300005 19685 300035
rect 19715 300005 19845 300035
rect 19875 300005 19880 300035
rect 19680 300000 19880 300005
rect 19680 299955 19880 299960
rect 19680 299925 19685 299955
rect 19715 299925 19845 299955
rect 19875 299925 19880 299955
rect 19680 299920 19880 299925
rect 19680 299875 19880 299880
rect 19680 299845 19685 299875
rect 19715 299845 19845 299875
rect 19875 299845 19880 299875
rect 19680 299840 19880 299845
rect 19680 299795 19880 299800
rect 19680 299765 19685 299795
rect 19715 299765 19845 299795
rect 19875 299765 19880 299795
rect 19680 299760 19880 299765
rect 19680 299715 19880 299720
rect 19680 299685 19685 299715
rect 19715 299685 19845 299715
rect 19875 299685 19880 299715
rect 19680 299680 19880 299685
rect 19680 299635 19880 299640
rect 19680 299605 19685 299635
rect 19715 299605 19845 299635
rect 19875 299605 19880 299635
rect 19680 299600 19880 299605
rect 19680 299555 19880 299560
rect 19680 299525 19685 299555
rect 19715 299525 19845 299555
rect 19875 299525 19880 299555
rect 19680 299520 19880 299525
rect 19680 299475 19880 299480
rect 19680 299445 19685 299475
rect 19715 299445 19845 299475
rect 19875 299445 19880 299475
rect 19680 299440 19880 299445
rect 19680 299395 19880 299400
rect 19680 299365 19685 299395
rect 19715 299365 19845 299395
rect 19875 299365 19880 299395
rect 19680 299360 19880 299365
rect 19680 299315 19880 299320
rect 19680 299285 19685 299315
rect 19715 299285 19845 299315
rect 19875 299285 19880 299315
rect 19680 299280 19880 299285
rect 19680 299235 19880 299240
rect 19680 299205 19685 299235
rect 19715 299205 19845 299235
rect 19875 299205 19880 299235
rect 19680 299200 19880 299205
rect 19680 299155 19880 299160
rect 19680 299125 19685 299155
rect 19715 299125 19845 299155
rect 19875 299125 19880 299155
rect 19680 299120 19880 299125
rect 19680 299075 19880 299080
rect 19680 299045 19685 299075
rect 19715 299045 19845 299075
rect 19875 299045 19880 299075
rect 19680 299040 19880 299045
rect 19680 298995 19880 299000
rect 19680 298965 19685 298995
rect 19715 298965 19845 298995
rect 19875 298965 19880 298995
rect 19680 298960 19880 298965
rect 19680 298915 19880 298920
rect 19680 298885 19685 298915
rect 19715 298885 19845 298915
rect 19875 298885 19880 298915
rect 19680 298880 19880 298885
rect 19680 298835 19880 298840
rect 19680 298805 19685 298835
rect 19715 298805 19845 298835
rect 19875 298805 19880 298835
rect 19680 298800 19880 298805
rect 19680 298755 19880 298760
rect 19680 298725 19685 298755
rect 19715 298725 19845 298755
rect 19875 298725 19880 298755
rect 19680 298720 19880 298725
rect 19680 298675 19880 298680
rect 19680 298645 19685 298675
rect 19715 298645 19845 298675
rect 19875 298645 19880 298675
rect 19680 298640 19880 298645
rect 19680 298595 19880 298600
rect 19680 298565 19685 298595
rect 19715 298565 19845 298595
rect 19875 298565 19880 298595
rect 19680 298560 19880 298565
rect 19680 298515 19880 298520
rect 19680 298485 19685 298515
rect 19715 298485 19845 298515
rect 19875 298485 19880 298515
rect 19680 298480 19880 298485
rect 19680 298435 19880 298440
rect 19680 298405 19685 298435
rect 19715 298405 19845 298435
rect 19875 298405 19880 298435
rect 19680 298400 19880 298405
rect 19680 298355 19880 298360
rect 19680 298325 19685 298355
rect 19715 298325 19845 298355
rect 19875 298325 19880 298355
rect 19680 298320 19880 298325
rect 19680 298275 19880 298280
rect 19680 298245 19685 298275
rect 19715 298245 19845 298275
rect 19875 298245 19880 298275
rect 19680 298240 19880 298245
rect 19680 298195 19880 298200
rect 19680 298165 19685 298195
rect 19715 298165 19845 298195
rect 19875 298165 19880 298195
rect 19680 298160 19880 298165
rect 19680 298115 19880 298120
rect 19680 298085 19685 298115
rect 19715 298085 19845 298115
rect 19875 298085 19880 298115
rect 19680 298080 19880 298085
rect 19680 298035 19880 298040
rect 19680 298005 19685 298035
rect 19715 298005 19845 298035
rect 19875 298005 19880 298035
rect 19680 298000 19880 298005
rect 19680 297955 19880 297960
rect 19680 297925 19685 297955
rect 19715 297925 19845 297955
rect 19875 297925 19880 297955
rect 19680 297920 19880 297925
rect 19680 297875 19880 297880
rect 19680 297845 19685 297875
rect 19715 297845 19845 297875
rect 19875 297845 19880 297875
rect 19680 297840 19880 297845
rect 19680 297795 19880 297800
rect 19680 297765 19685 297795
rect 19715 297765 19845 297795
rect 19875 297765 19880 297795
rect 19680 297760 19880 297765
rect 19680 297715 19880 297720
rect 19680 297685 19685 297715
rect 19715 297685 19845 297715
rect 19875 297685 19880 297715
rect 19680 297680 19880 297685
rect 19680 297635 19880 297640
rect 19680 297605 19685 297635
rect 19715 297605 19845 297635
rect 19875 297605 19880 297635
rect 19680 297600 19880 297605
rect 19680 297555 19880 297560
rect 19680 297525 19685 297555
rect 19715 297525 19845 297555
rect 19875 297525 19880 297555
rect 19680 297520 19880 297525
rect 19680 297475 19880 297480
rect 19680 297445 19685 297475
rect 19715 297445 19845 297475
rect 19875 297445 19880 297475
rect 19680 297440 19880 297445
rect 19680 297395 19880 297400
rect 19680 297365 19685 297395
rect 19715 297365 19845 297395
rect 19875 297365 19880 297395
rect 19680 297360 19880 297365
rect 19680 297315 19880 297320
rect 19680 297285 19685 297315
rect 19715 297285 19845 297315
rect 19875 297285 19880 297315
rect 19680 297280 19880 297285
rect 19680 297235 19880 297240
rect 19680 297205 19685 297235
rect 19715 297205 19845 297235
rect 19875 297205 19880 297235
rect 19680 297200 19880 297205
rect 19680 297155 19880 297160
rect 19680 297125 19685 297155
rect 19715 297125 19845 297155
rect 19875 297125 19880 297155
rect 19680 297120 19880 297125
rect 19680 297075 19880 297080
rect 19680 297045 19685 297075
rect 19715 297045 19845 297075
rect 19875 297045 19880 297075
rect 19680 297040 19880 297045
rect 19680 296995 19880 297000
rect 19680 296965 19685 296995
rect 19715 296965 19845 296995
rect 19875 296965 19880 296995
rect 19680 296960 19880 296965
rect 19680 296915 19880 296920
rect 19680 296885 19685 296915
rect 19715 296885 19845 296915
rect 19875 296885 19880 296915
rect 19680 296880 19880 296885
rect 19680 296835 19880 296840
rect 19680 296805 19685 296835
rect 19715 296805 19845 296835
rect 19875 296805 19880 296835
rect 19680 296800 19880 296805
rect 19680 296755 19880 296760
rect 19680 296725 19685 296755
rect 19715 296725 19845 296755
rect 19875 296725 19880 296755
rect 19680 296720 19880 296725
rect 19680 296675 19880 296680
rect 19680 296645 19685 296675
rect 19715 296645 19845 296675
rect 19875 296645 19880 296675
rect 19680 296640 19880 296645
rect 19680 296595 19880 296600
rect 19680 296565 19685 296595
rect 19715 296565 19845 296595
rect 19875 296565 19880 296595
rect 19680 296560 19880 296565
rect 19680 296515 19880 296520
rect 19680 296485 19685 296515
rect 19715 296485 19845 296515
rect 19875 296485 19880 296515
rect 19680 296480 19880 296485
rect 19680 296435 19880 296440
rect 19680 296405 19685 296435
rect 19715 296405 19845 296435
rect 19875 296405 19880 296435
rect 19680 296400 19880 296405
rect 19680 296355 19880 296360
rect 19680 296325 19685 296355
rect 19715 296325 19845 296355
rect 19875 296325 19880 296355
rect 19680 296320 19880 296325
rect 19680 296275 19880 296280
rect 19680 296245 19685 296275
rect 19715 296245 19845 296275
rect 19875 296245 19880 296275
rect 19680 296240 19880 296245
rect 19680 296195 19880 296200
rect 19680 296165 19685 296195
rect 19715 296165 19845 296195
rect 19875 296165 19880 296195
rect 19680 296160 19880 296165
rect 19680 296115 19880 296120
rect 19680 296085 19685 296115
rect 19715 296085 19845 296115
rect 19875 296085 19880 296115
rect 19680 296080 19880 296085
rect 19680 296035 19880 296040
rect 19680 296005 19685 296035
rect 19715 296005 19845 296035
rect 19875 296005 19880 296035
rect 19680 296000 19880 296005
rect 19680 295955 19880 295960
rect 19680 295925 19685 295955
rect 19715 295925 19845 295955
rect 19875 295925 19880 295955
rect 19680 295920 19880 295925
rect 19680 295875 19880 295880
rect 19680 295845 19685 295875
rect 19715 295845 19845 295875
rect 19875 295845 19880 295875
rect 19680 295840 19880 295845
rect 19680 295795 19880 295800
rect 19680 295765 19685 295795
rect 19715 295765 19845 295795
rect 19875 295765 19880 295795
rect 19680 295760 19880 295765
rect 19680 295715 19880 295720
rect 19680 295685 19685 295715
rect 19715 295685 19845 295715
rect 19875 295685 19880 295715
rect 19680 295680 19880 295685
rect 19680 295635 19880 295640
rect 19680 295605 19685 295635
rect 19715 295605 19845 295635
rect 19875 295605 19880 295635
rect 19680 295600 19880 295605
rect 19680 295555 19880 295560
rect 19680 295525 19685 295555
rect 19715 295525 19845 295555
rect 19875 295525 19880 295555
rect 19680 295520 19880 295525
rect 19680 295475 19880 295480
rect 19680 295445 19685 295475
rect 19715 295445 19845 295475
rect 19875 295445 19880 295475
rect 19680 295440 19880 295445
rect 19680 295395 19880 295400
rect 19680 295365 19685 295395
rect 19715 295365 19845 295395
rect 19875 295365 19880 295395
rect 19680 295360 19880 295365
rect 19680 295315 19880 295320
rect 19680 295285 19685 295315
rect 19715 295285 19845 295315
rect 19875 295285 19880 295315
rect 19680 295280 19880 295285
rect 19680 295235 19880 295240
rect 19680 295205 19685 295235
rect 19715 295205 19845 295235
rect 19875 295205 19880 295235
rect 19680 295200 19880 295205
rect 19680 295155 19880 295160
rect 19680 295125 19685 295155
rect 19715 295125 19845 295155
rect 19875 295125 19880 295155
rect 19680 295120 19880 295125
rect 19680 295075 19880 295080
rect 19680 295045 19685 295075
rect 19715 295045 19845 295075
rect 19875 295045 19880 295075
rect 19680 295040 19880 295045
rect 19680 294995 19880 295000
rect 19680 294965 19685 294995
rect 19715 294965 19845 294995
rect 19875 294965 19880 294995
rect 19680 294960 19880 294965
rect 19680 294915 19880 294920
rect 19680 294885 19685 294915
rect 19715 294885 19845 294915
rect 19875 294885 19880 294915
rect 19680 294880 19880 294885
rect 19680 294835 19880 294840
rect 19680 294805 19685 294835
rect 19715 294805 19845 294835
rect 19875 294805 19880 294835
rect 19680 294800 19880 294805
rect 19680 294755 19880 294760
rect 19680 294725 19685 294755
rect 19715 294725 19845 294755
rect 19875 294725 19880 294755
rect 19680 294720 19880 294725
rect 19680 294675 19880 294680
rect 19680 294645 19685 294675
rect 19715 294645 19845 294675
rect 19875 294645 19880 294675
rect 19680 294640 19880 294645
rect 19680 294595 19880 294600
rect 19680 294565 19685 294595
rect 19715 294565 19845 294595
rect 19875 294565 19880 294595
rect 19680 294560 19880 294565
rect 19680 294515 19880 294520
rect 19680 294485 19685 294515
rect 19715 294485 19845 294515
rect 19875 294485 19880 294515
rect 19680 294480 19880 294485
rect 19680 294435 19880 294440
rect 19680 294405 19685 294435
rect 19715 294405 19845 294435
rect 19875 294405 19880 294435
rect 19680 294400 19880 294405
rect 19680 294355 19880 294360
rect 19680 294325 19685 294355
rect 19715 294325 19845 294355
rect 19875 294325 19880 294355
rect 19680 294320 19880 294325
rect 19680 294275 19880 294280
rect 19680 294245 19685 294275
rect 19715 294245 19845 294275
rect 19875 294245 19880 294275
rect 19680 294240 19880 294245
rect 19680 294195 19880 294200
rect 19680 294165 19685 294195
rect 19715 294165 19845 294195
rect 19875 294165 19880 294195
rect 19680 294160 19880 294165
rect 19680 294115 19880 294120
rect 19680 294085 19685 294115
rect 19715 294085 19845 294115
rect 19875 294085 19880 294115
rect 19680 294080 19880 294085
rect 19680 294035 19880 294040
rect 19680 294005 19685 294035
rect 19715 294005 19845 294035
rect 19875 294005 19880 294035
rect 19680 294000 19880 294005
rect 19680 293955 19880 293960
rect 19680 293925 19685 293955
rect 19715 293925 19845 293955
rect 19875 293925 19880 293955
rect 19680 293920 19880 293925
rect 19680 293875 19880 293880
rect 19680 293845 19685 293875
rect 19715 293845 19845 293875
rect 19875 293845 19880 293875
rect 19680 293840 19880 293845
rect 19680 293795 19880 293800
rect 19680 293765 19685 293795
rect 19715 293765 19845 293795
rect 19875 293765 19880 293795
rect 19680 293760 19880 293765
rect 19680 293715 19880 293720
rect 19680 293685 19685 293715
rect 19715 293685 19845 293715
rect 19875 293685 19880 293715
rect 19680 293680 19880 293685
rect 19680 293635 19880 293640
rect 19680 293605 19685 293635
rect 19715 293605 19845 293635
rect 19875 293605 19880 293635
rect 19680 293600 19880 293605
rect 19680 293555 19880 293560
rect 19680 293525 19685 293555
rect 19715 293525 19845 293555
rect 19875 293525 19880 293555
rect 19680 293520 19880 293525
rect 19680 293475 19880 293480
rect 19680 293445 19685 293475
rect 19715 293445 19845 293475
rect 19875 293445 19880 293475
rect 19680 293440 19880 293445
rect 19680 293395 19880 293400
rect 19680 293365 19685 293395
rect 19715 293365 19845 293395
rect 19875 293365 19880 293395
rect 19680 293360 19880 293365
rect 19680 293315 19880 293320
rect 19680 293285 19685 293315
rect 19715 293285 19845 293315
rect 19875 293285 19880 293315
rect 19680 293280 19880 293285
rect 19680 293235 19880 293240
rect 19680 293205 19685 293235
rect 19715 293205 19845 293235
rect 19875 293205 19880 293235
rect 19680 293200 19880 293205
rect 19680 293155 19880 293160
rect 19680 293125 19685 293155
rect 19715 293125 19845 293155
rect 19875 293125 19880 293155
rect 19680 293120 19880 293125
rect 19680 293075 19880 293080
rect 19680 293045 19685 293075
rect 19715 293045 19845 293075
rect 19875 293045 19880 293075
rect 19680 293040 19880 293045
rect 19680 292995 19880 293000
rect 19680 292965 19685 292995
rect 19715 292965 19845 292995
rect 19875 292965 19880 292995
rect 19680 292960 19880 292965
rect 19680 292915 19880 292920
rect 19680 292885 19685 292915
rect 19715 292885 19845 292915
rect 19875 292885 19880 292915
rect 19680 292880 19880 292885
rect 19680 292835 19880 292840
rect 19680 292805 19685 292835
rect 19715 292805 19845 292835
rect 19875 292805 19880 292835
rect 19680 292800 19880 292805
rect 19680 292755 19880 292760
rect 19680 292725 19685 292755
rect 19715 292725 19845 292755
rect 19875 292725 19880 292755
rect 19680 292720 19880 292725
rect 19680 292675 19880 292680
rect 19680 292645 19685 292675
rect 19715 292645 19845 292675
rect 19875 292645 19880 292675
rect 19680 292640 19880 292645
rect 19680 292595 19880 292600
rect 19680 292565 19685 292595
rect 19715 292565 19845 292595
rect 19875 292565 19880 292595
rect 19680 292560 19880 292565
rect 19680 292515 19880 292520
rect 19680 292485 19685 292515
rect 19715 292485 19845 292515
rect 19875 292485 19880 292515
rect 19680 292480 19880 292485
rect 19680 292435 19880 292440
rect 19680 292405 19685 292435
rect 19715 292405 19845 292435
rect 19875 292405 19880 292435
rect 19680 292400 19880 292405
rect 19680 292355 19880 292360
rect 19680 292325 19685 292355
rect 19715 292325 19845 292355
rect 19875 292325 19880 292355
rect 19680 292320 19880 292325
rect 19680 292275 19880 292280
rect 19680 292245 19685 292275
rect 19715 292245 19845 292275
rect 19875 292245 19880 292275
rect 19680 292240 19880 292245
rect 19680 292195 19880 292200
rect 19680 292165 19685 292195
rect 19715 292165 19845 292195
rect 19875 292165 19880 292195
rect 19680 292160 19880 292165
rect 19680 292115 19880 292120
rect 19680 292085 19685 292115
rect 19715 292085 19845 292115
rect 19875 292085 19880 292115
rect 19680 292080 19880 292085
rect 19680 292035 19880 292040
rect 19680 292005 19685 292035
rect 19715 292005 19845 292035
rect 19875 292005 19880 292035
rect 19680 292000 19880 292005
rect 19680 291955 19880 291960
rect 19680 291925 19685 291955
rect 19715 291925 19845 291955
rect 19875 291925 19880 291955
rect 19680 291920 19880 291925
rect 19680 291875 19880 291880
rect 19680 291845 19685 291875
rect 19715 291845 19845 291875
rect 19875 291845 19880 291875
rect 19680 291840 19880 291845
rect 19680 291795 19880 291800
rect 19680 291765 19685 291795
rect 19715 291765 19845 291795
rect 19875 291765 19880 291795
rect 19680 291760 19880 291765
rect 19680 291715 19880 291720
rect 19680 291685 19685 291715
rect 19715 291685 19845 291715
rect 19875 291685 19880 291715
rect 19680 291680 19880 291685
rect 19680 291635 19880 291640
rect 19680 291605 19685 291635
rect 19715 291605 19845 291635
rect 19875 291605 19880 291635
rect 19680 291600 19880 291605
rect 19680 291555 19880 291560
rect 19680 291525 19685 291555
rect 19715 291525 19845 291555
rect 19875 291525 19880 291555
rect 19680 291520 19880 291525
rect 19680 291475 19880 291480
rect 19680 291445 19685 291475
rect 19715 291445 19845 291475
rect 19875 291445 19880 291475
rect 19680 291440 19880 291445
rect 19680 291395 19880 291400
rect 19680 291365 19685 291395
rect 19715 291365 19845 291395
rect 19875 291365 19880 291395
rect 19680 291360 19880 291365
rect 19680 291315 19880 291320
rect 19680 291285 19685 291315
rect 19715 291285 19845 291315
rect 19875 291285 19880 291315
rect 19680 291280 19880 291285
rect 19680 291235 19880 291240
rect 19680 291205 19685 291235
rect 19715 291205 19845 291235
rect 19875 291205 19880 291235
rect 19680 291200 19880 291205
rect 19680 291155 19880 291160
rect 19680 291125 19685 291155
rect 19715 291125 19845 291155
rect 19875 291125 19880 291155
rect 19680 291120 19880 291125
rect 19680 291075 19880 291080
rect 19680 291045 19685 291075
rect 19715 291045 19845 291075
rect 19875 291045 19880 291075
rect 19680 291040 19880 291045
rect 19680 290995 19880 291000
rect 19680 290965 19685 290995
rect 19715 290965 19845 290995
rect 19875 290965 19880 290995
rect 19680 290960 19880 290965
rect 19680 290915 19880 290920
rect 19680 290885 19685 290915
rect 19715 290885 19845 290915
rect 19875 290885 19880 290915
rect 19680 290880 19880 290885
rect 19680 290835 19880 290840
rect 19680 290805 19685 290835
rect 19715 290805 19845 290835
rect 19875 290805 19880 290835
rect 19680 290800 19880 290805
rect 19680 290755 19880 290760
rect 19680 290725 19685 290755
rect 19715 290725 19845 290755
rect 19875 290725 19880 290755
rect 19680 290720 19880 290725
rect 19680 290675 19880 290680
rect 19680 290645 19685 290675
rect 19715 290645 19845 290675
rect 19875 290645 19880 290675
rect 19680 290640 19880 290645
rect 19680 290595 19880 290600
rect 19680 290565 19685 290595
rect 19715 290565 19845 290595
rect 19875 290565 19880 290595
rect 19680 290560 19880 290565
rect 19680 290515 19880 290520
rect 19680 290485 19685 290515
rect 19715 290485 19845 290515
rect 19875 290485 19880 290515
rect 19680 290480 19880 290485
rect 19680 290435 19880 290440
rect 19680 290405 19685 290435
rect 19715 290405 19845 290435
rect 19875 290405 19880 290435
rect 19680 290400 19880 290405
rect 19680 290355 19880 290360
rect 19680 290325 19685 290355
rect 19715 290325 19845 290355
rect 19875 290325 19880 290355
rect 19680 290320 19880 290325
rect 19680 290275 19880 290280
rect 19680 290245 19685 290275
rect 19715 290245 19845 290275
rect 19875 290245 19880 290275
rect 19680 290240 19880 290245
rect 19680 290195 19880 290200
rect 19680 290165 19685 290195
rect 19715 290165 19845 290195
rect 19875 290165 19880 290195
rect 19680 290160 19880 290165
rect 19680 290115 19880 290120
rect 19680 290085 19685 290115
rect 19715 290085 19845 290115
rect 19875 290085 19880 290115
rect 19680 290080 19880 290085
rect 19680 290035 19880 290040
rect 19680 290005 19685 290035
rect 19715 290005 19845 290035
rect 19875 290005 19880 290035
rect 19680 290000 19880 290005
rect 19680 289955 19880 289960
rect 19680 289925 19685 289955
rect 19715 289925 19845 289955
rect 19875 289925 19880 289955
rect 19680 289920 19880 289925
rect 19680 289875 19880 289880
rect 19680 289845 19685 289875
rect 19715 289845 19845 289875
rect 19875 289845 19880 289875
rect 19680 289840 19880 289845
rect 19680 289795 19880 289800
rect 19680 289765 19685 289795
rect 19715 289765 19845 289795
rect 19875 289765 19880 289795
rect 19680 289760 19880 289765
rect 19680 289715 19880 289720
rect 19680 289685 19685 289715
rect 19715 289685 19845 289715
rect 19875 289685 19880 289715
rect 19680 289680 19880 289685
rect 19680 289635 19880 289640
rect 19680 289605 19685 289635
rect 19715 289605 19845 289635
rect 19875 289605 19880 289635
rect 19680 289600 19880 289605
rect 19680 289555 19880 289560
rect 19680 289525 19685 289555
rect 19715 289525 19845 289555
rect 19875 289525 19880 289555
rect 19680 289520 19880 289525
rect 19680 289475 19880 289480
rect 19680 289445 19685 289475
rect 19715 289445 19845 289475
rect 19875 289445 19880 289475
rect 19680 289440 19880 289445
rect 19680 289395 19880 289400
rect 19680 289365 19685 289395
rect 19715 289365 19845 289395
rect 19875 289365 19880 289395
rect 19680 289360 19880 289365
rect 19680 289315 19880 289320
rect 19680 289285 19685 289315
rect 19715 289285 19845 289315
rect 19875 289285 19880 289315
rect 19680 289280 19880 289285
rect 19680 289235 19880 289240
rect 19680 289205 19685 289235
rect 19715 289205 19845 289235
rect 19875 289205 19880 289235
rect 19680 289200 19880 289205
rect 19680 289155 19880 289160
rect 19680 289125 19685 289155
rect 19715 289125 19845 289155
rect 19875 289125 19880 289155
rect 19680 289120 19880 289125
rect 19680 289075 19880 289080
rect 19680 289045 19685 289075
rect 19715 289045 19845 289075
rect 19875 289045 19880 289075
rect 19680 289040 19880 289045
rect 19680 288995 19880 289000
rect 19680 288965 19685 288995
rect 19715 288965 19845 288995
rect 19875 288965 19880 288995
rect 19680 288960 19880 288965
rect 19680 288915 19880 288920
rect 19680 288885 19685 288915
rect 19715 288885 19845 288915
rect 19875 288885 19880 288915
rect 19680 288880 19880 288885
rect 19680 288835 19880 288840
rect 19680 288805 19685 288835
rect 19715 288805 19845 288835
rect 19875 288805 19880 288835
rect 19680 288800 19880 288805
rect 19680 288755 19880 288760
rect 19680 288725 19685 288755
rect 19715 288725 19845 288755
rect 19875 288725 19880 288755
rect 19680 288720 19880 288725
rect 19680 288675 19880 288680
rect 19680 288645 19685 288675
rect 19715 288645 19845 288675
rect 19875 288645 19880 288675
rect 19680 288640 19880 288645
rect 19680 288595 19880 288600
rect 19680 288565 19685 288595
rect 19715 288565 19845 288595
rect 19875 288565 19880 288595
rect 19680 288560 19880 288565
rect 19680 288515 19880 288520
rect 19680 288485 19685 288515
rect 19715 288485 19845 288515
rect 19875 288485 19880 288515
rect 19680 288480 19880 288485
rect 19680 288435 19880 288440
rect 19680 288405 19685 288435
rect 19715 288405 19845 288435
rect 19875 288405 19880 288435
rect 19680 288400 19880 288405
rect 19680 288355 19880 288360
rect 19680 288325 19685 288355
rect 19715 288325 19845 288355
rect 19875 288325 19880 288355
rect 19680 288320 19880 288325
rect 19680 288275 19880 288280
rect 19680 288245 19685 288275
rect 19715 288245 19845 288275
rect 19875 288245 19880 288275
rect 19680 288240 19880 288245
rect 19680 288195 19880 288200
rect 19680 288165 19685 288195
rect 19715 288165 19845 288195
rect 19875 288165 19880 288195
rect 19680 288160 19880 288165
rect 19680 288115 19880 288120
rect 19680 288085 19685 288115
rect 19715 288085 19845 288115
rect 19875 288085 19880 288115
rect 19680 288080 19880 288085
rect 19680 288035 19880 288040
rect 19680 288005 19685 288035
rect 19715 288005 19845 288035
rect 19875 288005 19880 288035
rect 19680 288000 19880 288005
rect 19680 287955 19880 287960
rect 19680 287925 19685 287955
rect 19715 287925 19845 287955
rect 19875 287925 19880 287955
rect 19680 287920 19880 287925
rect 19680 287875 19880 287880
rect 19680 287845 19685 287875
rect 19715 287845 19845 287875
rect 19875 287845 19880 287875
rect 19680 287840 19880 287845
rect 19680 287795 19880 287800
rect 19680 287765 19685 287795
rect 19715 287765 19845 287795
rect 19875 287765 19880 287795
rect 19680 287760 19880 287765
rect 19680 287715 19880 287720
rect 19680 287685 19685 287715
rect 19715 287685 19845 287715
rect 19875 287685 19880 287715
rect 19680 287680 19880 287685
rect 19680 287635 19880 287640
rect 19680 287605 19685 287635
rect 19715 287605 19845 287635
rect 19875 287605 19880 287635
rect 19680 287600 19880 287605
rect 19680 287555 19880 287560
rect 19680 287525 19685 287555
rect 19715 287525 19845 287555
rect 19875 287525 19880 287555
rect 19680 287520 19880 287525
rect 19680 287475 19880 287480
rect 19680 287445 19685 287475
rect 19715 287445 19845 287475
rect 19875 287445 19880 287475
rect 19680 287440 19880 287445
rect 19680 287395 19880 287400
rect 19680 287365 19685 287395
rect 19715 287365 19845 287395
rect 19875 287365 19880 287395
rect 19680 287360 19880 287365
rect 19680 287315 19880 287320
rect 19680 287285 19685 287315
rect 19715 287285 19845 287315
rect 19875 287285 19880 287315
rect 19680 287280 19880 287285
rect 19680 287235 19880 287240
rect 19680 287205 19685 287235
rect 19715 287205 19845 287235
rect 19875 287205 19880 287235
rect 19680 287200 19880 287205
rect 19680 287155 19880 287160
rect 19680 287125 19685 287155
rect 19715 287125 19845 287155
rect 19875 287125 19880 287155
rect 19680 287120 19880 287125
rect 19680 287075 19880 287080
rect 19680 287045 19685 287075
rect 19715 287045 19845 287075
rect 19875 287045 19880 287075
rect 19680 287040 19880 287045
rect 19680 286995 19880 287000
rect 19680 286965 19685 286995
rect 19715 286965 19845 286995
rect 19875 286965 19880 286995
rect 19680 286960 19880 286965
rect 19680 286915 19880 286920
rect 19680 286885 19685 286915
rect 19715 286885 19845 286915
rect 19875 286885 19880 286915
rect 19680 286880 19880 286885
rect 19680 286835 19880 286840
rect 19680 286805 19685 286835
rect 19715 286805 19845 286835
rect 19875 286805 19880 286835
rect 19680 286800 19880 286805
rect 19680 286755 19880 286760
rect 19680 286725 19685 286755
rect 19715 286725 19845 286755
rect 19875 286725 19880 286755
rect 19680 286720 19880 286725
rect 19680 286675 19880 286680
rect 19680 286645 19685 286675
rect 19715 286645 19845 286675
rect 19875 286645 19880 286675
rect 19680 286640 19880 286645
rect 19680 286595 19880 286600
rect 19680 286565 19685 286595
rect 19715 286565 19845 286595
rect 19875 286565 19880 286595
rect 19680 286560 19880 286565
rect 19680 286515 19880 286520
rect 19680 286485 19685 286515
rect 19715 286485 19845 286515
rect 19875 286485 19880 286515
rect 19680 286480 19880 286485
rect 19680 286435 19880 286440
rect 19680 286405 19685 286435
rect 19715 286405 19845 286435
rect 19875 286405 19880 286435
rect 19680 286400 19880 286405
rect 19680 286355 19880 286360
rect 19680 286325 19685 286355
rect 19715 286325 19845 286355
rect 19875 286325 19880 286355
rect 19680 286320 19880 286325
rect 19680 286275 19880 286280
rect 19680 286245 19685 286275
rect 19715 286245 19845 286275
rect 19875 286245 19880 286275
rect 19680 286240 19880 286245
rect 19680 286195 19880 286200
rect 19680 286165 19685 286195
rect 19715 286165 19845 286195
rect 19875 286165 19880 286195
rect 19680 286160 19880 286165
rect 19680 286115 19880 286120
rect 19680 286085 19685 286115
rect 19715 286085 19845 286115
rect 19875 286085 19880 286115
rect 19680 286080 19880 286085
rect 19680 286035 19880 286040
rect 19680 286005 19685 286035
rect 19715 286005 19845 286035
rect 19875 286005 19880 286035
rect 19680 286000 19880 286005
rect 19680 285955 19880 285960
rect 19680 285925 19685 285955
rect 19715 285925 19845 285955
rect 19875 285925 19880 285955
rect 19680 285920 19880 285925
rect 19680 285875 19880 285880
rect 19680 285845 19685 285875
rect 19715 285845 19845 285875
rect 19875 285845 19880 285875
rect 19680 285840 19880 285845
rect 19680 285795 19880 285800
rect 19680 285765 19685 285795
rect 19715 285765 19845 285795
rect 19875 285765 19880 285795
rect 19680 285760 19880 285765
rect 19680 285715 19880 285720
rect 19680 285685 19685 285715
rect 19715 285685 19845 285715
rect 19875 285685 19880 285715
rect 19680 285680 19880 285685
rect 19680 285635 19880 285640
rect 19680 285605 19685 285635
rect 19715 285605 19845 285635
rect 19875 285605 19880 285635
rect 19680 285600 19880 285605
rect 19680 285555 19880 285560
rect 19680 285525 19685 285555
rect 19715 285525 19845 285555
rect 19875 285525 19880 285555
rect 19680 285520 19880 285525
rect 19680 285475 19880 285480
rect 19680 285445 19685 285475
rect 19715 285445 19845 285475
rect 19875 285445 19880 285475
rect 19680 285440 19880 285445
rect 19680 285395 19880 285400
rect 19680 285365 19685 285395
rect 19715 285365 19845 285395
rect 19875 285365 19880 285395
rect 19680 285360 19880 285365
rect 19680 285315 19880 285320
rect 19680 285285 19685 285315
rect 19715 285285 19845 285315
rect 19875 285285 19880 285315
rect 19680 285280 19880 285285
rect 19680 285235 19880 285240
rect 19680 285205 19685 285235
rect 19715 285205 19845 285235
rect 19875 285205 19880 285235
rect 19680 285200 19880 285205
rect 19680 285155 19880 285160
rect 19680 285125 19685 285155
rect 19715 285125 19845 285155
rect 19875 285125 19880 285155
rect 19680 285120 19880 285125
rect 19680 285075 19880 285080
rect 19680 285045 19685 285075
rect 19715 285045 19845 285075
rect 19875 285045 19880 285075
rect 19680 285040 19880 285045
rect 19680 284995 19880 285000
rect 19680 284965 19685 284995
rect 19715 284965 19845 284995
rect 19875 284965 19880 284995
rect 19680 284960 19880 284965
rect 19680 284915 19880 284920
rect 19680 284885 19685 284915
rect 19715 284885 19845 284915
rect 19875 284885 19880 284915
rect 19680 284880 19880 284885
rect 19680 284835 19880 284840
rect 19680 284805 19685 284835
rect 19715 284805 19845 284835
rect 19875 284805 19880 284835
rect 19680 284800 19880 284805
rect 19680 284755 19880 284760
rect 19680 284725 19685 284755
rect 19715 284725 19845 284755
rect 19875 284725 19880 284755
rect 19680 284720 19880 284725
rect 19680 284675 19880 284680
rect 19680 284645 19685 284675
rect 19715 284645 19845 284675
rect 19875 284645 19880 284675
rect 19680 284640 19880 284645
rect 19680 284595 19880 284600
rect 19680 284565 19685 284595
rect 19715 284565 19845 284595
rect 19875 284565 19880 284595
rect 19680 284560 19880 284565
rect 19680 284515 19880 284520
rect 19680 284485 19685 284515
rect 19715 284485 19845 284515
rect 19875 284485 19880 284515
rect 19680 284480 19880 284485
rect 19680 284435 19880 284440
rect 19680 284405 19685 284435
rect 19715 284405 19845 284435
rect 19875 284405 19880 284435
rect 19680 284400 19880 284405
rect 19680 284355 19880 284360
rect 19680 284325 19685 284355
rect 19715 284325 19845 284355
rect 19875 284325 19880 284355
rect 19680 284320 19880 284325
rect 19680 284275 19880 284280
rect 19680 284245 19685 284275
rect 19715 284245 19845 284275
rect 19875 284245 19880 284275
rect 19680 284240 19880 284245
rect 19680 284195 19880 284200
rect 19680 284165 19685 284195
rect 19715 284165 19845 284195
rect 19875 284165 19880 284195
rect 19680 284160 19880 284165
rect 19680 284115 19880 284120
rect 19680 284085 19685 284115
rect 19715 284085 19845 284115
rect 19875 284085 19880 284115
rect 19680 284080 19880 284085
rect 19680 284035 19880 284040
rect 19680 284005 19685 284035
rect 19715 284005 19845 284035
rect 19875 284005 19880 284035
rect 19680 284000 19880 284005
rect 19680 283955 19880 283960
rect 19680 283925 19685 283955
rect 19715 283925 19845 283955
rect 19875 283925 19880 283955
rect 19680 283920 19880 283925
rect 19680 283875 19880 283880
rect 19680 283845 19685 283875
rect 19715 283845 19845 283875
rect 19875 283845 19880 283875
rect 19680 283840 19880 283845
rect 19680 283795 19880 283800
rect 19680 283765 19685 283795
rect 19715 283765 19845 283795
rect 19875 283765 19880 283795
rect 19680 283760 19880 283765
rect 19680 283715 19880 283720
rect 19680 283685 19685 283715
rect 19715 283685 19845 283715
rect 19875 283685 19880 283715
rect 19680 283680 19880 283685
rect 19680 283635 19880 283640
rect 19680 283605 19685 283635
rect 19715 283605 19845 283635
rect 19875 283605 19880 283635
rect 19680 283600 19880 283605
rect 19680 283555 19880 283560
rect 19680 283525 19685 283555
rect 19715 283525 19845 283555
rect 19875 283525 19880 283555
rect 19680 283520 19880 283525
rect 19680 283475 19880 283480
rect 19680 283445 19685 283475
rect 19715 283445 19845 283475
rect 19875 283445 19880 283475
rect 19680 283440 19880 283445
rect 19680 283395 19880 283400
rect 19680 283365 19685 283395
rect 19715 283365 19845 283395
rect 19875 283365 19880 283395
rect 19680 283360 19880 283365
rect 19680 283315 19880 283320
rect 19680 283285 19685 283315
rect 19715 283285 19845 283315
rect 19875 283285 19880 283315
rect 19680 283280 19880 283285
rect 19680 283235 19880 283240
rect 19680 283205 19685 283235
rect 19715 283205 19845 283235
rect 19875 283205 19880 283235
rect 19680 283200 19880 283205
rect 19680 283155 19880 283160
rect 19680 283125 19685 283155
rect 19715 283125 19845 283155
rect 19875 283125 19880 283155
rect 19680 283120 19880 283125
rect 19680 283075 19880 283080
rect 19680 283045 19685 283075
rect 19715 283045 19845 283075
rect 19875 283045 19880 283075
rect 19680 283040 19880 283045
rect 19680 282995 19880 283000
rect 19680 282965 19685 282995
rect 19715 282965 19845 282995
rect 19875 282965 19880 282995
rect 19680 282960 19880 282965
rect 19680 282915 19880 282920
rect 19680 282885 19685 282915
rect 19715 282885 19845 282915
rect 19875 282885 19880 282915
rect 19680 282880 19880 282885
rect 19680 282835 19880 282840
rect 19680 282805 19685 282835
rect 19715 282805 19845 282835
rect 19875 282805 19880 282835
rect 19680 282800 19880 282805
rect 19680 282755 19880 282760
rect 19680 282725 19685 282755
rect 19715 282725 19845 282755
rect 19875 282725 19880 282755
rect 19680 282720 19880 282725
rect 19680 282675 19880 282680
rect 19680 282645 19685 282675
rect 19715 282645 19845 282675
rect 19875 282645 19880 282675
rect 19680 282640 19880 282645
rect 19680 282595 19880 282600
rect 19680 282565 19685 282595
rect 19715 282565 19845 282595
rect 19875 282565 19880 282595
rect 19680 282560 19880 282565
rect 19680 282515 19880 282520
rect 19680 282485 19685 282515
rect 19715 282485 19845 282515
rect 19875 282485 19880 282515
rect 19680 282480 19880 282485
rect 19680 282435 19880 282440
rect 19680 282405 19685 282435
rect 19715 282405 19845 282435
rect 19875 282405 19880 282435
rect 19680 282400 19880 282405
rect 19680 282355 19880 282360
rect 19680 282325 19685 282355
rect 19715 282325 19845 282355
rect 19875 282325 19880 282355
rect 19680 282320 19880 282325
rect 19680 282275 19880 282280
rect 19680 282245 19685 282275
rect 19715 282245 19845 282275
rect 19875 282245 19880 282275
rect 19680 282240 19880 282245
rect 19680 282195 19880 282200
rect 19680 282165 19685 282195
rect 19715 282165 19845 282195
rect 19875 282165 19880 282195
rect 19680 282160 19880 282165
rect 19680 282115 19880 282120
rect 19680 282085 19685 282115
rect 19715 282085 19845 282115
rect 19875 282085 19880 282115
rect 19680 282080 19880 282085
rect 19680 282035 19880 282040
rect 19680 282005 19685 282035
rect 19715 282005 19845 282035
rect 19875 282005 19880 282035
rect 19680 282000 19880 282005
rect 19680 281955 19880 281960
rect 19680 281925 19685 281955
rect 19715 281925 19845 281955
rect 19875 281925 19880 281955
rect 19680 281920 19880 281925
rect 19680 281875 19880 281880
rect 19680 281845 19685 281875
rect 19715 281845 19845 281875
rect 19875 281845 19880 281875
rect 19680 281840 19880 281845
rect 19680 281795 19880 281800
rect 19680 281765 19685 281795
rect 19715 281765 19845 281795
rect 19875 281765 19880 281795
rect 19680 281760 19880 281765
rect 19680 281715 19880 281720
rect 19680 281685 19685 281715
rect 19715 281685 19845 281715
rect 19875 281685 19880 281715
rect 19680 281680 19880 281685
rect 19680 281635 19880 281640
rect 19680 281605 19685 281635
rect 19715 281605 19845 281635
rect 19875 281605 19880 281635
rect 19680 281600 19880 281605
rect 19680 281555 19880 281560
rect 19680 281525 19685 281555
rect 19715 281525 19845 281555
rect 19875 281525 19880 281555
rect 19680 281520 19880 281525
rect 19680 281475 19880 281480
rect 19680 281445 19685 281475
rect 19715 281445 19845 281475
rect 19875 281445 19880 281475
rect 19680 281440 19880 281445
rect 19680 281395 19880 281400
rect 19680 281365 19685 281395
rect 19715 281365 19845 281395
rect 19875 281365 19880 281395
rect 19680 281360 19880 281365
rect 19680 281315 19880 281320
rect 19680 281285 19685 281315
rect 19715 281285 19845 281315
rect 19875 281285 19880 281315
rect 19680 281280 19880 281285
rect 19680 281235 19880 281240
rect 19680 281205 19685 281235
rect 19715 281205 19845 281235
rect 19875 281205 19880 281235
rect 19680 281200 19880 281205
rect 19680 281155 19880 281160
rect 19680 281125 19685 281155
rect 19715 281125 19845 281155
rect 19875 281125 19880 281155
rect 19680 281120 19880 281125
rect 19680 281075 19880 281080
rect 19680 281045 19685 281075
rect 19715 281045 19845 281075
rect 19875 281045 19880 281075
rect 19680 281040 19880 281045
rect 19680 280995 19880 281000
rect 19680 280965 19685 280995
rect 19715 280965 19845 280995
rect 19875 280965 19880 280995
rect 19680 280960 19880 280965
rect 19680 280915 19880 280920
rect 19680 280885 19685 280915
rect 19715 280885 19845 280915
rect 19875 280885 19880 280915
rect 19680 280880 19880 280885
rect 19680 280835 19880 280840
rect 19680 280805 19685 280835
rect 19715 280805 19845 280835
rect 19875 280805 19880 280835
rect 19680 280800 19880 280805
rect 19680 280755 19880 280760
rect 19680 280725 19685 280755
rect 19715 280725 19845 280755
rect 19875 280725 19880 280755
rect 19680 280720 19880 280725
rect 19680 280675 19880 280680
rect 19680 280645 19685 280675
rect 19715 280645 19845 280675
rect 19875 280645 19880 280675
rect 19680 280640 19880 280645
rect 19680 280595 19880 280600
rect 19680 280565 19685 280595
rect 19715 280565 19845 280595
rect 19875 280565 19880 280595
rect 19680 280560 19880 280565
rect 19680 280515 19880 280520
rect 19680 280485 19685 280515
rect 19715 280485 19845 280515
rect 19875 280485 19880 280515
rect 19680 280480 19880 280485
rect 19680 280435 19880 280440
rect 19680 280405 19685 280435
rect 19715 280405 19845 280435
rect 19875 280405 19880 280435
rect 19680 280400 19880 280405
rect 19680 280355 19880 280360
rect 19680 280325 19685 280355
rect 19715 280325 19845 280355
rect 19875 280325 19880 280355
rect 19680 280320 19880 280325
rect 19680 280275 19880 280280
rect 19680 280245 19685 280275
rect 19715 280245 19845 280275
rect 19875 280245 19880 280275
rect 19680 280240 19880 280245
rect 19680 280195 19880 280200
rect 19680 280165 19685 280195
rect 19715 280165 19845 280195
rect 19875 280165 19880 280195
rect 19680 280160 19880 280165
rect 19680 280115 19880 280120
rect 19680 280085 19685 280115
rect 19715 280085 19845 280115
rect 19875 280085 19880 280115
rect 19680 280080 19880 280085
rect 19680 280035 19880 280040
rect 19680 280005 19685 280035
rect 19715 280005 19845 280035
rect 19875 280005 19880 280035
rect 19680 280000 19880 280005
rect 19680 279955 19880 279960
rect 19680 279925 19685 279955
rect 19715 279925 19845 279955
rect 19875 279925 19880 279955
rect 19680 279920 19880 279925
rect 19680 279875 19880 279880
rect 19680 279845 19685 279875
rect 19715 279845 19845 279875
rect 19875 279845 19880 279875
rect 19680 279840 19880 279845
rect 19680 279795 19880 279800
rect 19680 279765 19685 279795
rect 19715 279765 19845 279795
rect 19875 279765 19880 279795
rect 19680 279760 19880 279765
rect 19680 279715 19880 279720
rect 19680 279685 19685 279715
rect 19715 279685 19845 279715
rect 19875 279685 19880 279715
rect 19680 279680 19880 279685
rect 19680 279635 19880 279640
rect 19680 279605 19685 279635
rect 19715 279605 19845 279635
rect 19875 279605 19880 279635
rect 19680 279600 19880 279605
rect 19680 279555 19880 279560
rect 19680 279525 19685 279555
rect 19715 279525 19845 279555
rect 19875 279525 19880 279555
rect 19680 279520 19880 279525
rect 19680 279475 19880 279480
rect 19680 279445 19685 279475
rect 19715 279445 19845 279475
rect 19875 279445 19880 279475
rect 19680 279440 19880 279445
rect 19680 279395 19880 279400
rect 19680 279365 19685 279395
rect 19715 279365 19845 279395
rect 19875 279365 19880 279395
rect 19680 279360 19880 279365
rect 19680 279315 19880 279320
rect 19680 279285 19685 279315
rect 19715 279285 19845 279315
rect 19875 279285 19880 279315
rect 19680 279280 19880 279285
rect 19680 279235 19880 279240
rect 19680 279205 19685 279235
rect 19715 279205 19845 279235
rect 19875 279205 19880 279235
rect 19680 279200 19880 279205
rect 19680 279155 19880 279160
rect 19680 279125 19685 279155
rect 19715 279125 19845 279155
rect 19875 279125 19880 279155
rect 19680 279120 19880 279125
rect 19680 279075 19880 279080
rect 19680 279045 19685 279075
rect 19715 279045 19845 279075
rect 19875 279045 19880 279075
rect 19680 279040 19880 279045
rect 19680 278995 19880 279000
rect 19680 278965 19685 278995
rect 19715 278965 19845 278995
rect 19875 278965 19880 278995
rect 19680 278960 19880 278965
rect 19680 278915 19880 278920
rect 19680 278885 19685 278915
rect 19715 278885 19845 278915
rect 19875 278885 19880 278915
rect 19680 278880 19880 278885
rect 19680 278835 19880 278840
rect 19680 278805 19685 278835
rect 19715 278805 19845 278835
rect 19875 278805 19880 278835
rect 19680 278800 19880 278805
rect 19680 278755 19880 278760
rect 19680 278725 19685 278755
rect 19715 278725 19845 278755
rect 19875 278725 19880 278755
rect 19680 278720 19880 278725
rect 17040 278675 17800 278680
rect 17040 278645 17045 278675
rect 17075 278645 17205 278675
rect 17235 278645 17285 278675
rect 17315 278645 17365 278675
rect 17395 278645 17445 278675
rect 17475 278645 17525 278675
rect 17555 278645 17605 278675
rect 17635 278645 17685 278675
rect 17715 278645 17765 278675
rect 17795 278645 17800 278675
rect 17040 278640 17800 278645
rect 19520 278675 19880 278680
rect 19520 278645 19525 278675
rect 19555 278645 19605 278675
rect 19635 278645 19685 278675
rect 19715 278645 19845 278675
rect 19875 278645 19880 278675
rect 19520 278640 19880 278645
rect 17040 278560 17080 278600
rect 17120 278595 17800 278600
rect 17120 278565 17125 278595
rect 17155 278565 17800 278595
rect 17120 278560 17800 278565
rect 19520 278595 19800 278600
rect 19520 278565 19765 278595
rect 19795 278565 19800 278595
rect 19520 278560 19800 278565
rect 17040 278515 17800 278520
rect 17040 278485 17045 278515
rect 17075 278485 17205 278515
rect 17235 278485 17285 278515
rect 17315 278485 17365 278515
rect 17395 278485 17445 278515
rect 17475 278485 17525 278515
rect 17555 278485 17605 278515
rect 17635 278485 17685 278515
rect 17715 278485 17765 278515
rect 17795 278485 17800 278515
rect 17040 278480 17800 278485
rect 19520 278515 19880 278520
rect 19520 278485 19525 278515
rect 19555 278485 19605 278515
rect 19635 278485 19685 278515
rect 19715 278485 19845 278515
rect 19875 278485 19880 278515
rect 19520 278480 19880 278485
rect 17040 278435 17240 278440
rect 17040 278405 17045 278435
rect 17075 278405 17205 278435
rect 17235 278405 17240 278435
rect 17040 278400 17240 278405
rect 17040 278355 17240 278360
rect 17040 278325 17045 278355
rect 17075 278325 17205 278355
rect 17235 278325 17240 278355
rect 17040 278320 17240 278325
rect 17040 278275 17240 278280
rect 17040 278245 17045 278275
rect 17075 278245 17205 278275
rect 17235 278245 17240 278275
rect 17040 278240 17240 278245
rect 17040 278195 17240 278200
rect 17040 278165 17045 278195
rect 17075 278165 17205 278195
rect 17235 278165 17240 278195
rect 17040 278160 17240 278165
rect 17040 278115 17240 278120
rect 17040 278085 17045 278115
rect 17075 278085 17205 278115
rect 17235 278085 17240 278115
rect 17040 278080 17240 278085
rect 17040 278035 17240 278040
rect 17040 278005 17045 278035
rect 17075 278005 17205 278035
rect 17235 278005 17240 278035
rect 17040 278000 17240 278005
rect 17040 277955 17240 277960
rect 17040 277925 17045 277955
rect 17075 277925 17205 277955
rect 17235 277925 17240 277955
rect 17040 277920 17240 277925
rect 17040 277875 17240 277880
rect 17040 277845 17045 277875
rect 17075 277845 17205 277875
rect 17235 277845 17240 277875
rect 17040 277840 17240 277845
rect 28400 275355 28760 275360
rect 28400 275325 28405 275355
rect 28435 275325 28565 275355
rect 28595 275325 28725 275355
rect 28755 275325 28760 275355
rect 28400 275320 28760 275325
rect 28400 275275 28760 275280
rect 28400 275245 28405 275275
rect 28435 275245 28565 275275
rect 28595 275245 28725 275275
rect 28755 275245 28760 275275
rect 28400 275240 28760 275245
rect 1000 275195 28760 275200
rect 1000 275160 13525 275195
rect 1000 275040 1040 275160
rect 1160 275040 13525 275160
rect 1000 275005 13525 275040
rect 13555 275005 13685 275195
rect 13715 275005 13845 275195
rect 13875 275005 14005 275195
rect 14035 275005 14165 275195
rect 14195 275005 14325 275195
rect 14355 275005 27925 275195
rect 27955 275005 28085 275195
rect 28115 275005 28245 275195
rect 28275 275005 28405 275195
rect 28435 275005 28565 275195
rect 28595 275005 28725 275195
rect 28755 275005 28760 275195
rect 1000 275000 28760 275005
rect 262 -400 318 240
rect 853 -400 909 240
rect 1444 -400 1500 240
rect 2035 -400 2091 240
rect 2626 -400 2682 240
rect 3217 -400 3273 240
rect 3808 -400 3864 240
rect 4399 -400 4455 240
rect 4990 -400 5046 240
rect 5581 -400 5637 240
rect 6172 -400 6228 240
rect 6763 -400 6819 240
rect 7354 -400 7410 240
rect 7945 -400 8001 240
rect 8536 -400 8592 240
rect 9127 -400 9183 240
rect 9718 -400 9774 240
rect 10309 -400 10365 240
rect 10900 -400 10956 240
rect 11491 -400 11547 240
rect 12082 -400 12138 240
rect 12673 -400 12729 240
rect 13264 -400 13320 240
rect 13855 -400 13911 240
rect 14446 -400 14502 240
rect 15037 -400 15093 240
rect 15628 -400 15684 240
rect 16219 -400 16275 240
rect 16810 -400 16866 240
rect 17401 -400 17457 240
rect 17992 -400 18048 240
rect 18583 -400 18639 240
rect 19174 -400 19230 240
rect 19765 -400 19821 240
rect 20356 -400 20412 240
rect 20947 -400 21003 240
rect 21538 -400 21594 240
rect 22129 -400 22185 240
rect 22720 -400 22776 240
rect 23311 -400 23367 240
rect 23902 -400 23958 240
rect 24493 -400 24549 240
rect 25084 -400 25140 240
rect 25675 -400 25731 240
rect 26266 -400 26322 240
rect 26857 -400 26913 240
rect 27448 -400 27504 240
rect 28039 -400 28095 240
rect 28630 -400 28686 240
rect 29221 -400 29277 240
rect 29812 -400 29868 240
rect 30403 -400 30459 240
rect 30994 -400 31050 240
rect 31585 -400 31641 240
rect 32176 -400 32232 240
rect 32767 -400 32823 240
rect 33358 -400 33414 240
rect 33949 -400 34005 240
rect 34540 -400 34596 240
rect 35131 -400 35187 240
rect 35722 -400 35778 240
rect 36313 -400 36369 240
rect 36904 -400 36960 240
rect 37495 -400 37551 240
rect 38086 -400 38142 240
rect 38677 -400 38733 240
rect 39268 -400 39324 240
rect 39859 -400 39915 240
rect 40450 -400 40506 240
rect 41041 -400 41097 240
rect 41632 -400 41688 240
rect 42223 -400 42279 240
rect 42814 -400 42870 240
rect 43405 -400 43461 240
rect 43996 -400 44052 240
rect 44587 -400 44643 240
rect 45178 -400 45234 240
rect 45769 -400 45825 240
rect 46360 -400 46416 240
rect 46951 -400 47007 240
rect 47542 -400 47598 240
rect 48133 -400 48189 240
rect 48724 -400 48780 240
rect 49315 -400 49371 240
rect 49906 -400 49962 240
rect 50497 -400 50553 240
rect 51088 -400 51144 240
rect 51679 -400 51735 240
rect 52270 -400 52326 240
rect 52861 -400 52917 240
rect 53452 -400 53508 240
rect 54043 -400 54099 240
rect 54634 -400 54690 240
rect 55225 -400 55281 240
rect 55816 -400 55872 240
rect 56407 -400 56463 240
rect 56998 -400 57054 240
rect 57589 -400 57645 240
rect 58180 -400 58236 240
rect 58771 -400 58827 240
rect 59362 -400 59418 240
rect 59953 -400 60009 240
rect 60544 -400 60600 240
rect 61135 -400 61191 240
rect 61726 -400 61782 240
rect 62317 -400 62373 240
rect 62908 -400 62964 240
rect 63499 -400 63555 240
rect 64090 -400 64146 240
rect 64681 -400 64737 240
rect 65272 -400 65328 240
rect 65863 -400 65919 240
rect 66454 -400 66510 240
rect 67045 -400 67101 240
rect 67636 -400 67692 240
rect 68227 -400 68283 240
rect 68818 -400 68874 240
rect 69409 -400 69465 240
rect 70000 -400 70056 240
rect 70591 -400 70647 240
rect 71182 -400 71238 240
rect 71773 -400 71829 240
rect 72364 -400 72420 240
rect 72955 -400 73011 240
rect 73546 -400 73602 240
rect 74137 -400 74193 240
rect 74728 -400 74784 240
rect 75319 -400 75375 240
rect 75910 -400 75966 240
rect 76501 -400 76557 240
rect 77092 -400 77148 240
rect 77683 -400 77739 240
rect 78274 -400 78330 240
rect 78865 -400 78921 240
rect 79456 -400 79512 240
rect 80047 -400 80103 240
rect 80638 -400 80694 240
rect 81229 -400 81285 240
rect 81820 -400 81876 240
rect 82411 -400 82467 240
rect 83002 -400 83058 240
rect 83593 -400 83649 240
rect 84184 -400 84240 240
rect 84775 -400 84831 240
rect 85366 -400 85422 240
rect 85957 -400 86013 240
rect 86548 -400 86604 240
rect 87139 -400 87195 240
rect 87730 -400 87786 240
rect 88321 -400 88377 240
rect 88912 -400 88968 240
rect 89503 -400 89559 240
rect 90094 -400 90150 240
rect 90685 -400 90741 240
rect 91276 -400 91332 240
rect 91867 -400 91923 240
rect 92458 -400 92514 240
rect 93049 -400 93105 240
rect 93640 -400 93696 240
rect 94231 -400 94287 240
rect 94822 -400 94878 240
rect 95413 -400 95469 240
rect 96004 -400 96060 240
rect 96595 -400 96651 240
rect 97186 -400 97242 240
rect 97777 -400 97833 240
rect 98368 -400 98424 240
rect 98959 -400 99015 240
rect 99550 -400 99606 240
rect 100141 -400 100197 240
rect 100732 -400 100788 240
rect 101323 -400 101379 240
rect 101914 -400 101970 240
rect 102505 -400 102561 240
rect 103096 -400 103152 240
rect 103687 -400 103743 240
rect 104278 -400 104334 240
rect 104869 -400 104925 240
rect 105460 -400 105516 240
rect 106051 -400 106107 240
rect 106642 -400 106698 240
rect 107233 -400 107289 240
rect 107824 -400 107880 240
rect 108415 -400 108471 240
rect 109006 -400 109062 240
rect 109597 -400 109653 240
rect 110188 -400 110244 240
rect 110779 -400 110835 240
rect 111370 -400 111426 240
rect 111961 -400 112017 240
rect 112552 -400 112608 240
rect 113143 -400 113199 240
rect 113734 -400 113790 240
rect 114325 -400 114381 240
rect 114916 -400 114972 240
rect 115507 -400 115563 240
rect 116098 -400 116154 240
rect 116689 -400 116745 240
rect 117280 -400 117336 240
rect 117871 -400 117927 240
rect 118462 -400 118518 240
rect 119053 -400 119109 240
rect 119644 -400 119700 240
rect 120235 -400 120291 240
rect 120826 -400 120882 240
rect 121417 -400 121473 240
rect 122008 -400 122064 240
rect 122599 -400 122655 240
rect 123190 -400 123246 240
rect 123781 -400 123837 240
rect 124372 -400 124428 240
rect 124963 -400 125019 240
rect 125554 -400 125610 240
rect 126145 -400 126201 240
rect 126736 -400 126792 240
rect 127327 -400 127383 240
rect 127918 -400 127974 240
rect 128509 -400 128565 240
rect 129100 -400 129156 240
rect 129691 -400 129747 240
rect 130282 -400 130338 240
rect 130873 -400 130929 240
rect 131464 -400 131520 240
rect 132055 -400 132111 240
rect 132646 -400 132702 240
rect 133237 -400 133293 240
rect 133828 -400 133884 240
rect 134419 -400 134475 240
rect 135010 -400 135066 240
rect 135601 -400 135657 240
rect 136192 -400 136248 240
rect 136783 -400 136839 240
rect 137374 -400 137430 240
rect 137965 -400 138021 240
rect 138556 -400 138612 240
rect 139147 -400 139203 240
rect 139738 -400 139794 240
rect 140329 -400 140385 240
rect 140920 -400 140976 240
rect 141511 -400 141567 240
rect 142102 -400 142158 240
rect 142693 -400 142749 240
rect 143284 -400 143340 240
rect 143875 -400 143931 240
rect 144466 -400 144522 240
rect 145057 -400 145113 240
rect 145648 -400 145704 240
rect 146239 -400 146295 240
rect 146830 -400 146886 240
rect 147421 -400 147477 240
rect 148012 -400 148068 240
rect 148603 -400 148659 240
rect 149194 -400 149250 240
rect 149785 -400 149841 240
rect 150376 -400 150432 240
rect 150967 -400 151023 240
rect 151558 -400 151614 240
rect 152149 -400 152205 240
rect 152740 -400 152796 240
rect 153331 -400 153387 240
rect 153922 -400 153978 240
rect 154513 -400 154569 240
rect 155104 -400 155160 240
rect 155695 -400 155751 240
rect 156286 -400 156342 240
rect 156877 -400 156933 240
rect 157468 -400 157524 240
rect 158059 -400 158115 240
rect 158650 -400 158706 240
rect 159241 -400 159297 240
rect 159832 -400 159888 240
rect 160423 -400 160479 240
rect 161014 -400 161070 240
rect 161605 -400 161661 240
rect 162196 -400 162252 240
rect 162787 -400 162843 240
rect 163378 -400 163434 240
rect 163969 -400 164025 240
rect 164560 -400 164616 240
rect 165151 -400 165207 240
rect 165742 -400 165798 240
rect 166333 -400 166389 240
rect 166924 -400 166980 240
rect 167515 -400 167571 240
rect 168106 -400 168162 240
rect 168697 -400 168753 240
rect 169288 -400 169344 240
rect 169879 -400 169935 240
rect 170470 -400 170526 240
rect 171061 -400 171117 240
rect 171652 -400 171708 240
rect 172243 -400 172299 240
rect 172834 -400 172890 240
rect 173425 -400 173481 240
rect 174016 -400 174072 240
rect 174607 -400 174663 240
rect 175198 -400 175254 240
rect 175789 -400 175845 240
rect 176380 -400 176436 240
rect 176971 -400 177027 240
rect 177562 -400 177618 240
rect 178153 -400 178209 240
rect 178744 -400 178800 240
rect 179335 -400 179391 240
rect 179926 -400 179982 240
rect 180517 -400 180573 240
rect 181108 -400 181164 240
rect 181699 -400 181755 240
rect 182290 -400 182346 240
rect 182881 -400 182937 240
rect 183472 -400 183528 240
rect 184063 -400 184119 240
rect 184654 -400 184710 240
rect 185245 -400 185301 240
rect 185836 -400 185892 240
rect 186427 -400 186483 240
rect 187018 -400 187074 240
rect 187609 -400 187665 240
rect 188200 -400 188256 240
rect 188791 -400 188847 240
rect 189382 -400 189438 240
rect 189973 -400 190029 240
rect 190564 -400 190620 240
rect 191155 -400 191211 240
rect 191746 -400 191802 240
rect 192337 -400 192393 240
rect 192928 -400 192984 240
rect 193519 -400 193575 240
rect 194110 -400 194166 240
rect 194701 -400 194757 240
rect 195292 -400 195348 240
rect 195883 -400 195939 240
rect 196474 -400 196530 240
rect 197065 -400 197121 240
rect 197656 -400 197712 240
rect 198247 -400 198303 240
rect 198838 -400 198894 240
rect 199429 -400 199485 240
rect 200020 -400 200076 240
rect 200611 -400 200667 240
rect 201202 -400 201258 240
rect 201793 -400 201849 240
rect 202384 -400 202440 240
rect 202975 -400 203031 240
rect 203566 -400 203622 240
rect 204157 -400 204213 240
rect 204748 -400 204804 240
rect 205339 -400 205395 240
rect 205930 -400 205986 240
rect 206521 -400 206577 240
rect 207112 -400 207168 240
rect 207703 -400 207759 240
rect 208294 -400 208350 240
rect 208885 -400 208941 240
rect 209476 -400 209532 240
rect 210067 -400 210123 240
rect 210658 -400 210714 240
rect 211249 -400 211305 240
rect 211840 -400 211896 240
rect 212431 -400 212487 240
rect 213022 -400 213078 240
rect 213613 -400 213669 240
rect 214204 -400 214260 240
rect 214795 -400 214851 240
rect 215386 -400 215442 240
rect 215977 -400 216033 240
rect 216568 -400 216624 240
rect 217159 -400 217215 240
rect 217750 -400 217806 240
rect 218341 -400 218397 240
rect 218932 -400 218988 240
rect 219523 -400 219579 240
rect 220114 -400 220170 240
rect 220705 -400 220761 240
rect 221296 -400 221352 240
rect 221887 -400 221943 240
rect 222478 -400 222534 240
rect 223069 -400 223125 240
rect 223660 -400 223716 240
rect 224251 -400 224307 240
rect 224842 -400 224898 240
rect 225433 -400 225489 240
rect 226024 -400 226080 240
rect 226615 -400 226671 240
rect 227206 -400 227262 240
rect 227797 -400 227853 240
rect 228388 -400 228444 240
rect 228979 -400 229035 240
rect 229570 -400 229626 240
rect 230161 -400 230217 240
rect 230752 -400 230808 240
rect 231343 -400 231399 240
rect 231934 -400 231990 240
rect 232525 -400 232581 240
rect 233116 -400 233172 240
rect 233707 -400 233763 240
rect 234298 -400 234354 240
rect 234889 -400 234945 240
rect 235480 -400 235536 240
rect 236071 -400 236127 240
rect 236662 -400 236718 240
rect 237253 -400 237309 240
rect 237844 -400 237900 240
rect 238435 -400 238491 240
rect 239026 -400 239082 240
rect 239617 -400 239673 240
rect 240208 -400 240264 240
rect 240799 -400 240855 240
rect 241390 -400 241446 240
rect 241981 -400 242037 240
rect 242572 -400 242628 240
rect 243163 -400 243219 240
rect 243754 -400 243810 240
rect 244345 -400 244401 240
rect 244936 -400 244992 240
rect 245527 -400 245583 240
rect 246118 -400 246174 240
rect 246709 -400 246765 240
rect 247300 -400 247356 240
rect 247891 -400 247947 240
rect 248482 -400 248538 240
rect 249073 -400 249129 240
rect 249664 -400 249720 240
rect 250255 -400 250311 240
rect 250846 -400 250902 240
rect 251437 -400 251493 240
rect 252028 -400 252084 240
rect 252619 -400 252675 240
rect 253210 -400 253266 240
rect 253801 -400 253857 240
rect 254392 -400 254448 240
rect 254983 -400 255039 240
rect 255574 -400 255630 240
rect 256165 -400 256221 240
rect 256756 -400 256812 240
rect 257347 -400 257403 240
rect 257938 -400 257994 240
rect 258529 -400 258585 240
rect 259120 -400 259176 240
rect 259711 -400 259767 240
rect 260302 -400 260358 240
rect 260893 -400 260949 240
rect 261484 -400 261540 240
rect 262075 -400 262131 240
rect 262666 -400 262722 240
rect 263257 -400 263313 240
rect 263848 -400 263904 240
rect 264439 -400 264495 240
rect 265030 -400 265086 240
rect 265621 -400 265677 240
rect 266212 -400 266268 240
rect 266803 -400 266859 240
rect 267394 -400 267450 240
rect 267985 -400 268041 240
rect 268576 -400 268632 240
rect 269167 -400 269223 240
rect 269758 -400 269814 240
rect 270349 -400 270405 240
rect 270940 -400 270996 240
rect 271531 -400 271587 240
rect 272122 -400 272178 240
rect 272713 -400 272769 240
rect 273304 -400 273360 240
rect 273895 -400 273951 240
rect 274486 -400 274542 240
rect 275077 -400 275133 240
rect 275668 -400 275724 240
rect 276259 -400 276315 240
rect 276850 -400 276906 240
rect 277441 -400 277497 240
rect 278032 -400 278088 240
rect 278623 -400 278679 240
rect 279214 -400 279270 240
rect 279805 -400 279861 240
rect 280396 -400 280452 240
rect 280987 -400 281043 240
rect 281578 -400 281634 240
rect 282169 -400 282225 240
rect 282760 -400 282816 240
rect 283351 -400 283407 240
rect 283942 -400 283998 240
rect 284533 -400 284589 240
rect 285124 -400 285180 240
rect 285715 -400 285771 240
rect 286306 -400 286362 240
rect 286897 -400 286953 240
rect 287488 -400 287544 240
rect 288079 -400 288135 240
rect 288670 -400 288726 240
rect 289261 -400 289317 240
rect 289852 -400 289908 240
rect 290443 -400 290499 240
rect 291034 -400 291090 240
rect 291625 -400 291681 240
<< via2 >>
rect 10725 351365 10755 351395
rect 10805 351365 10835 351395
rect 10885 351365 10915 351395
rect 10965 351365 10995 351395
rect 11045 351365 11075 351395
rect 11125 351365 11155 351395
rect 11205 351365 11235 351395
rect 11285 351365 11315 351395
rect 11365 351365 11395 351395
rect 11445 351365 11475 351395
rect 11525 351365 11555 351395
rect 11605 351365 11635 351395
rect 11685 351365 11715 351395
rect 11765 351365 11795 351395
rect 11845 351365 11875 351395
rect 11925 351365 11955 351395
rect 12005 351365 12035 351395
rect 12085 351365 12115 351395
rect 12165 351365 12195 351395
rect 12245 351365 12275 351395
rect 12325 351365 12355 351395
rect 12405 351365 12435 351395
rect 12485 351365 12515 351395
rect 12565 351365 12595 351395
rect 12645 351365 12675 351395
rect 12725 351365 12755 351395
rect 12805 351365 12835 351395
rect 12885 351365 12915 351395
rect 12965 351365 12995 351395
rect 13045 351365 13075 351395
rect 13125 351365 13155 351395
rect 13205 351365 13235 351395
rect 13285 351365 13315 351395
rect 13365 351365 13395 351395
rect 13445 351365 13475 351395
rect 13525 351365 13555 351395
rect 13605 351365 13635 351395
rect 13685 351365 13715 351395
rect 13765 351365 13795 351395
rect 13845 351365 13875 351395
rect 13925 351365 13955 351395
rect 14005 351365 14035 351395
rect 14085 351365 14115 351395
rect 14165 351365 14195 351395
rect 14245 351365 14275 351395
rect 14325 351365 14355 351395
rect 14405 351365 14435 351395
rect 14485 351365 14515 351395
rect 14565 351365 14595 351395
rect 14645 351365 14675 351395
rect 14725 351365 14755 351395
rect 14805 351365 14835 351395
rect 14885 351365 14915 351395
rect 14965 351365 14995 351395
rect 15045 351365 15075 351395
rect 15125 351365 15155 351395
rect 15205 351365 15235 351395
rect 15285 351365 15315 351395
rect 15365 351365 15395 351395
rect 15445 351365 15475 351395
rect 15525 351365 15555 351395
rect 15605 351365 15635 351395
rect 15685 351365 15715 351395
rect 15765 351365 15795 351395
rect 15845 351365 15875 351395
rect 15925 351365 15955 351395
rect 16005 351365 16035 351395
rect 16085 351365 16115 351395
rect 16165 351365 16195 351395
rect 16245 351365 16275 351395
rect 16325 351365 16355 351395
rect 16405 351365 16435 351395
rect 16485 351365 16515 351395
rect 16565 351365 16595 351395
rect 16645 351365 16675 351395
rect 16725 351365 16755 351395
rect 16805 351365 16835 351395
rect 16885 351365 16915 351395
rect 16965 351365 16995 351395
rect 17045 351365 17075 351395
rect 17125 351365 17155 351395
rect 17205 351365 17235 351395
rect 17285 351365 17315 351395
rect 17365 351365 17395 351395
rect 17445 351365 17475 351395
rect 17525 351365 17555 351395
rect 17605 351365 17635 351395
rect 17685 351365 17715 351395
rect 17765 351365 17795 351395
rect 17845 351365 17875 351395
rect 17925 351365 17955 351395
rect 18005 351365 18035 351395
rect 18085 351365 18115 351395
rect 18165 351365 18195 351395
rect 18245 351365 18275 351395
rect 18325 351365 18355 351395
rect 18405 351365 18435 351395
rect 18485 351365 18515 351395
rect 18565 351365 18595 351395
rect 18645 351365 18675 351395
rect 18725 351365 18755 351395
rect 18805 351365 18835 351395
rect 18885 351365 18915 351395
rect 18965 351365 18995 351395
rect 19045 351365 19075 351395
rect 19125 351365 19155 351395
rect 19205 351365 19235 351395
rect 19285 351365 19315 351395
rect 19365 351365 19395 351395
rect 19445 351365 19475 351395
rect 19525 351365 19555 351395
rect 19605 351365 19635 351395
rect 19685 351365 19715 351395
rect 19845 351365 19875 351395
rect 10645 351285 10675 351315
rect 19765 351285 19795 351315
rect 10725 351205 10755 351235
rect 10805 351205 10835 351235
rect 10885 351205 10915 351235
rect 10965 351205 10995 351235
rect 11045 351205 11075 351235
rect 11125 351205 11155 351235
rect 11205 351205 11235 351235
rect 11285 351205 11315 351235
rect 11365 351205 11395 351235
rect 11445 351205 11475 351235
rect 11525 351205 11555 351235
rect 11605 351205 11635 351235
rect 11685 351205 11715 351235
rect 11765 351205 11795 351235
rect 11845 351205 11875 351235
rect 11925 351205 11955 351235
rect 12005 351205 12035 351235
rect 12085 351205 12115 351235
rect 12165 351205 12195 351235
rect 12245 351205 12275 351235
rect 12325 351205 12355 351235
rect 12405 351205 12435 351235
rect 12485 351205 12515 351235
rect 12565 351205 12595 351235
rect 12645 351205 12675 351235
rect 12725 351205 12755 351235
rect 12805 351205 12835 351235
rect 12885 351205 12915 351235
rect 12965 351205 12995 351235
rect 13045 351205 13075 351235
rect 13125 351205 13155 351235
rect 13205 351205 13235 351235
rect 13285 351205 13315 351235
rect 13365 351205 13395 351235
rect 13445 351205 13475 351235
rect 13525 351205 13555 351235
rect 13605 351205 13635 351235
rect 13685 351205 13715 351235
rect 13765 351205 13795 351235
rect 13845 351205 13875 351235
rect 13925 351205 13955 351235
rect 14005 351205 14035 351235
rect 14085 351205 14115 351235
rect 14165 351205 14195 351235
rect 14245 351205 14275 351235
rect 14325 351205 14355 351235
rect 14405 351205 14435 351235
rect 14485 351205 14515 351235
rect 14565 351205 14595 351235
rect 14645 351205 14675 351235
rect 14725 351205 14755 351235
rect 14805 351205 14835 351235
rect 14885 351205 14915 351235
rect 14965 351205 14995 351235
rect 15045 351205 15075 351235
rect 15125 351205 15155 351235
rect 15205 351205 15235 351235
rect 15285 351205 15315 351235
rect 15365 351205 15395 351235
rect 15445 351205 15475 351235
rect 15525 351205 15555 351235
rect 15605 351205 15635 351235
rect 15685 351205 15715 351235
rect 15765 351205 15795 351235
rect 15845 351205 15875 351235
rect 15925 351205 15955 351235
rect 16005 351205 16035 351235
rect 16085 351205 16115 351235
rect 16165 351205 16195 351235
rect 16245 351205 16275 351235
rect 16325 351205 16355 351235
rect 16405 351205 16435 351235
rect 16485 351205 16515 351235
rect 16565 351205 16595 351235
rect 16645 351205 16675 351235
rect 16725 351205 16755 351235
rect 16805 351205 16835 351235
rect 16885 351205 16915 351235
rect 16965 351205 16995 351235
rect 17045 351205 17075 351235
rect 17125 351205 17155 351235
rect 17205 351205 17235 351235
rect 17285 351205 17315 351235
rect 17365 351205 17395 351235
rect 17445 351205 17475 351235
rect 17525 351205 17555 351235
rect 17605 351205 17635 351235
rect 17685 351205 17715 351235
rect 17765 351205 17795 351235
rect 17845 351205 17875 351235
rect 17925 351205 17955 351235
rect 18005 351205 18035 351235
rect 18085 351205 18115 351235
rect 18165 351205 18195 351235
rect 18245 351205 18275 351235
rect 18325 351205 18355 351235
rect 18405 351205 18435 351235
rect 18485 351205 18515 351235
rect 18565 351205 18595 351235
rect 18645 351205 18675 351235
rect 18725 351205 18755 351235
rect 18805 351205 18835 351235
rect 18885 351205 18915 351235
rect 18965 351205 18995 351235
rect 19045 351205 19075 351235
rect 19125 351205 19155 351235
rect 19205 351205 19235 351235
rect 19285 351205 19315 351235
rect 19365 351205 19395 351235
rect 19445 351205 19475 351235
rect 19525 351205 19555 351235
rect 19605 351205 19635 351235
rect 19685 351205 19715 351235
rect 19845 351205 19875 351235
rect 19685 351125 19715 351155
rect 19845 351125 19875 351155
rect 19685 351045 19715 351075
rect 19845 351045 19875 351075
rect 19685 350965 19715 350995
rect 19845 350965 19875 350995
rect 19685 350885 19715 350915
rect 19845 350885 19875 350915
rect 19685 350805 19715 350835
rect 19845 350805 19875 350835
rect 19685 350725 19715 350755
rect 19845 350725 19875 350755
rect 19685 350645 19715 350675
rect 19845 350645 19875 350675
rect 19685 350565 19715 350595
rect 19845 350565 19875 350595
rect 19685 350485 19715 350515
rect 19845 350485 19875 350515
rect 19685 350405 19715 350435
rect 19845 350405 19875 350435
rect 19685 350325 19715 350355
rect 19845 350325 19875 350355
rect 19685 350245 19715 350275
rect 19845 350245 19875 350275
rect 19685 350165 19715 350195
rect 19845 350165 19875 350195
rect 19685 350085 19715 350115
rect 19845 350085 19875 350115
rect 19685 350005 19715 350035
rect 19845 350005 19875 350035
rect 19685 349925 19715 349955
rect 19845 349925 19875 349955
rect 19685 349845 19715 349875
rect 19845 349845 19875 349875
rect 19685 349765 19715 349795
rect 19845 349765 19875 349795
rect 19685 349685 19715 349715
rect 19845 349685 19875 349715
rect 19685 349605 19715 349635
rect 19845 349605 19875 349635
rect 19685 349525 19715 349555
rect 19845 349525 19875 349555
rect 19685 349445 19715 349475
rect 19845 349445 19875 349475
rect 19685 349365 19715 349395
rect 19845 349365 19875 349395
rect 19685 349285 19715 349315
rect 19845 349285 19875 349315
rect 19685 349205 19715 349235
rect 19845 349205 19875 349235
rect 19685 349125 19715 349155
rect 19845 349125 19875 349155
rect 19685 349045 19715 349075
rect 19845 349045 19875 349075
rect 19685 348965 19715 348995
rect 19845 348965 19875 348995
rect 19685 348885 19715 348915
rect 19845 348885 19875 348915
rect 19685 348805 19715 348835
rect 19845 348805 19875 348835
rect 19685 348725 19715 348755
rect 19845 348725 19875 348755
rect 19685 348645 19715 348675
rect 19845 348645 19875 348675
rect 19685 348565 19715 348595
rect 19845 348565 19875 348595
rect 19685 348485 19715 348515
rect 19845 348485 19875 348515
rect 19685 348405 19715 348435
rect 19845 348405 19875 348435
rect 19685 348325 19715 348355
rect 19845 348325 19875 348355
rect 19685 348245 19715 348275
rect 19845 348245 19875 348275
rect 19685 348165 19715 348195
rect 19845 348165 19875 348195
rect 19685 348085 19715 348115
rect 19845 348085 19875 348115
rect 19685 348005 19715 348035
rect 19845 348005 19875 348035
rect 19685 347925 19715 347955
rect 19845 347925 19875 347955
rect 19685 347845 19715 347875
rect 19845 347845 19875 347875
rect 19685 347765 19715 347795
rect 19845 347765 19875 347795
rect 19685 347685 19715 347715
rect 19845 347685 19875 347715
rect 19685 347605 19715 347635
rect 19845 347605 19875 347635
rect 19685 347525 19715 347555
rect 19845 347525 19875 347555
rect 19685 347445 19715 347475
rect 19845 347445 19875 347475
rect 19685 347365 19715 347395
rect 19845 347365 19875 347395
rect 19685 347285 19715 347315
rect 19845 347285 19875 347315
rect 19685 347205 19715 347235
rect 19845 347205 19875 347235
rect 19685 347125 19715 347155
rect 19845 347125 19875 347155
rect 19685 347045 19715 347075
rect 19845 347045 19875 347075
rect 19685 346965 19715 346995
rect 19845 346965 19875 346995
rect 19685 346885 19715 346915
rect 19845 346885 19875 346915
rect 19685 346805 19715 346835
rect 19845 346805 19875 346835
rect 19685 346725 19715 346755
rect 19845 346725 19875 346755
rect 19685 346645 19715 346675
rect 19845 346645 19875 346675
rect 19685 346565 19715 346595
rect 19845 346565 19875 346595
rect 19685 346485 19715 346515
rect 19845 346485 19875 346515
rect 19685 346405 19715 346435
rect 19845 346405 19875 346435
rect 19685 346325 19715 346355
rect 19845 346325 19875 346355
rect 19685 346245 19715 346275
rect 19845 346245 19875 346275
rect 19685 346165 19715 346195
rect 19845 346165 19875 346195
rect 19685 346085 19715 346115
rect 19845 346085 19875 346115
rect 19685 346005 19715 346035
rect 19845 346005 19875 346035
rect 19685 345925 19715 345955
rect 19845 345925 19875 345955
rect 19685 345845 19715 345875
rect 19845 345845 19875 345875
rect 19685 345765 19715 345795
rect 19845 345765 19875 345795
rect 19685 345685 19715 345715
rect 19845 345685 19875 345715
rect 19685 345605 19715 345635
rect 19845 345605 19875 345635
rect 19685 345525 19715 345555
rect 19845 345525 19875 345555
rect 19685 345445 19715 345475
rect 19845 345445 19875 345475
rect 19685 345365 19715 345395
rect 19845 345365 19875 345395
rect 19685 345285 19715 345315
rect 19845 345285 19875 345315
rect 19685 345205 19715 345235
rect 19845 345205 19875 345235
rect 19685 345125 19715 345155
rect 19845 345125 19875 345155
rect 19685 345045 19715 345075
rect 19845 345045 19875 345075
rect 19685 344965 19715 344995
rect 19845 344965 19875 344995
rect 19685 344885 19715 344915
rect 19845 344885 19875 344915
rect 19685 344805 19715 344835
rect 19845 344805 19875 344835
rect 19685 344725 19715 344755
rect 19845 344725 19875 344755
rect 19685 344645 19715 344675
rect 19845 344645 19875 344675
rect 19685 344565 19715 344595
rect 19845 344565 19875 344595
rect 19685 344485 19715 344515
rect 19845 344485 19875 344515
rect 19685 344405 19715 344435
rect 19845 344405 19875 344435
rect 19685 344325 19715 344355
rect 19845 344325 19875 344355
rect 19685 344245 19715 344275
rect 19845 344245 19875 344275
rect 19685 344165 19715 344195
rect 19845 344165 19875 344195
rect 19685 344085 19715 344115
rect 19845 344085 19875 344115
rect 19685 344005 19715 344035
rect 19845 344005 19875 344035
rect 19685 343925 19715 343955
rect 19845 343925 19875 343955
rect 19685 343845 19715 343875
rect 19845 343845 19875 343875
rect 19685 343765 19715 343795
rect 19845 343765 19875 343795
rect 19685 343685 19715 343715
rect 19845 343685 19875 343715
rect 19685 343605 19715 343635
rect 19845 343605 19875 343635
rect 19685 343525 19715 343555
rect 19845 343525 19875 343555
rect 19685 343445 19715 343475
rect 19845 343445 19875 343475
rect 19685 343365 19715 343395
rect 19845 343365 19875 343395
rect 19685 343285 19715 343315
rect 19845 343285 19875 343315
rect 19685 343205 19715 343235
rect 19845 343205 19875 343235
rect 19685 343125 19715 343155
rect 19845 343125 19875 343155
rect 19685 343045 19715 343075
rect 19845 343045 19875 343075
rect 19685 342965 19715 342995
rect 19845 342965 19875 342995
rect 19685 342885 19715 342915
rect 19845 342885 19875 342915
rect 19685 342805 19715 342835
rect 19845 342805 19875 342835
rect 19685 342725 19715 342755
rect 19845 342725 19875 342755
rect 19685 342645 19715 342675
rect 19845 342645 19875 342675
rect 19685 342565 19715 342595
rect 19845 342565 19875 342595
rect 19685 342485 19715 342515
rect 19845 342485 19875 342515
rect 19685 342405 19715 342435
rect 19845 342405 19875 342435
rect 19685 342325 19715 342355
rect 19845 342325 19875 342355
rect 19685 342245 19715 342275
rect 19845 342245 19875 342275
rect 19685 342165 19715 342195
rect 19845 342165 19875 342195
rect 19685 342085 19715 342115
rect 19845 342085 19875 342115
rect 19685 342005 19715 342035
rect 19845 342005 19875 342035
rect 19685 341925 19715 341955
rect 19845 341925 19875 341955
rect 19685 341845 19715 341875
rect 19845 341845 19875 341875
rect 19685 341765 19715 341795
rect 19845 341765 19875 341795
rect 19685 341685 19715 341715
rect 19845 341685 19875 341715
rect 19685 341605 19715 341635
rect 19845 341605 19875 341635
rect 19685 341525 19715 341555
rect 19845 341525 19875 341555
rect 19685 341445 19715 341475
rect 19845 341445 19875 341475
rect 19685 341365 19715 341395
rect 19845 341365 19875 341395
rect 19685 341285 19715 341315
rect 19845 341285 19875 341315
rect 19685 341205 19715 341235
rect 19845 341205 19875 341235
rect 19685 341125 19715 341155
rect 19845 341125 19875 341155
rect 19685 341045 19715 341075
rect 19845 341045 19875 341075
rect 19685 340965 19715 340995
rect 19845 340965 19875 340995
rect 19685 340885 19715 340915
rect 19845 340885 19875 340915
rect 19685 340805 19715 340835
rect 19845 340805 19875 340835
rect 19685 340725 19715 340755
rect 19845 340725 19875 340755
rect 19685 340645 19715 340675
rect 19845 340645 19875 340675
rect 19685 340565 19715 340595
rect 19845 340565 19875 340595
rect 19685 340485 19715 340515
rect 19845 340485 19875 340515
rect 19685 340405 19715 340435
rect 19845 340405 19875 340435
rect 19685 340325 19715 340355
rect 19845 340325 19875 340355
rect 19685 340245 19715 340275
rect 19845 340245 19875 340275
rect 19685 340165 19715 340195
rect 19845 340165 19875 340195
rect 19685 340085 19715 340115
rect 19845 340085 19875 340115
rect 19685 340005 19715 340035
rect 19845 340005 19875 340035
rect 19685 339925 19715 339955
rect 19845 339925 19875 339955
rect 19685 339845 19715 339875
rect 19845 339845 19875 339875
rect 19685 339765 19715 339795
rect 19845 339765 19875 339795
rect 19685 339685 19715 339715
rect 19845 339685 19875 339715
rect 19685 339605 19715 339635
rect 19845 339605 19875 339635
rect 19685 339525 19715 339555
rect 19845 339525 19875 339555
rect 19685 339445 19715 339475
rect 19845 339445 19875 339475
rect 19685 339365 19715 339395
rect 19845 339365 19875 339395
rect 19685 339285 19715 339315
rect 19845 339285 19875 339315
rect 19685 339205 19715 339235
rect 19845 339205 19875 339235
rect 19685 339125 19715 339155
rect 19845 339125 19875 339155
rect 19685 339045 19715 339075
rect 19845 339045 19875 339075
rect 19685 338965 19715 338995
rect 19845 338965 19875 338995
rect 19685 338885 19715 338915
rect 19845 338885 19875 338915
rect 19685 338805 19715 338835
rect 19845 338805 19875 338835
rect 19685 338725 19715 338755
rect 19845 338725 19875 338755
rect 19685 338645 19715 338675
rect 19845 338645 19875 338675
rect 19685 338565 19715 338595
rect 19845 338565 19875 338595
rect 19685 338485 19715 338515
rect 19845 338485 19875 338515
rect 19685 338405 19715 338435
rect 19845 338405 19875 338435
rect 19685 338325 19715 338355
rect 19845 338325 19875 338355
rect 19685 338245 19715 338275
rect 19845 338245 19875 338275
rect 19685 338165 19715 338195
rect 19845 338165 19875 338195
rect 19685 338085 19715 338115
rect 19845 338085 19875 338115
rect 19685 338005 19715 338035
rect 19845 338005 19875 338035
rect 19685 337925 19715 337955
rect 19845 337925 19875 337955
rect 19685 337845 19715 337875
rect 19845 337845 19875 337875
rect 19685 337765 19715 337795
rect 19845 337765 19875 337795
rect 19685 337685 19715 337715
rect 19845 337685 19875 337715
rect 19685 337605 19715 337635
rect 19845 337605 19875 337635
rect 19685 337525 19715 337555
rect 19845 337525 19875 337555
rect 19685 337445 19715 337475
rect 19845 337445 19875 337475
rect 19685 337365 19715 337395
rect 19845 337365 19875 337395
rect 19685 337285 19715 337315
rect 19845 337285 19875 337315
rect 19685 337205 19715 337235
rect 19845 337205 19875 337235
rect 19685 337125 19715 337155
rect 19845 337125 19875 337155
rect 19685 337045 19715 337075
rect 19845 337045 19875 337075
rect 19685 336965 19715 336995
rect 19845 336965 19875 336995
rect 19685 336885 19715 336915
rect 19845 336885 19875 336915
rect 19685 336805 19715 336835
rect 19845 336805 19875 336835
rect 19685 336725 19715 336755
rect 19845 336725 19875 336755
rect 19685 336645 19715 336675
rect 19845 336645 19875 336675
rect 19685 336565 19715 336595
rect 19845 336565 19875 336595
rect 19685 336485 19715 336515
rect 19845 336485 19875 336515
rect 19685 336405 19715 336435
rect 19845 336405 19875 336435
rect 19685 336325 19715 336355
rect 19845 336325 19875 336355
rect 19685 336245 19715 336275
rect 19845 336245 19875 336275
rect 19685 336165 19715 336195
rect 19845 336165 19875 336195
rect 19685 336085 19715 336115
rect 19845 336085 19875 336115
rect 19685 336005 19715 336035
rect 19845 336005 19875 336035
rect 19685 335925 19715 335955
rect 19845 335925 19875 335955
rect 19685 335845 19715 335875
rect 19845 335845 19875 335875
rect 19685 335765 19715 335795
rect 19845 335765 19875 335795
rect 19685 335685 19715 335715
rect 19845 335685 19875 335715
rect 19685 335605 19715 335635
rect 19845 335605 19875 335635
rect 19685 335525 19715 335555
rect 19845 335525 19875 335555
rect 19685 335445 19715 335475
rect 19845 335445 19875 335475
rect 19685 335365 19715 335395
rect 19845 335365 19875 335395
rect 19685 335285 19715 335315
rect 19845 335285 19875 335315
rect 19685 335205 19715 335235
rect 19845 335205 19875 335235
rect 19685 335125 19715 335155
rect 19845 335125 19875 335155
rect 19685 335045 19715 335075
rect 19845 335045 19875 335075
rect 19685 334965 19715 334995
rect 19845 334965 19875 334995
rect 19685 334885 19715 334915
rect 19845 334885 19875 334915
rect 19685 334805 19715 334835
rect 19845 334805 19875 334835
rect 19685 334725 19715 334755
rect 19845 334725 19875 334755
rect 19685 334645 19715 334675
rect 19845 334645 19875 334675
rect 19685 334565 19715 334595
rect 19845 334565 19875 334595
rect 19685 334485 19715 334515
rect 19845 334485 19875 334515
rect 19685 334405 19715 334435
rect 19845 334405 19875 334435
rect 19685 334325 19715 334355
rect 19845 334325 19875 334355
rect 19685 334245 19715 334275
rect 19845 334245 19875 334275
rect 19685 334165 19715 334195
rect 19845 334165 19875 334195
rect 19685 334085 19715 334115
rect 19845 334085 19875 334115
rect 19685 334005 19715 334035
rect 19845 334005 19875 334035
rect 19685 333925 19715 333955
rect 19845 333925 19875 333955
rect 19685 333845 19715 333875
rect 19845 333845 19875 333875
rect 19685 333765 19715 333795
rect 19845 333765 19875 333795
rect 19685 333685 19715 333715
rect 19845 333685 19875 333715
rect 19685 333605 19715 333635
rect 19845 333605 19875 333635
rect 19685 333525 19715 333555
rect 19845 333525 19875 333555
rect 19685 333445 19715 333475
rect 19845 333445 19875 333475
rect 19685 333365 19715 333395
rect 19845 333365 19875 333395
rect 19685 333285 19715 333315
rect 19845 333285 19875 333315
rect 19685 333205 19715 333235
rect 19845 333205 19875 333235
rect 19685 333125 19715 333155
rect 19845 333125 19875 333155
rect 19685 333045 19715 333075
rect 19845 333045 19875 333075
rect 19685 332965 19715 332995
rect 19845 332965 19875 332995
rect 19685 332885 19715 332915
rect 19845 332885 19875 332915
rect 19685 332805 19715 332835
rect 19845 332805 19875 332835
rect 19685 332725 19715 332755
rect 19845 332725 19875 332755
rect 19685 332645 19715 332675
rect 19845 332645 19875 332675
rect 19685 332565 19715 332595
rect 19845 332565 19875 332595
rect 19685 332485 19715 332515
rect 19845 332485 19875 332515
rect 19685 332405 19715 332435
rect 19845 332405 19875 332435
rect 19685 332325 19715 332355
rect 19845 332325 19875 332355
rect 19685 332245 19715 332275
rect 19845 332245 19875 332275
rect 19685 332165 19715 332195
rect 19845 332165 19875 332195
rect 19685 332085 19715 332115
rect 19845 332085 19875 332115
rect 19685 332005 19715 332035
rect 19845 332005 19875 332035
rect 19685 331925 19715 331955
rect 19845 331925 19875 331955
rect 19685 331845 19715 331875
rect 19845 331845 19875 331875
rect 19685 331765 19715 331795
rect 19845 331765 19875 331795
rect 19685 331685 19715 331715
rect 19845 331685 19875 331715
rect 19685 331605 19715 331635
rect 19845 331605 19875 331635
rect 19685 331525 19715 331555
rect 19845 331525 19875 331555
rect 19685 331445 19715 331475
rect 19845 331445 19875 331475
rect 19685 331365 19715 331395
rect 19845 331365 19875 331395
rect 19685 331285 19715 331315
rect 19845 331285 19875 331315
rect 19685 331205 19715 331235
rect 19845 331205 19875 331235
rect 19685 331125 19715 331155
rect 19845 331125 19875 331155
rect 19685 331045 19715 331075
rect 19845 331045 19875 331075
rect 19685 330965 19715 330995
rect 19845 330965 19875 330995
rect 19685 330885 19715 330915
rect 19845 330885 19875 330915
rect 19685 330805 19715 330835
rect 19845 330805 19875 330835
rect 19685 330725 19715 330755
rect 19845 330725 19875 330755
rect 19685 330645 19715 330675
rect 19845 330645 19875 330675
rect 19685 330565 19715 330595
rect 19845 330565 19875 330595
rect 19685 330485 19715 330515
rect 19845 330485 19875 330515
rect 19685 330405 19715 330435
rect 19845 330405 19875 330435
rect 19685 330325 19715 330355
rect 19845 330325 19875 330355
rect 19685 330245 19715 330275
rect 19845 330245 19875 330275
rect 19685 330165 19715 330195
rect 19845 330165 19875 330195
rect 19685 330085 19715 330115
rect 19845 330085 19875 330115
rect 19685 330005 19715 330035
rect 19845 330005 19875 330035
rect 19685 329925 19715 329955
rect 19845 329925 19875 329955
rect 19685 329845 19715 329875
rect 19845 329845 19875 329875
rect 19685 329765 19715 329795
rect 19845 329765 19875 329795
rect 19685 329685 19715 329715
rect 19845 329685 19875 329715
rect 19685 329605 19715 329635
rect 19845 329605 19875 329635
rect 19685 329525 19715 329555
rect 19845 329525 19875 329555
rect 19685 329445 19715 329475
rect 19845 329445 19875 329475
rect 19685 329365 19715 329395
rect 19845 329365 19875 329395
rect 19685 329285 19715 329315
rect 19845 329285 19875 329315
rect 19685 329205 19715 329235
rect 19845 329205 19875 329235
rect 19685 329125 19715 329155
rect 19845 329125 19875 329155
rect 19685 329045 19715 329075
rect 19845 329045 19875 329075
rect 19685 328965 19715 328995
rect 19845 328965 19875 328995
rect 19685 328885 19715 328915
rect 19845 328885 19875 328915
rect 19685 328805 19715 328835
rect 19845 328805 19875 328835
rect 19685 328725 19715 328755
rect 19845 328725 19875 328755
rect 19685 328645 19715 328675
rect 19845 328645 19875 328675
rect 19685 328565 19715 328595
rect 19845 328565 19875 328595
rect 19685 328485 19715 328515
rect 19845 328485 19875 328515
rect 19685 328405 19715 328435
rect 19845 328405 19875 328435
rect 19685 328325 19715 328355
rect 19845 328325 19875 328355
rect 19685 328245 19715 328275
rect 19845 328245 19875 328275
rect 19685 328165 19715 328195
rect 19845 328165 19875 328195
rect 19685 328085 19715 328115
rect 19845 328085 19875 328115
rect 19685 328005 19715 328035
rect 19845 328005 19875 328035
rect 19685 327925 19715 327955
rect 19845 327925 19875 327955
rect 19685 327845 19715 327875
rect 19845 327845 19875 327875
rect 19685 327765 19715 327795
rect 19845 327765 19875 327795
rect 19685 327685 19715 327715
rect 19845 327685 19875 327715
rect 19685 327605 19715 327635
rect 19845 327605 19875 327635
rect 19685 327525 19715 327555
rect 19845 327525 19875 327555
rect 19685 327445 19715 327475
rect 19845 327445 19875 327475
rect 19685 327365 19715 327395
rect 19845 327365 19875 327395
rect 19685 327285 19715 327315
rect 19845 327285 19875 327315
rect 19685 327205 19715 327235
rect 19845 327205 19875 327235
rect 19685 327125 19715 327155
rect 19845 327125 19875 327155
rect 19685 327045 19715 327075
rect 19845 327045 19875 327075
rect 19685 326965 19715 326995
rect 19845 326965 19875 326995
rect 19685 326885 19715 326915
rect 19845 326885 19875 326915
rect 19685 326805 19715 326835
rect 19845 326805 19875 326835
rect 19685 326725 19715 326755
rect 19845 326725 19875 326755
rect 19685 326645 19715 326675
rect 19845 326645 19875 326675
rect 19685 326565 19715 326595
rect 19845 326565 19875 326595
rect 19685 326485 19715 326515
rect 19845 326485 19875 326515
rect 19685 326405 19715 326435
rect 19845 326405 19875 326435
rect 19685 326325 19715 326355
rect 19845 326325 19875 326355
rect 19685 326245 19715 326275
rect 19845 326245 19875 326275
rect 19685 326165 19715 326195
rect 19845 326165 19875 326195
rect 19685 326085 19715 326115
rect 19845 326085 19875 326115
rect 19685 326005 19715 326035
rect 19845 326005 19875 326035
rect 19685 325925 19715 325955
rect 19845 325925 19875 325955
rect 19685 325845 19715 325875
rect 19845 325845 19875 325875
rect 19685 325765 19715 325795
rect 19845 325765 19875 325795
rect 19685 325685 19715 325715
rect 19845 325685 19875 325715
rect 19685 325605 19715 325635
rect 19845 325605 19875 325635
rect 19685 325525 19715 325555
rect 19845 325525 19875 325555
rect 19685 325445 19715 325475
rect 19845 325445 19875 325475
rect 19685 325365 19715 325395
rect 19845 325365 19875 325395
rect 19685 325285 19715 325315
rect 19845 325285 19875 325315
rect 19685 325205 19715 325235
rect 19845 325205 19875 325235
rect 19685 325125 19715 325155
rect 19845 325125 19875 325155
rect 19685 325045 19715 325075
rect 19845 325045 19875 325075
rect 19685 324965 19715 324995
rect 19845 324965 19875 324995
rect 19685 324885 19715 324915
rect 19845 324885 19875 324915
rect 19685 324805 19715 324835
rect 19845 324805 19875 324835
rect 19685 324725 19715 324755
rect 19845 324725 19875 324755
rect 19685 324645 19715 324675
rect 19845 324645 19875 324675
rect 19685 324565 19715 324595
rect 19845 324565 19875 324595
rect 19685 324485 19715 324515
rect 19845 324485 19875 324515
rect 19685 324405 19715 324435
rect 19845 324405 19875 324435
rect 19685 324325 19715 324355
rect 19845 324325 19875 324355
rect 19685 324245 19715 324275
rect 19845 324245 19875 324275
rect 19685 324165 19715 324195
rect 19845 324165 19875 324195
rect 19685 324085 19715 324115
rect 19845 324085 19875 324115
rect 19685 324005 19715 324035
rect 19845 324005 19875 324035
rect 19685 323925 19715 323955
rect 19845 323925 19875 323955
rect 19685 323845 19715 323875
rect 19845 323845 19875 323875
rect 19685 323765 19715 323795
rect 19845 323765 19875 323795
rect 19685 323685 19715 323715
rect 19845 323685 19875 323715
rect 19685 323605 19715 323635
rect 19845 323605 19875 323635
rect 19685 323525 19715 323555
rect 19845 323525 19875 323555
rect 19685 323445 19715 323475
rect 19845 323445 19875 323475
rect 19685 323365 19715 323395
rect 19845 323365 19875 323395
rect 19685 323285 19715 323315
rect 19845 323285 19875 323315
rect 19685 323205 19715 323235
rect 19845 323205 19875 323235
rect 19685 323125 19715 323155
rect 19845 323125 19875 323155
rect 19685 323045 19715 323075
rect 19845 323045 19875 323075
rect 19685 322965 19715 322995
rect 19845 322965 19875 322995
rect 19685 322885 19715 322915
rect 19845 322885 19875 322915
rect 19685 322805 19715 322835
rect 19845 322805 19875 322835
rect 19685 322725 19715 322755
rect 19845 322725 19875 322755
rect 19685 322645 19715 322675
rect 19845 322645 19875 322675
rect 19685 322565 19715 322595
rect 19845 322565 19875 322595
rect 19685 322485 19715 322515
rect 19845 322485 19875 322515
rect 19685 322405 19715 322435
rect 19845 322405 19875 322435
rect 19685 322325 19715 322355
rect 19845 322325 19875 322355
rect 19685 322245 19715 322275
rect 19845 322245 19875 322275
rect 19685 322165 19715 322195
rect 19845 322165 19875 322195
rect 19685 322085 19715 322115
rect 19845 322085 19875 322115
rect 19685 322005 19715 322035
rect 19845 322005 19875 322035
rect 19685 321925 19715 321955
rect 19845 321925 19875 321955
rect 19685 321845 19715 321875
rect 19845 321845 19875 321875
rect 19685 321765 19715 321795
rect 19845 321765 19875 321795
rect 19685 321685 19715 321715
rect 19845 321685 19875 321715
rect 19685 321605 19715 321635
rect 19845 321605 19875 321635
rect 19685 321525 19715 321555
rect 19845 321525 19875 321555
rect 19685 321445 19715 321475
rect 19845 321445 19875 321475
rect 19685 321365 19715 321395
rect 19845 321365 19875 321395
rect 19685 321285 19715 321315
rect 19845 321285 19875 321315
rect 19685 321205 19715 321235
rect 19845 321205 19875 321235
rect 19685 321125 19715 321155
rect 19845 321125 19875 321155
rect 19685 321045 19715 321075
rect 19845 321045 19875 321075
rect 19685 320965 19715 320995
rect 19845 320965 19875 320995
rect 19685 320885 19715 320915
rect 19845 320885 19875 320915
rect 19685 320805 19715 320835
rect 19845 320805 19875 320835
rect 19685 320725 19715 320755
rect 19845 320725 19875 320755
rect 19685 320645 19715 320675
rect 19845 320645 19875 320675
rect 19685 320565 19715 320595
rect 19845 320565 19875 320595
rect 19685 320485 19715 320515
rect 19845 320485 19875 320515
rect 19685 320405 19715 320435
rect 19845 320405 19875 320435
rect 19685 320325 19715 320355
rect 19845 320325 19875 320355
rect 19685 320245 19715 320275
rect 19845 320245 19875 320275
rect 19685 320165 19715 320195
rect 19845 320165 19875 320195
rect 19685 320085 19715 320115
rect 19845 320085 19875 320115
rect 19685 320005 19715 320035
rect 19845 320005 19875 320035
rect 19685 319925 19715 319955
rect 19845 319925 19875 319955
rect 19685 319845 19715 319875
rect 19845 319845 19875 319875
rect 19685 319765 19715 319795
rect 19845 319765 19875 319795
rect 19685 319685 19715 319715
rect 19845 319685 19875 319715
rect 19685 319605 19715 319635
rect 19845 319605 19875 319635
rect 19685 319525 19715 319555
rect 19845 319525 19875 319555
rect 19685 319445 19715 319475
rect 19845 319445 19875 319475
rect 19685 319365 19715 319395
rect 19845 319365 19875 319395
rect 19685 319285 19715 319315
rect 19845 319285 19875 319315
rect 19685 319205 19715 319235
rect 19845 319205 19875 319235
rect 19685 319125 19715 319155
rect 19845 319125 19875 319155
rect 19685 319045 19715 319075
rect 19845 319045 19875 319075
rect 19685 318965 19715 318995
rect 19845 318965 19875 318995
rect 19685 318885 19715 318915
rect 19845 318885 19875 318915
rect 19685 318805 19715 318835
rect 19845 318805 19875 318835
rect 19685 318725 19715 318755
rect 19845 318725 19875 318755
rect 19685 318645 19715 318675
rect 19845 318645 19875 318675
rect 19685 318565 19715 318595
rect 19845 318565 19875 318595
rect 19685 318485 19715 318515
rect 19845 318485 19875 318515
rect 19685 318405 19715 318435
rect 19845 318405 19875 318435
rect 19685 318325 19715 318355
rect 19845 318325 19875 318355
rect 19685 318245 19715 318275
rect 19845 318245 19875 318275
rect 19685 318165 19715 318195
rect 19845 318165 19875 318195
rect 19685 318085 19715 318115
rect 19845 318085 19875 318115
rect 19685 318005 19715 318035
rect 19845 318005 19875 318035
rect 19685 317925 19715 317955
rect 19845 317925 19875 317955
rect 19685 317845 19715 317875
rect 19845 317845 19875 317875
rect 19685 317765 19715 317795
rect 19845 317765 19875 317795
rect 19685 317685 19715 317715
rect 19845 317685 19875 317715
rect 19685 317605 19715 317635
rect 19845 317605 19875 317635
rect 19685 317525 19715 317555
rect 19845 317525 19875 317555
rect 19685 317445 19715 317475
rect 19845 317445 19875 317475
rect 19685 317365 19715 317395
rect 19845 317365 19875 317395
rect 19685 317285 19715 317315
rect 19845 317285 19875 317315
rect 19685 317205 19715 317235
rect 19845 317205 19875 317235
rect 19685 317125 19715 317155
rect 19845 317125 19875 317155
rect 19685 317045 19715 317075
rect 19845 317045 19875 317075
rect 19685 316965 19715 316995
rect 19845 316965 19875 316995
rect 19685 316885 19715 316915
rect 19845 316885 19875 316915
rect 19685 316805 19715 316835
rect 19845 316805 19875 316835
rect 19685 316725 19715 316755
rect 19845 316725 19875 316755
rect 19685 316645 19715 316675
rect 19845 316645 19875 316675
rect 19685 316565 19715 316595
rect 19845 316565 19875 316595
rect 19685 316485 19715 316515
rect 19845 316485 19875 316515
rect 19685 316405 19715 316435
rect 19845 316405 19875 316435
rect 19685 316325 19715 316355
rect 19845 316325 19875 316355
rect 19685 316245 19715 316275
rect 19845 316245 19875 316275
rect 19685 316165 19715 316195
rect 19845 316165 19875 316195
rect 19685 316085 19715 316115
rect 19845 316085 19875 316115
rect 19685 316005 19715 316035
rect 19845 316005 19875 316035
rect 19685 315925 19715 315955
rect 19845 315925 19875 315955
rect 19685 315845 19715 315875
rect 19845 315845 19875 315875
rect 19685 315765 19715 315795
rect 19845 315765 19875 315795
rect 19685 315685 19715 315715
rect 19845 315685 19875 315715
rect 19685 315605 19715 315635
rect 19845 315605 19875 315635
rect 19685 315525 19715 315555
rect 19845 315525 19875 315555
rect 19685 315445 19715 315475
rect 19845 315445 19875 315475
rect 19685 315365 19715 315395
rect 19845 315365 19875 315395
rect 19685 315285 19715 315315
rect 19845 315285 19875 315315
rect 19685 315205 19715 315235
rect 19845 315205 19875 315235
rect 19685 315125 19715 315155
rect 19845 315125 19875 315155
rect 19685 315045 19715 315075
rect 19845 315045 19875 315075
rect 19685 314965 19715 314995
rect 19845 314965 19875 314995
rect 19685 314885 19715 314915
rect 19845 314885 19875 314915
rect 19685 314805 19715 314835
rect 19845 314805 19875 314835
rect 19685 314725 19715 314755
rect 19845 314725 19875 314755
rect 19685 314645 19715 314675
rect 19845 314645 19875 314675
rect 19685 314565 19715 314595
rect 19845 314565 19875 314595
rect 19685 314485 19715 314515
rect 19845 314485 19875 314515
rect 19685 314405 19715 314435
rect 19845 314405 19875 314435
rect 19685 314325 19715 314355
rect 19845 314325 19875 314355
rect 19685 314245 19715 314275
rect 19845 314245 19875 314275
rect 19685 314165 19715 314195
rect 19845 314165 19875 314195
rect 19685 314085 19715 314115
rect 19845 314085 19875 314115
rect 19685 314005 19715 314035
rect 19845 314005 19875 314035
rect 19685 313925 19715 313955
rect 19845 313925 19875 313955
rect 19685 313845 19715 313875
rect 19845 313845 19875 313875
rect 19685 313765 19715 313795
rect 19845 313765 19875 313795
rect 19685 313685 19715 313715
rect 19845 313685 19875 313715
rect 19685 313605 19715 313635
rect 19845 313605 19875 313635
rect 19685 313525 19715 313555
rect 19845 313525 19875 313555
rect 19685 313445 19715 313475
rect 19845 313445 19875 313475
rect 19685 313365 19715 313395
rect 19845 313365 19875 313395
rect 19685 313285 19715 313315
rect 19845 313285 19875 313315
rect 19685 313205 19715 313235
rect 19845 313205 19875 313235
rect 19685 313125 19715 313155
rect 19845 313125 19875 313155
rect 19685 313045 19715 313075
rect 19845 313045 19875 313075
rect 19685 312965 19715 312995
rect 19845 312965 19875 312995
rect 19685 312885 19715 312915
rect 19845 312885 19875 312915
rect 19685 312805 19715 312835
rect 19845 312805 19875 312835
rect 19685 312725 19715 312755
rect 19845 312725 19875 312755
rect 19685 312645 19715 312675
rect 19845 312645 19875 312675
rect 19685 312565 19715 312595
rect 19845 312565 19875 312595
rect 19685 312485 19715 312515
rect 19845 312485 19875 312515
rect 19685 312405 19715 312435
rect 19845 312405 19875 312435
rect 19685 312325 19715 312355
rect 19845 312325 19875 312355
rect 19685 312245 19715 312275
rect 19845 312245 19875 312275
rect 19685 312165 19715 312195
rect 19845 312165 19875 312195
rect 19685 312085 19715 312115
rect 19845 312085 19875 312115
rect 19685 312005 19715 312035
rect 19845 312005 19875 312035
rect 19685 311925 19715 311955
rect 19845 311925 19875 311955
rect 19685 311845 19715 311875
rect 19845 311845 19875 311875
rect 19685 311765 19715 311795
rect 19845 311765 19875 311795
rect 19685 311685 19715 311715
rect 19845 311685 19875 311715
rect 19685 311605 19715 311635
rect 19845 311605 19875 311635
rect 19685 311525 19715 311555
rect 19845 311525 19875 311555
rect 19685 311445 19715 311475
rect 19845 311445 19875 311475
rect 19685 311365 19715 311395
rect 19845 311365 19875 311395
rect 19685 311285 19715 311315
rect 19845 311285 19875 311315
rect 19685 311205 19715 311235
rect 19845 311205 19875 311235
rect 19685 311125 19715 311155
rect 19845 311125 19875 311155
rect 19685 311045 19715 311075
rect 19845 311045 19875 311075
rect 19685 310965 19715 310995
rect 19845 310965 19875 310995
rect 19685 310885 19715 310915
rect 19845 310885 19875 310915
rect 19685 310805 19715 310835
rect 19845 310805 19875 310835
rect 19685 310725 19715 310755
rect 19845 310725 19875 310755
rect 19685 310645 19715 310675
rect 19845 310645 19875 310675
rect 19685 310565 19715 310595
rect 19845 310565 19875 310595
rect 19685 310485 19715 310515
rect 19845 310485 19875 310515
rect 19685 310405 19715 310435
rect 19845 310405 19875 310435
rect 19685 310325 19715 310355
rect 19845 310325 19875 310355
rect 19685 310245 19715 310275
rect 19845 310245 19875 310275
rect 19685 310165 19715 310195
rect 19845 310165 19875 310195
rect 19685 310085 19715 310115
rect 19845 310085 19875 310115
rect 19685 310005 19715 310035
rect 19845 310005 19875 310035
rect 19685 309925 19715 309955
rect 19845 309925 19875 309955
rect 19685 309845 19715 309875
rect 19845 309845 19875 309875
rect 19685 309765 19715 309795
rect 19845 309765 19875 309795
rect 19685 309685 19715 309715
rect 19845 309685 19875 309715
rect 19685 309605 19715 309635
rect 19845 309605 19875 309635
rect 19685 309525 19715 309555
rect 19845 309525 19875 309555
rect 19685 309445 19715 309475
rect 19845 309445 19875 309475
rect 19685 309365 19715 309395
rect 19845 309365 19875 309395
rect 19685 309285 19715 309315
rect 19845 309285 19875 309315
rect 19685 309205 19715 309235
rect 19845 309205 19875 309235
rect 19685 309125 19715 309155
rect 19845 309125 19875 309155
rect 19685 309045 19715 309075
rect 19845 309045 19875 309075
rect 19685 308965 19715 308995
rect 19845 308965 19875 308995
rect 19685 308885 19715 308915
rect 19845 308885 19875 308915
rect 19685 308805 19715 308835
rect 19845 308805 19875 308835
rect 19685 308725 19715 308755
rect 19845 308725 19875 308755
rect 19685 308645 19715 308675
rect 19845 308645 19875 308675
rect 19685 308565 19715 308595
rect 19845 308565 19875 308595
rect 19685 308485 19715 308515
rect 19845 308485 19875 308515
rect 19685 308405 19715 308435
rect 19845 308405 19875 308435
rect 19685 308325 19715 308355
rect 19845 308325 19875 308355
rect 19685 308245 19715 308275
rect 19845 308245 19875 308275
rect 19685 308165 19715 308195
rect 19845 308165 19875 308195
rect 19685 308085 19715 308115
rect 19845 308085 19875 308115
rect 19685 308005 19715 308035
rect 19845 308005 19875 308035
rect 19685 307925 19715 307955
rect 19845 307925 19875 307955
rect 19685 307845 19715 307875
rect 19845 307845 19875 307875
rect 19685 307765 19715 307795
rect 19845 307765 19875 307795
rect 19685 307685 19715 307715
rect 19845 307685 19875 307715
rect 19685 307605 19715 307635
rect 19845 307605 19875 307635
rect 19685 307525 19715 307555
rect 19845 307525 19875 307555
rect 19685 307445 19715 307475
rect 19845 307445 19875 307475
rect 19685 307365 19715 307395
rect 19845 307365 19875 307395
rect 19685 307285 19715 307315
rect 19845 307285 19875 307315
rect 19685 307205 19715 307235
rect 19845 307205 19875 307235
rect 19685 307125 19715 307155
rect 19845 307125 19875 307155
rect 19685 307045 19715 307075
rect 19845 307045 19875 307075
rect 19685 306965 19715 306995
rect 19845 306965 19875 306995
rect 19685 306885 19715 306915
rect 19845 306885 19875 306915
rect 19685 306805 19715 306835
rect 19845 306805 19875 306835
rect 19685 306725 19715 306755
rect 19845 306725 19875 306755
rect 19685 306645 19715 306675
rect 19845 306645 19875 306675
rect 19685 306565 19715 306595
rect 19845 306565 19875 306595
rect 19685 306485 19715 306515
rect 19845 306485 19875 306515
rect 19685 306405 19715 306435
rect 19845 306405 19875 306435
rect 19685 306325 19715 306355
rect 19845 306325 19875 306355
rect 19685 306245 19715 306275
rect 19845 306245 19875 306275
rect 19685 306165 19715 306195
rect 19845 306165 19875 306195
rect 19685 306085 19715 306115
rect 19845 306085 19875 306115
rect 19685 306005 19715 306035
rect 19845 306005 19875 306035
rect 19685 305925 19715 305955
rect 19845 305925 19875 305955
rect 19685 305845 19715 305875
rect 19845 305845 19875 305875
rect 19685 305765 19715 305795
rect 19845 305765 19875 305795
rect 19685 305685 19715 305715
rect 19845 305685 19875 305715
rect 19685 305605 19715 305635
rect 19845 305605 19875 305635
rect 19685 305525 19715 305555
rect 19845 305525 19875 305555
rect 19685 305445 19715 305475
rect 19845 305445 19875 305475
rect 19685 305365 19715 305395
rect 19845 305365 19875 305395
rect 19685 305285 19715 305315
rect 19845 305285 19875 305315
rect 19685 305205 19715 305235
rect 19845 305205 19875 305235
rect 19685 305125 19715 305155
rect 19845 305125 19875 305155
rect 19685 305045 19715 305075
rect 19845 305045 19875 305075
rect 19685 304965 19715 304995
rect 19845 304965 19875 304995
rect 19685 304885 19715 304915
rect 19845 304885 19875 304915
rect 19685 304805 19715 304835
rect 19845 304805 19875 304835
rect 19685 304725 19715 304755
rect 19845 304725 19875 304755
rect 19685 304645 19715 304675
rect 19845 304645 19875 304675
rect 19685 304565 19715 304595
rect 19845 304565 19875 304595
rect 19685 304485 19715 304515
rect 19845 304485 19875 304515
rect 19685 304405 19715 304435
rect 19845 304405 19875 304435
rect 19685 304325 19715 304355
rect 19845 304325 19875 304355
rect 19685 304245 19715 304275
rect 19845 304245 19875 304275
rect 19685 304165 19715 304195
rect 19845 304165 19875 304195
rect 19685 304085 19715 304115
rect 19845 304085 19875 304115
rect 19685 304005 19715 304035
rect 19845 304005 19875 304035
rect 19685 303925 19715 303955
rect 19845 303925 19875 303955
rect 19685 303845 19715 303875
rect 19845 303845 19875 303875
rect 19685 303765 19715 303795
rect 19845 303765 19875 303795
rect 19685 303685 19715 303715
rect 19845 303685 19875 303715
rect 19685 303605 19715 303635
rect 19845 303605 19875 303635
rect 19685 303525 19715 303555
rect 19845 303525 19875 303555
rect 19685 303445 19715 303475
rect 19845 303445 19875 303475
rect 19685 303365 19715 303395
rect 19845 303365 19875 303395
rect 19685 303285 19715 303315
rect 19845 303285 19875 303315
rect 19685 303205 19715 303235
rect 19845 303205 19875 303235
rect 19685 303125 19715 303155
rect 19845 303125 19875 303155
rect 19685 303045 19715 303075
rect 19845 303045 19875 303075
rect 19685 302965 19715 302995
rect 19845 302965 19875 302995
rect 19685 302885 19715 302915
rect 19845 302885 19875 302915
rect 19685 302805 19715 302835
rect 19845 302805 19875 302835
rect 19685 302725 19715 302755
rect 19845 302725 19875 302755
rect 19685 302645 19715 302675
rect 19845 302645 19875 302675
rect 19685 302565 19715 302595
rect 19845 302565 19875 302595
rect 19685 302485 19715 302515
rect 19845 302485 19875 302515
rect 19685 302405 19715 302435
rect 19845 302405 19875 302435
rect 19685 302325 19715 302355
rect 19845 302325 19875 302355
rect 19685 302245 19715 302275
rect 19845 302245 19875 302275
rect 19685 302165 19715 302195
rect 19845 302165 19875 302195
rect 19685 302085 19715 302115
rect 19845 302085 19875 302115
rect 19685 302005 19715 302035
rect 19845 302005 19875 302035
rect 19685 301925 19715 301955
rect 19845 301925 19875 301955
rect 19685 301845 19715 301875
rect 19845 301845 19875 301875
rect 19685 301765 19715 301795
rect 19845 301765 19875 301795
rect 19685 301685 19715 301715
rect 19845 301685 19875 301715
rect 19685 301605 19715 301635
rect 19845 301605 19875 301635
rect 19685 301525 19715 301555
rect 19845 301525 19875 301555
rect 19685 301445 19715 301475
rect 19845 301445 19875 301475
rect 19685 301365 19715 301395
rect 19845 301365 19875 301395
rect 19685 301285 19715 301315
rect 19845 301285 19875 301315
rect 19685 301205 19715 301235
rect 19845 301205 19875 301235
rect 19685 301125 19715 301155
rect 19845 301125 19875 301155
rect 19685 301045 19715 301075
rect 19845 301045 19875 301075
rect 19685 300965 19715 300995
rect 19845 300965 19875 300995
rect 19685 300885 19715 300915
rect 19845 300885 19875 300915
rect 19685 300805 19715 300835
rect 19845 300805 19875 300835
rect 19685 300725 19715 300755
rect 19845 300725 19875 300755
rect 19685 300645 19715 300675
rect 19845 300645 19875 300675
rect 19685 300565 19715 300595
rect 19845 300565 19875 300595
rect 19685 300485 19715 300515
rect 19845 300485 19875 300515
rect 19685 300405 19715 300435
rect 19845 300405 19875 300435
rect 19685 300325 19715 300355
rect 19845 300325 19875 300355
rect 19685 300245 19715 300275
rect 19845 300245 19875 300275
rect 19685 300165 19715 300195
rect 19845 300165 19875 300195
rect 19685 300085 19715 300115
rect 19845 300085 19875 300115
rect 19685 300005 19715 300035
rect 19845 300005 19875 300035
rect 19685 299925 19715 299955
rect 19845 299925 19875 299955
rect 19685 299845 19715 299875
rect 19845 299845 19875 299875
rect 19685 299765 19715 299795
rect 19845 299765 19875 299795
rect 19685 299685 19715 299715
rect 19845 299685 19875 299715
rect 19685 299605 19715 299635
rect 19845 299605 19875 299635
rect 19685 299525 19715 299555
rect 19845 299525 19875 299555
rect 19685 299445 19715 299475
rect 19845 299445 19875 299475
rect 19685 299365 19715 299395
rect 19845 299365 19875 299395
rect 19685 299285 19715 299315
rect 19845 299285 19875 299315
rect 19685 299205 19715 299235
rect 19845 299205 19875 299235
rect 19685 299125 19715 299155
rect 19845 299125 19875 299155
rect 19685 299045 19715 299075
rect 19845 299045 19875 299075
rect 19685 298965 19715 298995
rect 19845 298965 19875 298995
rect 19685 298885 19715 298915
rect 19845 298885 19875 298915
rect 19685 298805 19715 298835
rect 19845 298805 19875 298835
rect 19685 298725 19715 298755
rect 19845 298725 19875 298755
rect 19685 298645 19715 298675
rect 19845 298645 19875 298675
rect 19685 298565 19715 298595
rect 19845 298565 19875 298595
rect 19685 298485 19715 298515
rect 19845 298485 19875 298515
rect 19685 298405 19715 298435
rect 19845 298405 19875 298435
rect 19685 298325 19715 298355
rect 19845 298325 19875 298355
rect 19685 298245 19715 298275
rect 19845 298245 19875 298275
rect 19685 298165 19715 298195
rect 19845 298165 19875 298195
rect 19685 298085 19715 298115
rect 19845 298085 19875 298115
rect 19685 298005 19715 298035
rect 19845 298005 19875 298035
rect 19685 297925 19715 297955
rect 19845 297925 19875 297955
rect 19685 297845 19715 297875
rect 19845 297845 19875 297875
rect 19685 297765 19715 297795
rect 19845 297765 19875 297795
rect 19685 297685 19715 297715
rect 19845 297685 19875 297715
rect 19685 297605 19715 297635
rect 19845 297605 19875 297635
rect 19685 297525 19715 297555
rect 19845 297525 19875 297555
rect 19685 297445 19715 297475
rect 19845 297445 19875 297475
rect 19685 297365 19715 297395
rect 19845 297365 19875 297395
rect 19685 297285 19715 297315
rect 19845 297285 19875 297315
rect 19685 297205 19715 297235
rect 19845 297205 19875 297235
rect 19685 297125 19715 297155
rect 19845 297125 19875 297155
rect 19685 297045 19715 297075
rect 19845 297045 19875 297075
rect 19685 296965 19715 296995
rect 19845 296965 19875 296995
rect 19685 296885 19715 296915
rect 19845 296885 19875 296915
rect 19685 296805 19715 296835
rect 19845 296805 19875 296835
rect 19685 296725 19715 296755
rect 19845 296725 19875 296755
rect 19685 296645 19715 296675
rect 19845 296645 19875 296675
rect 19685 296565 19715 296595
rect 19845 296565 19875 296595
rect 19685 296485 19715 296515
rect 19845 296485 19875 296515
rect 19685 296405 19715 296435
rect 19845 296405 19875 296435
rect 19685 296325 19715 296355
rect 19845 296325 19875 296355
rect 19685 296245 19715 296275
rect 19845 296245 19875 296275
rect 19685 296165 19715 296195
rect 19845 296165 19875 296195
rect 19685 296085 19715 296115
rect 19845 296085 19875 296115
rect 19685 296005 19715 296035
rect 19845 296005 19875 296035
rect 19685 295925 19715 295955
rect 19845 295925 19875 295955
rect 19685 295845 19715 295875
rect 19845 295845 19875 295875
rect 19685 295765 19715 295795
rect 19845 295765 19875 295795
rect 19685 295685 19715 295715
rect 19845 295685 19875 295715
rect 19685 295605 19715 295635
rect 19845 295605 19875 295635
rect 19685 295525 19715 295555
rect 19845 295525 19875 295555
rect 19685 295445 19715 295475
rect 19845 295445 19875 295475
rect 19685 295365 19715 295395
rect 19845 295365 19875 295395
rect 19685 295285 19715 295315
rect 19845 295285 19875 295315
rect 19685 295205 19715 295235
rect 19845 295205 19875 295235
rect 19685 295125 19715 295155
rect 19845 295125 19875 295155
rect 19685 295045 19715 295075
rect 19845 295045 19875 295075
rect 19685 294965 19715 294995
rect 19845 294965 19875 294995
rect 19685 294885 19715 294915
rect 19845 294885 19875 294915
rect 19685 294805 19715 294835
rect 19845 294805 19875 294835
rect 19685 294725 19715 294755
rect 19845 294725 19875 294755
rect 19685 294645 19715 294675
rect 19845 294645 19875 294675
rect 19685 294565 19715 294595
rect 19845 294565 19875 294595
rect 19685 294485 19715 294515
rect 19845 294485 19875 294515
rect 19685 294405 19715 294435
rect 19845 294405 19875 294435
rect 19685 294325 19715 294355
rect 19845 294325 19875 294355
rect 19685 294245 19715 294275
rect 19845 294245 19875 294275
rect 19685 294165 19715 294195
rect 19845 294165 19875 294195
rect 19685 294085 19715 294115
rect 19845 294085 19875 294115
rect 19685 294005 19715 294035
rect 19845 294005 19875 294035
rect 19685 293925 19715 293955
rect 19845 293925 19875 293955
rect 19685 293845 19715 293875
rect 19845 293845 19875 293875
rect 19685 293765 19715 293795
rect 19845 293765 19875 293795
rect 19685 293685 19715 293715
rect 19845 293685 19875 293715
rect 19685 293605 19715 293635
rect 19845 293605 19875 293635
rect 19685 293525 19715 293555
rect 19845 293525 19875 293555
rect 19685 293445 19715 293475
rect 19845 293445 19875 293475
rect 19685 293365 19715 293395
rect 19845 293365 19875 293395
rect 19685 293285 19715 293315
rect 19845 293285 19875 293315
rect 19685 293205 19715 293235
rect 19845 293205 19875 293235
rect 19685 293125 19715 293155
rect 19845 293125 19875 293155
rect 19685 293045 19715 293075
rect 19845 293045 19875 293075
rect 19685 292965 19715 292995
rect 19845 292965 19875 292995
rect 19685 292885 19715 292915
rect 19845 292885 19875 292915
rect 19685 292805 19715 292835
rect 19845 292805 19875 292835
rect 19685 292725 19715 292755
rect 19845 292725 19875 292755
rect 19685 292645 19715 292675
rect 19845 292645 19875 292675
rect 19685 292565 19715 292595
rect 19845 292565 19875 292595
rect 19685 292485 19715 292515
rect 19845 292485 19875 292515
rect 19685 292405 19715 292435
rect 19845 292405 19875 292435
rect 19685 292325 19715 292355
rect 19845 292325 19875 292355
rect 19685 292245 19715 292275
rect 19845 292245 19875 292275
rect 19685 292165 19715 292195
rect 19845 292165 19875 292195
rect 19685 292085 19715 292115
rect 19845 292085 19875 292115
rect 19685 292005 19715 292035
rect 19845 292005 19875 292035
rect 19685 291925 19715 291955
rect 19845 291925 19875 291955
rect 19685 291845 19715 291875
rect 19845 291845 19875 291875
rect 19685 291765 19715 291795
rect 19845 291765 19875 291795
rect 19685 291685 19715 291715
rect 19845 291685 19875 291715
rect 19685 291605 19715 291635
rect 19845 291605 19875 291635
rect 19685 291525 19715 291555
rect 19845 291525 19875 291555
rect 19685 291445 19715 291475
rect 19845 291445 19875 291475
rect 19685 291365 19715 291395
rect 19845 291365 19875 291395
rect 19685 291285 19715 291315
rect 19845 291285 19875 291315
rect 19685 291205 19715 291235
rect 19845 291205 19875 291235
rect 19685 291125 19715 291155
rect 19845 291125 19875 291155
rect 19685 291045 19715 291075
rect 19845 291045 19875 291075
rect 19685 290965 19715 290995
rect 19845 290965 19875 290995
rect 19685 290885 19715 290915
rect 19845 290885 19875 290915
rect 19685 290805 19715 290835
rect 19845 290805 19875 290835
rect 19685 290725 19715 290755
rect 19845 290725 19875 290755
rect 19685 290645 19715 290675
rect 19845 290645 19875 290675
rect 19685 290565 19715 290595
rect 19845 290565 19875 290595
rect 19685 290485 19715 290515
rect 19845 290485 19875 290515
rect 19685 290405 19715 290435
rect 19845 290405 19875 290435
rect 19685 290325 19715 290355
rect 19845 290325 19875 290355
rect 19685 290245 19715 290275
rect 19845 290245 19875 290275
rect 19685 290165 19715 290195
rect 19845 290165 19875 290195
rect 19685 290085 19715 290115
rect 19845 290085 19875 290115
rect 19685 290005 19715 290035
rect 19845 290005 19875 290035
rect 19685 289925 19715 289955
rect 19845 289925 19875 289955
rect 19685 289845 19715 289875
rect 19845 289845 19875 289875
rect 19685 289765 19715 289795
rect 19845 289765 19875 289795
rect 19685 289685 19715 289715
rect 19845 289685 19875 289715
rect 19685 289605 19715 289635
rect 19845 289605 19875 289635
rect 19685 289525 19715 289555
rect 19845 289525 19875 289555
rect 19685 289445 19715 289475
rect 19845 289445 19875 289475
rect 19685 289365 19715 289395
rect 19845 289365 19875 289395
rect 19685 289285 19715 289315
rect 19845 289285 19875 289315
rect 19685 289205 19715 289235
rect 19845 289205 19875 289235
rect 19685 289125 19715 289155
rect 19845 289125 19875 289155
rect 19685 289045 19715 289075
rect 19845 289045 19875 289075
rect 19685 288965 19715 288995
rect 19845 288965 19875 288995
rect 19685 288885 19715 288915
rect 19845 288885 19875 288915
rect 19685 288805 19715 288835
rect 19845 288805 19875 288835
rect 19685 288725 19715 288755
rect 19845 288725 19875 288755
rect 19685 288645 19715 288675
rect 19845 288645 19875 288675
rect 19685 288565 19715 288595
rect 19845 288565 19875 288595
rect 19685 288485 19715 288515
rect 19845 288485 19875 288515
rect 19685 288405 19715 288435
rect 19845 288405 19875 288435
rect 19685 288325 19715 288355
rect 19845 288325 19875 288355
rect 19685 288245 19715 288275
rect 19845 288245 19875 288275
rect 19685 288165 19715 288195
rect 19845 288165 19875 288195
rect 19685 288085 19715 288115
rect 19845 288085 19875 288115
rect 19685 288005 19715 288035
rect 19845 288005 19875 288035
rect 19685 287925 19715 287955
rect 19845 287925 19875 287955
rect 19685 287845 19715 287875
rect 19845 287845 19875 287875
rect 19685 287765 19715 287795
rect 19845 287765 19875 287795
rect 19685 287685 19715 287715
rect 19845 287685 19875 287715
rect 19685 287605 19715 287635
rect 19845 287605 19875 287635
rect 19685 287525 19715 287555
rect 19845 287525 19875 287555
rect 19685 287445 19715 287475
rect 19845 287445 19875 287475
rect 19685 287365 19715 287395
rect 19845 287365 19875 287395
rect 19685 287285 19715 287315
rect 19845 287285 19875 287315
rect 19685 287205 19715 287235
rect 19845 287205 19875 287235
rect 19685 287125 19715 287155
rect 19845 287125 19875 287155
rect 19685 287045 19715 287075
rect 19845 287045 19875 287075
rect 19685 286965 19715 286995
rect 19845 286965 19875 286995
rect 19685 286885 19715 286915
rect 19845 286885 19875 286915
rect 19685 286805 19715 286835
rect 19845 286805 19875 286835
rect 19685 286725 19715 286755
rect 19845 286725 19875 286755
rect 19685 286645 19715 286675
rect 19845 286645 19875 286675
rect 19685 286565 19715 286595
rect 19845 286565 19875 286595
rect 19685 286485 19715 286515
rect 19845 286485 19875 286515
rect 19685 286405 19715 286435
rect 19845 286405 19875 286435
rect 19685 286325 19715 286355
rect 19845 286325 19875 286355
rect 19685 286245 19715 286275
rect 19845 286245 19875 286275
rect 19685 286165 19715 286195
rect 19845 286165 19875 286195
rect 19685 286085 19715 286115
rect 19845 286085 19875 286115
rect 19685 286005 19715 286035
rect 19845 286005 19875 286035
rect 19685 285925 19715 285955
rect 19845 285925 19875 285955
rect 19685 285845 19715 285875
rect 19845 285845 19875 285875
rect 19685 285765 19715 285795
rect 19845 285765 19875 285795
rect 19685 285685 19715 285715
rect 19845 285685 19875 285715
rect 19685 285605 19715 285635
rect 19845 285605 19875 285635
rect 19685 285525 19715 285555
rect 19845 285525 19875 285555
rect 19685 285445 19715 285475
rect 19845 285445 19875 285475
rect 19685 285365 19715 285395
rect 19845 285365 19875 285395
rect 19685 285285 19715 285315
rect 19845 285285 19875 285315
rect 19685 285205 19715 285235
rect 19845 285205 19875 285235
rect 19685 285125 19715 285155
rect 19845 285125 19875 285155
rect 19685 285045 19715 285075
rect 19845 285045 19875 285075
rect 19685 284965 19715 284995
rect 19845 284965 19875 284995
rect 19685 284885 19715 284915
rect 19845 284885 19875 284915
rect 19685 284805 19715 284835
rect 19845 284805 19875 284835
rect 19685 284725 19715 284755
rect 19845 284725 19875 284755
rect 19685 284645 19715 284675
rect 19845 284645 19875 284675
rect 19685 284565 19715 284595
rect 19845 284565 19875 284595
rect 19685 284485 19715 284515
rect 19845 284485 19875 284515
rect 19685 284405 19715 284435
rect 19845 284405 19875 284435
rect 19685 284325 19715 284355
rect 19845 284325 19875 284355
rect 19685 284245 19715 284275
rect 19845 284245 19875 284275
rect 19685 284165 19715 284195
rect 19845 284165 19875 284195
rect 19685 284085 19715 284115
rect 19845 284085 19875 284115
rect 19685 284005 19715 284035
rect 19845 284005 19875 284035
rect 19685 283925 19715 283955
rect 19845 283925 19875 283955
rect 19685 283845 19715 283875
rect 19845 283845 19875 283875
rect 19685 283765 19715 283795
rect 19845 283765 19875 283795
rect 19685 283685 19715 283715
rect 19845 283685 19875 283715
rect 19685 283605 19715 283635
rect 19845 283605 19875 283635
rect 19685 283525 19715 283555
rect 19845 283525 19875 283555
rect 19685 283445 19715 283475
rect 19845 283445 19875 283475
rect 19685 283365 19715 283395
rect 19845 283365 19875 283395
rect 19685 283285 19715 283315
rect 19845 283285 19875 283315
rect 19685 283205 19715 283235
rect 19845 283205 19875 283235
rect 19685 283125 19715 283155
rect 19845 283125 19875 283155
rect 19685 283045 19715 283075
rect 19845 283045 19875 283075
rect 19685 282965 19715 282995
rect 19845 282965 19875 282995
rect 19685 282885 19715 282915
rect 19845 282885 19875 282915
rect 19685 282805 19715 282835
rect 19845 282805 19875 282835
rect 19685 282725 19715 282755
rect 19845 282725 19875 282755
rect 19685 282645 19715 282675
rect 19845 282645 19875 282675
rect 19685 282565 19715 282595
rect 19845 282565 19875 282595
rect 19685 282485 19715 282515
rect 19845 282485 19875 282515
rect 19685 282405 19715 282435
rect 19845 282405 19875 282435
rect 19685 282325 19715 282355
rect 19845 282325 19875 282355
rect 19685 282245 19715 282275
rect 19845 282245 19875 282275
rect 19685 282165 19715 282195
rect 19845 282165 19875 282195
rect 19685 282085 19715 282115
rect 19845 282085 19875 282115
rect 19685 282005 19715 282035
rect 19845 282005 19875 282035
rect 19685 281925 19715 281955
rect 19845 281925 19875 281955
rect 19685 281845 19715 281875
rect 19845 281845 19875 281875
rect 19685 281765 19715 281795
rect 19845 281765 19875 281795
rect 19685 281685 19715 281715
rect 19845 281685 19875 281715
rect 19685 281605 19715 281635
rect 19845 281605 19875 281635
rect 19685 281525 19715 281555
rect 19845 281525 19875 281555
rect 19685 281445 19715 281475
rect 19845 281445 19875 281475
rect 19685 281365 19715 281395
rect 19845 281365 19875 281395
rect 19685 281285 19715 281315
rect 19845 281285 19875 281315
rect 19685 281205 19715 281235
rect 19845 281205 19875 281235
rect 19685 281125 19715 281155
rect 19845 281125 19875 281155
rect 19685 281045 19715 281075
rect 19845 281045 19875 281075
rect 19685 280965 19715 280995
rect 19845 280965 19875 280995
rect 19685 280885 19715 280915
rect 19845 280885 19875 280915
rect 19685 280805 19715 280835
rect 19845 280805 19875 280835
rect 19685 280725 19715 280755
rect 19845 280725 19875 280755
rect 19685 280645 19715 280675
rect 19845 280645 19875 280675
rect 19685 280565 19715 280595
rect 19845 280565 19875 280595
rect 19685 280485 19715 280515
rect 19845 280485 19875 280515
rect 19685 280405 19715 280435
rect 19845 280405 19875 280435
rect 19685 280325 19715 280355
rect 19845 280325 19875 280355
rect 19685 280245 19715 280275
rect 19845 280245 19875 280275
rect 19685 280165 19715 280195
rect 19845 280165 19875 280195
rect 19685 280085 19715 280115
rect 19845 280085 19875 280115
rect 19685 280005 19715 280035
rect 19845 280005 19875 280035
rect 19685 279925 19715 279955
rect 19845 279925 19875 279955
rect 19685 279845 19715 279875
rect 19845 279845 19875 279875
rect 19685 279765 19715 279795
rect 19845 279765 19875 279795
rect 19685 279685 19715 279715
rect 19845 279685 19875 279715
rect 19685 279605 19715 279635
rect 19845 279605 19875 279635
rect 19685 279525 19715 279555
rect 19845 279525 19875 279555
rect 19685 279445 19715 279475
rect 19845 279445 19875 279475
rect 19685 279365 19715 279395
rect 19845 279365 19875 279395
rect 19685 279285 19715 279315
rect 19845 279285 19875 279315
rect 19685 279205 19715 279235
rect 19845 279205 19875 279235
rect 19685 279125 19715 279155
rect 19845 279125 19875 279155
rect 19685 279045 19715 279075
rect 19845 279045 19875 279075
rect 19685 278965 19715 278995
rect 19845 278965 19875 278995
rect 19685 278885 19715 278915
rect 19845 278885 19875 278915
rect 19685 278805 19715 278835
rect 19845 278805 19875 278835
rect 19685 278725 19715 278755
rect 19845 278725 19875 278755
rect 17045 278645 17075 278675
rect 17205 278645 17235 278675
rect 17285 278645 17315 278675
rect 17365 278645 17395 278675
rect 17445 278645 17475 278675
rect 17525 278645 17555 278675
rect 17605 278645 17635 278675
rect 17685 278645 17715 278675
rect 17765 278645 17795 278675
rect 19525 278645 19555 278675
rect 19605 278645 19635 278675
rect 19685 278645 19715 278675
rect 19845 278645 19875 278675
rect 17125 278565 17155 278595
rect 19765 278565 19795 278595
rect 17045 278485 17075 278515
rect 17205 278485 17235 278515
rect 17285 278485 17315 278515
rect 17365 278485 17395 278515
rect 17445 278485 17475 278515
rect 17525 278485 17555 278515
rect 17605 278485 17635 278515
rect 17685 278485 17715 278515
rect 17765 278485 17795 278515
rect 19525 278485 19555 278515
rect 19605 278485 19635 278515
rect 19685 278485 19715 278515
rect 19845 278485 19875 278515
rect 17045 278405 17075 278435
rect 17205 278405 17235 278435
rect 17045 278325 17075 278355
rect 17205 278325 17235 278355
rect 17045 278245 17075 278275
rect 17205 278245 17235 278275
rect 17045 278165 17075 278195
rect 17205 278165 17235 278195
rect 17045 278085 17075 278115
rect 17205 278085 17235 278115
rect 17045 278005 17075 278035
rect 17205 278005 17235 278035
rect 17045 277925 17075 277955
rect 17205 277925 17235 277955
rect 17045 277845 17075 277875
rect 17205 277845 17235 277875
rect 28405 275325 28435 275355
rect 28565 275325 28595 275355
rect 28725 275325 28755 275355
rect 28405 275245 28435 275275
rect 28565 275245 28595 275275
rect 28725 275245 28755 275275
rect 1040 275040 1160 275160
rect 13525 275005 13555 275195
rect 13685 275005 13715 275195
rect 13845 275005 13875 275195
rect 14005 275005 14035 275195
rect 14165 275005 14195 275195
rect 14325 275005 14355 275195
rect 27925 275005 27955 275195
rect 28085 275005 28115 275195
rect 28245 275005 28275 275195
rect 28405 275005 28435 275195
rect 28565 275005 28595 275195
rect 28725 275005 28755 275195
<< metal3 >>
rect 8097 351400 10597 352400
rect 8097 351320 10600 351400
rect 10720 351396 10760 351400
rect 10720 351364 10724 351396
rect 10756 351364 10760 351396
rect 8097 351315 10680 351320
rect 8097 351285 10645 351315
rect 10675 351285 10680 351315
rect 8097 351280 10680 351285
rect 10720 351316 10760 351364
rect 10720 351284 10724 351316
rect 10756 351284 10760 351316
rect 8097 351200 10600 351280
rect 10720 351236 10760 351284
rect 10720 351204 10724 351236
rect 10756 351204 10760 351236
rect 10720 351200 10760 351204
rect 10800 351396 10840 351400
rect 10800 351364 10804 351396
rect 10836 351364 10840 351396
rect 10800 351316 10840 351364
rect 10800 351284 10804 351316
rect 10836 351284 10840 351316
rect 10800 351236 10840 351284
rect 10800 351204 10804 351236
rect 10836 351204 10840 351236
rect 10800 351200 10840 351204
rect 10880 351396 10920 351400
rect 10880 351364 10884 351396
rect 10916 351364 10920 351396
rect 10880 351316 10920 351364
rect 10880 351284 10884 351316
rect 10916 351284 10920 351316
rect 10880 351236 10920 351284
rect 10880 351204 10884 351236
rect 10916 351204 10920 351236
rect 10880 351200 10920 351204
rect 10960 351396 11000 351400
rect 10960 351364 10964 351396
rect 10996 351364 11000 351396
rect 10960 351316 11000 351364
rect 10960 351284 10964 351316
rect 10996 351284 11000 351316
rect 10960 351236 11000 351284
rect 10960 351204 10964 351236
rect 10996 351204 11000 351236
rect 10960 351200 11000 351204
rect 11040 351396 11080 351400
rect 11040 351364 11044 351396
rect 11076 351364 11080 351396
rect 11040 351316 11080 351364
rect 11040 351284 11044 351316
rect 11076 351284 11080 351316
rect 11040 351236 11080 351284
rect 11040 351204 11044 351236
rect 11076 351204 11080 351236
rect 11040 351200 11080 351204
rect 11120 351396 11160 351400
rect 11120 351364 11124 351396
rect 11156 351364 11160 351396
rect 11120 351316 11160 351364
rect 11120 351284 11124 351316
rect 11156 351284 11160 351316
rect 11120 351236 11160 351284
rect 11120 351204 11124 351236
rect 11156 351204 11160 351236
rect 11120 351200 11160 351204
rect 11200 351396 11240 351400
rect 11200 351364 11204 351396
rect 11236 351364 11240 351396
rect 11200 351316 11240 351364
rect 11200 351284 11204 351316
rect 11236 351284 11240 351316
rect 11200 351236 11240 351284
rect 11200 351204 11204 351236
rect 11236 351204 11240 351236
rect 11200 351200 11240 351204
rect 11280 351396 11320 351400
rect 11280 351364 11284 351396
rect 11316 351364 11320 351396
rect 11280 351316 11320 351364
rect 11280 351284 11284 351316
rect 11316 351284 11320 351316
rect 11280 351236 11320 351284
rect 11280 351204 11284 351236
rect 11316 351204 11320 351236
rect 11280 351200 11320 351204
rect 11360 351396 11400 351400
rect 11360 351364 11364 351396
rect 11396 351364 11400 351396
rect 11360 351316 11400 351364
rect 11360 351284 11364 351316
rect 11396 351284 11400 351316
rect 11360 351236 11400 351284
rect 11360 351204 11364 351236
rect 11396 351204 11400 351236
rect 11360 351200 11400 351204
rect 11440 351396 11480 351400
rect 11440 351364 11444 351396
rect 11476 351364 11480 351396
rect 11440 351316 11480 351364
rect 11440 351284 11444 351316
rect 11476 351284 11480 351316
rect 11440 351236 11480 351284
rect 11440 351204 11444 351236
rect 11476 351204 11480 351236
rect 11440 351200 11480 351204
rect 11520 351396 11560 351400
rect 11520 351364 11524 351396
rect 11556 351364 11560 351396
rect 11520 351316 11560 351364
rect 11520 351284 11524 351316
rect 11556 351284 11560 351316
rect 11520 351236 11560 351284
rect 11520 351204 11524 351236
rect 11556 351204 11560 351236
rect 11520 351200 11560 351204
rect 11600 351396 11640 351400
rect 11600 351364 11604 351396
rect 11636 351364 11640 351396
rect 11600 351316 11640 351364
rect 11600 351284 11604 351316
rect 11636 351284 11640 351316
rect 11600 351236 11640 351284
rect 11600 351204 11604 351236
rect 11636 351204 11640 351236
rect 11600 351200 11640 351204
rect 11680 351396 11720 351400
rect 11680 351364 11684 351396
rect 11716 351364 11720 351396
rect 11680 351316 11720 351364
rect 11680 351284 11684 351316
rect 11716 351284 11720 351316
rect 11680 351236 11720 351284
rect 11680 351204 11684 351236
rect 11716 351204 11720 351236
rect 11680 351200 11720 351204
rect 11760 351396 11800 351400
rect 11760 351364 11764 351396
rect 11796 351364 11800 351396
rect 11760 351316 11800 351364
rect 11760 351284 11764 351316
rect 11796 351284 11800 351316
rect 11760 351236 11800 351284
rect 11760 351204 11764 351236
rect 11796 351204 11800 351236
rect 11760 351200 11800 351204
rect 11840 351396 11880 351400
rect 11840 351364 11844 351396
rect 11876 351364 11880 351396
rect 11840 351316 11880 351364
rect 11840 351284 11844 351316
rect 11876 351284 11880 351316
rect 11840 351236 11880 351284
rect 11840 351204 11844 351236
rect 11876 351204 11880 351236
rect 11840 351200 11880 351204
rect 11920 351396 11960 351400
rect 11920 351364 11924 351396
rect 11956 351364 11960 351396
rect 11920 351316 11960 351364
rect 11920 351284 11924 351316
rect 11956 351284 11960 351316
rect 11920 351236 11960 351284
rect 11920 351204 11924 351236
rect 11956 351204 11960 351236
rect 11920 351200 11960 351204
rect 12000 351396 12040 351400
rect 12000 351364 12004 351396
rect 12036 351364 12040 351396
rect 12000 351316 12040 351364
rect 12000 351284 12004 351316
rect 12036 351284 12040 351316
rect 12000 351236 12040 351284
rect 12000 351204 12004 351236
rect 12036 351204 12040 351236
rect 12000 351200 12040 351204
rect 12080 351396 12120 351400
rect 12080 351364 12084 351396
rect 12116 351364 12120 351396
rect 12080 351316 12120 351364
rect 12080 351284 12084 351316
rect 12116 351284 12120 351316
rect 12080 351236 12120 351284
rect 12080 351204 12084 351236
rect 12116 351204 12120 351236
rect 12080 351200 12120 351204
rect 12160 351396 12200 351400
rect 12160 351364 12164 351396
rect 12196 351364 12200 351396
rect 12160 351316 12200 351364
rect 12160 351284 12164 351316
rect 12196 351284 12200 351316
rect 12160 351236 12200 351284
rect 12160 351204 12164 351236
rect 12196 351204 12200 351236
rect 12160 351200 12200 351204
rect 12240 351396 12280 351400
rect 12240 351364 12244 351396
rect 12276 351364 12280 351396
rect 12240 351316 12280 351364
rect 12240 351284 12244 351316
rect 12276 351284 12280 351316
rect 12240 351236 12280 351284
rect 12240 351204 12244 351236
rect 12276 351204 12280 351236
rect 12240 351200 12280 351204
rect 12320 351396 12360 351400
rect 12320 351364 12324 351396
rect 12356 351364 12360 351396
rect 12320 351316 12360 351364
rect 12320 351284 12324 351316
rect 12356 351284 12360 351316
rect 12320 351236 12360 351284
rect 12320 351204 12324 351236
rect 12356 351204 12360 351236
rect 12320 351200 12360 351204
rect 12400 351396 12440 351400
rect 12400 351364 12404 351396
rect 12436 351364 12440 351396
rect 12400 351316 12440 351364
rect 12400 351284 12404 351316
rect 12436 351284 12440 351316
rect 12400 351236 12440 351284
rect 12400 351204 12404 351236
rect 12436 351204 12440 351236
rect 12400 351200 12440 351204
rect 12480 351396 12520 351400
rect 12480 351364 12484 351396
rect 12516 351364 12520 351396
rect 12480 351316 12520 351364
rect 12480 351284 12484 351316
rect 12516 351284 12520 351316
rect 12480 351236 12520 351284
rect 12480 351204 12484 351236
rect 12516 351204 12520 351236
rect 12480 351200 12520 351204
rect 12560 351396 12600 351400
rect 12560 351364 12564 351396
rect 12596 351364 12600 351396
rect 12560 351316 12600 351364
rect 12560 351284 12564 351316
rect 12596 351284 12600 351316
rect 12560 351236 12600 351284
rect 12560 351204 12564 351236
rect 12596 351204 12600 351236
rect 12560 351200 12600 351204
rect 12640 351396 12680 351400
rect 12640 351364 12644 351396
rect 12676 351364 12680 351396
rect 12640 351316 12680 351364
rect 12640 351284 12644 351316
rect 12676 351284 12680 351316
rect 12640 351236 12680 351284
rect 12640 351204 12644 351236
rect 12676 351204 12680 351236
rect 12640 351200 12680 351204
rect 12720 351396 12760 351400
rect 12720 351364 12724 351396
rect 12756 351364 12760 351396
rect 12720 351316 12760 351364
rect 12720 351284 12724 351316
rect 12756 351284 12760 351316
rect 12720 351236 12760 351284
rect 12720 351204 12724 351236
rect 12756 351204 12760 351236
rect 12720 351200 12760 351204
rect 12800 351396 12840 351400
rect 12800 351364 12804 351396
rect 12836 351364 12840 351396
rect 12800 351316 12840 351364
rect 12800 351284 12804 351316
rect 12836 351284 12840 351316
rect 12800 351236 12840 351284
rect 12800 351204 12804 351236
rect 12836 351204 12840 351236
rect 12800 351200 12840 351204
rect 12880 351396 12920 351400
rect 12880 351364 12884 351396
rect 12916 351364 12920 351396
rect 12880 351316 12920 351364
rect 12880 351284 12884 351316
rect 12916 351284 12920 351316
rect 12880 351236 12920 351284
rect 12880 351204 12884 351236
rect 12916 351204 12920 351236
rect 12880 351200 12920 351204
rect 12960 351396 13000 351400
rect 12960 351364 12964 351396
rect 12996 351364 13000 351396
rect 12960 351316 13000 351364
rect 12960 351284 12964 351316
rect 12996 351284 13000 351316
rect 12960 351236 13000 351284
rect 12960 351204 12964 351236
rect 12996 351204 13000 351236
rect 12960 351200 13000 351204
rect 13040 351396 13080 351400
rect 13040 351364 13044 351396
rect 13076 351364 13080 351396
rect 13040 351316 13080 351364
rect 13040 351284 13044 351316
rect 13076 351284 13080 351316
rect 13040 351236 13080 351284
rect 13040 351204 13044 351236
rect 13076 351204 13080 351236
rect 13040 351200 13080 351204
rect 13120 351396 13160 351400
rect 13120 351364 13124 351396
rect 13156 351364 13160 351396
rect 13120 351316 13160 351364
rect 13120 351284 13124 351316
rect 13156 351284 13160 351316
rect 13120 351236 13160 351284
rect 13120 351204 13124 351236
rect 13156 351204 13160 351236
rect 13120 351200 13160 351204
rect 13200 351396 13240 351400
rect 13200 351364 13204 351396
rect 13236 351364 13240 351396
rect 13200 351316 13240 351364
rect 13200 351284 13204 351316
rect 13236 351284 13240 351316
rect 13200 351236 13240 351284
rect 13200 351204 13204 351236
rect 13236 351204 13240 351236
rect 13200 351200 13240 351204
rect 13280 351396 13320 351400
rect 13280 351364 13284 351396
rect 13316 351364 13320 351396
rect 13280 351316 13320 351364
rect 13280 351284 13284 351316
rect 13316 351284 13320 351316
rect 13280 351236 13320 351284
rect 13280 351204 13284 351236
rect 13316 351204 13320 351236
rect 13280 351200 13320 351204
rect 13360 351396 13400 351400
rect 13360 351364 13364 351396
rect 13396 351364 13400 351396
rect 13360 351316 13400 351364
rect 13360 351284 13364 351316
rect 13396 351284 13400 351316
rect 13360 351236 13400 351284
rect 13360 351204 13364 351236
rect 13396 351204 13400 351236
rect 13360 351200 13400 351204
rect 13440 351396 13480 351400
rect 13440 351364 13444 351396
rect 13476 351364 13480 351396
rect 13440 351316 13480 351364
rect 13440 351284 13444 351316
rect 13476 351284 13480 351316
rect 13440 351236 13480 351284
rect 13440 351204 13444 351236
rect 13476 351204 13480 351236
rect 13440 351200 13480 351204
rect 13520 351396 13560 351400
rect 13520 351364 13524 351396
rect 13556 351364 13560 351396
rect 13520 351316 13560 351364
rect 13520 351284 13524 351316
rect 13556 351284 13560 351316
rect 13520 351236 13560 351284
rect 13520 351204 13524 351236
rect 13556 351204 13560 351236
rect 13520 351200 13560 351204
rect 13600 351396 13640 351400
rect 13600 351364 13604 351396
rect 13636 351364 13640 351396
rect 13600 351316 13640 351364
rect 13600 351284 13604 351316
rect 13636 351284 13640 351316
rect 13600 351236 13640 351284
rect 13600 351204 13604 351236
rect 13636 351204 13640 351236
rect 13600 351200 13640 351204
rect 13680 351396 13720 351400
rect 13680 351364 13684 351396
rect 13716 351364 13720 351396
rect 13680 351316 13720 351364
rect 13680 351284 13684 351316
rect 13716 351284 13720 351316
rect 13680 351236 13720 351284
rect 13680 351204 13684 351236
rect 13716 351204 13720 351236
rect 13680 351200 13720 351204
rect 13760 351396 13800 351400
rect 13760 351364 13764 351396
rect 13796 351364 13800 351396
rect 13760 351316 13800 351364
rect 13760 351284 13764 351316
rect 13796 351284 13800 351316
rect 13760 351236 13800 351284
rect 13760 351204 13764 351236
rect 13796 351204 13800 351236
rect 13760 351200 13800 351204
rect 13840 351396 13880 351400
rect 13840 351364 13844 351396
rect 13876 351364 13880 351396
rect 13840 351316 13880 351364
rect 13840 351284 13844 351316
rect 13876 351284 13880 351316
rect 13840 351236 13880 351284
rect 13840 351204 13844 351236
rect 13876 351204 13880 351236
rect 13840 351200 13880 351204
rect 13920 351396 13960 351400
rect 13920 351364 13924 351396
rect 13956 351364 13960 351396
rect 13920 351316 13960 351364
rect 13920 351284 13924 351316
rect 13956 351284 13960 351316
rect 13920 351236 13960 351284
rect 13920 351204 13924 351236
rect 13956 351204 13960 351236
rect 13920 351200 13960 351204
rect 14000 351396 14040 351400
rect 14000 351364 14004 351396
rect 14036 351364 14040 351396
rect 14000 351316 14040 351364
rect 14000 351284 14004 351316
rect 14036 351284 14040 351316
rect 14000 351236 14040 351284
rect 14000 351204 14004 351236
rect 14036 351204 14040 351236
rect 14000 351200 14040 351204
rect 14080 351396 14120 351400
rect 14080 351364 14084 351396
rect 14116 351364 14120 351396
rect 14080 351316 14120 351364
rect 14080 351284 14084 351316
rect 14116 351284 14120 351316
rect 14080 351236 14120 351284
rect 14080 351204 14084 351236
rect 14116 351204 14120 351236
rect 14080 351200 14120 351204
rect 14160 351396 14200 351400
rect 14160 351364 14164 351396
rect 14196 351364 14200 351396
rect 14160 351316 14200 351364
rect 14160 351284 14164 351316
rect 14196 351284 14200 351316
rect 14160 351236 14200 351284
rect 14160 351204 14164 351236
rect 14196 351204 14200 351236
rect 14160 351200 14200 351204
rect 14240 351396 14280 351400
rect 14240 351364 14244 351396
rect 14276 351364 14280 351396
rect 14240 351316 14280 351364
rect 14240 351284 14244 351316
rect 14276 351284 14280 351316
rect 14240 351236 14280 351284
rect 14240 351204 14244 351236
rect 14276 351204 14280 351236
rect 14240 351200 14280 351204
rect 14320 351396 14360 351400
rect 14320 351364 14324 351396
rect 14356 351364 14360 351396
rect 14320 351316 14360 351364
rect 14320 351284 14324 351316
rect 14356 351284 14360 351316
rect 14320 351236 14360 351284
rect 14320 351204 14324 351236
rect 14356 351204 14360 351236
rect 14320 351200 14360 351204
rect 14400 351396 14440 351400
rect 14400 351364 14404 351396
rect 14436 351364 14440 351396
rect 14400 351316 14440 351364
rect 14400 351284 14404 351316
rect 14436 351284 14440 351316
rect 14400 351236 14440 351284
rect 14400 351204 14404 351236
rect 14436 351204 14440 351236
rect 14400 351200 14440 351204
rect 14480 351396 14520 351400
rect 14480 351364 14484 351396
rect 14516 351364 14520 351396
rect 14480 351316 14520 351364
rect 14480 351284 14484 351316
rect 14516 351284 14520 351316
rect 14480 351236 14520 351284
rect 14480 351204 14484 351236
rect 14516 351204 14520 351236
rect 14480 351200 14520 351204
rect 14560 351396 14600 351400
rect 14560 351364 14564 351396
rect 14596 351364 14600 351396
rect 14560 351316 14600 351364
rect 14560 351284 14564 351316
rect 14596 351284 14600 351316
rect 14560 351236 14600 351284
rect 14560 351204 14564 351236
rect 14596 351204 14600 351236
rect 14560 351200 14600 351204
rect 14640 351396 14680 351400
rect 14640 351364 14644 351396
rect 14676 351364 14680 351396
rect 14640 351316 14680 351364
rect 14640 351284 14644 351316
rect 14676 351284 14680 351316
rect 14640 351236 14680 351284
rect 14640 351204 14644 351236
rect 14676 351204 14680 351236
rect 14640 351200 14680 351204
rect 14720 351396 14760 351400
rect 14720 351364 14724 351396
rect 14756 351364 14760 351396
rect 14720 351316 14760 351364
rect 14720 351284 14724 351316
rect 14756 351284 14760 351316
rect 14720 351236 14760 351284
rect 14720 351204 14724 351236
rect 14756 351204 14760 351236
rect 14720 351200 14760 351204
rect 14800 351396 14840 351400
rect 14800 351364 14804 351396
rect 14836 351364 14840 351396
rect 14800 351316 14840 351364
rect 14800 351284 14804 351316
rect 14836 351284 14840 351316
rect 14800 351236 14840 351284
rect 14800 351204 14804 351236
rect 14836 351204 14840 351236
rect 14800 351200 14840 351204
rect 14880 351396 14920 351400
rect 14880 351364 14884 351396
rect 14916 351364 14920 351396
rect 14880 351316 14920 351364
rect 14880 351284 14884 351316
rect 14916 351284 14920 351316
rect 14880 351236 14920 351284
rect 14880 351204 14884 351236
rect 14916 351204 14920 351236
rect 14880 351200 14920 351204
rect 14960 351396 15000 351400
rect 14960 351364 14964 351396
rect 14996 351364 15000 351396
rect 14960 351316 15000 351364
rect 14960 351284 14964 351316
rect 14996 351284 15000 351316
rect 14960 351236 15000 351284
rect 14960 351204 14964 351236
rect 14996 351204 15000 351236
rect 14960 351200 15000 351204
rect 15040 351396 15080 351400
rect 15040 351364 15044 351396
rect 15076 351364 15080 351396
rect 15040 351316 15080 351364
rect 15040 351284 15044 351316
rect 15076 351284 15080 351316
rect 15040 351236 15080 351284
rect 15040 351204 15044 351236
rect 15076 351204 15080 351236
rect 15040 351200 15080 351204
rect 15120 351396 15160 351400
rect 15120 351364 15124 351396
rect 15156 351364 15160 351396
rect 15120 351316 15160 351364
rect 15120 351284 15124 351316
rect 15156 351284 15160 351316
rect 15120 351236 15160 351284
rect 15120 351204 15124 351236
rect 15156 351204 15160 351236
rect 15120 351200 15160 351204
rect 15200 351396 15240 351400
rect 15200 351364 15204 351396
rect 15236 351364 15240 351396
rect 15200 351316 15240 351364
rect 15200 351284 15204 351316
rect 15236 351284 15240 351316
rect 15200 351236 15240 351284
rect 15200 351204 15204 351236
rect 15236 351204 15240 351236
rect 15200 351200 15240 351204
rect 15280 351396 15320 351400
rect 15280 351364 15284 351396
rect 15316 351364 15320 351396
rect 15280 351316 15320 351364
rect 15280 351284 15284 351316
rect 15316 351284 15320 351316
rect 15280 351236 15320 351284
rect 15280 351204 15284 351236
rect 15316 351204 15320 351236
rect 15280 351200 15320 351204
rect 15360 351396 15400 351400
rect 15360 351364 15364 351396
rect 15396 351364 15400 351396
rect 15360 351316 15400 351364
rect 15360 351284 15364 351316
rect 15396 351284 15400 351316
rect 15360 351236 15400 351284
rect 15360 351204 15364 351236
rect 15396 351204 15400 351236
rect 15360 351200 15400 351204
rect 15440 351396 15480 351400
rect 15440 351364 15444 351396
rect 15476 351364 15480 351396
rect 15440 351316 15480 351364
rect 15440 351284 15444 351316
rect 15476 351284 15480 351316
rect 15440 351236 15480 351284
rect 15440 351204 15444 351236
rect 15476 351204 15480 351236
rect 15440 351200 15480 351204
rect 15520 351396 15560 351400
rect 15520 351364 15524 351396
rect 15556 351364 15560 351396
rect 15520 351316 15560 351364
rect 15520 351284 15524 351316
rect 15556 351284 15560 351316
rect 15520 351236 15560 351284
rect 15520 351204 15524 351236
rect 15556 351204 15560 351236
rect 15520 351200 15560 351204
rect 15600 351396 15640 351400
rect 15600 351364 15604 351396
rect 15636 351364 15640 351396
rect 15600 351316 15640 351364
rect 15600 351284 15604 351316
rect 15636 351284 15640 351316
rect 15600 351236 15640 351284
rect 15600 351204 15604 351236
rect 15636 351204 15640 351236
rect 15600 351200 15640 351204
rect 15680 351396 15720 351400
rect 15680 351364 15684 351396
rect 15716 351364 15720 351396
rect 15680 351316 15720 351364
rect 15680 351284 15684 351316
rect 15716 351284 15720 351316
rect 15680 351236 15720 351284
rect 15680 351204 15684 351236
rect 15716 351204 15720 351236
rect 15680 351200 15720 351204
rect 15760 351396 15800 351400
rect 15760 351364 15764 351396
rect 15796 351364 15800 351396
rect 15760 351316 15800 351364
rect 15760 351284 15764 351316
rect 15796 351284 15800 351316
rect 15760 351236 15800 351284
rect 15760 351204 15764 351236
rect 15796 351204 15800 351236
rect 15760 351200 15800 351204
rect 15840 351396 15880 351400
rect 15840 351364 15844 351396
rect 15876 351364 15880 351396
rect 15840 351316 15880 351364
rect 15840 351284 15844 351316
rect 15876 351284 15880 351316
rect 15840 351236 15880 351284
rect 15840 351204 15844 351236
rect 15876 351204 15880 351236
rect 15840 351200 15880 351204
rect 15920 351396 15960 351400
rect 15920 351364 15924 351396
rect 15956 351364 15960 351396
rect 15920 351316 15960 351364
rect 15920 351284 15924 351316
rect 15956 351284 15960 351316
rect 15920 351236 15960 351284
rect 15920 351204 15924 351236
rect 15956 351204 15960 351236
rect 15920 351200 15960 351204
rect 16000 351396 16040 351400
rect 16000 351364 16004 351396
rect 16036 351364 16040 351396
rect 16000 351316 16040 351364
rect 16000 351284 16004 351316
rect 16036 351284 16040 351316
rect 16000 351236 16040 351284
rect 16000 351204 16004 351236
rect 16036 351204 16040 351236
rect 16000 351200 16040 351204
rect 16080 351396 16120 351400
rect 16080 351364 16084 351396
rect 16116 351364 16120 351396
rect 16080 351316 16120 351364
rect 16080 351284 16084 351316
rect 16116 351284 16120 351316
rect 16080 351236 16120 351284
rect 16080 351204 16084 351236
rect 16116 351204 16120 351236
rect 16080 351200 16120 351204
rect 16160 351396 16200 351400
rect 16160 351364 16164 351396
rect 16196 351364 16200 351396
rect 16160 351316 16200 351364
rect 16160 351284 16164 351316
rect 16196 351284 16200 351316
rect 16160 351236 16200 351284
rect 16160 351204 16164 351236
rect 16196 351204 16200 351236
rect 16160 351200 16200 351204
rect 16240 351396 16280 351400
rect 16240 351364 16244 351396
rect 16276 351364 16280 351396
rect 16240 351316 16280 351364
rect 16240 351284 16244 351316
rect 16276 351284 16280 351316
rect 16240 351236 16280 351284
rect 16240 351204 16244 351236
rect 16276 351204 16280 351236
rect 16240 351200 16280 351204
rect 16320 351396 16360 351400
rect 16320 351364 16324 351396
rect 16356 351364 16360 351396
rect 16320 351316 16360 351364
rect 16320 351284 16324 351316
rect 16356 351284 16360 351316
rect 16320 351236 16360 351284
rect 16320 351204 16324 351236
rect 16356 351204 16360 351236
rect 16320 351200 16360 351204
rect 16400 351396 16440 351400
rect 16400 351364 16404 351396
rect 16436 351364 16440 351396
rect 16400 351316 16440 351364
rect 16400 351284 16404 351316
rect 16436 351284 16440 351316
rect 16400 351236 16440 351284
rect 16400 351204 16404 351236
rect 16436 351204 16440 351236
rect 16400 351200 16440 351204
rect 16480 351396 16520 351400
rect 16480 351364 16484 351396
rect 16516 351364 16520 351396
rect 16480 351316 16520 351364
rect 16480 351284 16484 351316
rect 16516 351284 16520 351316
rect 16480 351236 16520 351284
rect 16480 351204 16484 351236
rect 16516 351204 16520 351236
rect 16480 351200 16520 351204
rect 16560 351396 16600 351400
rect 16560 351364 16564 351396
rect 16596 351364 16600 351396
rect 16560 351316 16600 351364
rect 16560 351284 16564 351316
rect 16596 351284 16600 351316
rect 16560 351236 16600 351284
rect 16560 351204 16564 351236
rect 16596 351204 16600 351236
rect 16560 351200 16600 351204
rect 16640 351396 16680 351400
rect 16640 351364 16644 351396
rect 16676 351364 16680 351396
rect 16640 351316 16680 351364
rect 16640 351284 16644 351316
rect 16676 351284 16680 351316
rect 16640 351236 16680 351284
rect 16640 351204 16644 351236
rect 16676 351204 16680 351236
rect 16640 351200 16680 351204
rect 16720 351396 16760 351400
rect 16720 351364 16724 351396
rect 16756 351364 16760 351396
rect 16720 351316 16760 351364
rect 16720 351284 16724 351316
rect 16756 351284 16760 351316
rect 16720 351236 16760 351284
rect 16720 351204 16724 351236
rect 16756 351204 16760 351236
rect 16720 351200 16760 351204
rect 16800 351396 16840 351400
rect 16800 351364 16804 351396
rect 16836 351364 16840 351396
rect 16800 351316 16840 351364
rect 16800 351284 16804 351316
rect 16836 351284 16840 351316
rect 16800 351236 16840 351284
rect 16800 351204 16804 351236
rect 16836 351204 16840 351236
rect 16800 351200 16840 351204
rect 16880 351396 16920 351400
rect 16880 351364 16884 351396
rect 16916 351364 16920 351396
rect 16880 351316 16920 351364
rect 16880 351284 16884 351316
rect 16916 351284 16920 351316
rect 16880 351236 16920 351284
rect 16880 351204 16884 351236
rect 16916 351204 16920 351236
rect 16880 351200 16920 351204
rect 16960 351396 17000 351400
rect 16960 351364 16964 351396
rect 16996 351364 17000 351396
rect 16960 351316 17000 351364
rect 16960 351284 16964 351316
rect 16996 351284 17000 351316
rect 16960 351236 17000 351284
rect 16960 351204 16964 351236
rect 16996 351204 17000 351236
rect 16960 351200 17000 351204
rect 17040 351396 17080 351400
rect 17040 351364 17044 351396
rect 17076 351364 17080 351396
rect 17040 351316 17080 351364
rect 17040 351284 17044 351316
rect 17076 351284 17080 351316
rect 17040 351236 17080 351284
rect 17040 351204 17044 351236
rect 17076 351204 17080 351236
rect 17040 351200 17080 351204
rect 17120 351396 17160 351400
rect 17120 351364 17124 351396
rect 17156 351364 17160 351396
rect 17120 351316 17160 351364
rect 17120 351284 17124 351316
rect 17156 351284 17160 351316
rect 17120 351236 17160 351284
rect 17120 351204 17124 351236
rect 17156 351204 17160 351236
rect 17120 351200 17160 351204
rect 17200 351396 17240 351400
rect 17200 351364 17204 351396
rect 17236 351364 17240 351396
rect 17200 351316 17240 351364
rect 17200 351284 17204 351316
rect 17236 351284 17240 351316
rect 17200 351236 17240 351284
rect 17200 351204 17204 351236
rect 17236 351204 17240 351236
rect 17200 351200 17240 351204
rect 17280 351396 17320 351400
rect 17280 351364 17284 351396
rect 17316 351364 17320 351396
rect 17280 351316 17320 351364
rect 17280 351284 17284 351316
rect 17316 351284 17320 351316
rect 17280 351236 17320 351284
rect 17280 351204 17284 351236
rect 17316 351204 17320 351236
rect 17280 351200 17320 351204
rect 17360 351396 17400 351400
rect 17360 351364 17364 351396
rect 17396 351364 17400 351396
rect 17360 351316 17400 351364
rect 17360 351284 17364 351316
rect 17396 351284 17400 351316
rect 17360 351236 17400 351284
rect 17360 351204 17364 351236
rect 17396 351204 17400 351236
rect 17360 351200 17400 351204
rect 17440 351396 17480 351400
rect 17440 351364 17444 351396
rect 17476 351364 17480 351396
rect 17440 351316 17480 351364
rect 17440 351284 17444 351316
rect 17476 351284 17480 351316
rect 17440 351236 17480 351284
rect 17440 351204 17444 351236
rect 17476 351204 17480 351236
rect 17440 351200 17480 351204
rect 17520 351396 17560 351400
rect 17520 351364 17524 351396
rect 17556 351364 17560 351396
rect 17520 351316 17560 351364
rect 17520 351284 17524 351316
rect 17556 351284 17560 351316
rect 17520 351236 17560 351284
rect 17520 351204 17524 351236
rect 17556 351204 17560 351236
rect 17520 351200 17560 351204
rect 17600 351396 17640 351400
rect 17600 351364 17604 351396
rect 17636 351364 17640 351396
rect 17600 351316 17640 351364
rect 17600 351284 17604 351316
rect 17636 351284 17640 351316
rect 17600 351236 17640 351284
rect 17600 351204 17604 351236
rect 17636 351204 17640 351236
rect 17600 351200 17640 351204
rect 17680 351396 17720 351400
rect 17680 351364 17684 351396
rect 17716 351364 17720 351396
rect 17680 351316 17720 351364
rect 17680 351284 17684 351316
rect 17716 351284 17720 351316
rect 17680 351236 17720 351284
rect 17680 351204 17684 351236
rect 17716 351204 17720 351236
rect 17680 351200 17720 351204
rect 17760 351396 17800 351400
rect 17760 351364 17764 351396
rect 17796 351364 17800 351396
rect 17760 351316 17800 351364
rect 17760 351284 17764 351316
rect 17796 351284 17800 351316
rect 17760 351236 17800 351284
rect 17760 351204 17764 351236
rect 17796 351204 17800 351236
rect 17760 351200 17800 351204
rect 17840 351396 17880 351400
rect 17840 351364 17844 351396
rect 17876 351364 17880 351396
rect 17840 351316 17880 351364
rect 17840 351284 17844 351316
rect 17876 351284 17880 351316
rect 17840 351236 17880 351284
rect 17840 351204 17844 351236
rect 17876 351204 17880 351236
rect 17840 351200 17880 351204
rect 17920 351396 17960 351400
rect 17920 351364 17924 351396
rect 17956 351364 17960 351396
rect 17920 351316 17960 351364
rect 17920 351284 17924 351316
rect 17956 351284 17960 351316
rect 17920 351236 17960 351284
rect 17920 351204 17924 351236
rect 17956 351204 17960 351236
rect 17920 351200 17960 351204
rect 18000 351396 18040 351400
rect 18000 351364 18004 351396
rect 18036 351364 18040 351396
rect 18000 351316 18040 351364
rect 18000 351284 18004 351316
rect 18036 351284 18040 351316
rect 18000 351236 18040 351284
rect 18000 351204 18004 351236
rect 18036 351204 18040 351236
rect 18000 351200 18040 351204
rect 18080 351396 18120 351400
rect 18080 351364 18084 351396
rect 18116 351364 18120 351396
rect 18080 351316 18120 351364
rect 18080 351284 18084 351316
rect 18116 351284 18120 351316
rect 18080 351236 18120 351284
rect 18080 351204 18084 351236
rect 18116 351204 18120 351236
rect 18080 351200 18120 351204
rect 18160 351396 18200 351400
rect 18160 351364 18164 351396
rect 18196 351364 18200 351396
rect 18160 351316 18200 351364
rect 18160 351284 18164 351316
rect 18196 351284 18200 351316
rect 18160 351236 18200 351284
rect 18160 351204 18164 351236
rect 18196 351204 18200 351236
rect 18160 351200 18200 351204
rect 18240 351396 18280 351400
rect 18240 351364 18244 351396
rect 18276 351364 18280 351396
rect 18240 351316 18280 351364
rect 18240 351284 18244 351316
rect 18276 351284 18280 351316
rect 18240 351236 18280 351284
rect 18240 351204 18244 351236
rect 18276 351204 18280 351236
rect 18240 351200 18280 351204
rect 18320 351396 18360 351400
rect 18320 351364 18324 351396
rect 18356 351364 18360 351396
rect 18320 351316 18360 351364
rect 18320 351284 18324 351316
rect 18356 351284 18360 351316
rect 18320 351236 18360 351284
rect 18320 351204 18324 351236
rect 18356 351204 18360 351236
rect 18320 351200 18360 351204
rect 18400 351396 18440 351400
rect 18400 351364 18404 351396
rect 18436 351364 18440 351396
rect 18400 351316 18440 351364
rect 18400 351284 18404 351316
rect 18436 351284 18440 351316
rect 18400 351236 18440 351284
rect 18400 351204 18404 351236
rect 18436 351204 18440 351236
rect 18400 351200 18440 351204
rect 18480 351396 18520 351400
rect 18480 351364 18484 351396
rect 18516 351364 18520 351396
rect 18480 351316 18520 351364
rect 18480 351284 18484 351316
rect 18516 351284 18520 351316
rect 18480 351236 18520 351284
rect 18480 351204 18484 351236
rect 18516 351204 18520 351236
rect 18480 351200 18520 351204
rect 18560 351396 18600 351400
rect 18560 351364 18564 351396
rect 18596 351364 18600 351396
rect 18560 351316 18600 351364
rect 18560 351284 18564 351316
rect 18596 351284 18600 351316
rect 18560 351236 18600 351284
rect 18560 351204 18564 351236
rect 18596 351204 18600 351236
rect 18560 351200 18600 351204
rect 18640 351396 18680 351400
rect 18640 351364 18644 351396
rect 18676 351364 18680 351396
rect 18640 351316 18680 351364
rect 18640 351284 18644 351316
rect 18676 351284 18680 351316
rect 18640 351236 18680 351284
rect 18640 351204 18644 351236
rect 18676 351204 18680 351236
rect 18640 351200 18680 351204
rect 18720 351396 18760 351400
rect 18720 351364 18724 351396
rect 18756 351364 18760 351396
rect 18720 351316 18760 351364
rect 18720 351284 18724 351316
rect 18756 351284 18760 351316
rect 18720 351236 18760 351284
rect 18720 351204 18724 351236
rect 18756 351204 18760 351236
rect 18720 351200 18760 351204
rect 18800 351396 18840 351400
rect 18800 351364 18804 351396
rect 18836 351364 18840 351396
rect 18800 351316 18840 351364
rect 18800 351284 18804 351316
rect 18836 351284 18840 351316
rect 18800 351236 18840 351284
rect 18800 351204 18804 351236
rect 18836 351204 18840 351236
rect 18800 351200 18840 351204
rect 18880 351396 18920 351400
rect 18880 351364 18884 351396
rect 18916 351364 18920 351396
rect 18880 351316 18920 351364
rect 18880 351284 18884 351316
rect 18916 351284 18920 351316
rect 18880 351236 18920 351284
rect 18880 351204 18884 351236
rect 18916 351204 18920 351236
rect 18880 351200 18920 351204
rect 18960 351396 19000 351400
rect 18960 351364 18964 351396
rect 18996 351364 19000 351396
rect 18960 351316 19000 351364
rect 18960 351284 18964 351316
rect 18996 351284 19000 351316
rect 18960 351236 19000 351284
rect 18960 351204 18964 351236
rect 18996 351204 19000 351236
rect 18960 351200 19000 351204
rect 19040 351396 19080 351400
rect 19040 351364 19044 351396
rect 19076 351364 19080 351396
rect 19040 351316 19080 351364
rect 19040 351284 19044 351316
rect 19076 351284 19080 351316
rect 19040 351236 19080 351284
rect 19040 351204 19044 351236
rect 19076 351204 19080 351236
rect 19040 351200 19080 351204
rect 19120 351396 19160 351400
rect 19120 351364 19124 351396
rect 19156 351364 19160 351396
rect 19120 351316 19160 351364
rect 19120 351284 19124 351316
rect 19156 351284 19160 351316
rect 19120 351236 19160 351284
rect 19120 351204 19124 351236
rect 19156 351204 19160 351236
rect 19120 351200 19160 351204
rect 19200 351396 19240 351400
rect 19200 351364 19204 351396
rect 19236 351364 19240 351396
rect 19200 351316 19240 351364
rect 19200 351284 19204 351316
rect 19236 351284 19240 351316
rect 19200 351236 19240 351284
rect 19200 351204 19204 351236
rect 19236 351204 19240 351236
rect 19200 351200 19240 351204
rect 19280 351396 19320 351400
rect 19280 351364 19284 351396
rect 19316 351364 19320 351396
rect 19280 351316 19320 351364
rect 19280 351284 19284 351316
rect 19316 351284 19320 351316
rect 19280 351236 19320 351284
rect 19280 351204 19284 351236
rect 19316 351204 19320 351236
rect 19280 351200 19320 351204
rect 19360 351396 19400 351400
rect 19360 351364 19364 351396
rect 19396 351364 19400 351396
rect 19360 351316 19400 351364
rect 19360 351284 19364 351316
rect 19396 351284 19400 351316
rect 19360 351236 19400 351284
rect 19360 351204 19364 351236
rect 19396 351204 19400 351236
rect 19360 351200 19400 351204
rect 19440 351396 19480 351400
rect 19440 351364 19444 351396
rect 19476 351364 19480 351396
rect 19440 351316 19480 351364
rect 19440 351284 19444 351316
rect 19476 351284 19480 351316
rect 19440 351236 19480 351284
rect 19440 351204 19444 351236
rect 19476 351204 19480 351236
rect 19440 351200 19480 351204
rect 19520 351396 19560 351400
rect 19520 351364 19524 351396
rect 19556 351364 19560 351396
rect 19520 351316 19560 351364
rect 19520 351284 19524 351316
rect 19556 351284 19560 351316
rect 19520 351236 19560 351284
rect 19520 351204 19524 351236
rect 19556 351204 19560 351236
rect 19520 351200 19560 351204
rect 19600 351396 19640 351400
rect 19600 351364 19604 351396
rect 19636 351364 19640 351396
rect 19600 351316 19640 351364
rect 19600 351284 19604 351316
rect 19636 351284 19640 351316
rect 19600 351236 19640 351284
rect 19600 351204 19604 351236
rect 19636 351204 19640 351236
rect 19600 351200 19640 351204
rect 19680 351396 19720 351400
rect 19680 351364 19684 351396
rect 19716 351364 19720 351396
rect 19680 351316 19720 351364
rect 19840 351396 19880 351400
rect 19840 351364 19844 351396
rect 19876 351364 19880 351396
rect 19680 351284 19684 351316
rect 19716 351284 19720 351316
rect 19680 351236 19720 351284
rect 19680 351204 19684 351236
rect 19716 351204 19720 351236
rect 8097 351150 10597 351200
rect 19680 351156 19720 351204
rect 19680 351124 19684 351156
rect 19716 351124 19720 351156
rect 19680 351076 19720 351124
rect 19680 351044 19684 351076
rect 19716 351044 19720 351076
rect 19680 350996 19720 351044
rect 19680 350964 19684 350996
rect 19716 350964 19720 350996
rect 19680 350916 19720 350964
rect 19680 350884 19684 350916
rect 19716 350884 19720 350916
rect 19680 350836 19720 350884
rect 19680 350804 19684 350836
rect 19716 350804 19720 350836
rect 19680 350756 19720 350804
rect 19680 350724 19684 350756
rect 19716 350724 19720 350756
rect 19680 350676 19720 350724
rect 19680 350644 19684 350676
rect 19716 350644 19720 350676
rect 19680 350596 19720 350644
rect 19680 350564 19684 350596
rect 19716 350564 19720 350596
rect 19680 350516 19720 350564
rect 19680 350484 19684 350516
rect 19716 350484 19720 350516
rect 19680 350436 19720 350484
rect 19680 350404 19684 350436
rect 19716 350404 19720 350436
rect 19680 350356 19720 350404
rect 19680 350324 19684 350356
rect 19716 350324 19720 350356
rect 19680 350276 19720 350324
rect 19680 350244 19684 350276
rect 19716 350244 19720 350276
rect 19680 350196 19720 350244
rect 19680 350164 19684 350196
rect 19716 350164 19720 350196
rect 19680 350116 19720 350164
rect 19680 350084 19684 350116
rect 19716 350084 19720 350116
rect 19680 350036 19720 350084
rect 19680 350004 19684 350036
rect 19716 350004 19720 350036
rect 19680 349956 19720 350004
rect 19680 349924 19684 349956
rect 19716 349924 19720 349956
rect 19680 349876 19720 349924
rect 19680 349844 19684 349876
rect 19716 349844 19720 349876
rect 19680 349796 19720 349844
rect 19680 349764 19684 349796
rect 19716 349764 19720 349796
rect 19680 349716 19720 349764
rect 19680 349684 19684 349716
rect 19716 349684 19720 349716
rect 19680 349636 19720 349684
rect 19680 349604 19684 349636
rect 19716 349604 19720 349636
rect 19680 349556 19720 349604
rect 19680 349524 19684 349556
rect 19716 349524 19720 349556
rect 19680 349476 19720 349524
rect 19680 349444 19684 349476
rect 19716 349444 19720 349476
rect 19680 349396 19720 349444
rect 19680 349364 19684 349396
rect 19716 349364 19720 349396
rect 19680 349316 19720 349364
rect 19680 349284 19684 349316
rect 19716 349284 19720 349316
rect 19680 349236 19720 349284
rect 19680 349204 19684 349236
rect 19716 349204 19720 349236
rect 19680 349156 19720 349204
rect 19680 349124 19684 349156
rect 19716 349124 19720 349156
rect 19680 349076 19720 349124
rect 19680 349044 19684 349076
rect 19716 349044 19720 349076
rect 19680 348996 19720 349044
rect 19680 348964 19684 348996
rect 19716 348964 19720 348996
rect 19680 348916 19720 348964
rect 19680 348884 19684 348916
rect 19716 348884 19720 348916
rect 19680 348836 19720 348884
rect 19680 348804 19684 348836
rect 19716 348804 19720 348836
rect 19680 348756 19720 348804
rect 19680 348724 19684 348756
rect 19716 348724 19720 348756
rect 19680 348676 19720 348724
rect 19680 348644 19684 348676
rect 19716 348644 19720 348676
rect 19680 348596 19720 348644
rect 19680 348564 19684 348596
rect 19716 348564 19720 348596
rect 19680 348516 19720 348564
rect 19680 348484 19684 348516
rect 19716 348484 19720 348516
rect 19680 348436 19720 348484
rect 19680 348404 19684 348436
rect 19716 348404 19720 348436
rect 19680 348356 19720 348404
rect 19680 348324 19684 348356
rect 19716 348324 19720 348356
rect 19680 348276 19720 348324
rect 19680 348244 19684 348276
rect 19716 348244 19720 348276
rect 19680 348196 19720 348244
rect 19680 348164 19684 348196
rect 19716 348164 19720 348196
rect 19680 348116 19720 348164
rect 19680 348084 19684 348116
rect 19716 348084 19720 348116
rect 19680 348036 19720 348084
rect 19680 348004 19684 348036
rect 19716 348004 19720 348036
rect 19680 347956 19720 348004
rect 19680 347924 19684 347956
rect 19716 347924 19720 347956
rect 19680 347876 19720 347924
rect 19680 347844 19684 347876
rect 19716 347844 19720 347876
rect 19680 347796 19720 347844
rect 19680 347764 19684 347796
rect 19716 347764 19720 347796
rect 19680 347716 19720 347764
rect 19680 347684 19684 347716
rect 19716 347684 19720 347716
rect 19680 347636 19720 347684
rect 19680 347604 19684 347636
rect 19716 347604 19720 347636
rect 19680 347556 19720 347604
rect 19680 347524 19684 347556
rect 19716 347524 19720 347556
rect 19680 347476 19720 347524
rect 19680 347444 19684 347476
rect 19716 347444 19720 347476
rect 19680 347396 19720 347444
rect 19680 347364 19684 347396
rect 19716 347364 19720 347396
rect 19680 347316 19720 347364
rect 19680 347284 19684 347316
rect 19716 347284 19720 347316
rect 19680 347236 19720 347284
rect 19680 347204 19684 347236
rect 19716 347204 19720 347236
rect 19680 347156 19720 347204
rect 19680 347124 19684 347156
rect 19716 347124 19720 347156
rect 19680 347076 19720 347124
rect 19680 347044 19684 347076
rect 19716 347044 19720 347076
rect 19680 346996 19720 347044
rect 19680 346964 19684 346996
rect 19716 346964 19720 346996
rect 19680 346916 19720 346964
rect 19680 346884 19684 346916
rect 19716 346884 19720 346916
rect 19680 346836 19720 346884
rect 19680 346804 19684 346836
rect 19716 346804 19720 346836
rect 19680 346756 19720 346804
rect 19680 346724 19684 346756
rect 19716 346724 19720 346756
rect 19680 346676 19720 346724
rect 19680 346644 19684 346676
rect 19716 346644 19720 346676
rect 19680 346596 19720 346644
rect 19680 346564 19684 346596
rect 19716 346564 19720 346596
rect 19680 346516 19720 346564
rect 19680 346484 19684 346516
rect 19716 346484 19720 346516
rect 19680 346436 19720 346484
rect 19680 346404 19684 346436
rect 19716 346404 19720 346436
rect 19680 346356 19720 346404
rect 19680 346324 19684 346356
rect 19716 346324 19720 346356
rect 19680 346276 19720 346324
rect 19680 346244 19684 346276
rect 19716 346244 19720 346276
rect 19680 346196 19720 346244
rect 19680 346164 19684 346196
rect 19716 346164 19720 346196
rect 19680 346116 19720 346164
rect 19680 346084 19684 346116
rect 19716 346084 19720 346116
rect 19680 346036 19720 346084
rect 19680 346004 19684 346036
rect 19716 346004 19720 346036
rect 19680 345956 19720 346004
rect 19680 345924 19684 345956
rect 19716 345924 19720 345956
rect 19680 345876 19720 345924
rect 19680 345844 19684 345876
rect 19716 345844 19720 345876
rect 19680 345796 19720 345844
rect 19680 345764 19684 345796
rect 19716 345764 19720 345796
rect 19680 345716 19720 345764
rect 19680 345684 19684 345716
rect 19716 345684 19720 345716
rect 19680 345636 19720 345684
rect 19680 345604 19684 345636
rect 19716 345604 19720 345636
rect 19680 345556 19720 345604
rect 19680 345524 19684 345556
rect 19716 345524 19720 345556
rect 19680 345476 19720 345524
rect 19680 345444 19684 345476
rect 19716 345444 19720 345476
rect 19680 345396 19720 345444
rect 19680 345364 19684 345396
rect 19716 345364 19720 345396
rect 19680 345316 19720 345364
rect 19680 345284 19684 345316
rect 19716 345284 19720 345316
rect 19680 345236 19720 345284
rect 19680 345204 19684 345236
rect 19716 345204 19720 345236
rect 19680 345156 19720 345204
rect 19680 345124 19684 345156
rect 19716 345124 19720 345156
rect 19680 345076 19720 345124
rect 19680 345044 19684 345076
rect 19716 345044 19720 345076
rect 19680 344996 19720 345044
rect 19680 344964 19684 344996
rect 19716 344964 19720 344996
rect 19680 344916 19720 344964
rect 19680 344884 19684 344916
rect 19716 344884 19720 344916
rect 19680 344836 19720 344884
rect 19680 344804 19684 344836
rect 19716 344804 19720 344836
rect 19680 344756 19720 344804
rect 19680 344724 19684 344756
rect 19716 344724 19720 344756
rect 19680 344676 19720 344724
rect 19680 344644 19684 344676
rect 19716 344644 19720 344676
rect 19680 344596 19720 344644
rect 19680 344564 19684 344596
rect 19716 344564 19720 344596
rect 19680 344516 19720 344564
rect 19680 344484 19684 344516
rect 19716 344484 19720 344516
rect 19680 344436 19720 344484
rect 19680 344404 19684 344436
rect 19716 344404 19720 344436
rect 19680 344356 19720 344404
rect 19680 344324 19684 344356
rect 19716 344324 19720 344356
rect 19680 344276 19720 344324
rect 19680 344244 19684 344276
rect 19716 344244 19720 344276
rect 19680 344196 19720 344244
rect 19680 344164 19684 344196
rect 19716 344164 19720 344196
rect 19680 344116 19720 344164
rect 19680 344084 19684 344116
rect 19716 344084 19720 344116
rect 19680 344036 19720 344084
rect 19680 344004 19684 344036
rect 19716 344004 19720 344036
rect 19680 343956 19720 344004
rect 19680 343924 19684 343956
rect 19716 343924 19720 343956
rect 19680 343876 19720 343924
rect 19680 343844 19684 343876
rect 19716 343844 19720 343876
rect 19680 343796 19720 343844
rect 19680 343764 19684 343796
rect 19716 343764 19720 343796
rect 19680 343716 19720 343764
rect 19680 343684 19684 343716
rect 19716 343684 19720 343716
rect 19680 343636 19720 343684
rect 19680 343604 19684 343636
rect 19716 343604 19720 343636
rect 19680 343556 19720 343604
rect 19680 343524 19684 343556
rect 19716 343524 19720 343556
rect 19680 343476 19720 343524
rect 19680 343444 19684 343476
rect 19716 343444 19720 343476
rect 19680 343396 19720 343444
rect 19680 343364 19684 343396
rect 19716 343364 19720 343396
rect 19680 343316 19720 343364
rect 19680 343284 19684 343316
rect 19716 343284 19720 343316
rect 19680 343236 19720 343284
rect 19680 343204 19684 343236
rect 19716 343204 19720 343236
rect 19680 343156 19720 343204
rect 19680 343124 19684 343156
rect 19716 343124 19720 343156
rect 19680 343076 19720 343124
rect 19680 343044 19684 343076
rect 19716 343044 19720 343076
rect 19680 342996 19720 343044
rect 19680 342964 19684 342996
rect 19716 342964 19720 342996
rect 19680 342916 19720 342964
rect 19680 342884 19684 342916
rect 19716 342884 19720 342916
rect 19680 342836 19720 342884
rect 19680 342804 19684 342836
rect 19716 342804 19720 342836
rect 19680 342756 19720 342804
rect 19680 342724 19684 342756
rect 19716 342724 19720 342756
rect 19680 342676 19720 342724
rect 19680 342644 19684 342676
rect 19716 342644 19720 342676
rect -400 340400 850 342621
rect 19680 342596 19720 342644
rect 19680 342564 19684 342596
rect 19716 342564 19720 342596
rect 19680 342516 19720 342564
rect 19680 342484 19684 342516
rect 19716 342484 19720 342516
rect 19680 342436 19720 342484
rect 19680 342404 19684 342436
rect 19716 342404 19720 342436
rect 19680 342356 19720 342404
rect 19680 342324 19684 342356
rect 19716 342324 19720 342356
rect 19680 342276 19720 342324
rect 19680 342244 19684 342276
rect 19716 342244 19720 342276
rect 19680 342196 19720 342244
rect 19680 342164 19684 342196
rect 19716 342164 19720 342196
rect 19680 342116 19720 342164
rect 19680 342084 19684 342116
rect 19716 342084 19720 342116
rect 19680 342036 19720 342084
rect 19680 342004 19684 342036
rect 19716 342004 19720 342036
rect 19680 341956 19720 342004
rect 19680 341924 19684 341956
rect 19716 341924 19720 341956
rect 19680 341876 19720 341924
rect 19680 341844 19684 341876
rect 19716 341844 19720 341876
rect 19680 341796 19720 341844
rect 19680 341764 19684 341796
rect 19716 341764 19720 341796
rect 19680 341716 19720 341764
rect 19680 341684 19684 341716
rect 19716 341684 19720 341716
rect 19680 341636 19720 341684
rect 19680 341604 19684 341636
rect 19716 341604 19720 341636
rect 19680 341556 19720 341604
rect 19680 341524 19684 341556
rect 19716 341524 19720 341556
rect 19680 341476 19720 341524
rect 19680 341444 19684 341476
rect 19716 341444 19720 341476
rect 19680 341396 19720 341444
rect 19680 341364 19684 341396
rect 19716 341364 19720 341396
rect 19680 341316 19720 341364
rect 19680 341284 19684 341316
rect 19716 341284 19720 341316
rect 19680 341236 19720 341284
rect 19680 341204 19684 341236
rect 19716 341204 19720 341236
rect 19680 341156 19720 341204
rect 19680 341124 19684 341156
rect 19716 341124 19720 341156
rect 19680 341076 19720 341124
rect 19680 341044 19684 341076
rect 19716 341044 19720 341076
rect 19680 340996 19720 341044
rect 19680 340964 19684 340996
rect 19716 340964 19720 340996
rect 19680 340916 19720 340964
rect 19680 340884 19684 340916
rect 19716 340884 19720 340916
rect 19680 340836 19720 340884
rect 19680 340804 19684 340836
rect 19716 340804 19720 340836
rect 19680 340756 19720 340804
rect 19680 340724 19684 340756
rect 19716 340724 19720 340756
rect 19680 340676 19720 340724
rect 19680 340644 19684 340676
rect 19716 340644 19720 340676
rect 19680 340596 19720 340644
rect 19680 340564 19684 340596
rect 19716 340564 19720 340596
rect 19680 340516 19720 340564
rect 19680 340484 19684 340516
rect 19716 340484 19720 340516
rect 19680 340436 19720 340484
rect 19680 340404 19684 340436
rect 19716 340404 19720 340436
rect -400 340200 14400 340400
rect -400 340121 850 340200
rect -400 321921 830 324321
rect -400 316921 830 319321
rect 3200 287160 3280 287200
rect 3240 287120 3280 287160
rect -400 279721 830 282121
rect 14200 279400 14400 340200
rect 19680 340356 19720 340404
rect 19680 340324 19684 340356
rect 19716 340324 19720 340356
rect 19680 340276 19720 340324
rect 19680 340244 19684 340276
rect 19716 340244 19720 340276
rect 19680 340196 19720 340244
rect 19680 340164 19684 340196
rect 19716 340164 19720 340196
rect 19680 340116 19720 340164
rect 19680 340084 19684 340116
rect 19716 340084 19720 340116
rect 19680 340036 19720 340084
rect 19680 340004 19684 340036
rect 19716 340004 19720 340036
rect 19680 339956 19720 340004
rect 19680 339924 19684 339956
rect 19716 339924 19720 339956
rect 19680 339876 19720 339924
rect 19680 339844 19684 339876
rect 19716 339844 19720 339876
rect 19680 339796 19720 339844
rect 19680 339764 19684 339796
rect 19716 339764 19720 339796
rect 19680 339716 19720 339764
rect 19680 339684 19684 339716
rect 19716 339684 19720 339716
rect 19680 339636 19720 339684
rect 19680 339604 19684 339636
rect 19716 339604 19720 339636
rect 19680 339556 19720 339604
rect 19680 339524 19684 339556
rect 19716 339524 19720 339556
rect 19680 339476 19720 339524
rect 19680 339444 19684 339476
rect 19716 339444 19720 339476
rect 19680 339396 19720 339444
rect 19680 339364 19684 339396
rect 19716 339364 19720 339396
rect 19680 339316 19720 339364
rect 19680 339284 19684 339316
rect 19716 339284 19720 339316
rect 19680 339236 19720 339284
rect 19680 339204 19684 339236
rect 19716 339204 19720 339236
rect 19680 339156 19720 339204
rect 19680 339124 19684 339156
rect 19716 339124 19720 339156
rect 19680 339076 19720 339124
rect 19680 339044 19684 339076
rect 19716 339044 19720 339076
rect 19680 338996 19720 339044
rect 19680 338964 19684 338996
rect 19716 338964 19720 338996
rect 19680 338916 19720 338964
rect 19680 338884 19684 338916
rect 19716 338884 19720 338916
rect 19680 338836 19720 338884
rect 19680 338804 19684 338836
rect 19716 338804 19720 338836
rect 19680 338756 19720 338804
rect 19680 338724 19684 338756
rect 19716 338724 19720 338756
rect 19680 338676 19720 338724
rect 19680 338644 19684 338676
rect 19716 338644 19720 338676
rect 19680 338596 19720 338644
rect 19680 338564 19684 338596
rect 19716 338564 19720 338596
rect 19680 338516 19720 338564
rect 19680 338484 19684 338516
rect 19716 338484 19720 338516
rect 19680 338436 19720 338484
rect 19680 338404 19684 338436
rect 19716 338404 19720 338436
rect 19680 338356 19720 338404
rect 19680 338324 19684 338356
rect 19716 338324 19720 338356
rect 19680 338276 19720 338324
rect 19680 338244 19684 338276
rect 19716 338244 19720 338276
rect 19680 338196 19720 338244
rect 19680 338164 19684 338196
rect 19716 338164 19720 338196
rect 19680 338116 19720 338164
rect 19680 338084 19684 338116
rect 19716 338084 19720 338116
rect 19680 338036 19720 338084
rect 19680 338004 19684 338036
rect 19716 338004 19720 338036
rect 19680 337956 19720 338004
rect 19680 337924 19684 337956
rect 19716 337924 19720 337956
rect 19680 337876 19720 337924
rect 19680 337844 19684 337876
rect 19716 337844 19720 337876
rect 19680 337796 19720 337844
rect 19680 337764 19684 337796
rect 19716 337764 19720 337796
rect 19680 337716 19720 337764
rect 19680 337684 19684 337716
rect 19716 337684 19720 337716
rect 19680 337636 19720 337684
rect 19680 337604 19684 337636
rect 19716 337604 19720 337636
rect 19680 337556 19720 337604
rect 19680 337524 19684 337556
rect 19716 337524 19720 337556
rect 19680 337476 19720 337524
rect 19680 337444 19684 337476
rect 19716 337444 19720 337476
rect 19680 337396 19720 337444
rect 19680 337364 19684 337396
rect 19716 337364 19720 337396
rect 19680 337316 19720 337364
rect 19680 337284 19684 337316
rect 19716 337284 19720 337316
rect 19680 337236 19720 337284
rect 19680 337204 19684 337236
rect 19716 337204 19720 337236
rect 19680 337156 19720 337204
rect 19680 337124 19684 337156
rect 19716 337124 19720 337156
rect 19680 337076 19720 337124
rect 19680 337044 19684 337076
rect 19716 337044 19720 337076
rect 19680 336996 19720 337044
rect 19680 336964 19684 336996
rect 19716 336964 19720 336996
rect 19680 336916 19720 336964
rect 19680 336884 19684 336916
rect 19716 336884 19720 336916
rect 19680 336836 19720 336884
rect 19680 336804 19684 336836
rect 19716 336804 19720 336836
rect 19680 336756 19720 336804
rect 19680 336724 19684 336756
rect 19716 336724 19720 336756
rect 19680 336676 19720 336724
rect 19680 336644 19684 336676
rect 19716 336644 19720 336676
rect 19680 336596 19720 336644
rect 19680 336564 19684 336596
rect 19716 336564 19720 336596
rect 19680 336516 19720 336564
rect 19680 336484 19684 336516
rect 19716 336484 19720 336516
rect 19680 336436 19720 336484
rect 19680 336404 19684 336436
rect 19716 336404 19720 336436
rect 19680 336356 19720 336404
rect 19680 336324 19684 336356
rect 19716 336324 19720 336356
rect 19680 336276 19720 336324
rect 19680 336244 19684 336276
rect 19716 336244 19720 336276
rect 19680 336196 19720 336244
rect 19680 336164 19684 336196
rect 19716 336164 19720 336196
rect 19680 336116 19720 336164
rect 19680 336084 19684 336116
rect 19716 336084 19720 336116
rect 19680 336036 19720 336084
rect 19680 336004 19684 336036
rect 19716 336004 19720 336036
rect 19680 335956 19720 336004
rect 19680 335924 19684 335956
rect 19716 335924 19720 335956
rect 19680 335876 19720 335924
rect 19680 335844 19684 335876
rect 19716 335844 19720 335876
rect 19680 335796 19720 335844
rect 19680 335764 19684 335796
rect 19716 335764 19720 335796
rect 19680 335716 19720 335764
rect 19680 335684 19684 335716
rect 19716 335684 19720 335716
rect 19680 335636 19720 335684
rect 19680 335604 19684 335636
rect 19716 335604 19720 335636
rect 19680 335556 19720 335604
rect 19680 335524 19684 335556
rect 19716 335524 19720 335556
rect 19680 335476 19720 335524
rect 19680 335444 19684 335476
rect 19716 335444 19720 335476
rect 19680 335396 19720 335444
rect 19680 335364 19684 335396
rect 19716 335364 19720 335396
rect 19680 335316 19720 335364
rect 19680 335284 19684 335316
rect 19716 335284 19720 335316
rect 19680 335236 19720 335284
rect 19680 335204 19684 335236
rect 19716 335204 19720 335236
rect 19680 335156 19720 335204
rect 19680 335124 19684 335156
rect 19716 335124 19720 335156
rect 19680 335076 19720 335124
rect 19680 335044 19684 335076
rect 19716 335044 19720 335076
rect 19680 334996 19720 335044
rect 19680 334964 19684 334996
rect 19716 334964 19720 334996
rect 19680 334916 19720 334964
rect 19680 334884 19684 334916
rect 19716 334884 19720 334916
rect 19680 334836 19720 334884
rect 19680 334804 19684 334836
rect 19716 334804 19720 334836
rect 19680 334756 19720 334804
rect 19680 334724 19684 334756
rect 19716 334724 19720 334756
rect 19680 334676 19720 334724
rect 19680 334644 19684 334676
rect 19716 334644 19720 334676
rect 19680 334596 19720 334644
rect 19680 334564 19684 334596
rect 19716 334564 19720 334596
rect 19680 334516 19720 334564
rect 19680 334484 19684 334516
rect 19716 334484 19720 334516
rect 19680 334436 19720 334484
rect 19680 334404 19684 334436
rect 19716 334404 19720 334436
rect 19680 334356 19720 334404
rect 19680 334324 19684 334356
rect 19716 334324 19720 334356
rect 19680 334276 19720 334324
rect 19680 334244 19684 334276
rect 19716 334244 19720 334276
rect 19680 334196 19720 334244
rect 19680 334164 19684 334196
rect 19716 334164 19720 334196
rect 19680 334116 19720 334164
rect 19680 334084 19684 334116
rect 19716 334084 19720 334116
rect 19680 334036 19720 334084
rect 19680 334004 19684 334036
rect 19716 334004 19720 334036
rect 19680 333956 19720 334004
rect 19680 333924 19684 333956
rect 19716 333924 19720 333956
rect 19680 333876 19720 333924
rect 19680 333844 19684 333876
rect 19716 333844 19720 333876
rect 19680 333796 19720 333844
rect 19680 333764 19684 333796
rect 19716 333764 19720 333796
rect 19680 333716 19720 333764
rect 19680 333684 19684 333716
rect 19716 333684 19720 333716
rect 19680 333636 19720 333684
rect 19680 333604 19684 333636
rect 19716 333604 19720 333636
rect 19680 333556 19720 333604
rect 19680 333524 19684 333556
rect 19716 333524 19720 333556
rect 19680 333476 19720 333524
rect 19680 333444 19684 333476
rect 19716 333444 19720 333476
rect 19680 333396 19720 333444
rect 19680 333364 19684 333396
rect 19716 333364 19720 333396
rect 19680 333316 19720 333364
rect 19680 333284 19684 333316
rect 19716 333284 19720 333316
rect 19680 333236 19720 333284
rect 19680 333204 19684 333236
rect 19716 333204 19720 333236
rect 19680 333156 19720 333204
rect 19680 333124 19684 333156
rect 19716 333124 19720 333156
rect 19680 333076 19720 333124
rect 19680 333044 19684 333076
rect 19716 333044 19720 333076
rect 19680 332996 19720 333044
rect 19680 332964 19684 332996
rect 19716 332964 19720 332996
rect 19680 332916 19720 332964
rect 19680 332884 19684 332916
rect 19716 332884 19720 332916
rect 19680 332836 19720 332884
rect 19680 332804 19684 332836
rect 19716 332804 19720 332836
rect 19680 332756 19720 332804
rect 19680 332724 19684 332756
rect 19716 332724 19720 332756
rect 19680 332676 19720 332724
rect 19680 332644 19684 332676
rect 19716 332644 19720 332676
rect 19680 332596 19720 332644
rect 19680 332564 19684 332596
rect 19716 332564 19720 332596
rect 19680 332516 19720 332564
rect 19680 332484 19684 332516
rect 19716 332484 19720 332516
rect 19680 332436 19720 332484
rect 19680 332404 19684 332436
rect 19716 332404 19720 332436
rect 19680 332356 19720 332404
rect 19680 332324 19684 332356
rect 19716 332324 19720 332356
rect 19680 332276 19720 332324
rect 19680 332244 19684 332276
rect 19716 332244 19720 332276
rect 19680 332196 19720 332244
rect 19680 332164 19684 332196
rect 19716 332164 19720 332196
rect 19680 332116 19720 332164
rect 19680 332084 19684 332116
rect 19716 332084 19720 332116
rect 19680 332036 19720 332084
rect 19680 332004 19684 332036
rect 19716 332004 19720 332036
rect 19680 331956 19720 332004
rect 19680 331924 19684 331956
rect 19716 331924 19720 331956
rect 19680 331876 19720 331924
rect 19680 331844 19684 331876
rect 19716 331844 19720 331876
rect 19680 331796 19720 331844
rect 19680 331764 19684 331796
rect 19716 331764 19720 331796
rect 19680 331716 19720 331764
rect 19680 331684 19684 331716
rect 19716 331684 19720 331716
rect 19680 331636 19720 331684
rect 19680 331604 19684 331636
rect 19716 331604 19720 331636
rect 19680 331556 19720 331604
rect 19680 331524 19684 331556
rect 19716 331524 19720 331556
rect 19680 331476 19720 331524
rect 19680 331444 19684 331476
rect 19716 331444 19720 331476
rect 19680 331396 19720 331444
rect 19680 331364 19684 331396
rect 19716 331364 19720 331396
rect 19680 331316 19720 331364
rect 19680 331284 19684 331316
rect 19716 331284 19720 331316
rect 19680 331236 19720 331284
rect 19680 331204 19684 331236
rect 19716 331204 19720 331236
rect 19680 331156 19720 331204
rect 19680 331124 19684 331156
rect 19716 331124 19720 331156
rect 19680 331076 19720 331124
rect 19680 331044 19684 331076
rect 19716 331044 19720 331076
rect 19680 330996 19720 331044
rect 19680 330964 19684 330996
rect 19716 330964 19720 330996
rect 19680 330916 19720 330964
rect 19680 330884 19684 330916
rect 19716 330884 19720 330916
rect 19680 330836 19720 330884
rect 19680 330804 19684 330836
rect 19716 330804 19720 330836
rect 19680 330756 19720 330804
rect 19680 330724 19684 330756
rect 19716 330724 19720 330756
rect 19680 330676 19720 330724
rect 19680 330644 19684 330676
rect 19716 330644 19720 330676
rect 19680 330596 19720 330644
rect 19680 330564 19684 330596
rect 19716 330564 19720 330596
rect 19680 330516 19720 330564
rect 19680 330484 19684 330516
rect 19716 330484 19720 330516
rect 19680 330436 19720 330484
rect 19680 330404 19684 330436
rect 19716 330404 19720 330436
rect 19680 330356 19720 330404
rect 19680 330324 19684 330356
rect 19716 330324 19720 330356
rect 19680 330276 19720 330324
rect 19680 330244 19684 330276
rect 19716 330244 19720 330276
rect 19680 330196 19720 330244
rect 19680 330164 19684 330196
rect 19716 330164 19720 330196
rect 19680 330116 19720 330164
rect 19680 330084 19684 330116
rect 19716 330084 19720 330116
rect 19680 330036 19720 330084
rect 19680 330004 19684 330036
rect 19716 330004 19720 330036
rect 19680 329956 19720 330004
rect 19680 329924 19684 329956
rect 19716 329924 19720 329956
rect 19680 329876 19720 329924
rect 19680 329844 19684 329876
rect 19716 329844 19720 329876
rect 19680 329796 19720 329844
rect 19680 329764 19684 329796
rect 19716 329764 19720 329796
rect 19680 329716 19720 329764
rect 19680 329684 19684 329716
rect 19716 329684 19720 329716
rect 19680 329636 19720 329684
rect 19680 329604 19684 329636
rect 19716 329604 19720 329636
rect 19680 329556 19720 329604
rect 19680 329524 19684 329556
rect 19716 329524 19720 329556
rect 19680 329476 19720 329524
rect 19680 329444 19684 329476
rect 19716 329444 19720 329476
rect 19680 329396 19720 329444
rect 19680 329364 19684 329396
rect 19716 329364 19720 329396
rect 19680 329316 19720 329364
rect 19680 329284 19684 329316
rect 19716 329284 19720 329316
rect 19680 329236 19720 329284
rect 19680 329204 19684 329236
rect 19716 329204 19720 329236
rect 19680 329156 19720 329204
rect 19680 329124 19684 329156
rect 19716 329124 19720 329156
rect 19680 329076 19720 329124
rect 19680 329044 19684 329076
rect 19716 329044 19720 329076
rect 19680 328996 19720 329044
rect 19680 328964 19684 328996
rect 19716 328964 19720 328996
rect 19680 328916 19720 328964
rect 19680 328884 19684 328916
rect 19716 328884 19720 328916
rect 19680 328836 19720 328884
rect 19680 328804 19684 328836
rect 19716 328804 19720 328836
rect 19680 328756 19720 328804
rect 19680 328724 19684 328756
rect 19716 328724 19720 328756
rect 19680 328676 19720 328724
rect 19680 328644 19684 328676
rect 19716 328644 19720 328676
rect 19680 328596 19720 328644
rect 19680 328564 19684 328596
rect 19716 328564 19720 328596
rect 19680 328516 19720 328564
rect 19680 328484 19684 328516
rect 19716 328484 19720 328516
rect 19680 328436 19720 328484
rect 19680 328404 19684 328436
rect 19716 328404 19720 328436
rect 19680 328356 19720 328404
rect 19680 328324 19684 328356
rect 19716 328324 19720 328356
rect 19680 328276 19720 328324
rect 19680 328244 19684 328276
rect 19716 328244 19720 328276
rect 19680 328196 19720 328244
rect 19680 328164 19684 328196
rect 19716 328164 19720 328196
rect 19680 328116 19720 328164
rect 19680 328084 19684 328116
rect 19716 328084 19720 328116
rect 19680 328036 19720 328084
rect 19680 328004 19684 328036
rect 19716 328004 19720 328036
rect 19680 327956 19720 328004
rect 19680 327924 19684 327956
rect 19716 327924 19720 327956
rect 19680 327876 19720 327924
rect 19680 327844 19684 327876
rect 19716 327844 19720 327876
rect 19680 327796 19720 327844
rect 19680 327764 19684 327796
rect 19716 327764 19720 327796
rect 19680 327716 19720 327764
rect 19680 327684 19684 327716
rect 19716 327684 19720 327716
rect 19680 327636 19720 327684
rect 19680 327604 19684 327636
rect 19716 327604 19720 327636
rect 19680 327556 19720 327604
rect 19680 327524 19684 327556
rect 19716 327524 19720 327556
rect 19680 327476 19720 327524
rect 19680 327444 19684 327476
rect 19716 327444 19720 327476
rect 19680 327396 19720 327444
rect 19680 327364 19684 327396
rect 19716 327364 19720 327396
rect 19680 327316 19720 327364
rect 19680 327284 19684 327316
rect 19716 327284 19720 327316
rect 19680 327236 19720 327284
rect 19680 327204 19684 327236
rect 19716 327204 19720 327236
rect 19680 327156 19720 327204
rect 19680 327124 19684 327156
rect 19716 327124 19720 327156
rect 19680 327076 19720 327124
rect 19680 327044 19684 327076
rect 19716 327044 19720 327076
rect 19680 326996 19720 327044
rect 19680 326964 19684 326996
rect 19716 326964 19720 326996
rect 19680 326916 19720 326964
rect 19680 326884 19684 326916
rect 19716 326884 19720 326916
rect 19680 326836 19720 326884
rect 19680 326804 19684 326836
rect 19716 326804 19720 326836
rect 19680 326756 19720 326804
rect 19680 326724 19684 326756
rect 19716 326724 19720 326756
rect 19680 326676 19720 326724
rect 19680 326644 19684 326676
rect 19716 326644 19720 326676
rect 19680 326596 19720 326644
rect 19680 326564 19684 326596
rect 19716 326564 19720 326596
rect 19680 326516 19720 326564
rect 19680 326484 19684 326516
rect 19716 326484 19720 326516
rect 19680 326436 19720 326484
rect 19680 326404 19684 326436
rect 19716 326404 19720 326436
rect 19680 326356 19720 326404
rect 19680 326324 19684 326356
rect 19716 326324 19720 326356
rect 19680 326276 19720 326324
rect 19680 326244 19684 326276
rect 19716 326244 19720 326276
rect 19680 326196 19720 326244
rect 19680 326164 19684 326196
rect 19716 326164 19720 326196
rect 19680 326116 19720 326164
rect 19680 326084 19684 326116
rect 19716 326084 19720 326116
rect 19680 326036 19720 326084
rect 19680 326004 19684 326036
rect 19716 326004 19720 326036
rect 19680 325956 19720 326004
rect 19680 325924 19684 325956
rect 19716 325924 19720 325956
rect 19680 325876 19720 325924
rect 19680 325844 19684 325876
rect 19716 325844 19720 325876
rect 19680 325796 19720 325844
rect 19680 325764 19684 325796
rect 19716 325764 19720 325796
rect 19680 325716 19720 325764
rect 19680 325684 19684 325716
rect 19716 325684 19720 325716
rect 19680 325636 19720 325684
rect 19680 325604 19684 325636
rect 19716 325604 19720 325636
rect 19680 325556 19720 325604
rect 19680 325524 19684 325556
rect 19716 325524 19720 325556
rect 19680 325476 19720 325524
rect 19680 325444 19684 325476
rect 19716 325444 19720 325476
rect 19680 325396 19720 325444
rect 19680 325364 19684 325396
rect 19716 325364 19720 325396
rect 19680 325316 19720 325364
rect 19680 325284 19684 325316
rect 19716 325284 19720 325316
rect 19680 325236 19720 325284
rect 19680 325204 19684 325236
rect 19716 325204 19720 325236
rect 19680 325156 19720 325204
rect 19680 325124 19684 325156
rect 19716 325124 19720 325156
rect 19680 325076 19720 325124
rect 19680 325044 19684 325076
rect 19716 325044 19720 325076
rect 19680 324996 19720 325044
rect 19680 324964 19684 324996
rect 19716 324964 19720 324996
rect 19680 324916 19720 324964
rect 19680 324884 19684 324916
rect 19716 324884 19720 324916
rect 19680 324836 19720 324884
rect 19680 324804 19684 324836
rect 19716 324804 19720 324836
rect 19680 324756 19720 324804
rect 19680 324724 19684 324756
rect 19716 324724 19720 324756
rect 19680 324676 19720 324724
rect 19680 324644 19684 324676
rect 19716 324644 19720 324676
rect 19680 324596 19720 324644
rect 19680 324564 19684 324596
rect 19716 324564 19720 324596
rect 19680 324516 19720 324564
rect 19680 324484 19684 324516
rect 19716 324484 19720 324516
rect 19680 324436 19720 324484
rect 19680 324404 19684 324436
rect 19716 324404 19720 324436
rect 19680 324356 19720 324404
rect 19680 324324 19684 324356
rect 19716 324324 19720 324356
rect 19680 324276 19720 324324
rect 19680 324244 19684 324276
rect 19716 324244 19720 324276
rect 19680 324196 19720 324244
rect 19680 324164 19684 324196
rect 19716 324164 19720 324196
rect 19680 324116 19720 324164
rect 19680 324084 19684 324116
rect 19716 324084 19720 324116
rect 19680 324036 19720 324084
rect 19680 324004 19684 324036
rect 19716 324004 19720 324036
rect 19680 323956 19720 324004
rect 19680 323924 19684 323956
rect 19716 323924 19720 323956
rect 19680 323876 19720 323924
rect 19680 323844 19684 323876
rect 19716 323844 19720 323876
rect 19680 323796 19720 323844
rect 19680 323764 19684 323796
rect 19716 323764 19720 323796
rect 19680 323716 19720 323764
rect 19680 323684 19684 323716
rect 19716 323684 19720 323716
rect 19680 323636 19720 323684
rect 19680 323604 19684 323636
rect 19716 323604 19720 323636
rect 19680 323556 19720 323604
rect 19680 323524 19684 323556
rect 19716 323524 19720 323556
rect 19680 323476 19720 323524
rect 19680 323444 19684 323476
rect 19716 323444 19720 323476
rect 19680 323396 19720 323444
rect 19680 323364 19684 323396
rect 19716 323364 19720 323396
rect 19680 323316 19720 323364
rect 19680 323284 19684 323316
rect 19716 323284 19720 323316
rect 19680 323236 19720 323284
rect 19680 323204 19684 323236
rect 19716 323204 19720 323236
rect 19680 323156 19720 323204
rect 19680 323124 19684 323156
rect 19716 323124 19720 323156
rect 19680 323076 19720 323124
rect 19680 323044 19684 323076
rect 19716 323044 19720 323076
rect 19680 322996 19720 323044
rect 19680 322964 19684 322996
rect 19716 322964 19720 322996
rect 19680 322916 19720 322964
rect 19680 322884 19684 322916
rect 19716 322884 19720 322916
rect 19680 322836 19720 322884
rect 19680 322804 19684 322836
rect 19716 322804 19720 322836
rect 19680 322756 19720 322804
rect 19680 322724 19684 322756
rect 19716 322724 19720 322756
rect 19680 322676 19720 322724
rect 19680 322644 19684 322676
rect 19716 322644 19720 322676
rect 19680 322596 19720 322644
rect 19680 322564 19684 322596
rect 19716 322564 19720 322596
rect 19680 322516 19720 322564
rect 19680 322484 19684 322516
rect 19716 322484 19720 322516
rect 19680 322436 19720 322484
rect 19680 322404 19684 322436
rect 19716 322404 19720 322436
rect 19680 322356 19720 322404
rect 19680 322324 19684 322356
rect 19716 322324 19720 322356
rect 19680 322276 19720 322324
rect 19680 322244 19684 322276
rect 19716 322244 19720 322276
rect 19680 322196 19720 322244
rect 19680 322164 19684 322196
rect 19716 322164 19720 322196
rect 19680 322116 19720 322164
rect 19680 322084 19684 322116
rect 19716 322084 19720 322116
rect 19680 322036 19720 322084
rect 19680 322004 19684 322036
rect 19716 322004 19720 322036
rect 19680 321956 19720 322004
rect 19680 321924 19684 321956
rect 19716 321924 19720 321956
rect 19680 321876 19720 321924
rect 19680 321844 19684 321876
rect 19716 321844 19720 321876
rect 19680 321796 19720 321844
rect 19680 321764 19684 321796
rect 19716 321764 19720 321796
rect 19680 321716 19720 321764
rect 19680 321684 19684 321716
rect 19716 321684 19720 321716
rect 19680 321636 19720 321684
rect 19680 321604 19684 321636
rect 19716 321604 19720 321636
rect 19680 321556 19720 321604
rect 19680 321524 19684 321556
rect 19716 321524 19720 321556
rect 19680 321476 19720 321524
rect 19680 321444 19684 321476
rect 19716 321444 19720 321476
rect 19680 321396 19720 321444
rect 19680 321364 19684 321396
rect 19716 321364 19720 321396
rect 19680 321316 19720 321364
rect 19680 321284 19684 321316
rect 19716 321284 19720 321316
rect 19680 321236 19720 321284
rect 19680 321204 19684 321236
rect 19716 321204 19720 321236
rect 19680 321156 19720 321204
rect 19680 321124 19684 321156
rect 19716 321124 19720 321156
rect 19680 321076 19720 321124
rect 19680 321044 19684 321076
rect 19716 321044 19720 321076
rect 19680 320996 19720 321044
rect 19680 320964 19684 320996
rect 19716 320964 19720 320996
rect 19680 320916 19720 320964
rect 19680 320884 19684 320916
rect 19716 320884 19720 320916
rect 19680 320836 19720 320884
rect 19680 320804 19684 320836
rect 19716 320804 19720 320836
rect 19680 320756 19720 320804
rect 19680 320724 19684 320756
rect 19716 320724 19720 320756
rect 19680 320676 19720 320724
rect 19680 320644 19684 320676
rect 19716 320644 19720 320676
rect 19680 320596 19720 320644
rect 19680 320564 19684 320596
rect 19716 320564 19720 320596
rect 19680 320516 19720 320564
rect 19680 320484 19684 320516
rect 19716 320484 19720 320516
rect 19680 320436 19720 320484
rect 19680 320404 19684 320436
rect 19716 320404 19720 320436
rect 19680 320356 19720 320404
rect 19680 320324 19684 320356
rect 19716 320324 19720 320356
rect 19680 320276 19720 320324
rect 19680 320244 19684 320276
rect 19716 320244 19720 320276
rect 19680 320196 19720 320244
rect 19680 320164 19684 320196
rect 19716 320164 19720 320196
rect 19680 320116 19720 320164
rect 19680 320084 19684 320116
rect 19716 320084 19720 320116
rect 19680 320036 19720 320084
rect 19680 320004 19684 320036
rect 19716 320004 19720 320036
rect 19680 319956 19720 320004
rect 19680 319924 19684 319956
rect 19716 319924 19720 319956
rect 19680 319876 19720 319924
rect 19680 319844 19684 319876
rect 19716 319844 19720 319876
rect 19680 319796 19720 319844
rect 19680 319764 19684 319796
rect 19716 319764 19720 319796
rect 19680 319716 19720 319764
rect 19680 319684 19684 319716
rect 19716 319684 19720 319716
rect 19680 319636 19720 319684
rect 19680 319604 19684 319636
rect 19716 319604 19720 319636
rect 19680 319556 19720 319604
rect 19680 319524 19684 319556
rect 19716 319524 19720 319556
rect 19680 319476 19720 319524
rect 19680 319444 19684 319476
rect 19716 319444 19720 319476
rect 19680 319396 19720 319444
rect 19680 319364 19684 319396
rect 19716 319364 19720 319396
rect 19680 319316 19720 319364
rect 19680 319284 19684 319316
rect 19716 319284 19720 319316
rect 19680 319236 19720 319284
rect 19680 319204 19684 319236
rect 19716 319204 19720 319236
rect 19680 319156 19720 319204
rect 19680 319124 19684 319156
rect 19716 319124 19720 319156
rect 19680 319076 19720 319124
rect 19680 319044 19684 319076
rect 19716 319044 19720 319076
rect 19680 318996 19720 319044
rect 19680 318964 19684 318996
rect 19716 318964 19720 318996
rect 19680 318916 19720 318964
rect 19680 318884 19684 318916
rect 19716 318884 19720 318916
rect 19680 318836 19720 318884
rect 19680 318804 19684 318836
rect 19716 318804 19720 318836
rect 19680 318756 19720 318804
rect 19680 318724 19684 318756
rect 19716 318724 19720 318756
rect 19680 318676 19720 318724
rect 19680 318644 19684 318676
rect 19716 318644 19720 318676
rect 19680 318596 19720 318644
rect 19680 318564 19684 318596
rect 19716 318564 19720 318596
rect 19680 318516 19720 318564
rect 19680 318484 19684 318516
rect 19716 318484 19720 318516
rect 19680 318436 19720 318484
rect 19680 318404 19684 318436
rect 19716 318404 19720 318436
rect 19680 318356 19720 318404
rect 19680 318324 19684 318356
rect 19716 318324 19720 318356
rect 19680 318276 19720 318324
rect 19680 318244 19684 318276
rect 19716 318244 19720 318276
rect 19680 318196 19720 318244
rect 19680 318164 19684 318196
rect 19716 318164 19720 318196
rect 19680 318116 19720 318164
rect 19680 318084 19684 318116
rect 19716 318084 19720 318116
rect 19680 318036 19720 318084
rect 19680 318004 19684 318036
rect 19716 318004 19720 318036
rect 19680 317956 19720 318004
rect 19680 317924 19684 317956
rect 19716 317924 19720 317956
rect 19680 317876 19720 317924
rect 19680 317844 19684 317876
rect 19716 317844 19720 317876
rect 19680 317796 19720 317844
rect 19680 317764 19684 317796
rect 19716 317764 19720 317796
rect 19680 317716 19720 317764
rect 19680 317684 19684 317716
rect 19716 317684 19720 317716
rect 19680 317636 19720 317684
rect 19680 317604 19684 317636
rect 19716 317604 19720 317636
rect 19680 317556 19720 317604
rect 19680 317524 19684 317556
rect 19716 317524 19720 317556
rect 19680 317476 19720 317524
rect 19680 317444 19684 317476
rect 19716 317444 19720 317476
rect 19680 317396 19720 317444
rect 19680 317364 19684 317396
rect 19716 317364 19720 317396
rect 19680 317316 19720 317364
rect 19680 317284 19684 317316
rect 19716 317284 19720 317316
rect 19680 317236 19720 317284
rect 19680 317204 19684 317236
rect 19716 317204 19720 317236
rect 19680 317156 19720 317204
rect 19680 317124 19684 317156
rect 19716 317124 19720 317156
rect 19680 317076 19720 317124
rect 19680 317044 19684 317076
rect 19716 317044 19720 317076
rect 19680 316996 19720 317044
rect 19680 316964 19684 316996
rect 19716 316964 19720 316996
rect 19680 316916 19720 316964
rect 19680 316884 19684 316916
rect 19716 316884 19720 316916
rect 19680 316836 19720 316884
rect 19680 316804 19684 316836
rect 19716 316804 19720 316836
rect 19680 316756 19720 316804
rect 19680 316724 19684 316756
rect 19716 316724 19720 316756
rect 19680 316676 19720 316724
rect 19680 316644 19684 316676
rect 19716 316644 19720 316676
rect 19680 316596 19720 316644
rect 19680 316564 19684 316596
rect 19716 316564 19720 316596
rect 19680 316516 19720 316564
rect 19680 316484 19684 316516
rect 19716 316484 19720 316516
rect 19680 316436 19720 316484
rect 19680 316404 19684 316436
rect 19716 316404 19720 316436
rect 19680 316356 19720 316404
rect 19680 316324 19684 316356
rect 19716 316324 19720 316356
rect 19680 316276 19720 316324
rect 19680 316244 19684 316276
rect 19716 316244 19720 316276
rect 19680 316196 19720 316244
rect 19680 316164 19684 316196
rect 19716 316164 19720 316196
rect 19680 316116 19720 316164
rect 19680 316084 19684 316116
rect 19716 316084 19720 316116
rect 19680 316036 19720 316084
rect 19680 316004 19684 316036
rect 19716 316004 19720 316036
rect 19680 315956 19720 316004
rect 19680 315924 19684 315956
rect 19716 315924 19720 315956
rect 19680 315876 19720 315924
rect 19680 315844 19684 315876
rect 19716 315844 19720 315876
rect 19680 315796 19720 315844
rect 19680 315764 19684 315796
rect 19716 315764 19720 315796
rect 19680 315716 19720 315764
rect 19680 315684 19684 315716
rect 19716 315684 19720 315716
rect 19680 315636 19720 315684
rect 19680 315604 19684 315636
rect 19716 315604 19720 315636
rect 19680 315556 19720 315604
rect 19680 315524 19684 315556
rect 19716 315524 19720 315556
rect 19680 315476 19720 315524
rect 19680 315444 19684 315476
rect 19716 315444 19720 315476
rect 19680 315396 19720 315444
rect 19680 315364 19684 315396
rect 19716 315364 19720 315396
rect 19680 315316 19720 315364
rect 19680 315284 19684 315316
rect 19716 315284 19720 315316
rect 19680 315236 19720 315284
rect 19680 315204 19684 315236
rect 19716 315204 19720 315236
rect 19680 315156 19720 315204
rect 19680 315124 19684 315156
rect 19716 315124 19720 315156
rect 19680 315076 19720 315124
rect 19680 315044 19684 315076
rect 19716 315044 19720 315076
rect 19680 314996 19720 315044
rect 19680 314964 19684 314996
rect 19716 314964 19720 314996
rect 19680 314916 19720 314964
rect 19680 314884 19684 314916
rect 19716 314884 19720 314916
rect 19680 314836 19720 314884
rect 19680 314804 19684 314836
rect 19716 314804 19720 314836
rect 19680 314756 19720 314804
rect 19680 314724 19684 314756
rect 19716 314724 19720 314756
rect 19680 314676 19720 314724
rect 19680 314644 19684 314676
rect 19716 314644 19720 314676
rect 19680 314596 19720 314644
rect 19680 314564 19684 314596
rect 19716 314564 19720 314596
rect 19680 314516 19720 314564
rect 19680 314484 19684 314516
rect 19716 314484 19720 314516
rect 19680 314436 19720 314484
rect 19680 314404 19684 314436
rect 19716 314404 19720 314436
rect 19680 314356 19720 314404
rect 19680 314324 19684 314356
rect 19716 314324 19720 314356
rect 19680 314276 19720 314324
rect 19680 314244 19684 314276
rect 19716 314244 19720 314276
rect 19680 314196 19720 314244
rect 19680 314164 19684 314196
rect 19716 314164 19720 314196
rect 19680 314116 19720 314164
rect 19680 314084 19684 314116
rect 19716 314084 19720 314116
rect 19680 314036 19720 314084
rect 19680 314004 19684 314036
rect 19716 314004 19720 314036
rect 19680 313956 19720 314004
rect 19680 313924 19684 313956
rect 19716 313924 19720 313956
rect 19680 313876 19720 313924
rect 19680 313844 19684 313876
rect 19716 313844 19720 313876
rect 19680 313796 19720 313844
rect 19680 313764 19684 313796
rect 19716 313764 19720 313796
rect 19680 313716 19720 313764
rect 19680 313684 19684 313716
rect 19716 313684 19720 313716
rect 19680 313636 19720 313684
rect 19680 313604 19684 313636
rect 19716 313604 19720 313636
rect 19680 313556 19720 313604
rect 19680 313524 19684 313556
rect 19716 313524 19720 313556
rect 19680 313476 19720 313524
rect 19680 313444 19684 313476
rect 19716 313444 19720 313476
rect 19680 313396 19720 313444
rect 19680 313364 19684 313396
rect 19716 313364 19720 313396
rect 19680 313316 19720 313364
rect 19680 313284 19684 313316
rect 19716 313284 19720 313316
rect 19680 313236 19720 313284
rect 19680 313204 19684 313236
rect 19716 313204 19720 313236
rect 19680 313156 19720 313204
rect 19680 313124 19684 313156
rect 19716 313124 19720 313156
rect 19680 313076 19720 313124
rect 19680 313044 19684 313076
rect 19716 313044 19720 313076
rect 19680 312996 19720 313044
rect 19680 312964 19684 312996
rect 19716 312964 19720 312996
rect 19680 312916 19720 312964
rect 19680 312884 19684 312916
rect 19716 312884 19720 312916
rect 19680 312836 19720 312884
rect 19680 312804 19684 312836
rect 19716 312804 19720 312836
rect 19680 312756 19720 312804
rect 19680 312724 19684 312756
rect 19716 312724 19720 312756
rect 19680 312676 19720 312724
rect 19680 312644 19684 312676
rect 19716 312644 19720 312676
rect 19680 312596 19720 312644
rect 19680 312564 19684 312596
rect 19716 312564 19720 312596
rect 19680 312516 19720 312564
rect 19680 312484 19684 312516
rect 19716 312484 19720 312516
rect 19680 312436 19720 312484
rect 19680 312404 19684 312436
rect 19716 312404 19720 312436
rect 19680 312356 19720 312404
rect 19680 312324 19684 312356
rect 19716 312324 19720 312356
rect 19680 312276 19720 312324
rect 19680 312244 19684 312276
rect 19716 312244 19720 312276
rect 19680 312196 19720 312244
rect 19680 312164 19684 312196
rect 19716 312164 19720 312196
rect 19680 312116 19720 312164
rect 19680 312084 19684 312116
rect 19716 312084 19720 312116
rect 19680 312036 19720 312084
rect 19680 312004 19684 312036
rect 19716 312004 19720 312036
rect 19680 311956 19720 312004
rect 19680 311924 19684 311956
rect 19716 311924 19720 311956
rect 19680 311876 19720 311924
rect 19680 311844 19684 311876
rect 19716 311844 19720 311876
rect 19680 311796 19720 311844
rect 19680 311764 19684 311796
rect 19716 311764 19720 311796
rect 19680 311716 19720 311764
rect 19680 311684 19684 311716
rect 19716 311684 19720 311716
rect 19680 311636 19720 311684
rect 19680 311604 19684 311636
rect 19716 311604 19720 311636
rect 19680 311556 19720 311604
rect 19680 311524 19684 311556
rect 19716 311524 19720 311556
rect 19680 311476 19720 311524
rect 19680 311444 19684 311476
rect 19716 311444 19720 311476
rect 19680 311396 19720 311444
rect 19680 311364 19684 311396
rect 19716 311364 19720 311396
rect 19680 311316 19720 311364
rect 19680 311284 19684 311316
rect 19716 311284 19720 311316
rect 19680 311236 19720 311284
rect 19680 311204 19684 311236
rect 19716 311204 19720 311236
rect 19680 311156 19720 311204
rect 19680 311124 19684 311156
rect 19716 311124 19720 311156
rect 19680 311076 19720 311124
rect 19680 311044 19684 311076
rect 19716 311044 19720 311076
rect 19680 310996 19720 311044
rect 19680 310964 19684 310996
rect 19716 310964 19720 310996
rect 19680 310916 19720 310964
rect 19680 310884 19684 310916
rect 19716 310884 19720 310916
rect 19680 310836 19720 310884
rect 19680 310804 19684 310836
rect 19716 310804 19720 310836
rect 19680 310756 19720 310804
rect 19680 310724 19684 310756
rect 19716 310724 19720 310756
rect 19680 310676 19720 310724
rect 19680 310644 19684 310676
rect 19716 310644 19720 310676
rect 19680 310596 19720 310644
rect 19680 310564 19684 310596
rect 19716 310564 19720 310596
rect 19680 310516 19720 310564
rect 19680 310484 19684 310516
rect 19716 310484 19720 310516
rect 19680 310436 19720 310484
rect 19680 310404 19684 310436
rect 19716 310404 19720 310436
rect 19680 310356 19720 310404
rect 19680 310324 19684 310356
rect 19716 310324 19720 310356
rect 19680 310276 19720 310324
rect 19680 310244 19684 310276
rect 19716 310244 19720 310276
rect 19680 310196 19720 310244
rect 19680 310164 19684 310196
rect 19716 310164 19720 310196
rect 19680 310116 19720 310164
rect 19680 310084 19684 310116
rect 19716 310084 19720 310116
rect 19680 310036 19720 310084
rect 19680 310004 19684 310036
rect 19716 310004 19720 310036
rect 19680 309956 19720 310004
rect 19680 309924 19684 309956
rect 19716 309924 19720 309956
rect 19680 309876 19720 309924
rect 19680 309844 19684 309876
rect 19716 309844 19720 309876
rect 19680 309796 19720 309844
rect 19680 309764 19684 309796
rect 19716 309764 19720 309796
rect 19680 309716 19720 309764
rect 19680 309684 19684 309716
rect 19716 309684 19720 309716
rect 19680 309636 19720 309684
rect 19680 309604 19684 309636
rect 19716 309604 19720 309636
rect 19680 309556 19720 309604
rect 19680 309524 19684 309556
rect 19716 309524 19720 309556
rect 19680 309476 19720 309524
rect 19680 309444 19684 309476
rect 19716 309444 19720 309476
rect 19680 309396 19720 309444
rect 19680 309364 19684 309396
rect 19716 309364 19720 309396
rect 19680 309316 19720 309364
rect 19680 309284 19684 309316
rect 19716 309284 19720 309316
rect 19680 309236 19720 309284
rect 19680 309204 19684 309236
rect 19716 309204 19720 309236
rect 19680 309156 19720 309204
rect 19680 309124 19684 309156
rect 19716 309124 19720 309156
rect 19680 309076 19720 309124
rect 19680 309044 19684 309076
rect 19716 309044 19720 309076
rect 19680 308996 19720 309044
rect 19680 308964 19684 308996
rect 19716 308964 19720 308996
rect 19680 308916 19720 308964
rect 19680 308884 19684 308916
rect 19716 308884 19720 308916
rect 19680 308836 19720 308884
rect 19680 308804 19684 308836
rect 19716 308804 19720 308836
rect 19680 308756 19720 308804
rect 19680 308724 19684 308756
rect 19716 308724 19720 308756
rect 19680 308676 19720 308724
rect 19680 308644 19684 308676
rect 19716 308644 19720 308676
rect 19680 308596 19720 308644
rect 19680 308564 19684 308596
rect 19716 308564 19720 308596
rect 19680 308516 19720 308564
rect 19680 308484 19684 308516
rect 19716 308484 19720 308516
rect 19680 308436 19720 308484
rect 19680 308404 19684 308436
rect 19716 308404 19720 308436
rect 19680 308356 19720 308404
rect 19680 308324 19684 308356
rect 19716 308324 19720 308356
rect 19680 308276 19720 308324
rect 19680 308244 19684 308276
rect 19716 308244 19720 308276
rect 19680 308196 19720 308244
rect 19680 308164 19684 308196
rect 19716 308164 19720 308196
rect 19680 308116 19720 308164
rect 19680 308084 19684 308116
rect 19716 308084 19720 308116
rect 19680 308036 19720 308084
rect 19680 308004 19684 308036
rect 19716 308004 19720 308036
rect 19680 307956 19720 308004
rect 19680 307924 19684 307956
rect 19716 307924 19720 307956
rect 19680 307876 19720 307924
rect 19680 307844 19684 307876
rect 19716 307844 19720 307876
rect 19680 307796 19720 307844
rect 19680 307764 19684 307796
rect 19716 307764 19720 307796
rect 19680 307716 19720 307764
rect 19680 307684 19684 307716
rect 19716 307684 19720 307716
rect 19680 307636 19720 307684
rect 19680 307604 19684 307636
rect 19716 307604 19720 307636
rect 19680 307556 19720 307604
rect 19680 307524 19684 307556
rect 19716 307524 19720 307556
rect 19680 307476 19720 307524
rect 19680 307444 19684 307476
rect 19716 307444 19720 307476
rect 19680 307396 19720 307444
rect 19680 307364 19684 307396
rect 19716 307364 19720 307396
rect 19680 307316 19720 307364
rect 19680 307284 19684 307316
rect 19716 307284 19720 307316
rect 19680 307236 19720 307284
rect 19680 307204 19684 307236
rect 19716 307204 19720 307236
rect 19680 307156 19720 307204
rect 19680 307124 19684 307156
rect 19716 307124 19720 307156
rect 19680 307076 19720 307124
rect 19680 307044 19684 307076
rect 19716 307044 19720 307076
rect 19680 306996 19720 307044
rect 19680 306964 19684 306996
rect 19716 306964 19720 306996
rect 19680 306916 19720 306964
rect 19680 306884 19684 306916
rect 19716 306884 19720 306916
rect 19680 306836 19720 306884
rect 19680 306804 19684 306836
rect 19716 306804 19720 306836
rect 19680 306756 19720 306804
rect 19680 306724 19684 306756
rect 19716 306724 19720 306756
rect 19680 306676 19720 306724
rect 19680 306644 19684 306676
rect 19716 306644 19720 306676
rect 19680 306596 19720 306644
rect 19680 306564 19684 306596
rect 19716 306564 19720 306596
rect 19680 306516 19720 306564
rect 19680 306484 19684 306516
rect 19716 306484 19720 306516
rect 19680 306436 19720 306484
rect 19680 306404 19684 306436
rect 19716 306404 19720 306436
rect 19680 306356 19720 306404
rect 19680 306324 19684 306356
rect 19716 306324 19720 306356
rect 19680 306276 19720 306324
rect 19680 306244 19684 306276
rect 19716 306244 19720 306276
rect 19680 306196 19720 306244
rect 19680 306164 19684 306196
rect 19716 306164 19720 306196
rect 19680 306116 19720 306164
rect 19680 306084 19684 306116
rect 19716 306084 19720 306116
rect 19680 306036 19720 306084
rect 19680 306004 19684 306036
rect 19716 306004 19720 306036
rect 19680 305956 19720 306004
rect 19680 305924 19684 305956
rect 19716 305924 19720 305956
rect 19680 305876 19720 305924
rect 19680 305844 19684 305876
rect 19716 305844 19720 305876
rect 19680 305796 19720 305844
rect 19680 305764 19684 305796
rect 19716 305764 19720 305796
rect 19680 305716 19720 305764
rect 19680 305684 19684 305716
rect 19716 305684 19720 305716
rect 19680 305636 19720 305684
rect 19680 305604 19684 305636
rect 19716 305604 19720 305636
rect 19680 305556 19720 305604
rect 19680 305524 19684 305556
rect 19716 305524 19720 305556
rect 19680 305476 19720 305524
rect 19680 305444 19684 305476
rect 19716 305444 19720 305476
rect 19680 305396 19720 305444
rect 19680 305364 19684 305396
rect 19716 305364 19720 305396
rect 19680 305316 19720 305364
rect 19680 305284 19684 305316
rect 19716 305284 19720 305316
rect 19680 305236 19720 305284
rect 19680 305204 19684 305236
rect 19716 305204 19720 305236
rect 19680 305156 19720 305204
rect 19680 305124 19684 305156
rect 19716 305124 19720 305156
rect 19680 305076 19720 305124
rect 19680 305044 19684 305076
rect 19716 305044 19720 305076
rect 19680 304996 19720 305044
rect 19680 304964 19684 304996
rect 19716 304964 19720 304996
rect 19680 304916 19720 304964
rect 19680 304884 19684 304916
rect 19716 304884 19720 304916
rect 19680 304836 19720 304884
rect 19680 304804 19684 304836
rect 19716 304804 19720 304836
rect 19680 304756 19720 304804
rect 19680 304724 19684 304756
rect 19716 304724 19720 304756
rect 19680 304676 19720 304724
rect 19680 304644 19684 304676
rect 19716 304644 19720 304676
rect 19680 304596 19720 304644
rect 19680 304564 19684 304596
rect 19716 304564 19720 304596
rect 19680 304516 19720 304564
rect 19680 304484 19684 304516
rect 19716 304484 19720 304516
rect 19680 304436 19720 304484
rect 19680 304404 19684 304436
rect 19716 304404 19720 304436
rect 19680 304356 19720 304404
rect 19680 304324 19684 304356
rect 19716 304324 19720 304356
rect 19680 304276 19720 304324
rect 19680 304244 19684 304276
rect 19716 304244 19720 304276
rect 19680 304196 19720 304244
rect 19680 304164 19684 304196
rect 19716 304164 19720 304196
rect 19680 304116 19720 304164
rect 19680 304084 19684 304116
rect 19716 304084 19720 304116
rect 19680 304036 19720 304084
rect 19680 304004 19684 304036
rect 19716 304004 19720 304036
rect 19680 303956 19720 304004
rect 19680 303924 19684 303956
rect 19716 303924 19720 303956
rect 19680 303876 19720 303924
rect 19680 303844 19684 303876
rect 19716 303844 19720 303876
rect 19680 303796 19720 303844
rect 19680 303764 19684 303796
rect 19716 303764 19720 303796
rect 19680 303716 19720 303764
rect 19680 303684 19684 303716
rect 19716 303684 19720 303716
rect 19680 303636 19720 303684
rect 19680 303604 19684 303636
rect 19716 303604 19720 303636
rect 19680 303556 19720 303604
rect 19680 303524 19684 303556
rect 19716 303524 19720 303556
rect 19680 303476 19720 303524
rect 19680 303444 19684 303476
rect 19716 303444 19720 303476
rect 19680 303396 19720 303444
rect 19680 303364 19684 303396
rect 19716 303364 19720 303396
rect 19680 303316 19720 303364
rect 19680 303284 19684 303316
rect 19716 303284 19720 303316
rect 19680 303236 19720 303284
rect 19680 303204 19684 303236
rect 19716 303204 19720 303236
rect 19680 303156 19720 303204
rect 19680 303124 19684 303156
rect 19716 303124 19720 303156
rect 19680 303076 19720 303124
rect 19680 303044 19684 303076
rect 19716 303044 19720 303076
rect 19680 302996 19720 303044
rect 19680 302964 19684 302996
rect 19716 302964 19720 302996
rect 19680 302916 19720 302964
rect 19680 302884 19684 302916
rect 19716 302884 19720 302916
rect 19680 302836 19720 302884
rect 19680 302804 19684 302836
rect 19716 302804 19720 302836
rect 19680 302756 19720 302804
rect 19680 302724 19684 302756
rect 19716 302724 19720 302756
rect 19680 302676 19720 302724
rect 19680 302644 19684 302676
rect 19716 302644 19720 302676
rect 19680 302596 19720 302644
rect 19680 302564 19684 302596
rect 19716 302564 19720 302596
rect 19680 302516 19720 302564
rect 19680 302484 19684 302516
rect 19716 302484 19720 302516
rect 19680 302436 19720 302484
rect 19680 302404 19684 302436
rect 19716 302404 19720 302436
rect 19680 302356 19720 302404
rect 19680 302324 19684 302356
rect 19716 302324 19720 302356
rect 19680 302276 19720 302324
rect 19680 302244 19684 302276
rect 19716 302244 19720 302276
rect 19680 302196 19720 302244
rect 19680 302164 19684 302196
rect 19716 302164 19720 302196
rect 19680 302116 19720 302164
rect 19680 302084 19684 302116
rect 19716 302084 19720 302116
rect 19680 302036 19720 302084
rect 19680 302004 19684 302036
rect 19716 302004 19720 302036
rect 19680 301956 19720 302004
rect 19680 301924 19684 301956
rect 19716 301924 19720 301956
rect 19680 301876 19720 301924
rect 19680 301844 19684 301876
rect 19716 301844 19720 301876
rect 19680 301796 19720 301844
rect 19680 301764 19684 301796
rect 19716 301764 19720 301796
rect 19680 301716 19720 301764
rect 19680 301684 19684 301716
rect 19716 301684 19720 301716
rect 19680 301636 19720 301684
rect 19680 301604 19684 301636
rect 19716 301604 19720 301636
rect 19680 301556 19720 301604
rect 19680 301524 19684 301556
rect 19716 301524 19720 301556
rect 19680 301476 19720 301524
rect 19680 301444 19684 301476
rect 19716 301444 19720 301476
rect 19680 301396 19720 301444
rect 19680 301364 19684 301396
rect 19716 301364 19720 301396
rect 19680 301316 19720 301364
rect 19680 301284 19684 301316
rect 19716 301284 19720 301316
rect 19680 301236 19720 301284
rect 19680 301204 19684 301236
rect 19716 301204 19720 301236
rect 19680 301156 19720 301204
rect 19680 301124 19684 301156
rect 19716 301124 19720 301156
rect 19680 301076 19720 301124
rect 19680 301044 19684 301076
rect 19716 301044 19720 301076
rect 19680 300996 19720 301044
rect 19680 300964 19684 300996
rect 19716 300964 19720 300996
rect 19680 300916 19720 300964
rect 19680 300884 19684 300916
rect 19716 300884 19720 300916
rect 19680 300836 19720 300884
rect 19680 300804 19684 300836
rect 19716 300804 19720 300836
rect 19680 300756 19720 300804
rect 19680 300724 19684 300756
rect 19716 300724 19720 300756
rect 19680 300676 19720 300724
rect 19680 300644 19684 300676
rect 19716 300644 19720 300676
rect 19680 300596 19720 300644
rect 19680 300564 19684 300596
rect 19716 300564 19720 300596
rect 19680 300516 19720 300564
rect 19680 300484 19684 300516
rect 19716 300484 19720 300516
rect 19680 300436 19720 300484
rect 19680 300404 19684 300436
rect 19716 300404 19720 300436
rect 19680 300356 19720 300404
rect 19680 300324 19684 300356
rect 19716 300324 19720 300356
rect 19680 300276 19720 300324
rect 19680 300244 19684 300276
rect 19716 300244 19720 300276
rect 19680 300196 19720 300244
rect 19680 300164 19684 300196
rect 19716 300164 19720 300196
rect 19680 300116 19720 300164
rect 19680 300084 19684 300116
rect 19716 300084 19720 300116
rect 19680 300036 19720 300084
rect 19680 300004 19684 300036
rect 19716 300004 19720 300036
rect 19680 299956 19720 300004
rect 19680 299924 19684 299956
rect 19716 299924 19720 299956
rect 19680 299876 19720 299924
rect 19680 299844 19684 299876
rect 19716 299844 19720 299876
rect 19680 299796 19720 299844
rect 19680 299764 19684 299796
rect 19716 299764 19720 299796
rect 19680 299716 19720 299764
rect 19680 299684 19684 299716
rect 19716 299684 19720 299716
rect 19680 299636 19720 299684
rect 19680 299604 19684 299636
rect 19716 299604 19720 299636
rect 19680 299556 19720 299604
rect 19680 299524 19684 299556
rect 19716 299524 19720 299556
rect 19680 299476 19720 299524
rect 19680 299444 19684 299476
rect 19716 299444 19720 299476
rect 19680 299396 19720 299444
rect 19680 299364 19684 299396
rect 19716 299364 19720 299396
rect 19680 299316 19720 299364
rect 19680 299284 19684 299316
rect 19716 299284 19720 299316
rect 19680 299236 19720 299284
rect 19680 299204 19684 299236
rect 19716 299204 19720 299236
rect 19680 299156 19720 299204
rect 19680 299124 19684 299156
rect 19716 299124 19720 299156
rect 19680 299076 19720 299124
rect 19680 299044 19684 299076
rect 19716 299044 19720 299076
rect 19680 298996 19720 299044
rect 19680 298964 19684 298996
rect 19716 298964 19720 298996
rect 19680 298916 19720 298964
rect 19680 298884 19684 298916
rect 19716 298884 19720 298916
rect 19680 298836 19720 298884
rect 19680 298804 19684 298836
rect 19716 298804 19720 298836
rect 19680 298756 19720 298804
rect 19680 298724 19684 298756
rect 19716 298724 19720 298756
rect 19680 298676 19720 298724
rect 19680 298644 19684 298676
rect 19716 298644 19720 298676
rect 19680 298596 19720 298644
rect 19680 298564 19684 298596
rect 19716 298564 19720 298596
rect 19680 298516 19720 298564
rect 19680 298484 19684 298516
rect 19716 298484 19720 298516
rect 19680 298436 19720 298484
rect 19680 298404 19684 298436
rect 19716 298404 19720 298436
rect 19680 298356 19720 298404
rect 19680 298324 19684 298356
rect 19716 298324 19720 298356
rect 19680 298276 19720 298324
rect 19680 298244 19684 298276
rect 19716 298244 19720 298276
rect 19680 298196 19720 298244
rect 19680 298164 19684 298196
rect 19716 298164 19720 298196
rect 19680 298116 19720 298164
rect 19680 298084 19684 298116
rect 19716 298084 19720 298116
rect 19680 298036 19720 298084
rect 19680 298004 19684 298036
rect 19716 298004 19720 298036
rect 19680 297956 19720 298004
rect 19680 297924 19684 297956
rect 19716 297924 19720 297956
rect 19680 297876 19720 297924
rect 19680 297844 19684 297876
rect 19716 297844 19720 297876
rect 19680 297796 19720 297844
rect 19680 297764 19684 297796
rect 19716 297764 19720 297796
rect 19680 297716 19720 297764
rect 19680 297684 19684 297716
rect 19716 297684 19720 297716
rect 19680 297636 19720 297684
rect 19680 297604 19684 297636
rect 19716 297604 19720 297636
rect 19680 297556 19720 297604
rect 19680 297524 19684 297556
rect 19716 297524 19720 297556
rect 19680 297476 19720 297524
rect 19680 297444 19684 297476
rect 19716 297444 19720 297476
rect 19680 297396 19720 297444
rect 19680 297364 19684 297396
rect 19716 297364 19720 297396
rect 19680 297316 19720 297364
rect 19680 297284 19684 297316
rect 19716 297284 19720 297316
rect 19680 297236 19720 297284
rect 19680 297204 19684 297236
rect 19716 297204 19720 297236
rect 19680 297156 19720 297204
rect 19680 297124 19684 297156
rect 19716 297124 19720 297156
rect 19680 297076 19720 297124
rect 19680 297044 19684 297076
rect 19716 297044 19720 297076
rect 19680 296996 19720 297044
rect 19680 296964 19684 296996
rect 19716 296964 19720 296996
rect 19680 296916 19720 296964
rect 19680 296884 19684 296916
rect 19716 296884 19720 296916
rect 19680 296836 19720 296884
rect 19680 296804 19684 296836
rect 19716 296804 19720 296836
rect 19680 296756 19720 296804
rect 19680 296724 19684 296756
rect 19716 296724 19720 296756
rect 19680 296676 19720 296724
rect 19680 296644 19684 296676
rect 19716 296644 19720 296676
rect 19680 296596 19720 296644
rect 19680 296564 19684 296596
rect 19716 296564 19720 296596
rect 19680 296516 19720 296564
rect 19680 296484 19684 296516
rect 19716 296484 19720 296516
rect 19680 296436 19720 296484
rect 19680 296404 19684 296436
rect 19716 296404 19720 296436
rect 19680 296356 19720 296404
rect 19680 296324 19684 296356
rect 19716 296324 19720 296356
rect 19680 296276 19720 296324
rect 19680 296244 19684 296276
rect 19716 296244 19720 296276
rect 19680 296196 19720 296244
rect 19680 296164 19684 296196
rect 19716 296164 19720 296196
rect 19680 296116 19720 296164
rect 19680 296084 19684 296116
rect 19716 296084 19720 296116
rect 19680 296036 19720 296084
rect 19680 296004 19684 296036
rect 19716 296004 19720 296036
rect 19680 295956 19720 296004
rect 19680 295924 19684 295956
rect 19716 295924 19720 295956
rect 19680 295876 19720 295924
rect 19680 295844 19684 295876
rect 19716 295844 19720 295876
rect 19680 295796 19720 295844
rect 19680 295764 19684 295796
rect 19716 295764 19720 295796
rect 19680 295716 19720 295764
rect 19680 295684 19684 295716
rect 19716 295684 19720 295716
rect 19680 295636 19720 295684
rect 19680 295604 19684 295636
rect 19716 295604 19720 295636
rect 19680 295556 19720 295604
rect 19680 295524 19684 295556
rect 19716 295524 19720 295556
rect 19680 295476 19720 295524
rect 19680 295444 19684 295476
rect 19716 295444 19720 295476
rect 19680 295396 19720 295444
rect 19680 295364 19684 295396
rect 19716 295364 19720 295396
rect 19680 295316 19720 295364
rect 19680 295284 19684 295316
rect 19716 295284 19720 295316
rect 19680 295236 19720 295284
rect 19680 295204 19684 295236
rect 19716 295204 19720 295236
rect 19680 295156 19720 295204
rect 19680 295124 19684 295156
rect 19716 295124 19720 295156
rect 19680 295076 19720 295124
rect 19680 295044 19684 295076
rect 19716 295044 19720 295076
rect 19680 294996 19720 295044
rect 19680 294964 19684 294996
rect 19716 294964 19720 294996
rect 19680 294916 19720 294964
rect 19680 294884 19684 294916
rect 19716 294884 19720 294916
rect 19680 294836 19720 294884
rect 19680 294804 19684 294836
rect 19716 294804 19720 294836
rect 19680 294756 19720 294804
rect 19680 294724 19684 294756
rect 19716 294724 19720 294756
rect 19680 294676 19720 294724
rect 19680 294644 19684 294676
rect 19716 294644 19720 294676
rect 19680 294596 19720 294644
rect 19680 294564 19684 294596
rect 19716 294564 19720 294596
rect 19680 294516 19720 294564
rect 19680 294484 19684 294516
rect 19716 294484 19720 294516
rect 19680 294436 19720 294484
rect 19680 294404 19684 294436
rect 19716 294404 19720 294436
rect 19680 294356 19720 294404
rect 19680 294324 19684 294356
rect 19716 294324 19720 294356
rect 19680 294276 19720 294324
rect 19680 294244 19684 294276
rect 19716 294244 19720 294276
rect 19680 294196 19720 294244
rect 19680 294164 19684 294196
rect 19716 294164 19720 294196
rect 19680 294116 19720 294164
rect 19680 294084 19684 294116
rect 19716 294084 19720 294116
rect 19680 294036 19720 294084
rect 19680 294004 19684 294036
rect 19716 294004 19720 294036
rect 19680 293956 19720 294004
rect 19680 293924 19684 293956
rect 19716 293924 19720 293956
rect 19680 293876 19720 293924
rect 19680 293844 19684 293876
rect 19716 293844 19720 293876
rect 19680 293796 19720 293844
rect 19680 293764 19684 293796
rect 19716 293764 19720 293796
rect 19680 293716 19720 293764
rect 19680 293684 19684 293716
rect 19716 293684 19720 293716
rect 19680 293636 19720 293684
rect 19680 293604 19684 293636
rect 19716 293604 19720 293636
rect 19680 293556 19720 293604
rect 19680 293524 19684 293556
rect 19716 293524 19720 293556
rect 19680 293476 19720 293524
rect 19680 293444 19684 293476
rect 19716 293444 19720 293476
rect 19680 293396 19720 293444
rect 19680 293364 19684 293396
rect 19716 293364 19720 293396
rect 19680 293316 19720 293364
rect 19680 293284 19684 293316
rect 19716 293284 19720 293316
rect 19680 293236 19720 293284
rect 19680 293204 19684 293236
rect 19716 293204 19720 293236
rect 19680 293156 19720 293204
rect 19680 293124 19684 293156
rect 19716 293124 19720 293156
rect 19680 293076 19720 293124
rect 19680 293044 19684 293076
rect 19716 293044 19720 293076
rect 19680 292996 19720 293044
rect 19680 292964 19684 292996
rect 19716 292964 19720 292996
rect 19680 292916 19720 292964
rect 19680 292884 19684 292916
rect 19716 292884 19720 292916
rect 19680 292836 19720 292884
rect 19680 292804 19684 292836
rect 19716 292804 19720 292836
rect 19680 292756 19720 292804
rect 19680 292724 19684 292756
rect 19716 292724 19720 292756
rect 19680 292676 19720 292724
rect 19680 292644 19684 292676
rect 19716 292644 19720 292676
rect 19680 292596 19720 292644
rect 19680 292564 19684 292596
rect 19716 292564 19720 292596
rect 19680 292516 19720 292564
rect 19680 292484 19684 292516
rect 19716 292484 19720 292516
rect 19680 292436 19720 292484
rect 19680 292404 19684 292436
rect 19716 292404 19720 292436
rect 19680 292356 19720 292404
rect 19680 292324 19684 292356
rect 19716 292324 19720 292356
rect 19680 292276 19720 292324
rect 19680 292244 19684 292276
rect 19716 292244 19720 292276
rect 19680 292196 19720 292244
rect 19680 292164 19684 292196
rect 19716 292164 19720 292196
rect 19680 292116 19720 292164
rect 19680 292084 19684 292116
rect 19716 292084 19720 292116
rect 19680 292036 19720 292084
rect 19680 292004 19684 292036
rect 19716 292004 19720 292036
rect 19680 291956 19720 292004
rect 19680 291924 19684 291956
rect 19716 291924 19720 291956
rect 19680 291876 19720 291924
rect 19680 291844 19684 291876
rect 19716 291844 19720 291876
rect 19680 291796 19720 291844
rect 19680 291764 19684 291796
rect 19716 291764 19720 291796
rect 19680 291716 19720 291764
rect 19680 291684 19684 291716
rect 19716 291684 19720 291716
rect 19680 291636 19720 291684
rect 19680 291604 19684 291636
rect 19716 291604 19720 291636
rect 19680 291556 19720 291604
rect 19680 291524 19684 291556
rect 19716 291524 19720 291556
rect 19680 291476 19720 291524
rect 19680 291444 19684 291476
rect 19716 291444 19720 291476
rect 19680 291396 19720 291444
rect 19680 291364 19684 291396
rect 19716 291364 19720 291396
rect 19680 291316 19720 291364
rect 19680 291284 19684 291316
rect 19716 291284 19720 291316
rect 19680 291236 19720 291284
rect 19680 291204 19684 291236
rect 19716 291204 19720 291236
rect 19680 291156 19720 291204
rect 19680 291124 19684 291156
rect 19716 291124 19720 291156
rect 19680 291076 19720 291124
rect 19680 291044 19684 291076
rect 19716 291044 19720 291076
rect 19680 290996 19720 291044
rect 19680 290964 19684 290996
rect 19716 290964 19720 290996
rect 19680 290916 19720 290964
rect 19680 290884 19684 290916
rect 19716 290884 19720 290916
rect 19680 290836 19720 290884
rect 19680 290804 19684 290836
rect 19716 290804 19720 290836
rect 19680 290756 19720 290804
rect 19680 290724 19684 290756
rect 19716 290724 19720 290756
rect 19680 290676 19720 290724
rect 19680 290644 19684 290676
rect 19716 290644 19720 290676
rect 19680 290596 19720 290644
rect 19680 290564 19684 290596
rect 19716 290564 19720 290596
rect 19680 290516 19720 290564
rect 19680 290484 19684 290516
rect 19716 290484 19720 290516
rect 19680 290436 19720 290484
rect 19680 290404 19684 290436
rect 19716 290404 19720 290436
rect 19680 290356 19720 290404
rect 19680 290324 19684 290356
rect 19716 290324 19720 290356
rect 19680 290276 19720 290324
rect 19680 290244 19684 290276
rect 19716 290244 19720 290276
rect 19680 290196 19720 290244
rect 19680 290164 19684 290196
rect 19716 290164 19720 290196
rect 19680 290116 19720 290164
rect 19680 290084 19684 290116
rect 19716 290084 19720 290116
rect 19680 290036 19720 290084
rect 19680 290004 19684 290036
rect 19716 290004 19720 290036
rect 19680 289956 19720 290004
rect 19680 289924 19684 289956
rect 19716 289924 19720 289956
rect 19680 289876 19720 289924
rect 19680 289844 19684 289876
rect 19716 289844 19720 289876
rect 19680 289796 19720 289844
rect 19680 289764 19684 289796
rect 19716 289764 19720 289796
rect 19680 289716 19720 289764
rect 19680 289684 19684 289716
rect 19716 289684 19720 289716
rect 19680 289636 19720 289684
rect 19680 289604 19684 289636
rect 19716 289604 19720 289636
rect 19680 289556 19720 289604
rect 19680 289524 19684 289556
rect 19716 289524 19720 289556
rect 19680 289476 19720 289524
rect 19680 289444 19684 289476
rect 19716 289444 19720 289476
rect 19680 289396 19720 289444
rect 19680 289364 19684 289396
rect 19716 289364 19720 289396
rect 19680 289316 19720 289364
rect 19680 289284 19684 289316
rect 19716 289284 19720 289316
rect 19680 289236 19720 289284
rect 19680 289204 19684 289236
rect 19716 289204 19720 289236
rect 19680 289156 19720 289204
rect 19680 289124 19684 289156
rect 19716 289124 19720 289156
rect 19680 289076 19720 289124
rect 19680 289044 19684 289076
rect 19716 289044 19720 289076
rect 19680 288996 19720 289044
rect 19680 288964 19684 288996
rect 19716 288964 19720 288996
rect 19680 288916 19720 288964
rect 19680 288884 19684 288916
rect 19716 288884 19720 288916
rect 19680 288836 19720 288884
rect 19680 288804 19684 288836
rect 19716 288804 19720 288836
rect 19680 288756 19720 288804
rect 19680 288724 19684 288756
rect 19716 288724 19720 288756
rect 19680 288676 19720 288724
rect 19680 288644 19684 288676
rect 19716 288644 19720 288676
rect 19680 288596 19720 288644
rect 19680 288564 19684 288596
rect 19716 288564 19720 288596
rect 19680 288516 19720 288564
rect 19680 288484 19684 288516
rect 19716 288484 19720 288516
rect 19680 288436 19720 288484
rect 19680 288404 19684 288436
rect 19716 288404 19720 288436
rect 19680 288356 19720 288404
rect 19680 288324 19684 288356
rect 19716 288324 19720 288356
rect 19680 288276 19720 288324
rect 19680 288244 19684 288276
rect 19716 288244 19720 288276
rect 19680 288196 19720 288244
rect 19680 288164 19684 288196
rect 19716 288164 19720 288196
rect 19680 288116 19720 288164
rect 19680 288084 19684 288116
rect 19716 288084 19720 288116
rect 19680 288036 19720 288084
rect 19680 288004 19684 288036
rect 19716 288004 19720 288036
rect 19680 287956 19720 288004
rect 19680 287924 19684 287956
rect 19716 287924 19720 287956
rect 19680 287876 19720 287924
rect 19680 287844 19684 287876
rect 19716 287844 19720 287876
rect 19680 287796 19720 287844
rect 19680 287764 19684 287796
rect 19716 287764 19720 287796
rect 19680 287716 19720 287764
rect 19680 287684 19684 287716
rect 19716 287684 19720 287716
rect 19680 287636 19720 287684
rect 19680 287604 19684 287636
rect 19716 287604 19720 287636
rect 19680 287556 19720 287604
rect 19680 287524 19684 287556
rect 19716 287524 19720 287556
rect 19680 287476 19720 287524
rect 19680 287444 19684 287476
rect 19716 287444 19720 287476
rect 19680 287396 19720 287444
rect 19680 287364 19684 287396
rect 19716 287364 19720 287396
rect 19680 287316 19720 287364
rect 19680 287284 19684 287316
rect 19716 287284 19720 287316
rect 19680 287236 19720 287284
rect 19680 287204 19684 287236
rect 19716 287204 19720 287236
rect 19680 287156 19720 287204
rect 19680 287124 19684 287156
rect 19716 287124 19720 287156
rect 19680 287076 19720 287124
rect 19680 287044 19684 287076
rect 19716 287044 19720 287076
rect 19680 286996 19720 287044
rect 19680 286964 19684 286996
rect 19716 286964 19720 286996
rect 19680 286916 19720 286964
rect 19680 286884 19684 286916
rect 19716 286884 19720 286916
rect 19680 286836 19720 286884
rect 19680 286804 19684 286836
rect 19716 286804 19720 286836
rect 19680 286756 19720 286804
rect 19680 286724 19684 286756
rect 19716 286724 19720 286756
rect 19680 286676 19720 286724
rect 19680 286644 19684 286676
rect 19716 286644 19720 286676
rect 19680 286596 19720 286644
rect 19680 286564 19684 286596
rect 19716 286564 19720 286596
rect 19680 286516 19720 286564
rect 19680 286484 19684 286516
rect 19716 286484 19720 286516
rect 19680 286436 19720 286484
rect 19680 286404 19684 286436
rect 19716 286404 19720 286436
rect 19680 286356 19720 286404
rect 19680 286324 19684 286356
rect 19716 286324 19720 286356
rect 19680 286276 19720 286324
rect 19680 286244 19684 286276
rect 19716 286244 19720 286276
rect 19680 286196 19720 286244
rect 19680 286164 19684 286196
rect 19716 286164 19720 286196
rect 19680 286116 19720 286164
rect 19680 286084 19684 286116
rect 19716 286084 19720 286116
rect 19680 286036 19720 286084
rect 19680 286004 19684 286036
rect 19716 286004 19720 286036
rect 19680 285956 19720 286004
rect 19680 285924 19684 285956
rect 19716 285924 19720 285956
rect 19680 285876 19720 285924
rect 19680 285844 19684 285876
rect 19716 285844 19720 285876
rect 19680 285796 19720 285844
rect 19680 285764 19684 285796
rect 19716 285764 19720 285796
rect 19680 285716 19720 285764
rect 19680 285684 19684 285716
rect 19716 285684 19720 285716
rect 19680 285636 19720 285684
rect 19680 285604 19684 285636
rect 19716 285604 19720 285636
rect 19680 285556 19720 285604
rect 19680 285524 19684 285556
rect 19716 285524 19720 285556
rect 19680 285476 19720 285524
rect 19680 285444 19684 285476
rect 19716 285444 19720 285476
rect 19680 285396 19720 285444
rect 19680 285364 19684 285396
rect 19716 285364 19720 285396
rect 19680 285316 19720 285364
rect 19680 285284 19684 285316
rect 19716 285284 19720 285316
rect 19680 285236 19720 285284
rect 19680 285204 19684 285236
rect 19716 285204 19720 285236
rect 19680 285156 19720 285204
rect 19680 285124 19684 285156
rect 19716 285124 19720 285156
rect 19680 285076 19720 285124
rect 19680 285044 19684 285076
rect 19716 285044 19720 285076
rect 19680 284996 19720 285044
rect 19680 284964 19684 284996
rect 19716 284964 19720 284996
rect 19680 284916 19720 284964
rect 19680 284884 19684 284916
rect 19716 284884 19720 284916
rect 19680 284836 19720 284884
rect 19680 284804 19684 284836
rect 19716 284804 19720 284836
rect 19680 284756 19720 284804
rect 19680 284724 19684 284756
rect 19716 284724 19720 284756
rect 19680 284676 19720 284724
rect 19680 284644 19684 284676
rect 19716 284644 19720 284676
rect 19680 284596 19720 284644
rect 19680 284564 19684 284596
rect 19716 284564 19720 284596
rect 19680 284516 19720 284564
rect 19680 284484 19684 284516
rect 19716 284484 19720 284516
rect 19680 284436 19720 284484
rect 19680 284404 19684 284436
rect 19716 284404 19720 284436
rect 19680 284356 19720 284404
rect 19680 284324 19684 284356
rect 19716 284324 19720 284356
rect 19680 284276 19720 284324
rect 19680 284244 19684 284276
rect 19716 284244 19720 284276
rect 19680 284196 19720 284244
rect 19680 284164 19684 284196
rect 19716 284164 19720 284196
rect 19680 284116 19720 284164
rect 19680 284084 19684 284116
rect 19716 284084 19720 284116
rect 19680 284036 19720 284084
rect 19680 284004 19684 284036
rect 19716 284004 19720 284036
rect 19680 283956 19720 284004
rect 19680 283924 19684 283956
rect 19716 283924 19720 283956
rect 19680 283876 19720 283924
rect 19680 283844 19684 283876
rect 19716 283844 19720 283876
rect 19680 283796 19720 283844
rect 19680 283764 19684 283796
rect 19716 283764 19720 283796
rect 19680 283716 19720 283764
rect 19680 283684 19684 283716
rect 19716 283684 19720 283716
rect 19680 283636 19720 283684
rect 19680 283604 19684 283636
rect 19716 283604 19720 283636
rect 19680 283556 19720 283604
rect 19680 283524 19684 283556
rect 19716 283524 19720 283556
rect 19680 283476 19720 283524
rect 19680 283444 19684 283476
rect 19716 283444 19720 283476
rect 19680 283396 19720 283444
rect 19680 283364 19684 283396
rect 19716 283364 19720 283396
rect 19680 283316 19720 283364
rect 19680 283284 19684 283316
rect 19716 283284 19720 283316
rect 19680 283236 19720 283284
rect 19680 283204 19684 283236
rect 19716 283204 19720 283236
rect 19680 283156 19720 283204
rect 19680 283124 19684 283156
rect 19716 283124 19720 283156
rect 19680 283076 19720 283124
rect 19680 283044 19684 283076
rect 19716 283044 19720 283076
rect 19680 282996 19720 283044
rect 19680 282964 19684 282996
rect 19716 282964 19720 282996
rect 19680 282916 19720 282964
rect 19680 282884 19684 282916
rect 19716 282884 19720 282916
rect 19680 282836 19720 282884
rect 19680 282804 19684 282836
rect 19716 282804 19720 282836
rect 19680 282756 19720 282804
rect 19680 282724 19684 282756
rect 19716 282724 19720 282756
rect 19680 282676 19720 282724
rect 19680 282644 19684 282676
rect 19716 282644 19720 282676
rect 19680 282596 19720 282644
rect 19680 282564 19684 282596
rect 19716 282564 19720 282596
rect 19680 282516 19720 282564
rect 19680 282484 19684 282516
rect 19716 282484 19720 282516
rect 19680 282436 19720 282484
rect 19680 282404 19684 282436
rect 19716 282404 19720 282436
rect 19680 282356 19720 282404
rect 19680 282324 19684 282356
rect 19716 282324 19720 282356
rect 19680 282276 19720 282324
rect 19680 282244 19684 282276
rect 19716 282244 19720 282276
rect 19680 282196 19720 282244
rect 19680 282164 19684 282196
rect 19716 282164 19720 282196
rect 19680 282116 19720 282164
rect 19680 282084 19684 282116
rect 19716 282084 19720 282116
rect 19680 282036 19720 282084
rect 19680 282004 19684 282036
rect 19716 282004 19720 282036
rect 19680 281956 19720 282004
rect 19680 281924 19684 281956
rect 19716 281924 19720 281956
rect 19680 281876 19720 281924
rect 19680 281844 19684 281876
rect 19716 281844 19720 281876
rect 19680 281796 19720 281844
rect 19680 281764 19684 281796
rect 19716 281764 19720 281796
rect 19680 281716 19720 281764
rect 19680 281684 19684 281716
rect 19716 281684 19720 281716
rect 19680 281636 19720 281684
rect 19680 281604 19684 281636
rect 19716 281604 19720 281636
rect 19680 281556 19720 281604
rect 19680 281524 19684 281556
rect 19716 281524 19720 281556
rect 19680 281476 19720 281524
rect 19680 281444 19684 281476
rect 19716 281444 19720 281476
rect 19680 281396 19720 281444
rect 19680 281364 19684 281396
rect 19716 281364 19720 281396
rect 19680 281316 19720 281364
rect 19680 281284 19684 281316
rect 19716 281284 19720 281316
rect 19680 281236 19720 281284
rect 19680 281204 19684 281236
rect 19716 281204 19720 281236
rect 19680 281156 19720 281204
rect 19680 281124 19684 281156
rect 19716 281124 19720 281156
rect 19680 281076 19720 281124
rect 19680 281044 19684 281076
rect 19716 281044 19720 281076
rect 19680 280996 19720 281044
rect 19680 280964 19684 280996
rect 19716 280964 19720 280996
rect 19680 280916 19720 280964
rect 19680 280884 19684 280916
rect 19716 280884 19720 280916
rect 19680 280836 19720 280884
rect 19680 280804 19684 280836
rect 19716 280804 19720 280836
rect 19680 280756 19720 280804
rect 19680 280724 19684 280756
rect 19716 280724 19720 280756
rect 19680 280676 19720 280724
rect 19680 280644 19684 280676
rect 19716 280644 19720 280676
rect 19680 280596 19720 280644
rect 19680 280564 19684 280596
rect 19716 280564 19720 280596
rect 19680 280516 19720 280564
rect 19680 280484 19684 280516
rect 19716 280484 19720 280516
rect 19680 280436 19720 280484
rect 19680 280404 19684 280436
rect 19716 280404 19720 280436
rect 19680 280356 19720 280404
rect 19680 280324 19684 280356
rect 19716 280324 19720 280356
rect 19680 280276 19720 280324
rect 19680 280244 19684 280276
rect 19716 280244 19720 280276
rect 19680 280196 19720 280244
rect 19680 280164 19684 280196
rect 19716 280164 19720 280196
rect 19680 280116 19720 280164
rect 19680 280084 19684 280116
rect 19716 280084 19720 280116
rect 19680 280036 19720 280084
rect 19680 280004 19684 280036
rect 19716 280004 19720 280036
rect 19680 279956 19720 280004
rect 19680 279924 19684 279956
rect 19716 279924 19720 279956
rect 19680 279876 19720 279924
rect 19680 279844 19684 279876
rect 19716 279844 19720 279876
rect 19680 279796 19720 279844
rect 19680 279764 19684 279796
rect 19716 279764 19720 279796
rect 19680 279716 19720 279764
rect 19680 279684 19684 279716
rect 19716 279684 19720 279716
rect 19680 279636 19720 279684
rect 19680 279604 19684 279636
rect 19716 279604 19720 279636
rect 19680 279556 19720 279604
rect 19680 279524 19684 279556
rect 19716 279524 19720 279556
rect 19680 279476 19720 279524
rect 19680 279444 19684 279476
rect 19716 279444 19720 279476
rect 2400 279350 2600 279400
rect 2400 279250 2450 279350
rect 2550 279250 2600 279350
rect -400 275500 830 277121
rect -400 275300 850 275500
rect -400 275200 830 275300
rect -400 275160 1200 275200
rect -400 275040 1040 275160
rect 1160 275040 1200 275160
rect -400 275000 1200 275040
rect -400 274721 830 275000
rect 2400 263200 2600 279250
rect 19680 279396 19720 279444
rect 19680 279364 19684 279396
rect 19716 279364 19720 279396
rect 19680 279316 19720 279364
rect 19680 279284 19684 279316
rect 19716 279284 19720 279316
rect 19680 279236 19720 279284
rect 19680 279204 19684 279236
rect 19716 279204 19720 279236
rect 14200 275800 14400 279200
rect 19680 279156 19720 279204
rect 19680 279124 19684 279156
rect 19716 279124 19720 279156
rect 19680 279076 19720 279124
rect 19680 279044 19684 279076
rect 19716 279044 19720 279076
rect 19680 278996 19720 279044
rect 19680 278964 19684 278996
rect 19716 278964 19720 278996
rect 19680 278916 19720 278964
rect 19680 278884 19684 278916
rect 19716 278884 19720 278916
rect 19680 278836 19720 278884
rect 19680 278804 19684 278836
rect 19716 278804 19720 278836
rect 19680 278756 19720 278804
rect 19680 278724 19684 278756
rect 19716 278724 19720 278756
rect 17040 278676 17080 278680
rect 17040 278644 17044 278676
rect 17076 278644 17080 278676
rect 17040 278596 17080 278644
rect 17200 278676 17240 278680
rect 17200 278644 17204 278676
rect 17236 278644 17240 278676
rect 17040 278564 17044 278596
rect 17076 278564 17080 278596
rect 17040 278516 17080 278564
rect 17040 278484 17044 278516
rect 17076 278484 17080 278516
rect 17040 278436 17080 278484
rect 17040 278404 17044 278436
rect 17076 278404 17080 278436
rect 17040 278356 17080 278404
rect 17040 278324 17044 278356
rect 17076 278324 17080 278356
rect 17040 278276 17080 278324
rect 17040 278244 17044 278276
rect 17076 278244 17080 278276
rect 17040 278196 17080 278244
rect 17040 278164 17044 278196
rect 17076 278164 17080 278196
rect 17040 278116 17080 278164
rect 17040 278084 17044 278116
rect 17076 278084 17080 278116
rect 17040 278036 17080 278084
rect 17040 278004 17044 278036
rect 17076 278004 17080 278036
rect 17040 277956 17080 278004
rect 17040 277924 17044 277956
rect 17076 277924 17080 277956
rect 17040 277876 17080 277924
rect 17040 277844 17044 277876
rect 17076 277844 17080 277876
rect 17040 277800 17080 277844
rect 17120 278595 17160 278600
rect 17120 278565 17125 278595
rect 17155 278565 17160 278595
rect 17120 277800 17160 278565
rect 17200 278596 17240 278644
rect 17200 278564 17204 278596
rect 17236 278564 17240 278596
rect 17200 278516 17240 278564
rect 17200 278484 17204 278516
rect 17236 278484 17240 278516
rect 17200 278436 17240 278484
rect 17280 278676 17320 278680
rect 17280 278644 17284 278676
rect 17316 278644 17320 278676
rect 17280 278596 17320 278644
rect 17280 278564 17284 278596
rect 17316 278564 17320 278596
rect 17280 278516 17320 278564
rect 17280 278484 17284 278516
rect 17316 278484 17320 278516
rect 17280 278480 17320 278484
rect 17360 278676 17400 278680
rect 17360 278644 17364 278676
rect 17396 278644 17400 278676
rect 17360 278596 17400 278644
rect 17360 278564 17364 278596
rect 17396 278564 17400 278596
rect 17360 278516 17400 278564
rect 17360 278484 17364 278516
rect 17396 278484 17400 278516
rect 17360 278480 17400 278484
rect 17440 278676 17480 278680
rect 17440 278644 17444 278676
rect 17476 278644 17480 278676
rect 17440 278596 17480 278644
rect 17440 278564 17444 278596
rect 17476 278564 17480 278596
rect 17440 278516 17480 278564
rect 17440 278484 17444 278516
rect 17476 278484 17480 278516
rect 17440 278480 17480 278484
rect 17520 278676 17560 278680
rect 17520 278644 17524 278676
rect 17556 278644 17560 278676
rect 17520 278596 17560 278644
rect 17520 278564 17524 278596
rect 17556 278564 17560 278596
rect 17520 278516 17560 278564
rect 17520 278484 17524 278516
rect 17556 278484 17560 278516
rect 17520 278480 17560 278484
rect 17600 278676 17640 278680
rect 17600 278644 17604 278676
rect 17636 278644 17640 278676
rect 17600 278596 17640 278644
rect 17600 278564 17604 278596
rect 17636 278564 17640 278596
rect 17600 278516 17640 278564
rect 17600 278484 17604 278516
rect 17636 278484 17640 278516
rect 17600 278480 17640 278484
rect 17680 278676 17720 278680
rect 17680 278644 17684 278676
rect 17716 278644 17720 278676
rect 17680 278596 17720 278644
rect 17680 278564 17684 278596
rect 17716 278564 17720 278596
rect 17680 278516 17720 278564
rect 17680 278484 17684 278516
rect 17716 278484 17720 278516
rect 17680 278480 17720 278484
rect 17760 278676 17800 278680
rect 17760 278644 17764 278676
rect 17796 278644 17800 278676
rect 17760 278596 17800 278644
rect 17760 278564 17764 278596
rect 17796 278564 17800 278596
rect 17760 278516 17800 278564
rect 17760 278484 17764 278516
rect 17796 278484 17800 278516
rect 17760 278480 17800 278484
rect 19520 278676 19560 278680
rect 19520 278644 19524 278676
rect 19556 278644 19560 278676
rect 19520 278596 19560 278644
rect 19520 278564 19524 278596
rect 19556 278564 19560 278596
rect 19520 278516 19560 278564
rect 19520 278484 19524 278516
rect 19556 278484 19560 278516
rect 19520 278480 19560 278484
rect 19600 278676 19640 278680
rect 19600 278644 19604 278676
rect 19636 278644 19640 278676
rect 19600 278596 19640 278644
rect 19600 278564 19604 278596
rect 19636 278564 19640 278596
rect 19600 278516 19640 278564
rect 19600 278484 19604 278516
rect 19636 278484 19640 278516
rect 19600 278480 19640 278484
rect 19680 278676 19720 278724
rect 19680 278644 19684 278676
rect 19716 278644 19720 278676
rect 19680 278596 19720 278644
rect 19680 278564 19684 278596
rect 19716 278564 19720 278596
rect 19680 278516 19720 278564
rect 19760 351315 19800 351320
rect 19760 351285 19765 351315
rect 19795 351285 19800 351315
rect 19760 278595 19800 351285
rect 19760 278565 19765 278595
rect 19795 278565 19800 278595
rect 19760 278560 19800 278565
rect 19840 351236 19880 351364
rect 19840 351204 19844 351236
rect 19876 351204 19880 351236
rect 19840 351156 19880 351204
rect 19840 351124 19844 351156
rect 19876 351124 19880 351156
rect 34097 351150 36597 352400
rect 60097 351150 62597 352400
rect 82797 351150 85297 352400
rect 85447 351150 86547 352400
rect 86697 351150 87797 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 111297 351150 112397 352400
rect 112547 351150 113647 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 162147 351150 163247 352400
rect 163397 351150 164497 352400
rect 164647 351150 167147 352400
rect 206697 351150 209197 352400
rect 232697 351150 235197 352400
rect 255297 351170 257697 352400
rect 260297 351170 262697 352400
rect 283297 351150 285797 352400
rect 19840 351076 19880 351124
rect 19840 351044 19844 351076
rect 19876 351044 19880 351076
rect 19840 350996 19880 351044
rect 19840 350964 19844 350996
rect 19876 350964 19880 350996
rect 19840 350916 19880 350964
rect 19840 350884 19844 350916
rect 19876 350884 19880 350916
rect 19840 350836 19880 350884
rect 19840 350804 19844 350836
rect 19876 350804 19880 350836
rect 19840 350756 19880 350804
rect 19840 350724 19844 350756
rect 19876 350724 19880 350756
rect 19840 350676 19880 350724
rect 19840 350644 19844 350676
rect 19876 350644 19880 350676
rect 19840 350596 19880 350644
rect 19840 350564 19844 350596
rect 19876 350564 19880 350596
rect 19840 350516 19880 350564
rect 19840 350484 19844 350516
rect 19876 350484 19880 350516
rect 19840 350436 19880 350484
rect 19840 350404 19844 350436
rect 19876 350404 19880 350436
rect 19840 350356 19880 350404
rect 19840 350324 19844 350356
rect 19876 350324 19880 350356
rect 19840 350276 19880 350324
rect 19840 350244 19844 350276
rect 19876 350244 19880 350276
rect 19840 350196 19880 350244
rect 19840 350164 19844 350196
rect 19876 350164 19880 350196
rect 19840 350116 19880 350164
rect 19840 350084 19844 350116
rect 19876 350084 19880 350116
rect 19840 350036 19880 350084
rect 19840 350004 19844 350036
rect 19876 350004 19880 350036
rect 19840 349956 19880 350004
rect 19840 349924 19844 349956
rect 19876 349924 19880 349956
rect 19840 349876 19880 349924
rect 19840 349844 19844 349876
rect 19876 349844 19880 349876
rect 19840 349796 19880 349844
rect 19840 349764 19844 349796
rect 19876 349764 19880 349796
rect 19840 349716 19880 349764
rect 19840 349684 19844 349716
rect 19876 349684 19880 349716
rect 19840 349636 19880 349684
rect 19840 349604 19844 349636
rect 19876 349604 19880 349636
rect 19840 349556 19880 349604
rect 19840 349524 19844 349556
rect 19876 349524 19880 349556
rect 19840 349476 19880 349524
rect 19840 349444 19844 349476
rect 19876 349444 19880 349476
rect 19840 349396 19880 349444
rect 19840 349364 19844 349396
rect 19876 349364 19880 349396
rect 19840 349316 19880 349364
rect 19840 349284 19844 349316
rect 19876 349284 19880 349316
rect 19840 349236 19880 349284
rect 19840 349204 19844 349236
rect 19876 349204 19880 349236
rect 19840 349156 19880 349204
rect 19840 349124 19844 349156
rect 19876 349124 19880 349156
rect 19840 349076 19880 349124
rect 19840 349044 19844 349076
rect 19876 349044 19880 349076
rect 19840 348996 19880 349044
rect 19840 348964 19844 348996
rect 19876 348964 19880 348996
rect 19840 348916 19880 348964
rect 19840 348884 19844 348916
rect 19876 348884 19880 348916
rect 19840 348836 19880 348884
rect 19840 348804 19844 348836
rect 19876 348804 19880 348836
rect 19840 348756 19880 348804
rect 19840 348724 19844 348756
rect 19876 348724 19880 348756
rect 19840 348676 19880 348724
rect 19840 348644 19844 348676
rect 19876 348644 19880 348676
rect 19840 348596 19880 348644
rect 19840 348564 19844 348596
rect 19876 348564 19880 348596
rect 19840 348516 19880 348564
rect 19840 348484 19844 348516
rect 19876 348484 19880 348516
rect 19840 348436 19880 348484
rect 19840 348404 19844 348436
rect 19876 348404 19880 348436
rect 19840 348356 19880 348404
rect 19840 348324 19844 348356
rect 19876 348324 19880 348356
rect 19840 348276 19880 348324
rect 19840 348244 19844 348276
rect 19876 348244 19880 348276
rect 19840 348196 19880 348244
rect 19840 348164 19844 348196
rect 19876 348164 19880 348196
rect 19840 348116 19880 348164
rect 19840 348084 19844 348116
rect 19876 348084 19880 348116
rect 19840 348036 19880 348084
rect 19840 348004 19844 348036
rect 19876 348004 19880 348036
rect 19840 347956 19880 348004
rect 19840 347924 19844 347956
rect 19876 347924 19880 347956
rect 19840 347876 19880 347924
rect 19840 347844 19844 347876
rect 19876 347844 19880 347876
rect 19840 347796 19880 347844
rect 19840 347764 19844 347796
rect 19876 347764 19880 347796
rect 19840 347716 19880 347764
rect 19840 347684 19844 347716
rect 19876 347684 19880 347716
rect 19840 347636 19880 347684
rect 19840 347604 19844 347636
rect 19876 347604 19880 347636
rect 19840 347556 19880 347604
rect 19840 347524 19844 347556
rect 19876 347524 19880 347556
rect 19840 347476 19880 347524
rect 19840 347444 19844 347476
rect 19876 347444 19880 347476
rect 19840 347396 19880 347444
rect 19840 347364 19844 347396
rect 19876 347364 19880 347396
rect 19840 347316 19880 347364
rect 19840 347284 19844 347316
rect 19876 347284 19880 347316
rect 19840 347236 19880 347284
rect 19840 347204 19844 347236
rect 19876 347204 19880 347236
rect 19840 347156 19880 347204
rect 19840 347124 19844 347156
rect 19876 347124 19880 347156
rect 19840 347076 19880 347124
rect 19840 347044 19844 347076
rect 19876 347044 19880 347076
rect 19840 346996 19880 347044
rect 19840 346964 19844 346996
rect 19876 346964 19880 346996
rect 19840 346916 19880 346964
rect 19840 346884 19844 346916
rect 19876 346884 19880 346916
rect 19840 346836 19880 346884
rect 19840 346804 19844 346836
rect 19876 346804 19880 346836
rect 19840 346756 19880 346804
rect 19840 346724 19844 346756
rect 19876 346724 19880 346756
rect 19840 346676 19880 346724
rect 19840 346644 19844 346676
rect 19876 346644 19880 346676
rect 19840 346596 19880 346644
rect 19840 346564 19844 346596
rect 19876 346564 19880 346596
rect 19840 346516 19880 346564
rect 19840 346484 19844 346516
rect 19876 346484 19880 346516
rect 19840 346436 19880 346484
rect 19840 346404 19844 346436
rect 19876 346404 19880 346436
rect 19840 346356 19880 346404
rect 19840 346324 19844 346356
rect 19876 346324 19880 346356
rect 19840 346276 19880 346324
rect 19840 346244 19844 346276
rect 19876 346244 19880 346276
rect 19840 346196 19880 346244
rect 19840 346164 19844 346196
rect 19876 346164 19880 346196
rect 19840 346116 19880 346164
rect 19840 346084 19844 346116
rect 19876 346084 19880 346116
rect 19840 346036 19880 346084
rect 19840 346004 19844 346036
rect 19876 346004 19880 346036
rect 19840 345956 19880 346004
rect 19840 345924 19844 345956
rect 19876 345924 19880 345956
rect 19840 345876 19880 345924
rect 19840 345844 19844 345876
rect 19876 345844 19880 345876
rect 19840 345796 19880 345844
rect 19840 345764 19844 345796
rect 19876 345764 19880 345796
rect 19840 345716 19880 345764
rect 19840 345684 19844 345716
rect 19876 345684 19880 345716
rect 19840 345636 19880 345684
rect 19840 345604 19844 345636
rect 19876 345604 19880 345636
rect 19840 345556 19880 345604
rect 19840 345524 19844 345556
rect 19876 345524 19880 345556
rect 19840 345476 19880 345524
rect 19840 345444 19844 345476
rect 19876 345444 19880 345476
rect 19840 345396 19880 345444
rect 19840 345364 19844 345396
rect 19876 345364 19880 345396
rect 19840 345316 19880 345364
rect 19840 345284 19844 345316
rect 19876 345284 19880 345316
rect 19840 345236 19880 345284
rect 19840 345204 19844 345236
rect 19876 345204 19880 345236
rect 19840 345156 19880 345204
rect 19840 345124 19844 345156
rect 19876 345124 19880 345156
rect 19840 345076 19880 345124
rect 19840 345044 19844 345076
rect 19876 345044 19880 345076
rect 19840 344996 19880 345044
rect 19840 344964 19844 344996
rect 19876 344964 19880 344996
rect 19840 344916 19880 344964
rect 19840 344884 19844 344916
rect 19876 344884 19880 344916
rect 19840 344836 19880 344884
rect 19840 344804 19844 344836
rect 19876 344804 19880 344836
rect 19840 344756 19880 344804
rect 19840 344724 19844 344756
rect 19876 344724 19880 344756
rect 19840 344676 19880 344724
rect 19840 344644 19844 344676
rect 19876 344644 19880 344676
rect 19840 344596 19880 344644
rect 19840 344564 19844 344596
rect 19876 344564 19880 344596
rect 19840 344516 19880 344564
rect 19840 344484 19844 344516
rect 19876 344484 19880 344516
rect 19840 344436 19880 344484
rect 19840 344404 19844 344436
rect 19876 344404 19880 344436
rect 19840 344356 19880 344404
rect 19840 344324 19844 344356
rect 19876 344324 19880 344356
rect 19840 344276 19880 344324
rect 19840 344244 19844 344276
rect 19876 344244 19880 344276
rect 19840 344196 19880 344244
rect 19840 344164 19844 344196
rect 19876 344164 19880 344196
rect 19840 344116 19880 344164
rect 19840 344084 19844 344116
rect 19876 344084 19880 344116
rect 19840 344036 19880 344084
rect 19840 344004 19844 344036
rect 19876 344004 19880 344036
rect 19840 343956 19880 344004
rect 19840 343924 19844 343956
rect 19876 343924 19880 343956
rect 19840 343876 19880 343924
rect 19840 343844 19844 343876
rect 19876 343844 19880 343876
rect 19840 343796 19880 343844
rect 19840 343764 19844 343796
rect 19876 343764 19880 343796
rect 19840 343716 19880 343764
rect 19840 343684 19844 343716
rect 19876 343684 19880 343716
rect 19840 343636 19880 343684
rect 19840 343604 19844 343636
rect 19876 343604 19880 343636
rect 19840 343556 19880 343604
rect 19840 343524 19844 343556
rect 19876 343524 19880 343556
rect 19840 343476 19880 343524
rect 19840 343444 19844 343476
rect 19876 343444 19880 343476
rect 19840 343396 19880 343444
rect 19840 343364 19844 343396
rect 19876 343364 19880 343396
rect 19840 343316 19880 343364
rect 19840 343284 19844 343316
rect 19876 343284 19880 343316
rect 19840 343236 19880 343284
rect 19840 343204 19844 343236
rect 19876 343204 19880 343236
rect 19840 343156 19880 343204
rect 19840 343124 19844 343156
rect 19876 343124 19880 343156
rect 19840 343076 19880 343124
rect 19840 343044 19844 343076
rect 19876 343044 19880 343076
rect 19840 342996 19880 343044
rect 19840 342964 19844 342996
rect 19876 342964 19880 342996
rect 19840 342916 19880 342964
rect 19840 342884 19844 342916
rect 19876 342884 19880 342916
rect 19840 342836 19880 342884
rect 19840 342804 19844 342836
rect 19876 342804 19880 342836
rect 19840 342756 19880 342804
rect 19840 342724 19844 342756
rect 19876 342724 19880 342756
rect 19840 342676 19880 342724
rect 19840 342644 19844 342676
rect 19876 342644 19880 342676
rect 19840 342596 19880 342644
rect 19840 342564 19844 342596
rect 19876 342564 19880 342596
rect 19840 342516 19880 342564
rect 19840 342484 19844 342516
rect 19876 342484 19880 342516
rect 19840 342436 19880 342484
rect 19840 342404 19844 342436
rect 19876 342404 19880 342436
rect 19840 342356 19880 342404
rect 19840 342324 19844 342356
rect 19876 342324 19880 342356
rect 19840 342276 19880 342324
rect 19840 342244 19844 342276
rect 19876 342244 19880 342276
rect 19840 342196 19880 342244
rect 19840 342164 19844 342196
rect 19876 342164 19880 342196
rect 19840 342116 19880 342164
rect 19840 342084 19844 342116
rect 19876 342084 19880 342116
rect 19840 342036 19880 342084
rect 19840 342004 19844 342036
rect 19876 342004 19880 342036
rect 19840 341956 19880 342004
rect 19840 341924 19844 341956
rect 19876 341924 19880 341956
rect 19840 341876 19880 341924
rect 19840 341844 19844 341876
rect 19876 341844 19880 341876
rect 19840 341796 19880 341844
rect 19840 341764 19844 341796
rect 19876 341764 19880 341796
rect 19840 341716 19880 341764
rect 19840 341684 19844 341716
rect 19876 341684 19880 341716
rect 19840 341636 19880 341684
rect 19840 341604 19844 341636
rect 19876 341604 19880 341636
rect 19840 341556 19880 341604
rect 19840 341524 19844 341556
rect 19876 341524 19880 341556
rect 19840 341476 19880 341524
rect 19840 341444 19844 341476
rect 19876 341444 19880 341476
rect 19840 341396 19880 341444
rect 19840 341364 19844 341396
rect 19876 341364 19880 341396
rect 19840 341316 19880 341364
rect 19840 341284 19844 341316
rect 19876 341284 19880 341316
rect 19840 341236 19880 341284
rect 19840 341204 19844 341236
rect 19876 341204 19880 341236
rect 19840 341156 19880 341204
rect 19840 341124 19844 341156
rect 19876 341124 19880 341156
rect 19840 341076 19880 341124
rect 19840 341044 19844 341076
rect 19876 341044 19880 341076
rect 19840 340996 19880 341044
rect 19840 340964 19844 340996
rect 19876 340964 19880 340996
rect 19840 340916 19880 340964
rect 19840 340884 19844 340916
rect 19876 340884 19880 340916
rect 19840 340836 19880 340884
rect 19840 340804 19844 340836
rect 19876 340804 19880 340836
rect 19840 340756 19880 340804
rect 19840 340724 19844 340756
rect 19876 340724 19880 340756
rect 19840 340676 19880 340724
rect 19840 340644 19844 340676
rect 19876 340644 19880 340676
rect 19840 340596 19880 340644
rect 19840 340564 19844 340596
rect 19876 340564 19880 340596
rect 19840 340516 19880 340564
rect 19840 340484 19844 340516
rect 19876 340484 19880 340516
rect 19840 340436 19880 340484
rect 19840 340404 19844 340436
rect 19876 340404 19880 340436
rect 19840 340356 19880 340404
rect 19840 340324 19844 340356
rect 19876 340324 19880 340356
rect 19840 340276 19880 340324
rect 19840 340244 19844 340276
rect 19876 340244 19880 340276
rect 19840 340196 19880 340244
rect 19840 340164 19844 340196
rect 19876 340164 19880 340196
rect 19840 340116 19880 340164
rect 19840 340084 19844 340116
rect 19876 340084 19880 340116
rect 19840 340036 19880 340084
rect 19840 340004 19844 340036
rect 19876 340004 19880 340036
rect 19840 339956 19880 340004
rect 19840 339924 19844 339956
rect 19876 339924 19880 339956
rect 19840 339876 19880 339924
rect 19840 339844 19844 339876
rect 19876 339844 19880 339876
rect 19840 339796 19880 339844
rect 19840 339764 19844 339796
rect 19876 339764 19880 339796
rect 19840 339716 19880 339764
rect 19840 339684 19844 339716
rect 19876 339684 19880 339716
rect 19840 339636 19880 339684
rect 19840 339604 19844 339636
rect 19876 339604 19880 339636
rect 19840 339556 19880 339604
rect 19840 339524 19844 339556
rect 19876 339524 19880 339556
rect 19840 339476 19880 339524
rect 19840 339444 19844 339476
rect 19876 339444 19880 339476
rect 19840 339396 19880 339444
rect 19840 339364 19844 339396
rect 19876 339364 19880 339396
rect 19840 339316 19880 339364
rect 19840 339284 19844 339316
rect 19876 339284 19880 339316
rect 19840 339236 19880 339284
rect 19840 339204 19844 339236
rect 19876 339204 19880 339236
rect 19840 339156 19880 339204
rect 19840 339124 19844 339156
rect 19876 339124 19880 339156
rect 19840 339076 19880 339124
rect 19840 339044 19844 339076
rect 19876 339044 19880 339076
rect 19840 338996 19880 339044
rect 19840 338964 19844 338996
rect 19876 338964 19880 338996
rect 291150 338992 292400 341492
rect 19840 338916 19880 338964
rect 19840 338884 19844 338916
rect 19876 338884 19880 338916
rect 19840 338836 19880 338884
rect 19840 338804 19844 338836
rect 19876 338804 19880 338836
rect 19840 338756 19880 338804
rect 19840 338724 19844 338756
rect 19876 338724 19880 338756
rect 19840 338676 19880 338724
rect 19840 338644 19844 338676
rect 19876 338644 19880 338676
rect 19840 338596 19880 338644
rect 19840 338564 19844 338596
rect 19876 338564 19880 338596
rect 19840 338516 19880 338564
rect 19840 338484 19844 338516
rect 19876 338484 19880 338516
rect 19840 338436 19880 338484
rect 19840 338404 19844 338436
rect 19876 338404 19880 338436
rect 19840 338356 19880 338404
rect 19840 338324 19844 338356
rect 19876 338324 19880 338356
rect 19840 338276 19880 338324
rect 19840 338244 19844 338276
rect 19876 338244 19880 338276
rect 19840 338196 19880 338244
rect 19840 338164 19844 338196
rect 19876 338164 19880 338196
rect 19840 338116 19880 338164
rect 19840 338084 19844 338116
rect 19876 338084 19880 338116
rect 19840 338036 19880 338084
rect 19840 338004 19844 338036
rect 19876 338004 19880 338036
rect 19840 337956 19880 338004
rect 19840 337924 19844 337956
rect 19876 337924 19880 337956
rect 19840 337876 19880 337924
rect 19840 337844 19844 337876
rect 19876 337844 19880 337876
rect 19840 337796 19880 337844
rect 19840 337764 19844 337796
rect 19876 337764 19880 337796
rect 19840 337716 19880 337764
rect 19840 337684 19844 337716
rect 19876 337684 19880 337716
rect 19840 337636 19880 337684
rect 19840 337604 19844 337636
rect 19876 337604 19880 337636
rect 19840 337556 19880 337604
rect 19840 337524 19844 337556
rect 19876 337524 19880 337556
rect 19840 337476 19880 337524
rect 19840 337444 19844 337476
rect 19876 337444 19880 337476
rect 19840 337396 19880 337444
rect 19840 337364 19844 337396
rect 19876 337364 19880 337396
rect 19840 337316 19880 337364
rect 19840 337284 19844 337316
rect 19876 337284 19880 337316
rect 19840 337236 19880 337284
rect 19840 337204 19844 337236
rect 19876 337204 19880 337236
rect 19840 337156 19880 337204
rect 19840 337124 19844 337156
rect 19876 337124 19880 337156
rect 19840 337076 19880 337124
rect 19840 337044 19844 337076
rect 19876 337044 19880 337076
rect 19840 336996 19880 337044
rect 19840 336964 19844 336996
rect 19876 336964 19880 336996
rect 19840 336916 19880 336964
rect 19840 336884 19844 336916
rect 19876 336884 19880 336916
rect 19840 336836 19880 336884
rect 19840 336804 19844 336836
rect 19876 336804 19880 336836
rect 19840 336756 19880 336804
rect 19840 336724 19844 336756
rect 19876 336724 19880 336756
rect 19840 336676 19880 336724
rect 19840 336644 19844 336676
rect 19876 336644 19880 336676
rect 19840 336596 19880 336644
rect 19840 336564 19844 336596
rect 19876 336564 19880 336596
rect 19840 336516 19880 336564
rect 19840 336484 19844 336516
rect 19876 336484 19880 336516
rect 19840 336436 19880 336484
rect 19840 336404 19844 336436
rect 19876 336404 19880 336436
rect 19840 336356 19880 336404
rect 19840 336324 19844 336356
rect 19876 336324 19880 336356
rect 19840 336276 19880 336324
rect 19840 336244 19844 336276
rect 19876 336244 19880 336276
rect 19840 336196 19880 336244
rect 19840 336164 19844 336196
rect 19876 336164 19880 336196
rect 19840 336116 19880 336164
rect 19840 336084 19844 336116
rect 19876 336084 19880 336116
rect 19840 336036 19880 336084
rect 19840 336004 19844 336036
rect 19876 336004 19880 336036
rect 19840 335956 19880 336004
rect 19840 335924 19844 335956
rect 19876 335924 19880 335956
rect 19840 335876 19880 335924
rect 19840 335844 19844 335876
rect 19876 335844 19880 335876
rect 19840 335796 19880 335844
rect 19840 335764 19844 335796
rect 19876 335764 19880 335796
rect 19840 335716 19880 335764
rect 19840 335684 19844 335716
rect 19876 335684 19880 335716
rect 19840 335636 19880 335684
rect 19840 335604 19844 335636
rect 19876 335604 19880 335636
rect 19840 335556 19880 335604
rect 19840 335524 19844 335556
rect 19876 335524 19880 335556
rect 19840 335476 19880 335524
rect 19840 335444 19844 335476
rect 19876 335444 19880 335476
rect 19840 335396 19880 335444
rect 19840 335364 19844 335396
rect 19876 335364 19880 335396
rect 19840 335316 19880 335364
rect 19840 335284 19844 335316
rect 19876 335284 19880 335316
rect 19840 335236 19880 335284
rect 19840 335204 19844 335236
rect 19876 335204 19880 335236
rect 19840 335156 19880 335204
rect 19840 335124 19844 335156
rect 19876 335124 19880 335156
rect 19840 335076 19880 335124
rect 19840 335044 19844 335076
rect 19876 335044 19880 335076
rect 19840 334996 19880 335044
rect 19840 334964 19844 334996
rect 19876 334964 19880 334996
rect 19840 334916 19880 334964
rect 19840 334884 19844 334916
rect 19876 334884 19880 334916
rect 19840 334836 19880 334884
rect 19840 334804 19844 334836
rect 19876 334804 19880 334836
rect 19840 334756 19880 334804
rect 19840 334724 19844 334756
rect 19876 334724 19880 334756
rect 19840 334676 19880 334724
rect 19840 334644 19844 334676
rect 19876 334644 19880 334676
rect 19840 334596 19880 334644
rect 19840 334564 19844 334596
rect 19876 334564 19880 334596
rect 19840 334516 19880 334564
rect 19840 334484 19844 334516
rect 19876 334484 19880 334516
rect 19840 334436 19880 334484
rect 19840 334404 19844 334436
rect 19876 334404 19880 334436
rect 19840 334356 19880 334404
rect 19840 334324 19844 334356
rect 19876 334324 19880 334356
rect 19840 334276 19880 334324
rect 19840 334244 19844 334276
rect 19876 334244 19880 334276
rect 19840 334196 19880 334244
rect 19840 334164 19844 334196
rect 19876 334164 19880 334196
rect 19840 334116 19880 334164
rect 19840 334084 19844 334116
rect 19876 334084 19880 334116
rect 19840 334036 19880 334084
rect 19840 334004 19844 334036
rect 19876 334004 19880 334036
rect 19840 333956 19880 334004
rect 19840 333924 19844 333956
rect 19876 333924 19880 333956
rect 19840 333876 19880 333924
rect 19840 333844 19844 333876
rect 19876 333844 19880 333876
rect 19840 333796 19880 333844
rect 19840 333764 19844 333796
rect 19876 333764 19880 333796
rect 19840 333716 19880 333764
rect 19840 333684 19844 333716
rect 19876 333684 19880 333716
rect 19840 333636 19880 333684
rect 19840 333604 19844 333636
rect 19876 333604 19880 333636
rect 19840 333556 19880 333604
rect 19840 333524 19844 333556
rect 19876 333524 19880 333556
rect 19840 333476 19880 333524
rect 19840 333444 19844 333476
rect 19876 333444 19880 333476
rect 19840 333396 19880 333444
rect 19840 333364 19844 333396
rect 19876 333364 19880 333396
rect 19840 333316 19880 333364
rect 19840 333284 19844 333316
rect 19876 333284 19880 333316
rect 19840 333236 19880 333284
rect 19840 333204 19844 333236
rect 19876 333204 19880 333236
rect 19840 333156 19880 333204
rect 19840 333124 19844 333156
rect 19876 333124 19880 333156
rect 19840 333076 19880 333124
rect 19840 333044 19844 333076
rect 19876 333044 19880 333076
rect 19840 332996 19880 333044
rect 19840 332964 19844 332996
rect 19876 332964 19880 332996
rect 19840 332916 19880 332964
rect 19840 332884 19844 332916
rect 19876 332884 19880 332916
rect 19840 332836 19880 332884
rect 19840 332804 19844 332836
rect 19876 332804 19880 332836
rect 19840 332756 19880 332804
rect 19840 332724 19844 332756
rect 19876 332724 19880 332756
rect 19840 332676 19880 332724
rect 19840 332644 19844 332676
rect 19876 332644 19880 332676
rect 19840 332596 19880 332644
rect 19840 332564 19844 332596
rect 19876 332564 19880 332596
rect 19840 332516 19880 332564
rect 19840 332484 19844 332516
rect 19876 332484 19880 332516
rect 19840 332436 19880 332484
rect 19840 332404 19844 332436
rect 19876 332404 19880 332436
rect 19840 332356 19880 332404
rect 19840 332324 19844 332356
rect 19876 332324 19880 332356
rect 19840 332276 19880 332324
rect 19840 332244 19844 332276
rect 19876 332244 19880 332276
rect 19840 332196 19880 332244
rect 19840 332164 19844 332196
rect 19876 332164 19880 332196
rect 19840 332116 19880 332164
rect 19840 332084 19844 332116
rect 19876 332084 19880 332116
rect 19840 332036 19880 332084
rect 19840 332004 19844 332036
rect 19876 332004 19880 332036
rect 19840 331956 19880 332004
rect 19840 331924 19844 331956
rect 19876 331924 19880 331956
rect 19840 331876 19880 331924
rect 19840 331844 19844 331876
rect 19876 331844 19880 331876
rect 19840 331796 19880 331844
rect 19840 331764 19844 331796
rect 19876 331764 19880 331796
rect 19840 331716 19880 331764
rect 19840 331684 19844 331716
rect 19876 331684 19880 331716
rect 19840 331636 19880 331684
rect 19840 331604 19844 331636
rect 19876 331604 19880 331636
rect 19840 331556 19880 331604
rect 19840 331524 19844 331556
rect 19876 331524 19880 331556
rect 19840 331476 19880 331524
rect 19840 331444 19844 331476
rect 19876 331444 19880 331476
rect 19840 331396 19880 331444
rect 19840 331364 19844 331396
rect 19876 331364 19880 331396
rect 19840 331316 19880 331364
rect 19840 331284 19844 331316
rect 19876 331284 19880 331316
rect 19840 331236 19880 331284
rect 19840 331204 19844 331236
rect 19876 331204 19880 331236
rect 19840 331156 19880 331204
rect 19840 331124 19844 331156
rect 19876 331124 19880 331156
rect 19840 331076 19880 331124
rect 19840 331044 19844 331076
rect 19876 331044 19880 331076
rect 19840 330996 19880 331044
rect 19840 330964 19844 330996
rect 19876 330964 19880 330996
rect 19840 330916 19880 330964
rect 19840 330884 19844 330916
rect 19876 330884 19880 330916
rect 19840 330836 19880 330884
rect 19840 330804 19844 330836
rect 19876 330804 19880 330836
rect 19840 330756 19880 330804
rect 19840 330724 19844 330756
rect 19876 330724 19880 330756
rect 19840 330676 19880 330724
rect 19840 330644 19844 330676
rect 19876 330644 19880 330676
rect 19840 330596 19880 330644
rect 19840 330564 19844 330596
rect 19876 330564 19880 330596
rect 19840 330516 19880 330564
rect 19840 330484 19844 330516
rect 19876 330484 19880 330516
rect 19840 330436 19880 330484
rect 19840 330404 19844 330436
rect 19876 330404 19880 330436
rect 19840 330356 19880 330404
rect 19840 330324 19844 330356
rect 19876 330324 19880 330356
rect 19840 330276 19880 330324
rect 19840 330244 19844 330276
rect 19876 330244 19880 330276
rect 19840 330196 19880 330244
rect 19840 330164 19844 330196
rect 19876 330164 19880 330196
rect 19840 330116 19880 330164
rect 19840 330084 19844 330116
rect 19876 330084 19880 330116
rect 19840 330036 19880 330084
rect 19840 330004 19844 330036
rect 19876 330004 19880 330036
rect 19840 329956 19880 330004
rect 19840 329924 19844 329956
rect 19876 329924 19880 329956
rect 19840 329876 19880 329924
rect 19840 329844 19844 329876
rect 19876 329844 19880 329876
rect 19840 329796 19880 329844
rect 19840 329764 19844 329796
rect 19876 329764 19880 329796
rect 19840 329716 19880 329764
rect 19840 329684 19844 329716
rect 19876 329684 19880 329716
rect 19840 329636 19880 329684
rect 19840 329604 19844 329636
rect 19876 329604 19880 329636
rect 19840 329556 19880 329604
rect 19840 329524 19844 329556
rect 19876 329524 19880 329556
rect 19840 329476 19880 329524
rect 19840 329444 19844 329476
rect 19876 329444 19880 329476
rect 19840 329396 19880 329444
rect 19840 329364 19844 329396
rect 19876 329364 19880 329396
rect 19840 329316 19880 329364
rect 19840 329284 19844 329316
rect 19876 329284 19880 329316
rect 19840 329236 19880 329284
rect 19840 329204 19844 329236
rect 19876 329204 19880 329236
rect 19840 329156 19880 329204
rect 19840 329124 19844 329156
rect 19876 329124 19880 329156
rect 19840 329076 19880 329124
rect 19840 329044 19844 329076
rect 19876 329044 19880 329076
rect 19840 328996 19880 329044
rect 19840 328964 19844 328996
rect 19876 328964 19880 328996
rect 19840 328916 19880 328964
rect 19840 328884 19844 328916
rect 19876 328884 19880 328916
rect 19840 328836 19880 328884
rect 19840 328804 19844 328836
rect 19876 328804 19880 328836
rect 19840 328756 19880 328804
rect 19840 328724 19844 328756
rect 19876 328724 19880 328756
rect 19840 328676 19880 328724
rect 19840 328644 19844 328676
rect 19876 328644 19880 328676
rect 19840 328596 19880 328644
rect 19840 328564 19844 328596
rect 19876 328564 19880 328596
rect 19840 328516 19880 328564
rect 19840 328484 19844 328516
rect 19876 328484 19880 328516
rect 19840 328436 19880 328484
rect 19840 328404 19844 328436
rect 19876 328404 19880 328436
rect 19840 328356 19880 328404
rect 19840 328324 19844 328356
rect 19876 328324 19880 328356
rect 19840 328276 19880 328324
rect 19840 328244 19844 328276
rect 19876 328244 19880 328276
rect 19840 328196 19880 328244
rect 19840 328164 19844 328196
rect 19876 328164 19880 328196
rect 19840 328116 19880 328164
rect 19840 328084 19844 328116
rect 19876 328084 19880 328116
rect 19840 328036 19880 328084
rect 19840 328004 19844 328036
rect 19876 328004 19880 328036
rect 19840 327956 19880 328004
rect 19840 327924 19844 327956
rect 19876 327924 19880 327956
rect 19840 327876 19880 327924
rect 19840 327844 19844 327876
rect 19876 327844 19880 327876
rect 19840 327796 19880 327844
rect 19840 327764 19844 327796
rect 19876 327764 19880 327796
rect 19840 327716 19880 327764
rect 19840 327684 19844 327716
rect 19876 327684 19880 327716
rect 19840 327636 19880 327684
rect 19840 327604 19844 327636
rect 19876 327604 19880 327636
rect 19840 327556 19880 327604
rect 19840 327524 19844 327556
rect 19876 327524 19880 327556
rect 19840 327476 19880 327524
rect 19840 327444 19844 327476
rect 19876 327444 19880 327476
rect 19840 327396 19880 327444
rect 19840 327364 19844 327396
rect 19876 327364 19880 327396
rect 19840 327316 19880 327364
rect 19840 327284 19844 327316
rect 19876 327284 19880 327316
rect 19840 327236 19880 327284
rect 19840 327204 19844 327236
rect 19876 327204 19880 327236
rect 19840 327156 19880 327204
rect 19840 327124 19844 327156
rect 19876 327124 19880 327156
rect 19840 327076 19880 327124
rect 19840 327044 19844 327076
rect 19876 327044 19880 327076
rect 19840 326996 19880 327044
rect 19840 326964 19844 326996
rect 19876 326964 19880 326996
rect 19840 326916 19880 326964
rect 19840 326884 19844 326916
rect 19876 326884 19880 326916
rect 19840 326836 19880 326884
rect 19840 326804 19844 326836
rect 19876 326804 19880 326836
rect 19840 326756 19880 326804
rect 19840 326724 19844 326756
rect 19876 326724 19880 326756
rect 19840 326676 19880 326724
rect 19840 326644 19844 326676
rect 19876 326644 19880 326676
rect 19840 326596 19880 326644
rect 19840 326564 19844 326596
rect 19876 326564 19880 326596
rect 19840 326516 19880 326564
rect 19840 326484 19844 326516
rect 19876 326484 19880 326516
rect 19840 326436 19880 326484
rect 19840 326404 19844 326436
rect 19876 326404 19880 326436
rect 19840 326356 19880 326404
rect 19840 326324 19844 326356
rect 19876 326324 19880 326356
rect 19840 326276 19880 326324
rect 19840 326244 19844 326276
rect 19876 326244 19880 326276
rect 19840 326196 19880 326244
rect 19840 326164 19844 326196
rect 19876 326164 19880 326196
rect 19840 326116 19880 326164
rect 19840 326084 19844 326116
rect 19876 326084 19880 326116
rect 19840 326036 19880 326084
rect 19840 326004 19844 326036
rect 19876 326004 19880 326036
rect 19840 325956 19880 326004
rect 19840 325924 19844 325956
rect 19876 325924 19880 325956
rect 19840 325876 19880 325924
rect 19840 325844 19844 325876
rect 19876 325844 19880 325876
rect 19840 325796 19880 325844
rect 19840 325764 19844 325796
rect 19876 325764 19880 325796
rect 19840 325716 19880 325764
rect 19840 325684 19844 325716
rect 19876 325684 19880 325716
rect 19840 325636 19880 325684
rect 19840 325604 19844 325636
rect 19876 325604 19880 325636
rect 19840 325556 19880 325604
rect 19840 325524 19844 325556
rect 19876 325524 19880 325556
rect 19840 325476 19880 325524
rect 19840 325444 19844 325476
rect 19876 325444 19880 325476
rect 19840 325396 19880 325444
rect 19840 325364 19844 325396
rect 19876 325364 19880 325396
rect 19840 325316 19880 325364
rect 19840 325284 19844 325316
rect 19876 325284 19880 325316
rect 19840 325236 19880 325284
rect 19840 325204 19844 325236
rect 19876 325204 19880 325236
rect 19840 325156 19880 325204
rect 19840 325124 19844 325156
rect 19876 325124 19880 325156
rect 19840 325076 19880 325124
rect 19840 325044 19844 325076
rect 19876 325044 19880 325076
rect 19840 324996 19880 325044
rect 19840 324964 19844 324996
rect 19876 324964 19880 324996
rect 19840 324916 19880 324964
rect 19840 324884 19844 324916
rect 19876 324884 19880 324916
rect 19840 324836 19880 324884
rect 19840 324804 19844 324836
rect 19876 324804 19880 324836
rect 19840 324756 19880 324804
rect 19840 324724 19844 324756
rect 19876 324724 19880 324756
rect 19840 324676 19880 324724
rect 19840 324644 19844 324676
rect 19876 324644 19880 324676
rect 19840 324596 19880 324644
rect 19840 324564 19844 324596
rect 19876 324564 19880 324596
rect 19840 324516 19880 324564
rect 19840 324484 19844 324516
rect 19876 324484 19880 324516
rect 19840 324436 19880 324484
rect 19840 324404 19844 324436
rect 19876 324404 19880 324436
rect 19840 324356 19880 324404
rect 19840 324324 19844 324356
rect 19876 324324 19880 324356
rect 19840 324276 19880 324324
rect 19840 324244 19844 324276
rect 19876 324244 19880 324276
rect 19840 324196 19880 324244
rect 19840 324164 19844 324196
rect 19876 324164 19880 324196
rect 19840 324116 19880 324164
rect 19840 324084 19844 324116
rect 19876 324084 19880 324116
rect 19840 324036 19880 324084
rect 19840 324004 19844 324036
rect 19876 324004 19880 324036
rect 19840 323956 19880 324004
rect 19840 323924 19844 323956
rect 19876 323924 19880 323956
rect 19840 323876 19880 323924
rect 19840 323844 19844 323876
rect 19876 323844 19880 323876
rect 19840 323796 19880 323844
rect 19840 323764 19844 323796
rect 19876 323764 19880 323796
rect 19840 323716 19880 323764
rect 19840 323684 19844 323716
rect 19876 323684 19880 323716
rect 19840 323636 19880 323684
rect 19840 323604 19844 323636
rect 19876 323604 19880 323636
rect 19840 323556 19880 323604
rect 19840 323524 19844 323556
rect 19876 323524 19880 323556
rect 19840 323476 19880 323524
rect 19840 323444 19844 323476
rect 19876 323444 19880 323476
rect 19840 323396 19880 323444
rect 19840 323364 19844 323396
rect 19876 323364 19880 323396
rect 19840 323316 19880 323364
rect 19840 323284 19844 323316
rect 19876 323284 19880 323316
rect 19840 323236 19880 323284
rect 19840 323204 19844 323236
rect 19876 323204 19880 323236
rect 19840 323156 19880 323204
rect 19840 323124 19844 323156
rect 19876 323124 19880 323156
rect 19840 323076 19880 323124
rect 19840 323044 19844 323076
rect 19876 323044 19880 323076
rect 19840 322996 19880 323044
rect 19840 322964 19844 322996
rect 19876 322964 19880 322996
rect 19840 322916 19880 322964
rect 19840 322884 19844 322916
rect 19876 322884 19880 322916
rect 19840 322836 19880 322884
rect 19840 322804 19844 322836
rect 19876 322804 19880 322836
rect 19840 322756 19880 322804
rect 19840 322724 19844 322756
rect 19876 322724 19880 322756
rect 19840 322676 19880 322724
rect 19840 322644 19844 322676
rect 19876 322644 19880 322676
rect 19840 322596 19880 322644
rect 19840 322564 19844 322596
rect 19876 322564 19880 322596
rect 19840 322516 19880 322564
rect 19840 322484 19844 322516
rect 19876 322484 19880 322516
rect 19840 322436 19880 322484
rect 19840 322404 19844 322436
rect 19876 322404 19880 322436
rect 19840 322356 19880 322404
rect 19840 322324 19844 322356
rect 19876 322324 19880 322356
rect 19840 322276 19880 322324
rect 19840 322244 19844 322276
rect 19876 322244 19880 322276
rect 19840 322196 19880 322244
rect 19840 322164 19844 322196
rect 19876 322164 19880 322196
rect 19840 322116 19880 322164
rect 19840 322084 19844 322116
rect 19876 322084 19880 322116
rect 19840 322036 19880 322084
rect 19840 322004 19844 322036
rect 19876 322004 19880 322036
rect 19840 321956 19880 322004
rect 19840 321924 19844 321956
rect 19876 321924 19880 321956
rect 19840 321876 19880 321924
rect 19840 321844 19844 321876
rect 19876 321844 19880 321876
rect 19840 321796 19880 321844
rect 19840 321764 19844 321796
rect 19876 321764 19880 321796
rect 19840 321716 19880 321764
rect 19840 321684 19844 321716
rect 19876 321684 19880 321716
rect 19840 321636 19880 321684
rect 19840 321604 19844 321636
rect 19876 321604 19880 321636
rect 19840 321556 19880 321604
rect 19840 321524 19844 321556
rect 19876 321524 19880 321556
rect 19840 321476 19880 321524
rect 19840 321444 19844 321476
rect 19876 321444 19880 321476
rect 19840 321396 19880 321444
rect 19840 321364 19844 321396
rect 19876 321364 19880 321396
rect 19840 321316 19880 321364
rect 19840 321284 19844 321316
rect 19876 321284 19880 321316
rect 19840 321236 19880 321284
rect 19840 321204 19844 321236
rect 19876 321204 19880 321236
rect 19840 321156 19880 321204
rect 19840 321124 19844 321156
rect 19876 321124 19880 321156
rect 19840 321076 19880 321124
rect 19840 321044 19844 321076
rect 19876 321044 19880 321076
rect 19840 320996 19880 321044
rect 19840 320964 19844 320996
rect 19876 320964 19880 320996
rect 19840 320916 19880 320964
rect 19840 320884 19844 320916
rect 19876 320884 19880 320916
rect 19840 320836 19880 320884
rect 19840 320804 19844 320836
rect 19876 320804 19880 320836
rect 19840 320756 19880 320804
rect 19840 320724 19844 320756
rect 19876 320724 19880 320756
rect 19840 320676 19880 320724
rect 19840 320644 19844 320676
rect 19876 320644 19880 320676
rect 19840 320596 19880 320644
rect 19840 320564 19844 320596
rect 19876 320564 19880 320596
rect 19840 320516 19880 320564
rect 19840 320484 19844 320516
rect 19876 320484 19880 320516
rect 19840 320436 19880 320484
rect 19840 320404 19844 320436
rect 19876 320404 19880 320436
rect 19840 320356 19880 320404
rect 19840 320324 19844 320356
rect 19876 320324 19880 320356
rect 19840 320276 19880 320324
rect 19840 320244 19844 320276
rect 19876 320244 19880 320276
rect 19840 320196 19880 320244
rect 19840 320164 19844 320196
rect 19876 320164 19880 320196
rect 19840 320116 19880 320164
rect 19840 320084 19844 320116
rect 19876 320084 19880 320116
rect 19840 320036 19880 320084
rect 19840 320004 19844 320036
rect 19876 320004 19880 320036
rect 19840 319956 19880 320004
rect 19840 319924 19844 319956
rect 19876 319924 19880 319956
rect 19840 319876 19880 319924
rect 291170 319892 292400 322292
rect 19840 319844 19844 319876
rect 19876 319844 19880 319876
rect 19840 319796 19880 319844
rect 19840 319764 19844 319796
rect 19876 319764 19880 319796
rect 19840 319716 19880 319764
rect 19840 319684 19844 319716
rect 19876 319684 19880 319716
rect 19840 319636 19880 319684
rect 19840 319604 19844 319636
rect 19876 319604 19880 319636
rect 19840 319556 19880 319604
rect 19840 319524 19844 319556
rect 19876 319524 19880 319556
rect 19840 319476 19880 319524
rect 19840 319444 19844 319476
rect 19876 319444 19880 319476
rect 19840 319396 19880 319444
rect 19840 319364 19844 319396
rect 19876 319364 19880 319396
rect 19840 319316 19880 319364
rect 19840 319284 19844 319316
rect 19876 319284 19880 319316
rect 19840 319236 19880 319284
rect 19840 319204 19844 319236
rect 19876 319204 19880 319236
rect 19840 319156 19880 319204
rect 19840 319124 19844 319156
rect 19876 319124 19880 319156
rect 19840 319076 19880 319124
rect 19840 319044 19844 319076
rect 19876 319044 19880 319076
rect 19840 318996 19880 319044
rect 19840 318964 19844 318996
rect 19876 318964 19880 318996
rect 19840 318916 19880 318964
rect 19840 318884 19844 318916
rect 19876 318884 19880 318916
rect 19840 318836 19880 318884
rect 19840 318804 19844 318836
rect 19876 318804 19880 318836
rect 19840 318756 19880 318804
rect 19840 318724 19844 318756
rect 19876 318724 19880 318756
rect 19840 318676 19880 318724
rect 19840 318644 19844 318676
rect 19876 318644 19880 318676
rect 19840 318596 19880 318644
rect 19840 318564 19844 318596
rect 19876 318564 19880 318596
rect 19840 318516 19880 318564
rect 19840 318484 19844 318516
rect 19876 318484 19880 318516
rect 19840 318436 19880 318484
rect 19840 318404 19844 318436
rect 19876 318404 19880 318436
rect 19840 318356 19880 318404
rect 19840 318324 19844 318356
rect 19876 318324 19880 318356
rect 19840 318276 19880 318324
rect 19840 318244 19844 318276
rect 19876 318244 19880 318276
rect 19840 318196 19880 318244
rect 19840 318164 19844 318196
rect 19876 318164 19880 318196
rect 19840 318116 19880 318164
rect 19840 318084 19844 318116
rect 19876 318084 19880 318116
rect 19840 318036 19880 318084
rect 19840 318004 19844 318036
rect 19876 318004 19880 318036
rect 19840 317956 19880 318004
rect 19840 317924 19844 317956
rect 19876 317924 19880 317956
rect 19840 317876 19880 317924
rect 19840 317844 19844 317876
rect 19876 317844 19880 317876
rect 19840 317796 19880 317844
rect 19840 317764 19844 317796
rect 19876 317764 19880 317796
rect 19840 317716 19880 317764
rect 19840 317684 19844 317716
rect 19876 317684 19880 317716
rect 19840 317636 19880 317684
rect 19840 317604 19844 317636
rect 19876 317604 19880 317636
rect 19840 317556 19880 317604
rect 19840 317524 19844 317556
rect 19876 317524 19880 317556
rect 19840 317476 19880 317524
rect 19840 317444 19844 317476
rect 19876 317444 19880 317476
rect 19840 317396 19880 317444
rect 19840 317364 19844 317396
rect 19876 317364 19880 317396
rect 19840 317316 19880 317364
rect 19840 317284 19844 317316
rect 19876 317284 19880 317316
rect 19840 317236 19880 317284
rect 19840 317204 19844 317236
rect 19876 317204 19880 317236
rect 19840 317156 19880 317204
rect 19840 317124 19844 317156
rect 19876 317124 19880 317156
rect 19840 317076 19880 317124
rect 19840 317044 19844 317076
rect 19876 317044 19880 317076
rect 19840 316996 19880 317044
rect 19840 316964 19844 316996
rect 19876 316964 19880 316996
rect 19840 316916 19880 316964
rect 19840 316884 19844 316916
rect 19876 316884 19880 316916
rect 19840 316836 19880 316884
rect 19840 316804 19844 316836
rect 19876 316804 19880 316836
rect 19840 316756 19880 316804
rect 19840 316724 19844 316756
rect 19876 316724 19880 316756
rect 19840 316676 19880 316724
rect 19840 316644 19844 316676
rect 19876 316644 19880 316676
rect 19840 316596 19880 316644
rect 19840 316564 19844 316596
rect 19876 316564 19880 316596
rect 19840 316516 19880 316564
rect 19840 316484 19844 316516
rect 19876 316484 19880 316516
rect 19840 316436 19880 316484
rect 19840 316404 19844 316436
rect 19876 316404 19880 316436
rect 19840 316356 19880 316404
rect 19840 316324 19844 316356
rect 19876 316324 19880 316356
rect 19840 316276 19880 316324
rect 19840 316244 19844 316276
rect 19876 316244 19880 316276
rect 19840 316196 19880 316244
rect 19840 316164 19844 316196
rect 19876 316164 19880 316196
rect 19840 316116 19880 316164
rect 19840 316084 19844 316116
rect 19876 316084 19880 316116
rect 19840 316036 19880 316084
rect 19840 316004 19844 316036
rect 19876 316004 19880 316036
rect 19840 315956 19880 316004
rect 19840 315924 19844 315956
rect 19876 315924 19880 315956
rect 19840 315876 19880 315924
rect 19840 315844 19844 315876
rect 19876 315844 19880 315876
rect 19840 315796 19880 315844
rect 19840 315764 19844 315796
rect 19876 315764 19880 315796
rect 19840 315716 19880 315764
rect 19840 315684 19844 315716
rect 19876 315684 19880 315716
rect 19840 315636 19880 315684
rect 19840 315604 19844 315636
rect 19876 315604 19880 315636
rect 19840 315556 19880 315604
rect 19840 315524 19844 315556
rect 19876 315524 19880 315556
rect 19840 315476 19880 315524
rect 19840 315444 19844 315476
rect 19876 315444 19880 315476
rect 19840 315396 19880 315444
rect 19840 315364 19844 315396
rect 19876 315364 19880 315396
rect 19840 315316 19880 315364
rect 19840 315284 19844 315316
rect 19876 315284 19880 315316
rect 19840 315236 19880 315284
rect 19840 315204 19844 315236
rect 19876 315204 19880 315236
rect 19840 315156 19880 315204
rect 19840 315124 19844 315156
rect 19876 315124 19880 315156
rect 19840 315076 19880 315124
rect 19840 315044 19844 315076
rect 19876 315044 19880 315076
rect 19840 314996 19880 315044
rect 19840 314964 19844 314996
rect 19876 314964 19880 314996
rect 19840 314916 19880 314964
rect 19840 314884 19844 314916
rect 19876 314884 19880 314916
rect 291170 314892 292400 317292
rect 19840 314836 19880 314884
rect 19840 314804 19844 314836
rect 19876 314804 19880 314836
rect 19840 314756 19880 314804
rect 19840 314724 19844 314756
rect 19876 314724 19880 314756
rect 19840 314676 19880 314724
rect 19840 314644 19844 314676
rect 19876 314644 19880 314676
rect 19840 314596 19880 314644
rect 19840 314564 19844 314596
rect 19876 314564 19880 314596
rect 19840 314516 19880 314564
rect 19840 314484 19844 314516
rect 19876 314484 19880 314516
rect 19840 314436 19880 314484
rect 19840 314404 19844 314436
rect 19876 314404 19880 314436
rect 19840 314356 19880 314404
rect 19840 314324 19844 314356
rect 19876 314324 19880 314356
rect 19840 314276 19880 314324
rect 19840 314244 19844 314276
rect 19876 314244 19880 314276
rect 19840 314196 19880 314244
rect 19840 314164 19844 314196
rect 19876 314164 19880 314196
rect 19840 314116 19880 314164
rect 19840 314084 19844 314116
rect 19876 314084 19880 314116
rect 19840 314036 19880 314084
rect 19840 314004 19844 314036
rect 19876 314004 19880 314036
rect 19840 313956 19880 314004
rect 19840 313924 19844 313956
rect 19876 313924 19880 313956
rect 19840 313876 19880 313924
rect 19840 313844 19844 313876
rect 19876 313844 19880 313876
rect 19840 313796 19880 313844
rect 19840 313764 19844 313796
rect 19876 313764 19880 313796
rect 19840 313716 19880 313764
rect 19840 313684 19844 313716
rect 19876 313684 19880 313716
rect 19840 313636 19880 313684
rect 19840 313604 19844 313636
rect 19876 313604 19880 313636
rect 19840 313556 19880 313604
rect 19840 313524 19844 313556
rect 19876 313524 19880 313556
rect 19840 313476 19880 313524
rect 19840 313444 19844 313476
rect 19876 313444 19880 313476
rect 19840 313396 19880 313444
rect 19840 313364 19844 313396
rect 19876 313364 19880 313396
rect 19840 313316 19880 313364
rect 19840 313284 19844 313316
rect 19876 313284 19880 313316
rect 19840 313236 19880 313284
rect 19840 313204 19844 313236
rect 19876 313204 19880 313236
rect 19840 313156 19880 313204
rect 19840 313124 19844 313156
rect 19876 313124 19880 313156
rect 19840 313076 19880 313124
rect 19840 313044 19844 313076
rect 19876 313044 19880 313076
rect 19840 312996 19880 313044
rect 19840 312964 19844 312996
rect 19876 312964 19880 312996
rect 19840 312916 19880 312964
rect 19840 312884 19844 312916
rect 19876 312884 19880 312916
rect 19840 312836 19880 312884
rect 19840 312804 19844 312836
rect 19876 312804 19880 312836
rect 19840 312756 19880 312804
rect 19840 312724 19844 312756
rect 19876 312724 19880 312756
rect 19840 312676 19880 312724
rect 19840 312644 19844 312676
rect 19876 312644 19880 312676
rect 19840 312596 19880 312644
rect 19840 312564 19844 312596
rect 19876 312564 19880 312596
rect 19840 312516 19880 312564
rect 19840 312484 19844 312516
rect 19876 312484 19880 312516
rect 19840 312436 19880 312484
rect 19840 312404 19844 312436
rect 19876 312404 19880 312436
rect 19840 312356 19880 312404
rect 19840 312324 19844 312356
rect 19876 312324 19880 312356
rect 19840 312276 19880 312324
rect 19840 312244 19844 312276
rect 19876 312244 19880 312276
rect 19840 312196 19880 312244
rect 19840 312164 19844 312196
rect 19876 312164 19880 312196
rect 19840 312116 19880 312164
rect 19840 312084 19844 312116
rect 19876 312084 19880 312116
rect 19840 312036 19880 312084
rect 19840 312004 19844 312036
rect 19876 312004 19880 312036
rect 19840 311956 19880 312004
rect 19840 311924 19844 311956
rect 19876 311924 19880 311956
rect 19840 311876 19880 311924
rect 19840 311844 19844 311876
rect 19876 311844 19880 311876
rect 19840 311796 19880 311844
rect 19840 311764 19844 311796
rect 19876 311764 19880 311796
rect 19840 311716 19880 311764
rect 19840 311684 19844 311716
rect 19876 311684 19880 311716
rect 19840 311636 19880 311684
rect 19840 311604 19844 311636
rect 19876 311604 19880 311636
rect 19840 311556 19880 311604
rect 19840 311524 19844 311556
rect 19876 311524 19880 311556
rect 19840 311476 19880 311524
rect 19840 311444 19844 311476
rect 19876 311444 19880 311476
rect 19840 311396 19880 311444
rect 19840 311364 19844 311396
rect 19876 311364 19880 311396
rect 19840 311316 19880 311364
rect 19840 311284 19844 311316
rect 19876 311284 19880 311316
rect 19840 311236 19880 311284
rect 19840 311204 19844 311236
rect 19876 311204 19880 311236
rect 19840 311156 19880 311204
rect 19840 311124 19844 311156
rect 19876 311124 19880 311156
rect 19840 311076 19880 311124
rect 19840 311044 19844 311076
rect 19876 311044 19880 311076
rect 19840 310996 19880 311044
rect 19840 310964 19844 310996
rect 19876 310964 19880 310996
rect 19840 310916 19880 310964
rect 19840 310884 19844 310916
rect 19876 310884 19880 310916
rect 19840 310836 19880 310884
rect 19840 310804 19844 310836
rect 19876 310804 19880 310836
rect 19840 310756 19880 310804
rect 19840 310724 19844 310756
rect 19876 310724 19880 310756
rect 19840 310676 19880 310724
rect 19840 310644 19844 310676
rect 19876 310644 19880 310676
rect 19840 310596 19880 310644
rect 19840 310564 19844 310596
rect 19876 310564 19880 310596
rect 19840 310516 19880 310564
rect 19840 310484 19844 310516
rect 19876 310484 19880 310516
rect 19840 310436 19880 310484
rect 19840 310404 19844 310436
rect 19876 310404 19880 310436
rect 19840 310356 19880 310404
rect 19840 310324 19844 310356
rect 19876 310324 19880 310356
rect 19840 310276 19880 310324
rect 19840 310244 19844 310276
rect 19876 310244 19880 310276
rect 19840 310196 19880 310244
rect 19840 310164 19844 310196
rect 19876 310164 19880 310196
rect 19840 310116 19880 310164
rect 19840 310084 19844 310116
rect 19876 310084 19880 310116
rect 19840 310036 19880 310084
rect 19840 310004 19844 310036
rect 19876 310004 19880 310036
rect 19840 309956 19880 310004
rect 19840 309924 19844 309956
rect 19876 309924 19880 309956
rect 19840 309876 19880 309924
rect 19840 309844 19844 309876
rect 19876 309844 19880 309876
rect 19840 309796 19880 309844
rect 19840 309764 19844 309796
rect 19876 309764 19880 309796
rect 19840 309716 19880 309764
rect 19840 309684 19844 309716
rect 19876 309684 19880 309716
rect 19840 309636 19880 309684
rect 19840 309604 19844 309636
rect 19876 309604 19880 309636
rect 19840 309556 19880 309604
rect 19840 309524 19844 309556
rect 19876 309524 19880 309556
rect 19840 309476 19880 309524
rect 19840 309444 19844 309476
rect 19876 309444 19880 309476
rect 19840 309396 19880 309444
rect 19840 309364 19844 309396
rect 19876 309364 19880 309396
rect 19840 309316 19880 309364
rect 19840 309284 19844 309316
rect 19876 309284 19880 309316
rect 19840 309236 19880 309284
rect 19840 309204 19844 309236
rect 19876 309204 19880 309236
rect 19840 309156 19880 309204
rect 19840 309124 19844 309156
rect 19876 309124 19880 309156
rect 19840 309076 19880 309124
rect 19840 309044 19844 309076
rect 19876 309044 19880 309076
rect 19840 308996 19880 309044
rect 19840 308964 19844 308996
rect 19876 308964 19880 308996
rect 19840 308916 19880 308964
rect 19840 308884 19844 308916
rect 19876 308884 19880 308916
rect 19840 308836 19880 308884
rect 19840 308804 19844 308836
rect 19876 308804 19880 308836
rect 19840 308756 19880 308804
rect 19840 308724 19844 308756
rect 19876 308724 19880 308756
rect 19840 308676 19880 308724
rect 19840 308644 19844 308676
rect 19876 308644 19880 308676
rect 19840 308596 19880 308644
rect 19840 308564 19844 308596
rect 19876 308564 19880 308596
rect 19840 308516 19880 308564
rect 19840 308484 19844 308516
rect 19876 308484 19880 308516
rect 19840 308436 19880 308484
rect 19840 308404 19844 308436
rect 19876 308404 19880 308436
rect 19840 308356 19880 308404
rect 19840 308324 19844 308356
rect 19876 308324 19880 308356
rect 19840 308276 19880 308324
rect 19840 308244 19844 308276
rect 19876 308244 19880 308276
rect 19840 308196 19880 308244
rect 19840 308164 19844 308196
rect 19876 308164 19880 308196
rect 19840 308116 19880 308164
rect 19840 308084 19844 308116
rect 19876 308084 19880 308116
rect 19840 308036 19880 308084
rect 19840 308004 19844 308036
rect 19876 308004 19880 308036
rect 19840 307956 19880 308004
rect 19840 307924 19844 307956
rect 19876 307924 19880 307956
rect 19840 307876 19880 307924
rect 19840 307844 19844 307876
rect 19876 307844 19880 307876
rect 19840 307796 19880 307844
rect 19840 307764 19844 307796
rect 19876 307764 19880 307796
rect 19840 307716 19880 307764
rect 19840 307684 19844 307716
rect 19876 307684 19880 307716
rect 19840 307636 19880 307684
rect 19840 307604 19844 307636
rect 19876 307604 19880 307636
rect 19840 307556 19880 307604
rect 19840 307524 19844 307556
rect 19876 307524 19880 307556
rect 19840 307476 19880 307524
rect 19840 307444 19844 307476
rect 19876 307444 19880 307476
rect 19840 307396 19880 307444
rect 19840 307364 19844 307396
rect 19876 307364 19880 307396
rect 19840 307316 19880 307364
rect 19840 307284 19844 307316
rect 19876 307284 19880 307316
rect 19840 307236 19880 307284
rect 19840 307204 19844 307236
rect 19876 307204 19880 307236
rect 19840 307156 19880 307204
rect 19840 307124 19844 307156
rect 19876 307124 19880 307156
rect 19840 307076 19880 307124
rect 19840 307044 19844 307076
rect 19876 307044 19880 307076
rect 19840 306996 19880 307044
rect 19840 306964 19844 306996
rect 19876 306964 19880 306996
rect 19840 306916 19880 306964
rect 19840 306884 19844 306916
rect 19876 306884 19880 306916
rect 19840 306836 19880 306884
rect 19840 306804 19844 306836
rect 19876 306804 19880 306836
rect 19840 306756 19880 306804
rect 19840 306724 19844 306756
rect 19876 306724 19880 306756
rect 19840 306676 19880 306724
rect 19840 306644 19844 306676
rect 19876 306644 19880 306676
rect 19840 306596 19880 306644
rect 19840 306564 19844 306596
rect 19876 306564 19880 306596
rect 19840 306516 19880 306564
rect 19840 306484 19844 306516
rect 19876 306484 19880 306516
rect 19840 306436 19880 306484
rect 19840 306404 19844 306436
rect 19876 306404 19880 306436
rect 19840 306356 19880 306404
rect 19840 306324 19844 306356
rect 19876 306324 19880 306356
rect 19840 306276 19880 306324
rect 19840 306244 19844 306276
rect 19876 306244 19880 306276
rect 19840 306196 19880 306244
rect 19840 306164 19844 306196
rect 19876 306164 19880 306196
rect 19840 306116 19880 306164
rect 19840 306084 19844 306116
rect 19876 306084 19880 306116
rect 19840 306036 19880 306084
rect 19840 306004 19844 306036
rect 19876 306004 19880 306036
rect 19840 305956 19880 306004
rect 19840 305924 19844 305956
rect 19876 305924 19880 305956
rect 19840 305876 19880 305924
rect 19840 305844 19844 305876
rect 19876 305844 19880 305876
rect 19840 305796 19880 305844
rect 19840 305764 19844 305796
rect 19876 305764 19880 305796
rect 19840 305716 19880 305764
rect 19840 305684 19844 305716
rect 19876 305684 19880 305716
rect 19840 305636 19880 305684
rect 19840 305604 19844 305636
rect 19876 305604 19880 305636
rect 19840 305556 19880 305604
rect 19840 305524 19844 305556
rect 19876 305524 19880 305556
rect 19840 305476 19880 305524
rect 19840 305444 19844 305476
rect 19876 305444 19880 305476
rect 19840 305396 19880 305444
rect 19840 305364 19844 305396
rect 19876 305364 19880 305396
rect 19840 305316 19880 305364
rect 19840 305284 19844 305316
rect 19876 305284 19880 305316
rect 19840 305236 19880 305284
rect 19840 305204 19844 305236
rect 19876 305204 19880 305236
rect 19840 305156 19880 305204
rect 19840 305124 19844 305156
rect 19876 305124 19880 305156
rect 19840 305076 19880 305124
rect 19840 305044 19844 305076
rect 19876 305044 19880 305076
rect 19840 304996 19880 305044
rect 19840 304964 19844 304996
rect 19876 304964 19880 304996
rect 19840 304916 19880 304964
rect 19840 304884 19844 304916
rect 19876 304884 19880 304916
rect 19840 304836 19880 304884
rect 19840 304804 19844 304836
rect 19876 304804 19880 304836
rect 19840 304756 19880 304804
rect 19840 304724 19844 304756
rect 19876 304724 19880 304756
rect 19840 304676 19880 304724
rect 19840 304644 19844 304676
rect 19876 304644 19880 304676
rect 19840 304596 19880 304644
rect 19840 304564 19844 304596
rect 19876 304564 19880 304596
rect 19840 304516 19880 304564
rect 19840 304484 19844 304516
rect 19876 304484 19880 304516
rect 19840 304436 19880 304484
rect 19840 304404 19844 304436
rect 19876 304404 19880 304436
rect 19840 304356 19880 304404
rect 19840 304324 19844 304356
rect 19876 304324 19880 304356
rect 19840 304276 19880 304324
rect 19840 304244 19844 304276
rect 19876 304244 19880 304276
rect 19840 304196 19880 304244
rect 19840 304164 19844 304196
rect 19876 304164 19880 304196
rect 19840 304116 19880 304164
rect 19840 304084 19844 304116
rect 19876 304084 19880 304116
rect 19840 304036 19880 304084
rect 19840 304004 19844 304036
rect 19876 304004 19880 304036
rect 19840 303956 19880 304004
rect 19840 303924 19844 303956
rect 19876 303924 19880 303956
rect 19840 303876 19880 303924
rect 19840 303844 19844 303876
rect 19876 303844 19880 303876
rect 19840 303796 19880 303844
rect 19840 303764 19844 303796
rect 19876 303764 19880 303796
rect 19840 303716 19880 303764
rect 19840 303684 19844 303716
rect 19876 303684 19880 303716
rect 19840 303636 19880 303684
rect 19840 303604 19844 303636
rect 19876 303604 19880 303636
rect 19840 303556 19880 303604
rect 19840 303524 19844 303556
rect 19876 303524 19880 303556
rect 19840 303476 19880 303524
rect 19840 303444 19844 303476
rect 19876 303444 19880 303476
rect 19840 303396 19880 303444
rect 19840 303364 19844 303396
rect 19876 303364 19880 303396
rect 19840 303316 19880 303364
rect 19840 303284 19844 303316
rect 19876 303284 19880 303316
rect 19840 303236 19880 303284
rect 19840 303204 19844 303236
rect 19876 303204 19880 303236
rect 19840 303156 19880 303204
rect 19840 303124 19844 303156
rect 19876 303124 19880 303156
rect 19840 303076 19880 303124
rect 19840 303044 19844 303076
rect 19876 303044 19880 303076
rect 19840 302996 19880 303044
rect 19840 302964 19844 302996
rect 19876 302964 19880 302996
rect 19840 302916 19880 302964
rect 19840 302884 19844 302916
rect 19876 302884 19880 302916
rect 19840 302836 19880 302884
rect 19840 302804 19844 302836
rect 19876 302804 19880 302836
rect 19840 302756 19880 302804
rect 19840 302724 19844 302756
rect 19876 302724 19880 302756
rect 19840 302676 19880 302724
rect 19840 302644 19844 302676
rect 19876 302644 19880 302676
rect 19840 302596 19880 302644
rect 19840 302564 19844 302596
rect 19876 302564 19880 302596
rect 19840 302516 19880 302564
rect 19840 302484 19844 302516
rect 19876 302484 19880 302516
rect 19840 302436 19880 302484
rect 19840 302404 19844 302436
rect 19876 302404 19880 302436
rect 19840 302356 19880 302404
rect 19840 302324 19844 302356
rect 19876 302324 19880 302356
rect 19840 302276 19880 302324
rect 19840 302244 19844 302276
rect 19876 302244 19880 302276
rect 19840 302196 19880 302244
rect 19840 302164 19844 302196
rect 19876 302164 19880 302196
rect 19840 302116 19880 302164
rect 19840 302084 19844 302116
rect 19876 302084 19880 302116
rect 19840 302036 19880 302084
rect 19840 302004 19844 302036
rect 19876 302004 19880 302036
rect 19840 301956 19880 302004
rect 19840 301924 19844 301956
rect 19876 301924 19880 301956
rect 19840 301876 19880 301924
rect 19840 301844 19844 301876
rect 19876 301844 19880 301876
rect 19840 301796 19880 301844
rect 19840 301764 19844 301796
rect 19876 301764 19880 301796
rect 19840 301716 19880 301764
rect 19840 301684 19844 301716
rect 19876 301684 19880 301716
rect 19840 301636 19880 301684
rect 19840 301604 19844 301636
rect 19876 301604 19880 301636
rect 19840 301556 19880 301604
rect 19840 301524 19844 301556
rect 19876 301524 19880 301556
rect 19840 301476 19880 301524
rect 19840 301444 19844 301476
rect 19876 301444 19880 301476
rect 19840 301396 19880 301444
rect 19840 301364 19844 301396
rect 19876 301364 19880 301396
rect 19840 301316 19880 301364
rect 19840 301284 19844 301316
rect 19876 301284 19880 301316
rect 19840 301236 19880 301284
rect 19840 301204 19844 301236
rect 19876 301204 19880 301236
rect 19840 301156 19880 301204
rect 19840 301124 19844 301156
rect 19876 301124 19880 301156
rect 19840 301076 19880 301124
rect 19840 301044 19844 301076
rect 19876 301044 19880 301076
rect 19840 300996 19880 301044
rect 19840 300964 19844 300996
rect 19876 300964 19880 300996
rect 19840 300916 19880 300964
rect 19840 300884 19844 300916
rect 19876 300884 19880 300916
rect 19840 300836 19880 300884
rect 19840 300804 19844 300836
rect 19876 300804 19880 300836
rect 19840 300756 19880 300804
rect 19840 300724 19844 300756
rect 19876 300724 19880 300756
rect 19840 300676 19880 300724
rect 19840 300644 19844 300676
rect 19876 300644 19880 300676
rect 19840 300596 19880 300644
rect 19840 300564 19844 300596
rect 19876 300564 19880 300596
rect 19840 300516 19880 300564
rect 19840 300484 19844 300516
rect 19876 300484 19880 300516
rect 19840 300436 19880 300484
rect 19840 300404 19844 300436
rect 19876 300404 19880 300436
rect 19840 300356 19880 300404
rect 19840 300324 19844 300356
rect 19876 300324 19880 300356
rect 19840 300276 19880 300324
rect 19840 300244 19844 300276
rect 19876 300244 19880 300276
rect 19840 300196 19880 300244
rect 19840 300164 19844 300196
rect 19876 300164 19880 300196
rect 19840 300116 19880 300164
rect 19840 300084 19844 300116
rect 19876 300084 19880 300116
rect 19840 300036 19880 300084
rect 19840 300004 19844 300036
rect 19876 300004 19880 300036
rect 19840 299956 19880 300004
rect 19840 299924 19844 299956
rect 19876 299924 19880 299956
rect 19840 299876 19880 299924
rect 19840 299844 19844 299876
rect 19876 299844 19880 299876
rect 19840 299796 19880 299844
rect 19840 299764 19844 299796
rect 19876 299764 19880 299796
rect 19840 299716 19880 299764
rect 19840 299684 19844 299716
rect 19876 299684 19880 299716
rect 19840 299636 19880 299684
rect 19840 299604 19844 299636
rect 19876 299604 19880 299636
rect 19840 299556 19880 299604
rect 19840 299524 19844 299556
rect 19876 299524 19880 299556
rect 19840 299476 19880 299524
rect 19840 299444 19844 299476
rect 19876 299444 19880 299476
rect 19840 299396 19880 299444
rect 19840 299364 19844 299396
rect 19876 299364 19880 299396
rect 19840 299316 19880 299364
rect 19840 299284 19844 299316
rect 19876 299284 19880 299316
rect 19840 299236 19880 299284
rect 19840 299204 19844 299236
rect 19876 299204 19880 299236
rect 19840 299156 19880 299204
rect 19840 299124 19844 299156
rect 19876 299124 19880 299156
rect 19840 299076 19880 299124
rect 19840 299044 19844 299076
rect 19876 299044 19880 299076
rect 19840 298996 19880 299044
rect 19840 298964 19844 298996
rect 19876 298964 19880 298996
rect 19840 298916 19880 298964
rect 19840 298884 19844 298916
rect 19876 298884 19880 298916
rect 19840 298836 19880 298884
rect 19840 298804 19844 298836
rect 19876 298804 19880 298836
rect 19840 298756 19880 298804
rect 19840 298724 19844 298756
rect 19876 298724 19880 298756
rect 19840 298676 19880 298724
rect 19840 298644 19844 298676
rect 19876 298644 19880 298676
rect 19840 298596 19880 298644
rect 19840 298564 19844 298596
rect 19876 298564 19880 298596
rect 19840 298516 19880 298564
rect 19840 298484 19844 298516
rect 19876 298484 19880 298516
rect 19840 298436 19880 298484
rect 19840 298404 19844 298436
rect 19876 298404 19880 298436
rect 19840 298356 19880 298404
rect 19840 298324 19844 298356
rect 19876 298324 19880 298356
rect 19840 298276 19880 298324
rect 19840 298244 19844 298276
rect 19876 298244 19880 298276
rect 19840 298196 19880 298244
rect 19840 298164 19844 298196
rect 19876 298164 19880 298196
rect 19840 298116 19880 298164
rect 19840 298084 19844 298116
rect 19876 298084 19880 298116
rect 19840 298036 19880 298084
rect 19840 298004 19844 298036
rect 19876 298004 19880 298036
rect 19840 297956 19880 298004
rect 19840 297924 19844 297956
rect 19876 297924 19880 297956
rect 19840 297876 19880 297924
rect 19840 297844 19844 297876
rect 19876 297844 19880 297876
rect 19840 297796 19880 297844
rect 19840 297764 19844 297796
rect 19876 297764 19880 297796
rect 19840 297716 19880 297764
rect 19840 297684 19844 297716
rect 19876 297684 19880 297716
rect 19840 297636 19880 297684
rect 19840 297604 19844 297636
rect 19876 297604 19880 297636
rect 19840 297556 19880 297604
rect 19840 297524 19844 297556
rect 19876 297524 19880 297556
rect 19840 297476 19880 297524
rect 19840 297444 19844 297476
rect 19876 297444 19880 297476
rect 19840 297396 19880 297444
rect 19840 297364 19844 297396
rect 19876 297364 19880 297396
rect 19840 297316 19880 297364
rect 19840 297284 19844 297316
rect 19876 297284 19880 297316
rect 19840 297236 19880 297284
rect 19840 297204 19844 297236
rect 19876 297204 19880 297236
rect 19840 297156 19880 297204
rect 19840 297124 19844 297156
rect 19876 297124 19880 297156
rect 19840 297076 19880 297124
rect 19840 297044 19844 297076
rect 19876 297044 19880 297076
rect 19840 296996 19880 297044
rect 19840 296964 19844 296996
rect 19876 296964 19880 296996
rect 19840 296916 19880 296964
rect 19840 296884 19844 296916
rect 19876 296884 19880 296916
rect 19840 296836 19880 296884
rect 19840 296804 19844 296836
rect 19876 296804 19880 296836
rect 19840 296756 19880 296804
rect 19840 296724 19844 296756
rect 19876 296724 19880 296756
rect 19840 296676 19880 296724
rect 19840 296644 19844 296676
rect 19876 296644 19880 296676
rect 19840 296596 19880 296644
rect 19840 296564 19844 296596
rect 19876 296564 19880 296596
rect 19840 296516 19880 296564
rect 19840 296484 19844 296516
rect 19876 296484 19880 296516
rect 19840 296436 19880 296484
rect 19840 296404 19844 296436
rect 19876 296404 19880 296436
rect 19840 296356 19880 296404
rect 19840 296324 19844 296356
rect 19876 296324 19880 296356
rect 19840 296276 19880 296324
rect 19840 296244 19844 296276
rect 19876 296244 19880 296276
rect 19840 296196 19880 296244
rect 19840 296164 19844 296196
rect 19876 296164 19880 296196
rect 19840 296116 19880 296164
rect 19840 296084 19844 296116
rect 19876 296084 19880 296116
rect 19840 296036 19880 296084
rect 19840 296004 19844 296036
rect 19876 296004 19880 296036
rect 19840 295956 19880 296004
rect 19840 295924 19844 295956
rect 19876 295924 19880 295956
rect 19840 295876 19880 295924
rect 19840 295844 19844 295876
rect 19876 295844 19880 295876
rect 19840 295796 19880 295844
rect 19840 295764 19844 295796
rect 19876 295764 19880 295796
rect 19840 295716 19880 295764
rect 19840 295684 19844 295716
rect 19876 295684 19880 295716
rect 19840 295636 19880 295684
rect 19840 295604 19844 295636
rect 19876 295604 19880 295636
rect 19840 295556 19880 295604
rect 19840 295524 19844 295556
rect 19876 295524 19880 295556
rect 19840 295476 19880 295524
rect 19840 295444 19844 295476
rect 19876 295444 19880 295476
rect 19840 295396 19880 295444
rect 19840 295364 19844 295396
rect 19876 295364 19880 295396
rect 19840 295316 19880 295364
rect 19840 295284 19844 295316
rect 19876 295284 19880 295316
rect 19840 295236 19880 295284
rect 19840 295204 19844 295236
rect 19876 295204 19880 295236
rect 19840 295156 19880 295204
rect 19840 295124 19844 295156
rect 19876 295124 19880 295156
rect 19840 295076 19880 295124
rect 19840 295044 19844 295076
rect 19876 295044 19880 295076
rect 19840 294996 19880 295044
rect 19840 294964 19844 294996
rect 19876 294964 19880 294996
rect 19840 294916 19880 294964
rect 19840 294884 19844 294916
rect 19876 294884 19880 294916
rect 19840 294836 19880 294884
rect 19840 294804 19844 294836
rect 19876 294804 19880 294836
rect 19840 294756 19880 294804
rect 19840 294724 19844 294756
rect 19876 294724 19880 294756
rect 291760 294736 292400 294792
rect 19840 294676 19880 294724
rect 19840 294644 19844 294676
rect 19876 294644 19880 294676
rect 19840 294596 19880 294644
rect 19840 294564 19844 294596
rect 19876 294564 19880 294596
rect 19840 294516 19880 294564
rect 19840 294484 19844 294516
rect 19876 294484 19880 294516
rect 19840 294436 19880 294484
rect 19840 294404 19844 294436
rect 19876 294404 19880 294436
rect 19840 294356 19880 294404
rect 19840 294324 19844 294356
rect 19876 294324 19880 294356
rect 19840 294276 19880 294324
rect 19840 294244 19844 294276
rect 19876 294244 19880 294276
rect 19840 294196 19880 294244
rect 19840 294164 19844 294196
rect 19876 294164 19880 294196
rect 19840 294116 19880 294164
rect 291760 294145 292400 294201
rect 19840 294084 19844 294116
rect 19876 294084 19880 294116
rect 19840 294036 19880 294084
rect 19840 294004 19844 294036
rect 19876 294004 19880 294036
rect 19840 293956 19880 294004
rect 19840 293924 19844 293956
rect 19876 293924 19880 293956
rect 19840 293876 19880 293924
rect 19840 293844 19844 293876
rect 19876 293844 19880 293876
rect 19840 293796 19880 293844
rect 19840 293764 19844 293796
rect 19876 293764 19880 293796
rect 19840 293716 19880 293764
rect 19840 293684 19844 293716
rect 19876 293684 19880 293716
rect 19840 293636 19880 293684
rect 19840 293604 19844 293636
rect 19876 293604 19880 293636
rect 19840 293556 19880 293604
rect 19840 293524 19844 293556
rect 19876 293524 19880 293556
rect 291760 293554 292400 293610
rect 19840 293476 19880 293524
rect 19840 293444 19844 293476
rect 19876 293444 19880 293476
rect 19840 293396 19880 293444
rect 19840 293364 19844 293396
rect 19876 293364 19880 293396
rect 19840 293316 19880 293364
rect 19840 293284 19844 293316
rect 19876 293284 19880 293316
rect 19840 293236 19880 293284
rect 19840 293204 19844 293236
rect 19876 293204 19880 293236
rect 19840 293156 19880 293204
rect 19840 293124 19844 293156
rect 19876 293124 19880 293156
rect 19840 293076 19880 293124
rect 19840 293044 19844 293076
rect 19876 293044 19880 293076
rect 19840 292996 19880 293044
rect 19840 292964 19844 292996
rect 19876 292964 19880 292996
rect 19840 292916 19880 292964
rect 291760 292963 292400 293019
rect 19840 292884 19844 292916
rect 19876 292884 19880 292916
rect 19840 292836 19880 292884
rect 19840 292804 19844 292836
rect 19876 292804 19880 292836
rect 19840 292756 19880 292804
rect 19840 292724 19844 292756
rect 19876 292724 19880 292756
rect 19840 292676 19880 292724
rect 19840 292644 19844 292676
rect 19876 292644 19880 292676
rect 19840 292596 19880 292644
rect 19840 292564 19844 292596
rect 19876 292564 19880 292596
rect 19840 292516 19880 292564
rect 19840 292484 19844 292516
rect 19876 292484 19880 292516
rect 19840 292436 19880 292484
rect 19840 292404 19844 292436
rect 19876 292404 19880 292436
rect 19840 292356 19880 292404
rect 291760 292372 292400 292428
rect 19840 292324 19844 292356
rect 19876 292324 19880 292356
rect 19840 292276 19880 292324
rect 19840 292244 19844 292276
rect 19876 292244 19880 292276
rect 19840 292196 19880 292244
rect 19840 292164 19844 292196
rect 19876 292164 19880 292196
rect 19840 292116 19880 292164
rect 19840 292084 19844 292116
rect 19876 292084 19880 292116
rect 19840 292036 19880 292084
rect 19840 292004 19844 292036
rect 19876 292004 19880 292036
rect 19840 291956 19880 292004
rect 19840 291924 19844 291956
rect 19876 291924 19880 291956
rect 19840 291876 19880 291924
rect 19840 291844 19844 291876
rect 19876 291844 19880 291876
rect 19840 291796 19880 291844
rect 19840 291764 19844 291796
rect 19876 291764 19880 291796
rect 291760 291781 292400 291837
rect 19840 291716 19880 291764
rect 19840 291684 19844 291716
rect 19876 291684 19880 291716
rect 19840 291636 19880 291684
rect 19840 291604 19844 291636
rect 19876 291604 19880 291636
rect 19840 291556 19880 291604
rect 19840 291524 19844 291556
rect 19876 291524 19880 291556
rect 19840 291476 19880 291524
rect 19840 291444 19844 291476
rect 19876 291444 19880 291476
rect 19840 291396 19880 291444
rect 19840 291364 19844 291396
rect 19876 291364 19880 291396
rect 19840 291316 19880 291364
rect 19840 291284 19844 291316
rect 19876 291284 19880 291316
rect 19840 291236 19880 291284
rect 19840 291204 19844 291236
rect 19876 291204 19880 291236
rect 19840 291156 19880 291204
rect 19840 291124 19844 291156
rect 19876 291124 19880 291156
rect 19840 291076 19880 291124
rect 19840 291044 19844 291076
rect 19876 291044 19880 291076
rect 19840 290996 19880 291044
rect 19840 290964 19844 290996
rect 19876 290964 19880 290996
rect 19840 290916 19880 290964
rect 19840 290884 19844 290916
rect 19876 290884 19880 290916
rect 19840 290836 19880 290884
rect 19840 290804 19844 290836
rect 19876 290804 19880 290836
rect 19840 290756 19880 290804
rect 19840 290724 19844 290756
rect 19876 290724 19880 290756
rect 19840 290676 19880 290724
rect 19840 290644 19844 290676
rect 19876 290644 19880 290676
rect 19840 290596 19880 290644
rect 19840 290564 19844 290596
rect 19876 290564 19880 290596
rect 19840 290516 19880 290564
rect 19840 290484 19844 290516
rect 19876 290484 19880 290516
rect 19840 290436 19880 290484
rect 19840 290404 19844 290436
rect 19876 290404 19880 290436
rect 19840 290356 19880 290404
rect 19840 290324 19844 290356
rect 19876 290324 19880 290356
rect 19840 290276 19880 290324
rect 19840 290244 19844 290276
rect 19876 290244 19880 290276
rect 19840 290196 19880 290244
rect 19840 290164 19844 290196
rect 19876 290164 19880 290196
rect 19840 290116 19880 290164
rect 19840 290084 19844 290116
rect 19876 290084 19880 290116
rect 19840 290036 19880 290084
rect 19840 290004 19844 290036
rect 19876 290004 19880 290036
rect 19840 289956 19880 290004
rect 19840 289924 19844 289956
rect 19876 289924 19880 289956
rect 19840 289876 19880 289924
rect 19840 289844 19844 289876
rect 19876 289844 19880 289876
rect 19840 289796 19880 289844
rect 19840 289764 19844 289796
rect 19876 289764 19880 289796
rect 19840 289716 19880 289764
rect 19840 289684 19844 289716
rect 19876 289684 19880 289716
rect 19840 289636 19880 289684
rect 19840 289604 19844 289636
rect 19876 289604 19880 289636
rect 19840 289556 19880 289604
rect 19840 289524 19844 289556
rect 19876 289524 19880 289556
rect 19840 289476 19880 289524
rect 19840 289444 19844 289476
rect 19876 289444 19880 289476
rect 19840 289396 19880 289444
rect 19840 289364 19844 289396
rect 19876 289364 19880 289396
rect 19840 289316 19880 289364
rect 19840 289284 19844 289316
rect 19876 289284 19880 289316
rect 19840 289236 19880 289284
rect 19840 289204 19844 289236
rect 19876 289204 19880 289236
rect 19840 289156 19880 289204
rect 19840 289124 19844 289156
rect 19876 289124 19880 289156
rect 19840 289076 19880 289124
rect 19840 289044 19844 289076
rect 19876 289044 19880 289076
rect 19840 288996 19880 289044
rect 19840 288964 19844 288996
rect 19876 288964 19880 288996
rect 19840 288916 19880 288964
rect 19840 288884 19844 288916
rect 19876 288884 19880 288916
rect 19840 288836 19880 288884
rect 19840 288804 19844 288836
rect 19876 288804 19880 288836
rect 19840 288756 19880 288804
rect 19840 288724 19844 288756
rect 19876 288724 19880 288756
rect 19840 288676 19880 288724
rect 19840 288644 19844 288676
rect 19876 288644 19880 288676
rect 19840 288596 19880 288644
rect 19840 288564 19844 288596
rect 19876 288564 19880 288596
rect 19840 288516 19880 288564
rect 19840 288484 19844 288516
rect 19876 288484 19880 288516
rect 19840 288436 19880 288484
rect 19840 288404 19844 288436
rect 19876 288404 19880 288436
rect 19840 288356 19880 288404
rect 19840 288324 19844 288356
rect 19876 288324 19880 288356
rect 19840 288276 19880 288324
rect 19840 288244 19844 288276
rect 19876 288244 19880 288276
rect 19840 288196 19880 288244
rect 19840 288164 19844 288196
rect 19876 288164 19880 288196
rect 19840 288116 19880 288164
rect 19840 288084 19844 288116
rect 19876 288084 19880 288116
rect 19840 288036 19880 288084
rect 19840 288004 19844 288036
rect 19876 288004 19880 288036
rect 19840 287956 19880 288004
rect 19840 287924 19844 287956
rect 19876 287924 19880 287956
rect 19840 287876 19880 287924
rect 19840 287844 19844 287876
rect 19876 287844 19880 287876
rect 19840 287796 19880 287844
rect 19840 287764 19844 287796
rect 19876 287764 19880 287796
rect 19840 287716 19880 287764
rect 19840 287684 19844 287716
rect 19876 287684 19880 287716
rect 19840 287636 19880 287684
rect 19840 287604 19844 287636
rect 19876 287604 19880 287636
rect 19840 287556 19880 287604
rect 19840 287524 19844 287556
rect 19876 287524 19880 287556
rect 19840 287476 19880 287524
rect 19840 287444 19844 287476
rect 19876 287444 19880 287476
rect 19840 287396 19880 287444
rect 19840 287364 19844 287396
rect 19876 287364 19880 287396
rect 19840 287316 19880 287364
rect 19840 287284 19844 287316
rect 19876 287284 19880 287316
rect 19840 287236 19880 287284
rect 19840 287204 19844 287236
rect 19876 287204 19880 287236
rect 19840 287156 19880 287204
rect 19840 287124 19844 287156
rect 19876 287124 19880 287156
rect 19840 287076 19880 287124
rect 19840 287044 19844 287076
rect 19876 287044 19880 287076
rect 19840 286996 19880 287044
rect 19840 286964 19844 286996
rect 19876 286964 19880 286996
rect 19840 286916 19880 286964
rect 19840 286884 19844 286916
rect 19876 286884 19880 286916
rect 19840 286836 19880 286884
rect 19840 286804 19844 286836
rect 19876 286804 19880 286836
rect 19840 286756 19880 286804
rect 19840 286724 19844 286756
rect 19876 286724 19880 286756
rect 19840 286676 19880 286724
rect 19840 286644 19844 286676
rect 19876 286644 19880 286676
rect 19840 286596 19880 286644
rect 19840 286564 19844 286596
rect 19876 286564 19880 286596
rect 19840 286516 19880 286564
rect 19840 286484 19844 286516
rect 19876 286484 19880 286516
rect 19840 286436 19880 286484
rect 19840 286404 19844 286436
rect 19876 286404 19880 286436
rect 19840 286356 19880 286404
rect 19840 286324 19844 286356
rect 19876 286324 19880 286356
rect 19840 286276 19880 286324
rect 19840 286244 19844 286276
rect 19876 286244 19880 286276
rect 19840 286196 19880 286244
rect 19840 286164 19844 286196
rect 19876 286164 19880 286196
rect 19840 286116 19880 286164
rect 19840 286084 19844 286116
rect 19876 286084 19880 286116
rect 19840 286036 19880 286084
rect 19840 286004 19844 286036
rect 19876 286004 19880 286036
rect 19840 285956 19880 286004
rect 19840 285924 19844 285956
rect 19876 285924 19880 285956
rect 19840 285876 19880 285924
rect 19840 285844 19844 285876
rect 19876 285844 19880 285876
rect 19840 285796 19880 285844
rect 19840 285764 19844 285796
rect 19876 285764 19880 285796
rect 19840 285716 19880 285764
rect 19840 285684 19844 285716
rect 19876 285684 19880 285716
rect 19840 285636 19880 285684
rect 19840 285604 19844 285636
rect 19876 285604 19880 285636
rect 19840 285556 19880 285604
rect 19840 285524 19844 285556
rect 19876 285524 19880 285556
rect 19840 285476 19880 285524
rect 19840 285444 19844 285476
rect 19876 285444 19880 285476
rect 19840 285396 19880 285444
rect 19840 285364 19844 285396
rect 19876 285364 19880 285396
rect 19840 285316 19880 285364
rect 19840 285284 19844 285316
rect 19876 285284 19880 285316
rect 19840 285236 19880 285284
rect 19840 285204 19844 285236
rect 19876 285204 19880 285236
rect 19840 285156 19880 285204
rect 19840 285124 19844 285156
rect 19876 285124 19880 285156
rect 19840 285076 19880 285124
rect 19840 285044 19844 285076
rect 19876 285044 19880 285076
rect 19840 284996 19880 285044
rect 19840 284964 19844 284996
rect 19876 284964 19880 284996
rect 19840 284916 19880 284964
rect 19840 284884 19844 284916
rect 19876 284884 19880 284916
rect 19840 284836 19880 284884
rect 19840 284804 19844 284836
rect 19876 284804 19880 284836
rect 19840 284756 19880 284804
rect 19840 284724 19844 284756
rect 19876 284724 19880 284756
rect 19840 284676 19880 284724
rect 19840 284644 19844 284676
rect 19876 284644 19880 284676
rect 19840 284596 19880 284644
rect 19840 284564 19844 284596
rect 19876 284564 19880 284596
rect 19840 284516 19880 284564
rect 19840 284484 19844 284516
rect 19876 284484 19880 284516
rect 19840 284436 19880 284484
rect 19840 284404 19844 284436
rect 19876 284404 19880 284436
rect 19840 284356 19880 284404
rect 19840 284324 19844 284356
rect 19876 284324 19880 284356
rect 19840 284276 19880 284324
rect 19840 284244 19844 284276
rect 19876 284244 19880 284276
rect 19840 284196 19880 284244
rect 19840 284164 19844 284196
rect 19876 284164 19880 284196
rect 19840 284116 19880 284164
rect 19840 284084 19844 284116
rect 19876 284084 19880 284116
rect 19840 284036 19880 284084
rect 19840 284004 19844 284036
rect 19876 284004 19880 284036
rect 19840 283956 19880 284004
rect 19840 283924 19844 283956
rect 19876 283924 19880 283956
rect 19840 283876 19880 283924
rect 19840 283844 19844 283876
rect 19876 283844 19880 283876
rect 19840 283796 19880 283844
rect 19840 283764 19844 283796
rect 19876 283764 19880 283796
rect 19840 283716 19880 283764
rect 19840 283684 19844 283716
rect 19876 283684 19880 283716
rect 19840 283636 19880 283684
rect 19840 283604 19844 283636
rect 19876 283604 19880 283636
rect 19840 283556 19880 283604
rect 19840 283524 19844 283556
rect 19876 283524 19880 283556
rect 19840 283476 19880 283524
rect 19840 283444 19844 283476
rect 19876 283444 19880 283476
rect 19840 283396 19880 283444
rect 19840 283364 19844 283396
rect 19876 283364 19880 283396
rect 19840 283316 19880 283364
rect 19840 283284 19844 283316
rect 19876 283284 19880 283316
rect 19840 283236 19880 283284
rect 19840 283204 19844 283236
rect 19876 283204 19880 283236
rect 19840 283156 19880 283204
rect 19840 283124 19844 283156
rect 19876 283124 19880 283156
rect 19840 283076 19880 283124
rect 19840 283044 19844 283076
rect 19876 283044 19880 283076
rect 19840 282996 19880 283044
rect 19840 282964 19844 282996
rect 19876 282964 19880 282996
rect 19840 282916 19880 282964
rect 19840 282884 19844 282916
rect 19876 282884 19880 282916
rect 19840 282836 19880 282884
rect 19840 282804 19844 282836
rect 19876 282804 19880 282836
rect 19840 282756 19880 282804
rect 19840 282724 19844 282756
rect 19876 282724 19880 282756
rect 19840 282676 19880 282724
rect 19840 282644 19844 282676
rect 19876 282644 19880 282676
rect 19840 282596 19880 282644
rect 19840 282564 19844 282596
rect 19876 282564 19880 282596
rect 19840 282516 19880 282564
rect 19840 282484 19844 282516
rect 19876 282484 19880 282516
rect 19840 282436 19880 282484
rect 19840 282404 19844 282436
rect 19876 282404 19880 282436
rect 19840 282356 19880 282404
rect 19840 282324 19844 282356
rect 19876 282324 19880 282356
rect 19840 282276 19880 282324
rect 19840 282244 19844 282276
rect 19876 282244 19880 282276
rect 19840 282196 19880 282244
rect 19840 282164 19844 282196
rect 19876 282164 19880 282196
rect 19840 282116 19880 282164
rect 19840 282084 19844 282116
rect 19876 282084 19880 282116
rect 19840 282036 19880 282084
rect 19840 282004 19844 282036
rect 19876 282004 19880 282036
rect 19840 281956 19880 282004
rect 19840 281924 19844 281956
rect 19876 281924 19880 281956
rect 19840 281876 19880 281924
rect 19840 281844 19844 281876
rect 19876 281844 19880 281876
rect 19840 281796 19880 281844
rect 19840 281764 19844 281796
rect 19876 281764 19880 281796
rect 19840 281716 19880 281764
rect 19840 281684 19844 281716
rect 19876 281684 19880 281716
rect 19840 281636 19880 281684
rect 19840 281604 19844 281636
rect 19876 281604 19880 281636
rect 19840 281556 19880 281604
rect 19840 281524 19844 281556
rect 19876 281524 19880 281556
rect 19840 281476 19880 281524
rect 19840 281444 19844 281476
rect 19876 281444 19880 281476
rect 19840 281396 19880 281444
rect 19840 281364 19844 281396
rect 19876 281364 19880 281396
rect 19840 281316 19880 281364
rect 19840 281284 19844 281316
rect 19876 281284 19880 281316
rect 19840 281236 19880 281284
rect 19840 281204 19844 281236
rect 19876 281204 19880 281236
rect 19840 281156 19880 281204
rect 19840 281124 19844 281156
rect 19876 281124 19880 281156
rect 19840 281076 19880 281124
rect 19840 281044 19844 281076
rect 19876 281044 19880 281076
rect 19840 280996 19880 281044
rect 19840 280964 19844 280996
rect 19876 280964 19880 280996
rect 19840 280916 19880 280964
rect 19840 280884 19844 280916
rect 19876 280884 19880 280916
rect 19840 280836 19880 280884
rect 19840 280804 19844 280836
rect 19876 280804 19880 280836
rect 19840 280756 19880 280804
rect 19840 280724 19844 280756
rect 19876 280724 19880 280756
rect 19840 280676 19880 280724
rect 19840 280644 19844 280676
rect 19876 280644 19880 280676
rect 19840 280596 19880 280644
rect 19840 280564 19844 280596
rect 19876 280564 19880 280596
rect 19840 280516 19880 280564
rect 19840 280484 19844 280516
rect 19876 280484 19880 280516
rect 19840 280436 19880 280484
rect 19840 280404 19844 280436
rect 19876 280404 19880 280436
rect 19840 280356 19880 280404
rect 19840 280324 19844 280356
rect 19876 280324 19880 280356
rect 19840 280276 19880 280324
rect 19840 280244 19844 280276
rect 19876 280244 19880 280276
rect 19840 280196 19880 280244
rect 19840 280164 19844 280196
rect 19876 280164 19880 280196
rect 19840 280116 19880 280164
rect 19840 280084 19844 280116
rect 19876 280084 19880 280116
rect 19840 280036 19880 280084
rect 19840 280004 19844 280036
rect 19876 280004 19880 280036
rect 19840 279956 19880 280004
rect 19840 279924 19844 279956
rect 19876 279924 19880 279956
rect 19840 279876 19880 279924
rect 19840 279844 19844 279876
rect 19876 279844 19880 279876
rect 19840 279796 19880 279844
rect 19840 279764 19844 279796
rect 19876 279764 19880 279796
rect 19840 279716 19880 279764
rect 19840 279684 19844 279716
rect 19876 279684 19880 279716
rect 19840 279636 19880 279684
rect 19840 279604 19844 279636
rect 19876 279604 19880 279636
rect 19840 279556 19880 279604
rect 19840 279524 19844 279556
rect 19876 279524 19880 279556
rect 19840 279476 19880 279524
rect 19840 279444 19844 279476
rect 19876 279444 19880 279476
rect 19840 279396 19880 279444
rect 19840 279364 19844 279396
rect 19876 279364 19880 279396
rect 19840 279316 19880 279364
rect 19840 279284 19844 279316
rect 19876 279284 19880 279316
rect 19840 279236 19880 279284
rect 19840 279204 19844 279236
rect 19876 279204 19880 279236
rect 19840 279156 19880 279204
rect 19840 279124 19844 279156
rect 19876 279124 19880 279156
rect 19840 279076 19880 279124
rect 19840 279044 19844 279076
rect 19876 279044 19880 279076
rect 19840 278996 19880 279044
rect 19840 278964 19844 278996
rect 19876 278964 19880 278996
rect 19840 278916 19880 278964
rect 19840 278884 19844 278916
rect 19876 278884 19880 278916
rect 19840 278836 19880 278884
rect 19840 278804 19844 278836
rect 19876 278804 19880 278836
rect 19840 278756 19880 278804
rect 19840 278724 19844 278756
rect 19876 278724 19880 278756
rect 19840 278676 19880 278724
rect 19840 278644 19844 278676
rect 19876 278644 19880 278676
rect 19680 278484 19684 278516
rect 19716 278484 19720 278516
rect 19680 278480 19720 278484
rect 19840 278516 19880 278644
rect 19840 278484 19844 278516
rect 19876 278484 19880 278516
rect 19840 278480 19880 278484
rect 17200 278404 17204 278436
rect 17236 278404 17240 278436
rect 17200 278356 17240 278404
rect 17200 278324 17204 278356
rect 17236 278324 17240 278356
rect 17200 278276 17240 278324
rect 17200 278244 17204 278276
rect 17236 278244 17240 278276
rect 17200 278196 17240 278244
rect 17200 278164 17204 278196
rect 17236 278164 17240 278196
rect 17200 278116 17240 278164
rect 17200 278084 17204 278116
rect 17236 278084 17240 278116
rect 17200 278036 17240 278084
rect 17200 278004 17204 278036
rect 17236 278004 17240 278036
rect 17200 277956 17240 278004
rect 17200 277924 17204 277956
rect 17236 277924 17240 277956
rect 17200 277876 17240 277924
rect 17200 277844 17204 277876
rect 17236 277844 17240 277876
rect 17200 277800 17240 277844
rect 17360 277800 17400 277840
rect 14220 275700 14300 275800
rect 13520 275195 13560 275200
rect 13520 275005 13525 275195
rect 13555 275005 13560 275195
rect 13520 274880 13560 275005
rect 13680 275195 13720 275200
rect 13680 275005 13685 275195
rect 13715 275005 13720 275195
rect 13680 274920 13720 275005
rect 13840 275195 13880 275200
rect 13840 275005 13845 275195
rect 13875 275005 13880 275195
rect 13840 274920 13880 275005
rect 14000 275195 14040 275200
rect 14000 275005 14005 275195
rect 14035 275005 14040 275195
rect 14000 274920 14040 275005
rect 14160 275195 14200 275200
rect 14160 275005 14165 275195
rect 14195 275005 14200 275195
rect 14160 274920 14200 275005
rect 14240 274920 14280 275700
rect 14320 275195 14360 275200
rect 14320 275005 14325 275195
rect 14355 275005 14360 275195
rect 14320 274920 14360 275005
rect 27920 275195 27960 275440
rect 27920 275005 27925 275195
rect 27955 275005 27960 275195
rect 27920 274880 27960 275005
rect 28080 275195 28120 275440
rect 28080 275005 28085 275195
rect 28115 275005 28120 275195
rect 28080 274920 28120 275005
rect 28240 275195 28280 275440
rect 28240 275005 28245 275195
rect 28275 275005 28280 275195
rect 28240 274920 28280 275005
rect 28400 275356 28440 275440
rect 28400 275324 28404 275356
rect 28436 275324 28440 275356
rect 28400 275276 28440 275324
rect 28400 275244 28404 275276
rect 28436 275244 28440 275276
rect 28400 275195 28440 275244
rect 28400 275005 28405 275195
rect 28435 275005 28440 275195
rect 28400 274920 28440 275005
rect 28480 274920 28520 275400
rect 28560 275356 28600 275440
rect 28560 275324 28564 275356
rect 28596 275324 28600 275356
rect 28560 275276 28600 275324
rect 28560 275244 28564 275276
rect 28596 275244 28600 275276
rect 28560 275195 28600 275244
rect 28560 275005 28565 275195
rect 28595 275005 28600 275195
rect 28560 274920 28600 275005
rect 28640 274920 28680 275400
rect 28720 275356 28760 275440
rect 28720 275324 28724 275356
rect 28756 275324 28760 275356
rect 28720 275276 28760 275324
rect 291170 275281 292400 277681
rect 28720 275244 28724 275276
rect 28756 275244 28760 275276
rect 28720 275195 28760 275244
rect 28720 275005 28725 275195
rect 28755 275005 28760 275195
rect 28720 274920 28760 275005
rect 291170 270281 292400 272681
rect 2800 263360 2840 263400
rect 2960 263360 3000 263400
rect 3120 263360 3160 263400
rect 3280 263360 3320 263400
rect 3440 263360 3480 263400
rect 2800 263320 3480 263360
rect 2800 263200 3000 263320
rect 17200 263200 17240 263400
rect 17360 263200 17400 263400
rect 17520 263200 17560 263400
rect 17680 263200 17720 263400
rect 17840 263200 17880 263400
rect 2400 263000 17880 263200
rect -400 255765 240 255821
rect -400 255174 240 255230
rect -400 254583 240 254639
rect -400 253992 240 254048
rect -400 253401 240 253457
rect -400 252810 240 252866
rect -400 234154 240 234210
rect -400 233563 240 233619
rect -400 232972 240 233028
rect -400 232381 240 232437
rect -400 231790 240 231846
rect -400 231199 240 231255
rect -400 212543 240 212599
rect -400 211952 240 212008
rect -400 211361 240 211417
rect -400 210770 240 210826
rect -400 210179 240 210235
rect -400 209588 240 209644
rect -400 190932 240 190988
rect -400 190341 240 190397
rect -400 189750 240 189806
rect -400 189159 240 189215
rect -400 188568 240 188624
rect -400 187977 240 188033
rect -400 169321 240 169377
rect -400 168730 240 168786
rect -400 168139 240 168195
rect -400 167548 240 167604
rect -400 166957 240 167013
rect -400 166366 240 166422
rect -400 147710 240 147766
rect -400 147119 240 147175
rect -400 146528 240 146584
rect -400 145937 240 145993
rect -400 145346 240 145402
rect -400 144755 240 144811
rect -400 126199 240 126255
rect -400 125608 240 125664
rect -400 125017 240 125073
rect -400 124426 240 124482
rect -400 123835 240 123891
rect -400 123244 240 123300
rect -400 109800 830 109844
rect 2800 109800 3000 263000
rect 291760 250025 292400 250081
rect 291760 249434 292400 249490
rect 291760 248843 292400 248899
rect 291760 248252 292400 248308
rect 291760 247661 292400 247717
rect 291760 247070 292400 247126
rect 291760 227814 292400 227870
rect 291760 227223 292400 227279
rect 291760 226632 292400 226688
rect 291760 226041 292400 226097
rect 291760 225450 292400 225506
rect 291760 224859 292400 224915
rect 291760 205603 292400 205659
rect 291760 205012 292400 205068
rect 291760 204421 292400 204477
rect 291760 203830 292400 203886
rect 291760 203239 292400 203295
rect 291760 202648 292400 202704
rect 291760 182392 292400 182448
rect 291760 181801 292400 181857
rect 291760 181210 292400 181266
rect 291760 180619 292400 180675
rect 291760 180028 292400 180084
rect 291760 179437 292400 179493
rect 291760 159781 292400 159837
rect 291760 159190 292400 159246
rect 291760 158599 292400 158655
rect 291760 158008 292400 158064
rect 291760 157417 292400 157473
rect 291760 156826 292400 156882
rect 291760 137570 292400 137626
rect 291760 136979 292400 137035
rect 291760 136388 292400 136444
rect 291760 135797 292400 135853
rect 291760 135206 292400 135262
rect 291760 134615 292400 134671
rect 291170 117615 292400 120015
rect 291170 112615 292400 115015
rect -400 109600 3000 109800
rect -400 107444 830 109600
rect -400 102444 830 104844
rect 291170 95715 292400 98115
rect 291170 90715 292400 93115
rect -400 86444 830 88844
rect -400 81444 830 83844
rect 291170 73415 292400 75815
rect 291170 68415 292400 70815
rect -400 62388 240 62444
rect -400 61797 240 61853
rect -400 61206 240 61262
rect -400 60615 240 60671
rect -400 60024 240 60080
rect -400 59433 240 59489
rect 291760 47559 292400 47615
rect 291760 46968 292400 47024
rect 291760 46377 292400 46433
rect 291760 45786 292400 45842
rect -400 40777 240 40833
rect -400 40186 240 40242
rect -400 39595 240 39651
rect -400 39004 240 39060
rect -400 38413 240 38469
rect -400 37822 240 37878
rect 291760 25230 292400 25286
rect 291760 24639 292400 24695
rect 291760 24048 292400 24104
rect 291760 23457 292400 23513
rect -400 19166 240 19222
rect -400 18575 240 18631
rect -400 17984 240 18040
rect -400 17393 240 17449
rect -400 16802 240 16858
rect -400 16211 240 16267
rect 291760 12001 292400 12057
rect 291760 11410 292400 11466
rect 291760 10819 292400 10875
rect 291760 10228 292400 10284
rect 291760 9637 292400 9693
rect 291760 9046 292400 9102
rect -400 8455 240 8511
rect 291760 8455 292400 8511
rect -400 7864 240 7920
rect 291760 7864 292400 7920
rect -400 7273 240 7329
rect 291760 7273 292400 7329
rect -400 6682 240 6738
rect 291760 6682 292400 6738
rect -400 6091 240 6147
rect 291760 6091 292400 6147
rect -400 5500 240 5556
rect 291760 5500 292400 5556
rect -400 4909 240 4965
rect 291760 4909 292400 4965
rect -400 4318 240 4374
rect 291760 4318 292400 4374
rect -400 3727 240 3783
rect 291760 3727 292400 3783
rect -400 3136 240 3192
rect 291760 3136 292400 3192
rect -400 2545 240 2601
rect 291760 2545 292400 2601
rect -400 1954 240 2010
rect 291760 1954 292400 2010
rect -400 1363 240 1419
rect 291760 1363 292400 1419
rect -400 772 240 828
rect 291760 772 292400 828
<< via3 >>
rect 10724 351395 10756 351396
rect 10724 351365 10725 351395
rect 10725 351365 10755 351395
rect 10755 351365 10756 351395
rect 10724 351364 10756 351365
rect 10724 351284 10756 351316
rect 10724 351235 10756 351236
rect 10724 351205 10725 351235
rect 10725 351205 10755 351235
rect 10755 351205 10756 351235
rect 10724 351204 10756 351205
rect 10804 351395 10836 351396
rect 10804 351365 10805 351395
rect 10805 351365 10835 351395
rect 10835 351365 10836 351395
rect 10804 351364 10836 351365
rect 10804 351284 10836 351316
rect 10804 351235 10836 351236
rect 10804 351205 10805 351235
rect 10805 351205 10835 351235
rect 10835 351205 10836 351235
rect 10804 351204 10836 351205
rect 10884 351395 10916 351396
rect 10884 351365 10885 351395
rect 10885 351365 10915 351395
rect 10915 351365 10916 351395
rect 10884 351364 10916 351365
rect 10884 351284 10916 351316
rect 10884 351235 10916 351236
rect 10884 351205 10885 351235
rect 10885 351205 10915 351235
rect 10915 351205 10916 351235
rect 10884 351204 10916 351205
rect 10964 351395 10996 351396
rect 10964 351365 10965 351395
rect 10965 351365 10995 351395
rect 10995 351365 10996 351395
rect 10964 351364 10996 351365
rect 10964 351284 10996 351316
rect 10964 351235 10996 351236
rect 10964 351205 10965 351235
rect 10965 351205 10995 351235
rect 10995 351205 10996 351235
rect 10964 351204 10996 351205
rect 11044 351395 11076 351396
rect 11044 351365 11045 351395
rect 11045 351365 11075 351395
rect 11075 351365 11076 351395
rect 11044 351364 11076 351365
rect 11044 351284 11076 351316
rect 11044 351235 11076 351236
rect 11044 351205 11045 351235
rect 11045 351205 11075 351235
rect 11075 351205 11076 351235
rect 11044 351204 11076 351205
rect 11124 351395 11156 351396
rect 11124 351365 11125 351395
rect 11125 351365 11155 351395
rect 11155 351365 11156 351395
rect 11124 351364 11156 351365
rect 11124 351284 11156 351316
rect 11124 351235 11156 351236
rect 11124 351205 11125 351235
rect 11125 351205 11155 351235
rect 11155 351205 11156 351235
rect 11124 351204 11156 351205
rect 11204 351395 11236 351396
rect 11204 351365 11205 351395
rect 11205 351365 11235 351395
rect 11235 351365 11236 351395
rect 11204 351364 11236 351365
rect 11204 351284 11236 351316
rect 11204 351235 11236 351236
rect 11204 351205 11205 351235
rect 11205 351205 11235 351235
rect 11235 351205 11236 351235
rect 11204 351204 11236 351205
rect 11284 351395 11316 351396
rect 11284 351365 11285 351395
rect 11285 351365 11315 351395
rect 11315 351365 11316 351395
rect 11284 351364 11316 351365
rect 11284 351284 11316 351316
rect 11284 351235 11316 351236
rect 11284 351205 11285 351235
rect 11285 351205 11315 351235
rect 11315 351205 11316 351235
rect 11284 351204 11316 351205
rect 11364 351395 11396 351396
rect 11364 351365 11365 351395
rect 11365 351365 11395 351395
rect 11395 351365 11396 351395
rect 11364 351364 11396 351365
rect 11364 351284 11396 351316
rect 11364 351235 11396 351236
rect 11364 351205 11365 351235
rect 11365 351205 11395 351235
rect 11395 351205 11396 351235
rect 11364 351204 11396 351205
rect 11444 351395 11476 351396
rect 11444 351365 11445 351395
rect 11445 351365 11475 351395
rect 11475 351365 11476 351395
rect 11444 351364 11476 351365
rect 11444 351284 11476 351316
rect 11444 351235 11476 351236
rect 11444 351205 11445 351235
rect 11445 351205 11475 351235
rect 11475 351205 11476 351235
rect 11444 351204 11476 351205
rect 11524 351395 11556 351396
rect 11524 351365 11525 351395
rect 11525 351365 11555 351395
rect 11555 351365 11556 351395
rect 11524 351364 11556 351365
rect 11524 351284 11556 351316
rect 11524 351235 11556 351236
rect 11524 351205 11525 351235
rect 11525 351205 11555 351235
rect 11555 351205 11556 351235
rect 11524 351204 11556 351205
rect 11604 351395 11636 351396
rect 11604 351365 11605 351395
rect 11605 351365 11635 351395
rect 11635 351365 11636 351395
rect 11604 351364 11636 351365
rect 11604 351284 11636 351316
rect 11604 351235 11636 351236
rect 11604 351205 11605 351235
rect 11605 351205 11635 351235
rect 11635 351205 11636 351235
rect 11604 351204 11636 351205
rect 11684 351395 11716 351396
rect 11684 351365 11685 351395
rect 11685 351365 11715 351395
rect 11715 351365 11716 351395
rect 11684 351364 11716 351365
rect 11684 351284 11716 351316
rect 11684 351235 11716 351236
rect 11684 351205 11685 351235
rect 11685 351205 11715 351235
rect 11715 351205 11716 351235
rect 11684 351204 11716 351205
rect 11764 351395 11796 351396
rect 11764 351365 11765 351395
rect 11765 351365 11795 351395
rect 11795 351365 11796 351395
rect 11764 351364 11796 351365
rect 11764 351284 11796 351316
rect 11764 351235 11796 351236
rect 11764 351205 11765 351235
rect 11765 351205 11795 351235
rect 11795 351205 11796 351235
rect 11764 351204 11796 351205
rect 11844 351395 11876 351396
rect 11844 351365 11845 351395
rect 11845 351365 11875 351395
rect 11875 351365 11876 351395
rect 11844 351364 11876 351365
rect 11844 351284 11876 351316
rect 11844 351235 11876 351236
rect 11844 351205 11845 351235
rect 11845 351205 11875 351235
rect 11875 351205 11876 351235
rect 11844 351204 11876 351205
rect 11924 351395 11956 351396
rect 11924 351365 11925 351395
rect 11925 351365 11955 351395
rect 11955 351365 11956 351395
rect 11924 351364 11956 351365
rect 11924 351284 11956 351316
rect 11924 351235 11956 351236
rect 11924 351205 11925 351235
rect 11925 351205 11955 351235
rect 11955 351205 11956 351235
rect 11924 351204 11956 351205
rect 12004 351395 12036 351396
rect 12004 351365 12005 351395
rect 12005 351365 12035 351395
rect 12035 351365 12036 351395
rect 12004 351364 12036 351365
rect 12004 351284 12036 351316
rect 12004 351235 12036 351236
rect 12004 351205 12005 351235
rect 12005 351205 12035 351235
rect 12035 351205 12036 351235
rect 12004 351204 12036 351205
rect 12084 351395 12116 351396
rect 12084 351365 12085 351395
rect 12085 351365 12115 351395
rect 12115 351365 12116 351395
rect 12084 351364 12116 351365
rect 12084 351284 12116 351316
rect 12084 351235 12116 351236
rect 12084 351205 12085 351235
rect 12085 351205 12115 351235
rect 12115 351205 12116 351235
rect 12084 351204 12116 351205
rect 12164 351395 12196 351396
rect 12164 351365 12165 351395
rect 12165 351365 12195 351395
rect 12195 351365 12196 351395
rect 12164 351364 12196 351365
rect 12164 351284 12196 351316
rect 12164 351235 12196 351236
rect 12164 351205 12165 351235
rect 12165 351205 12195 351235
rect 12195 351205 12196 351235
rect 12164 351204 12196 351205
rect 12244 351395 12276 351396
rect 12244 351365 12245 351395
rect 12245 351365 12275 351395
rect 12275 351365 12276 351395
rect 12244 351364 12276 351365
rect 12244 351284 12276 351316
rect 12244 351235 12276 351236
rect 12244 351205 12245 351235
rect 12245 351205 12275 351235
rect 12275 351205 12276 351235
rect 12244 351204 12276 351205
rect 12324 351395 12356 351396
rect 12324 351365 12325 351395
rect 12325 351365 12355 351395
rect 12355 351365 12356 351395
rect 12324 351364 12356 351365
rect 12324 351284 12356 351316
rect 12324 351235 12356 351236
rect 12324 351205 12325 351235
rect 12325 351205 12355 351235
rect 12355 351205 12356 351235
rect 12324 351204 12356 351205
rect 12404 351395 12436 351396
rect 12404 351365 12405 351395
rect 12405 351365 12435 351395
rect 12435 351365 12436 351395
rect 12404 351364 12436 351365
rect 12404 351284 12436 351316
rect 12404 351235 12436 351236
rect 12404 351205 12405 351235
rect 12405 351205 12435 351235
rect 12435 351205 12436 351235
rect 12404 351204 12436 351205
rect 12484 351395 12516 351396
rect 12484 351365 12485 351395
rect 12485 351365 12515 351395
rect 12515 351365 12516 351395
rect 12484 351364 12516 351365
rect 12484 351284 12516 351316
rect 12484 351235 12516 351236
rect 12484 351205 12485 351235
rect 12485 351205 12515 351235
rect 12515 351205 12516 351235
rect 12484 351204 12516 351205
rect 12564 351395 12596 351396
rect 12564 351365 12565 351395
rect 12565 351365 12595 351395
rect 12595 351365 12596 351395
rect 12564 351364 12596 351365
rect 12564 351284 12596 351316
rect 12564 351235 12596 351236
rect 12564 351205 12565 351235
rect 12565 351205 12595 351235
rect 12595 351205 12596 351235
rect 12564 351204 12596 351205
rect 12644 351395 12676 351396
rect 12644 351365 12645 351395
rect 12645 351365 12675 351395
rect 12675 351365 12676 351395
rect 12644 351364 12676 351365
rect 12644 351284 12676 351316
rect 12644 351235 12676 351236
rect 12644 351205 12645 351235
rect 12645 351205 12675 351235
rect 12675 351205 12676 351235
rect 12644 351204 12676 351205
rect 12724 351395 12756 351396
rect 12724 351365 12725 351395
rect 12725 351365 12755 351395
rect 12755 351365 12756 351395
rect 12724 351364 12756 351365
rect 12724 351284 12756 351316
rect 12724 351235 12756 351236
rect 12724 351205 12725 351235
rect 12725 351205 12755 351235
rect 12755 351205 12756 351235
rect 12724 351204 12756 351205
rect 12804 351395 12836 351396
rect 12804 351365 12805 351395
rect 12805 351365 12835 351395
rect 12835 351365 12836 351395
rect 12804 351364 12836 351365
rect 12804 351284 12836 351316
rect 12804 351235 12836 351236
rect 12804 351205 12805 351235
rect 12805 351205 12835 351235
rect 12835 351205 12836 351235
rect 12804 351204 12836 351205
rect 12884 351395 12916 351396
rect 12884 351365 12885 351395
rect 12885 351365 12915 351395
rect 12915 351365 12916 351395
rect 12884 351364 12916 351365
rect 12884 351284 12916 351316
rect 12884 351235 12916 351236
rect 12884 351205 12885 351235
rect 12885 351205 12915 351235
rect 12915 351205 12916 351235
rect 12884 351204 12916 351205
rect 12964 351395 12996 351396
rect 12964 351365 12965 351395
rect 12965 351365 12995 351395
rect 12995 351365 12996 351395
rect 12964 351364 12996 351365
rect 12964 351284 12996 351316
rect 12964 351235 12996 351236
rect 12964 351205 12965 351235
rect 12965 351205 12995 351235
rect 12995 351205 12996 351235
rect 12964 351204 12996 351205
rect 13044 351395 13076 351396
rect 13044 351365 13045 351395
rect 13045 351365 13075 351395
rect 13075 351365 13076 351395
rect 13044 351364 13076 351365
rect 13044 351284 13076 351316
rect 13044 351235 13076 351236
rect 13044 351205 13045 351235
rect 13045 351205 13075 351235
rect 13075 351205 13076 351235
rect 13044 351204 13076 351205
rect 13124 351395 13156 351396
rect 13124 351365 13125 351395
rect 13125 351365 13155 351395
rect 13155 351365 13156 351395
rect 13124 351364 13156 351365
rect 13124 351284 13156 351316
rect 13124 351235 13156 351236
rect 13124 351205 13125 351235
rect 13125 351205 13155 351235
rect 13155 351205 13156 351235
rect 13124 351204 13156 351205
rect 13204 351395 13236 351396
rect 13204 351365 13205 351395
rect 13205 351365 13235 351395
rect 13235 351365 13236 351395
rect 13204 351364 13236 351365
rect 13204 351284 13236 351316
rect 13204 351235 13236 351236
rect 13204 351205 13205 351235
rect 13205 351205 13235 351235
rect 13235 351205 13236 351235
rect 13204 351204 13236 351205
rect 13284 351395 13316 351396
rect 13284 351365 13285 351395
rect 13285 351365 13315 351395
rect 13315 351365 13316 351395
rect 13284 351364 13316 351365
rect 13284 351284 13316 351316
rect 13284 351235 13316 351236
rect 13284 351205 13285 351235
rect 13285 351205 13315 351235
rect 13315 351205 13316 351235
rect 13284 351204 13316 351205
rect 13364 351395 13396 351396
rect 13364 351365 13365 351395
rect 13365 351365 13395 351395
rect 13395 351365 13396 351395
rect 13364 351364 13396 351365
rect 13364 351284 13396 351316
rect 13364 351235 13396 351236
rect 13364 351205 13365 351235
rect 13365 351205 13395 351235
rect 13395 351205 13396 351235
rect 13364 351204 13396 351205
rect 13444 351395 13476 351396
rect 13444 351365 13445 351395
rect 13445 351365 13475 351395
rect 13475 351365 13476 351395
rect 13444 351364 13476 351365
rect 13444 351284 13476 351316
rect 13444 351235 13476 351236
rect 13444 351205 13445 351235
rect 13445 351205 13475 351235
rect 13475 351205 13476 351235
rect 13444 351204 13476 351205
rect 13524 351395 13556 351396
rect 13524 351365 13525 351395
rect 13525 351365 13555 351395
rect 13555 351365 13556 351395
rect 13524 351364 13556 351365
rect 13524 351284 13556 351316
rect 13524 351235 13556 351236
rect 13524 351205 13525 351235
rect 13525 351205 13555 351235
rect 13555 351205 13556 351235
rect 13524 351204 13556 351205
rect 13604 351395 13636 351396
rect 13604 351365 13605 351395
rect 13605 351365 13635 351395
rect 13635 351365 13636 351395
rect 13604 351364 13636 351365
rect 13604 351284 13636 351316
rect 13604 351235 13636 351236
rect 13604 351205 13605 351235
rect 13605 351205 13635 351235
rect 13635 351205 13636 351235
rect 13604 351204 13636 351205
rect 13684 351395 13716 351396
rect 13684 351365 13685 351395
rect 13685 351365 13715 351395
rect 13715 351365 13716 351395
rect 13684 351364 13716 351365
rect 13684 351284 13716 351316
rect 13684 351235 13716 351236
rect 13684 351205 13685 351235
rect 13685 351205 13715 351235
rect 13715 351205 13716 351235
rect 13684 351204 13716 351205
rect 13764 351395 13796 351396
rect 13764 351365 13765 351395
rect 13765 351365 13795 351395
rect 13795 351365 13796 351395
rect 13764 351364 13796 351365
rect 13764 351284 13796 351316
rect 13764 351235 13796 351236
rect 13764 351205 13765 351235
rect 13765 351205 13795 351235
rect 13795 351205 13796 351235
rect 13764 351204 13796 351205
rect 13844 351395 13876 351396
rect 13844 351365 13845 351395
rect 13845 351365 13875 351395
rect 13875 351365 13876 351395
rect 13844 351364 13876 351365
rect 13844 351284 13876 351316
rect 13844 351235 13876 351236
rect 13844 351205 13845 351235
rect 13845 351205 13875 351235
rect 13875 351205 13876 351235
rect 13844 351204 13876 351205
rect 13924 351395 13956 351396
rect 13924 351365 13925 351395
rect 13925 351365 13955 351395
rect 13955 351365 13956 351395
rect 13924 351364 13956 351365
rect 13924 351284 13956 351316
rect 13924 351235 13956 351236
rect 13924 351205 13925 351235
rect 13925 351205 13955 351235
rect 13955 351205 13956 351235
rect 13924 351204 13956 351205
rect 14004 351395 14036 351396
rect 14004 351365 14005 351395
rect 14005 351365 14035 351395
rect 14035 351365 14036 351395
rect 14004 351364 14036 351365
rect 14004 351284 14036 351316
rect 14004 351235 14036 351236
rect 14004 351205 14005 351235
rect 14005 351205 14035 351235
rect 14035 351205 14036 351235
rect 14004 351204 14036 351205
rect 14084 351395 14116 351396
rect 14084 351365 14085 351395
rect 14085 351365 14115 351395
rect 14115 351365 14116 351395
rect 14084 351364 14116 351365
rect 14084 351284 14116 351316
rect 14084 351235 14116 351236
rect 14084 351205 14085 351235
rect 14085 351205 14115 351235
rect 14115 351205 14116 351235
rect 14084 351204 14116 351205
rect 14164 351395 14196 351396
rect 14164 351365 14165 351395
rect 14165 351365 14195 351395
rect 14195 351365 14196 351395
rect 14164 351364 14196 351365
rect 14164 351284 14196 351316
rect 14164 351235 14196 351236
rect 14164 351205 14165 351235
rect 14165 351205 14195 351235
rect 14195 351205 14196 351235
rect 14164 351204 14196 351205
rect 14244 351395 14276 351396
rect 14244 351365 14245 351395
rect 14245 351365 14275 351395
rect 14275 351365 14276 351395
rect 14244 351364 14276 351365
rect 14244 351284 14276 351316
rect 14244 351235 14276 351236
rect 14244 351205 14245 351235
rect 14245 351205 14275 351235
rect 14275 351205 14276 351235
rect 14244 351204 14276 351205
rect 14324 351395 14356 351396
rect 14324 351365 14325 351395
rect 14325 351365 14355 351395
rect 14355 351365 14356 351395
rect 14324 351364 14356 351365
rect 14324 351284 14356 351316
rect 14324 351235 14356 351236
rect 14324 351205 14325 351235
rect 14325 351205 14355 351235
rect 14355 351205 14356 351235
rect 14324 351204 14356 351205
rect 14404 351395 14436 351396
rect 14404 351365 14405 351395
rect 14405 351365 14435 351395
rect 14435 351365 14436 351395
rect 14404 351364 14436 351365
rect 14404 351284 14436 351316
rect 14404 351235 14436 351236
rect 14404 351205 14405 351235
rect 14405 351205 14435 351235
rect 14435 351205 14436 351235
rect 14404 351204 14436 351205
rect 14484 351395 14516 351396
rect 14484 351365 14485 351395
rect 14485 351365 14515 351395
rect 14515 351365 14516 351395
rect 14484 351364 14516 351365
rect 14484 351284 14516 351316
rect 14484 351235 14516 351236
rect 14484 351205 14485 351235
rect 14485 351205 14515 351235
rect 14515 351205 14516 351235
rect 14484 351204 14516 351205
rect 14564 351395 14596 351396
rect 14564 351365 14565 351395
rect 14565 351365 14595 351395
rect 14595 351365 14596 351395
rect 14564 351364 14596 351365
rect 14564 351284 14596 351316
rect 14564 351235 14596 351236
rect 14564 351205 14565 351235
rect 14565 351205 14595 351235
rect 14595 351205 14596 351235
rect 14564 351204 14596 351205
rect 14644 351395 14676 351396
rect 14644 351365 14645 351395
rect 14645 351365 14675 351395
rect 14675 351365 14676 351395
rect 14644 351364 14676 351365
rect 14644 351284 14676 351316
rect 14644 351235 14676 351236
rect 14644 351205 14645 351235
rect 14645 351205 14675 351235
rect 14675 351205 14676 351235
rect 14644 351204 14676 351205
rect 14724 351395 14756 351396
rect 14724 351365 14725 351395
rect 14725 351365 14755 351395
rect 14755 351365 14756 351395
rect 14724 351364 14756 351365
rect 14724 351284 14756 351316
rect 14724 351235 14756 351236
rect 14724 351205 14725 351235
rect 14725 351205 14755 351235
rect 14755 351205 14756 351235
rect 14724 351204 14756 351205
rect 14804 351395 14836 351396
rect 14804 351365 14805 351395
rect 14805 351365 14835 351395
rect 14835 351365 14836 351395
rect 14804 351364 14836 351365
rect 14804 351284 14836 351316
rect 14804 351235 14836 351236
rect 14804 351205 14805 351235
rect 14805 351205 14835 351235
rect 14835 351205 14836 351235
rect 14804 351204 14836 351205
rect 14884 351395 14916 351396
rect 14884 351365 14885 351395
rect 14885 351365 14915 351395
rect 14915 351365 14916 351395
rect 14884 351364 14916 351365
rect 14884 351284 14916 351316
rect 14884 351235 14916 351236
rect 14884 351205 14885 351235
rect 14885 351205 14915 351235
rect 14915 351205 14916 351235
rect 14884 351204 14916 351205
rect 14964 351395 14996 351396
rect 14964 351365 14965 351395
rect 14965 351365 14995 351395
rect 14995 351365 14996 351395
rect 14964 351364 14996 351365
rect 14964 351284 14996 351316
rect 14964 351235 14996 351236
rect 14964 351205 14965 351235
rect 14965 351205 14995 351235
rect 14995 351205 14996 351235
rect 14964 351204 14996 351205
rect 15044 351395 15076 351396
rect 15044 351365 15045 351395
rect 15045 351365 15075 351395
rect 15075 351365 15076 351395
rect 15044 351364 15076 351365
rect 15044 351284 15076 351316
rect 15044 351235 15076 351236
rect 15044 351205 15045 351235
rect 15045 351205 15075 351235
rect 15075 351205 15076 351235
rect 15044 351204 15076 351205
rect 15124 351395 15156 351396
rect 15124 351365 15125 351395
rect 15125 351365 15155 351395
rect 15155 351365 15156 351395
rect 15124 351364 15156 351365
rect 15124 351284 15156 351316
rect 15124 351235 15156 351236
rect 15124 351205 15125 351235
rect 15125 351205 15155 351235
rect 15155 351205 15156 351235
rect 15124 351204 15156 351205
rect 15204 351395 15236 351396
rect 15204 351365 15205 351395
rect 15205 351365 15235 351395
rect 15235 351365 15236 351395
rect 15204 351364 15236 351365
rect 15204 351284 15236 351316
rect 15204 351235 15236 351236
rect 15204 351205 15205 351235
rect 15205 351205 15235 351235
rect 15235 351205 15236 351235
rect 15204 351204 15236 351205
rect 15284 351395 15316 351396
rect 15284 351365 15285 351395
rect 15285 351365 15315 351395
rect 15315 351365 15316 351395
rect 15284 351364 15316 351365
rect 15284 351284 15316 351316
rect 15284 351235 15316 351236
rect 15284 351205 15285 351235
rect 15285 351205 15315 351235
rect 15315 351205 15316 351235
rect 15284 351204 15316 351205
rect 15364 351395 15396 351396
rect 15364 351365 15365 351395
rect 15365 351365 15395 351395
rect 15395 351365 15396 351395
rect 15364 351364 15396 351365
rect 15364 351284 15396 351316
rect 15364 351235 15396 351236
rect 15364 351205 15365 351235
rect 15365 351205 15395 351235
rect 15395 351205 15396 351235
rect 15364 351204 15396 351205
rect 15444 351395 15476 351396
rect 15444 351365 15445 351395
rect 15445 351365 15475 351395
rect 15475 351365 15476 351395
rect 15444 351364 15476 351365
rect 15444 351284 15476 351316
rect 15444 351235 15476 351236
rect 15444 351205 15445 351235
rect 15445 351205 15475 351235
rect 15475 351205 15476 351235
rect 15444 351204 15476 351205
rect 15524 351395 15556 351396
rect 15524 351365 15525 351395
rect 15525 351365 15555 351395
rect 15555 351365 15556 351395
rect 15524 351364 15556 351365
rect 15524 351284 15556 351316
rect 15524 351235 15556 351236
rect 15524 351205 15525 351235
rect 15525 351205 15555 351235
rect 15555 351205 15556 351235
rect 15524 351204 15556 351205
rect 15604 351395 15636 351396
rect 15604 351365 15605 351395
rect 15605 351365 15635 351395
rect 15635 351365 15636 351395
rect 15604 351364 15636 351365
rect 15604 351284 15636 351316
rect 15604 351235 15636 351236
rect 15604 351205 15605 351235
rect 15605 351205 15635 351235
rect 15635 351205 15636 351235
rect 15604 351204 15636 351205
rect 15684 351395 15716 351396
rect 15684 351365 15685 351395
rect 15685 351365 15715 351395
rect 15715 351365 15716 351395
rect 15684 351364 15716 351365
rect 15684 351284 15716 351316
rect 15684 351235 15716 351236
rect 15684 351205 15685 351235
rect 15685 351205 15715 351235
rect 15715 351205 15716 351235
rect 15684 351204 15716 351205
rect 15764 351395 15796 351396
rect 15764 351365 15765 351395
rect 15765 351365 15795 351395
rect 15795 351365 15796 351395
rect 15764 351364 15796 351365
rect 15764 351284 15796 351316
rect 15764 351235 15796 351236
rect 15764 351205 15765 351235
rect 15765 351205 15795 351235
rect 15795 351205 15796 351235
rect 15764 351204 15796 351205
rect 15844 351395 15876 351396
rect 15844 351365 15845 351395
rect 15845 351365 15875 351395
rect 15875 351365 15876 351395
rect 15844 351364 15876 351365
rect 15844 351284 15876 351316
rect 15844 351235 15876 351236
rect 15844 351205 15845 351235
rect 15845 351205 15875 351235
rect 15875 351205 15876 351235
rect 15844 351204 15876 351205
rect 15924 351395 15956 351396
rect 15924 351365 15925 351395
rect 15925 351365 15955 351395
rect 15955 351365 15956 351395
rect 15924 351364 15956 351365
rect 15924 351284 15956 351316
rect 15924 351235 15956 351236
rect 15924 351205 15925 351235
rect 15925 351205 15955 351235
rect 15955 351205 15956 351235
rect 15924 351204 15956 351205
rect 16004 351395 16036 351396
rect 16004 351365 16005 351395
rect 16005 351365 16035 351395
rect 16035 351365 16036 351395
rect 16004 351364 16036 351365
rect 16004 351284 16036 351316
rect 16004 351235 16036 351236
rect 16004 351205 16005 351235
rect 16005 351205 16035 351235
rect 16035 351205 16036 351235
rect 16004 351204 16036 351205
rect 16084 351395 16116 351396
rect 16084 351365 16085 351395
rect 16085 351365 16115 351395
rect 16115 351365 16116 351395
rect 16084 351364 16116 351365
rect 16084 351284 16116 351316
rect 16084 351235 16116 351236
rect 16084 351205 16085 351235
rect 16085 351205 16115 351235
rect 16115 351205 16116 351235
rect 16084 351204 16116 351205
rect 16164 351395 16196 351396
rect 16164 351365 16165 351395
rect 16165 351365 16195 351395
rect 16195 351365 16196 351395
rect 16164 351364 16196 351365
rect 16164 351284 16196 351316
rect 16164 351235 16196 351236
rect 16164 351205 16165 351235
rect 16165 351205 16195 351235
rect 16195 351205 16196 351235
rect 16164 351204 16196 351205
rect 16244 351395 16276 351396
rect 16244 351365 16245 351395
rect 16245 351365 16275 351395
rect 16275 351365 16276 351395
rect 16244 351364 16276 351365
rect 16244 351284 16276 351316
rect 16244 351235 16276 351236
rect 16244 351205 16245 351235
rect 16245 351205 16275 351235
rect 16275 351205 16276 351235
rect 16244 351204 16276 351205
rect 16324 351395 16356 351396
rect 16324 351365 16325 351395
rect 16325 351365 16355 351395
rect 16355 351365 16356 351395
rect 16324 351364 16356 351365
rect 16324 351284 16356 351316
rect 16324 351235 16356 351236
rect 16324 351205 16325 351235
rect 16325 351205 16355 351235
rect 16355 351205 16356 351235
rect 16324 351204 16356 351205
rect 16404 351395 16436 351396
rect 16404 351365 16405 351395
rect 16405 351365 16435 351395
rect 16435 351365 16436 351395
rect 16404 351364 16436 351365
rect 16404 351284 16436 351316
rect 16404 351235 16436 351236
rect 16404 351205 16405 351235
rect 16405 351205 16435 351235
rect 16435 351205 16436 351235
rect 16404 351204 16436 351205
rect 16484 351395 16516 351396
rect 16484 351365 16485 351395
rect 16485 351365 16515 351395
rect 16515 351365 16516 351395
rect 16484 351364 16516 351365
rect 16484 351284 16516 351316
rect 16484 351235 16516 351236
rect 16484 351205 16485 351235
rect 16485 351205 16515 351235
rect 16515 351205 16516 351235
rect 16484 351204 16516 351205
rect 16564 351395 16596 351396
rect 16564 351365 16565 351395
rect 16565 351365 16595 351395
rect 16595 351365 16596 351395
rect 16564 351364 16596 351365
rect 16564 351284 16596 351316
rect 16564 351235 16596 351236
rect 16564 351205 16565 351235
rect 16565 351205 16595 351235
rect 16595 351205 16596 351235
rect 16564 351204 16596 351205
rect 16644 351395 16676 351396
rect 16644 351365 16645 351395
rect 16645 351365 16675 351395
rect 16675 351365 16676 351395
rect 16644 351364 16676 351365
rect 16644 351284 16676 351316
rect 16644 351235 16676 351236
rect 16644 351205 16645 351235
rect 16645 351205 16675 351235
rect 16675 351205 16676 351235
rect 16644 351204 16676 351205
rect 16724 351395 16756 351396
rect 16724 351365 16725 351395
rect 16725 351365 16755 351395
rect 16755 351365 16756 351395
rect 16724 351364 16756 351365
rect 16724 351284 16756 351316
rect 16724 351235 16756 351236
rect 16724 351205 16725 351235
rect 16725 351205 16755 351235
rect 16755 351205 16756 351235
rect 16724 351204 16756 351205
rect 16804 351395 16836 351396
rect 16804 351365 16805 351395
rect 16805 351365 16835 351395
rect 16835 351365 16836 351395
rect 16804 351364 16836 351365
rect 16804 351284 16836 351316
rect 16804 351235 16836 351236
rect 16804 351205 16805 351235
rect 16805 351205 16835 351235
rect 16835 351205 16836 351235
rect 16804 351204 16836 351205
rect 16884 351395 16916 351396
rect 16884 351365 16885 351395
rect 16885 351365 16915 351395
rect 16915 351365 16916 351395
rect 16884 351364 16916 351365
rect 16884 351284 16916 351316
rect 16884 351235 16916 351236
rect 16884 351205 16885 351235
rect 16885 351205 16915 351235
rect 16915 351205 16916 351235
rect 16884 351204 16916 351205
rect 16964 351395 16996 351396
rect 16964 351365 16965 351395
rect 16965 351365 16995 351395
rect 16995 351365 16996 351395
rect 16964 351364 16996 351365
rect 16964 351284 16996 351316
rect 16964 351235 16996 351236
rect 16964 351205 16965 351235
rect 16965 351205 16995 351235
rect 16995 351205 16996 351235
rect 16964 351204 16996 351205
rect 17044 351395 17076 351396
rect 17044 351365 17045 351395
rect 17045 351365 17075 351395
rect 17075 351365 17076 351395
rect 17044 351364 17076 351365
rect 17044 351284 17076 351316
rect 17044 351235 17076 351236
rect 17044 351205 17045 351235
rect 17045 351205 17075 351235
rect 17075 351205 17076 351235
rect 17044 351204 17076 351205
rect 17124 351395 17156 351396
rect 17124 351365 17125 351395
rect 17125 351365 17155 351395
rect 17155 351365 17156 351395
rect 17124 351364 17156 351365
rect 17124 351284 17156 351316
rect 17124 351235 17156 351236
rect 17124 351205 17125 351235
rect 17125 351205 17155 351235
rect 17155 351205 17156 351235
rect 17124 351204 17156 351205
rect 17204 351395 17236 351396
rect 17204 351365 17205 351395
rect 17205 351365 17235 351395
rect 17235 351365 17236 351395
rect 17204 351364 17236 351365
rect 17204 351284 17236 351316
rect 17204 351235 17236 351236
rect 17204 351205 17205 351235
rect 17205 351205 17235 351235
rect 17235 351205 17236 351235
rect 17204 351204 17236 351205
rect 17284 351395 17316 351396
rect 17284 351365 17285 351395
rect 17285 351365 17315 351395
rect 17315 351365 17316 351395
rect 17284 351364 17316 351365
rect 17284 351284 17316 351316
rect 17284 351235 17316 351236
rect 17284 351205 17285 351235
rect 17285 351205 17315 351235
rect 17315 351205 17316 351235
rect 17284 351204 17316 351205
rect 17364 351395 17396 351396
rect 17364 351365 17365 351395
rect 17365 351365 17395 351395
rect 17395 351365 17396 351395
rect 17364 351364 17396 351365
rect 17364 351284 17396 351316
rect 17364 351235 17396 351236
rect 17364 351205 17365 351235
rect 17365 351205 17395 351235
rect 17395 351205 17396 351235
rect 17364 351204 17396 351205
rect 17444 351395 17476 351396
rect 17444 351365 17445 351395
rect 17445 351365 17475 351395
rect 17475 351365 17476 351395
rect 17444 351364 17476 351365
rect 17444 351284 17476 351316
rect 17444 351235 17476 351236
rect 17444 351205 17445 351235
rect 17445 351205 17475 351235
rect 17475 351205 17476 351235
rect 17444 351204 17476 351205
rect 17524 351395 17556 351396
rect 17524 351365 17525 351395
rect 17525 351365 17555 351395
rect 17555 351365 17556 351395
rect 17524 351364 17556 351365
rect 17524 351284 17556 351316
rect 17524 351235 17556 351236
rect 17524 351205 17525 351235
rect 17525 351205 17555 351235
rect 17555 351205 17556 351235
rect 17524 351204 17556 351205
rect 17604 351395 17636 351396
rect 17604 351365 17605 351395
rect 17605 351365 17635 351395
rect 17635 351365 17636 351395
rect 17604 351364 17636 351365
rect 17604 351284 17636 351316
rect 17604 351235 17636 351236
rect 17604 351205 17605 351235
rect 17605 351205 17635 351235
rect 17635 351205 17636 351235
rect 17604 351204 17636 351205
rect 17684 351395 17716 351396
rect 17684 351365 17685 351395
rect 17685 351365 17715 351395
rect 17715 351365 17716 351395
rect 17684 351364 17716 351365
rect 17684 351284 17716 351316
rect 17684 351235 17716 351236
rect 17684 351205 17685 351235
rect 17685 351205 17715 351235
rect 17715 351205 17716 351235
rect 17684 351204 17716 351205
rect 17764 351395 17796 351396
rect 17764 351365 17765 351395
rect 17765 351365 17795 351395
rect 17795 351365 17796 351395
rect 17764 351364 17796 351365
rect 17764 351284 17796 351316
rect 17764 351235 17796 351236
rect 17764 351205 17765 351235
rect 17765 351205 17795 351235
rect 17795 351205 17796 351235
rect 17764 351204 17796 351205
rect 17844 351395 17876 351396
rect 17844 351365 17845 351395
rect 17845 351365 17875 351395
rect 17875 351365 17876 351395
rect 17844 351364 17876 351365
rect 17844 351284 17876 351316
rect 17844 351235 17876 351236
rect 17844 351205 17845 351235
rect 17845 351205 17875 351235
rect 17875 351205 17876 351235
rect 17844 351204 17876 351205
rect 17924 351395 17956 351396
rect 17924 351365 17925 351395
rect 17925 351365 17955 351395
rect 17955 351365 17956 351395
rect 17924 351364 17956 351365
rect 17924 351284 17956 351316
rect 17924 351235 17956 351236
rect 17924 351205 17925 351235
rect 17925 351205 17955 351235
rect 17955 351205 17956 351235
rect 17924 351204 17956 351205
rect 18004 351395 18036 351396
rect 18004 351365 18005 351395
rect 18005 351365 18035 351395
rect 18035 351365 18036 351395
rect 18004 351364 18036 351365
rect 18004 351284 18036 351316
rect 18004 351235 18036 351236
rect 18004 351205 18005 351235
rect 18005 351205 18035 351235
rect 18035 351205 18036 351235
rect 18004 351204 18036 351205
rect 18084 351395 18116 351396
rect 18084 351365 18085 351395
rect 18085 351365 18115 351395
rect 18115 351365 18116 351395
rect 18084 351364 18116 351365
rect 18084 351284 18116 351316
rect 18084 351235 18116 351236
rect 18084 351205 18085 351235
rect 18085 351205 18115 351235
rect 18115 351205 18116 351235
rect 18084 351204 18116 351205
rect 18164 351395 18196 351396
rect 18164 351365 18165 351395
rect 18165 351365 18195 351395
rect 18195 351365 18196 351395
rect 18164 351364 18196 351365
rect 18164 351284 18196 351316
rect 18164 351235 18196 351236
rect 18164 351205 18165 351235
rect 18165 351205 18195 351235
rect 18195 351205 18196 351235
rect 18164 351204 18196 351205
rect 18244 351395 18276 351396
rect 18244 351365 18245 351395
rect 18245 351365 18275 351395
rect 18275 351365 18276 351395
rect 18244 351364 18276 351365
rect 18244 351284 18276 351316
rect 18244 351235 18276 351236
rect 18244 351205 18245 351235
rect 18245 351205 18275 351235
rect 18275 351205 18276 351235
rect 18244 351204 18276 351205
rect 18324 351395 18356 351396
rect 18324 351365 18325 351395
rect 18325 351365 18355 351395
rect 18355 351365 18356 351395
rect 18324 351364 18356 351365
rect 18324 351284 18356 351316
rect 18324 351235 18356 351236
rect 18324 351205 18325 351235
rect 18325 351205 18355 351235
rect 18355 351205 18356 351235
rect 18324 351204 18356 351205
rect 18404 351395 18436 351396
rect 18404 351365 18405 351395
rect 18405 351365 18435 351395
rect 18435 351365 18436 351395
rect 18404 351364 18436 351365
rect 18404 351284 18436 351316
rect 18404 351235 18436 351236
rect 18404 351205 18405 351235
rect 18405 351205 18435 351235
rect 18435 351205 18436 351235
rect 18404 351204 18436 351205
rect 18484 351395 18516 351396
rect 18484 351365 18485 351395
rect 18485 351365 18515 351395
rect 18515 351365 18516 351395
rect 18484 351364 18516 351365
rect 18484 351284 18516 351316
rect 18484 351235 18516 351236
rect 18484 351205 18485 351235
rect 18485 351205 18515 351235
rect 18515 351205 18516 351235
rect 18484 351204 18516 351205
rect 18564 351395 18596 351396
rect 18564 351365 18565 351395
rect 18565 351365 18595 351395
rect 18595 351365 18596 351395
rect 18564 351364 18596 351365
rect 18564 351284 18596 351316
rect 18564 351235 18596 351236
rect 18564 351205 18565 351235
rect 18565 351205 18595 351235
rect 18595 351205 18596 351235
rect 18564 351204 18596 351205
rect 18644 351395 18676 351396
rect 18644 351365 18645 351395
rect 18645 351365 18675 351395
rect 18675 351365 18676 351395
rect 18644 351364 18676 351365
rect 18644 351284 18676 351316
rect 18644 351235 18676 351236
rect 18644 351205 18645 351235
rect 18645 351205 18675 351235
rect 18675 351205 18676 351235
rect 18644 351204 18676 351205
rect 18724 351395 18756 351396
rect 18724 351365 18725 351395
rect 18725 351365 18755 351395
rect 18755 351365 18756 351395
rect 18724 351364 18756 351365
rect 18724 351284 18756 351316
rect 18724 351235 18756 351236
rect 18724 351205 18725 351235
rect 18725 351205 18755 351235
rect 18755 351205 18756 351235
rect 18724 351204 18756 351205
rect 18804 351395 18836 351396
rect 18804 351365 18805 351395
rect 18805 351365 18835 351395
rect 18835 351365 18836 351395
rect 18804 351364 18836 351365
rect 18804 351284 18836 351316
rect 18804 351235 18836 351236
rect 18804 351205 18805 351235
rect 18805 351205 18835 351235
rect 18835 351205 18836 351235
rect 18804 351204 18836 351205
rect 18884 351395 18916 351396
rect 18884 351365 18885 351395
rect 18885 351365 18915 351395
rect 18915 351365 18916 351395
rect 18884 351364 18916 351365
rect 18884 351284 18916 351316
rect 18884 351235 18916 351236
rect 18884 351205 18885 351235
rect 18885 351205 18915 351235
rect 18915 351205 18916 351235
rect 18884 351204 18916 351205
rect 18964 351395 18996 351396
rect 18964 351365 18965 351395
rect 18965 351365 18995 351395
rect 18995 351365 18996 351395
rect 18964 351364 18996 351365
rect 18964 351284 18996 351316
rect 18964 351235 18996 351236
rect 18964 351205 18965 351235
rect 18965 351205 18995 351235
rect 18995 351205 18996 351235
rect 18964 351204 18996 351205
rect 19044 351395 19076 351396
rect 19044 351365 19045 351395
rect 19045 351365 19075 351395
rect 19075 351365 19076 351395
rect 19044 351364 19076 351365
rect 19044 351284 19076 351316
rect 19044 351235 19076 351236
rect 19044 351205 19045 351235
rect 19045 351205 19075 351235
rect 19075 351205 19076 351235
rect 19044 351204 19076 351205
rect 19124 351395 19156 351396
rect 19124 351365 19125 351395
rect 19125 351365 19155 351395
rect 19155 351365 19156 351395
rect 19124 351364 19156 351365
rect 19124 351284 19156 351316
rect 19124 351235 19156 351236
rect 19124 351205 19125 351235
rect 19125 351205 19155 351235
rect 19155 351205 19156 351235
rect 19124 351204 19156 351205
rect 19204 351395 19236 351396
rect 19204 351365 19205 351395
rect 19205 351365 19235 351395
rect 19235 351365 19236 351395
rect 19204 351364 19236 351365
rect 19204 351284 19236 351316
rect 19204 351235 19236 351236
rect 19204 351205 19205 351235
rect 19205 351205 19235 351235
rect 19235 351205 19236 351235
rect 19204 351204 19236 351205
rect 19284 351395 19316 351396
rect 19284 351365 19285 351395
rect 19285 351365 19315 351395
rect 19315 351365 19316 351395
rect 19284 351364 19316 351365
rect 19284 351284 19316 351316
rect 19284 351235 19316 351236
rect 19284 351205 19285 351235
rect 19285 351205 19315 351235
rect 19315 351205 19316 351235
rect 19284 351204 19316 351205
rect 19364 351395 19396 351396
rect 19364 351365 19365 351395
rect 19365 351365 19395 351395
rect 19395 351365 19396 351395
rect 19364 351364 19396 351365
rect 19364 351284 19396 351316
rect 19364 351235 19396 351236
rect 19364 351205 19365 351235
rect 19365 351205 19395 351235
rect 19395 351205 19396 351235
rect 19364 351204 19396 351205
rect 19444 351395 19476 351396
rect 19444 351365 19445 351395
rect 19445 351365 19475 351395
rect 19475 351365 19476 351395
rect 19444 351364 19476 351365
rect 19444 351284 19476 351316
rect 19444 351235 19476 351236
rect 19444 351205 19445 351235
rect 19445 351205 19475 351235
rect 19475 351205 19476 351235
rect 19444 351204 19476 351205
rect 19524 351395 19556 351396
rect 19524 351365 19525 351395
rect 19525 351365 19555 351395
rect 19555 351365 19556 351395
rect 19524 351364 19556 351365
rect 19524 351284 19556 351316
rect 19524 351235 19556 351236
rect 19524 351205 19525 351235
rect 19525 351205 19555 351235
rect 19555 351205 19556 351235
rect 19524 351204 19556 351205
rect 19604 351395 19636 351396
rect 19604 351365 19605 351395
rect 19605 351365 19635 351395
rect 19635 351365 19636 351395
rect 19604 351364 19636 351365
rect 19604 351284 19636 351316
rect 19604 351235 19636 351236
rect 19604 351205 19605 351235
rect 19605 351205 19635 351235
rect 19635 351205 19636 351235
rect 19604 351204 19636 351205
rect 19684 351395 19716 351396
rect 19684 351365 19685 351395
rect 19685 351365 19715 351395
rect 19715 351365 19716 351395
rect 19684 351364 19716 351365
rect 19844 351395 19876 351396
rect 19844 351365 19845 351395
rect 19845 351365 19875 351395
rect 19875 351365 19876 351395
rect 19844 351364 19876 351365
rect 19684 351284 19716 351316
rect 19684 351235 19716 351236
rect 19684 351205 19685 351235
rect 19685 351205 19715 351235
rect 19715 351205 19716 351235
rect 19684 351204 19716 351205
rect 19684 351155 19716 351156
rect 19684 351125 19685 351155
rect 19685 351125 19715 351155
rect 19715 351125 19716 351155
rect 19684 351124 19716 351125
rect 19684 351075 19716 351076
rect 19684 351045 19685 351075
rect 19685 351045 19715 351075
rect 19715 351045 19716 351075
rect 19684 351044 19716 351045
rect 19684 350995 19716 350996
rect 19684 350965 19685 350995
rect 19685 350965 19715 350995
rect 19715 350965 19716 350995
rect 19684 350964 19716 350965
rect 19684 350915 19716 350916
rect 19684 350885 19685 350915
rect 19685 350885 19715 350915
rect 19715 350885 19716 350915
rect 19684 350884 19716 350885
rect 19684 350835 19716 350836
rect 19684 350805 19685 350835
rect 19685 350805 19715 350835
rect 19715 350805 19716 350835
rect 19684 350804 19716 350805
rect 19684 350755 19716 350756
rect 19684 350725 19685 350755
rect 19685 350725 19715 350755
rect 19715 350725 19716 350755
rect 19684 350724 19716 350725
rect 19684 350675 19716 350676
rect 19684 350645 19685 350675
rect 19685 350645 19715 350675
rect 19715 350645 19716 350675
rect 19684 350644 19716 350645
rect 19684 350595 19716 350596
rect 19684 350565 19685 350595
rect 19685 350565 19715 350595
rect 19715 350565 19716 350595
rect 19684 350564 19716 350565
rect 19684 350515 19716 350516
rect 19684 350485 19685 350515
rect 19685 350485 19715 350515
rect 19715 350485 19716 350515
rect 19684 350484 19716 350485
rect 19684 350435 19716 350436
rect 19684 350405 19685 350435
rect 19685 350405 19715 350435
rect 19715 350405 19716 350435
rect 19684 350404 19716 350405
rect 19684 350355 19716 350356
rect 19684 350325 19685 350355
rect 19685 350325 19715 350355
rect 19715 350325 19716 350355
rect 19684 350324 19716 350325
rect 19684 350275 19716 350276
rect 19684 350245 19685 350275
rect 19685 350245 19715 350275
rect 19715 350245 19716 350275
rect 19684 350244 19716 350245
rect 19684 350195 19716 350196
rect 19684 350165 19685 350195
rect 19685 350165 19715 350195
rect 19715 350165 19716 350195
rect 19684 350164 19716 350165
rect 19684 350115 19716 350116
rect 19684 350085 19685 350115
rect 19685 350085 19715 350115
rect 19715 350085 19716 350115
rect 19684 350084 19716 350085
rect 19684 350035 19716 350036
rect 19684 350005 19685 350035
rect 19685 350005 19715 350035
rect 19715 350005 19716 350035
rect 19684 350004 19716 350005
rect 19684 349955 19716 349956
rect 19684 349925 19685 349955
rect 19685 349925 19715 349955
rect 19715 349925 19716 349955
rect 19684 349924 19716 349925
rect 19684 349875 19716 349876
rect 19684 349845 19685 349875
rect 19685 349845 19715 349875
rect 19715 349845 19716 349875
rect 19684 349844 19716 349845
rect 19684 349795 19716 349796
rect 19684 349765 19685 349795
rect 19685 349765 19715 349795
rect 19715 349765 19716 349795
rect 19684 349764 19716 349765
rect 19684 349715 19716 349716
rect 19684 349685 19685 349715
rect 19685 349685 19715 349715
rect 19715 349685 19716 349715
rect 19684 349684 19716 349685
rect 19684 349635 19716 349636
rect 19684 349605 19685 349635
rect 19685 349605 19715 349635
rect 19715 349605 19716 349635
rect 19684 349604 19716 349605
rect 19684 349555 19716 349556
rect 19684 349525 19685 349555
rect 19685 349525 19715 349555
rect 19715 349525 19716 349555
rect 19684 349524 19716 349525
rect 19684 349475 19716 349476
rect 19684 349445 19685 349475
rect 19685 349445 19715 349475
rect 19715 349445 19716 349475
rect 19684 349444 19716 349445
rect 19684 349395 19716 349396
rect 19684 349365 19685 349395
rect 19685 349365 19715 349395
rect 19715 349365 19716 349395
rect 19684 349364 19716 349365
rect 19684 349315 19716 349316
rect 19684 349285 19685 349315
rect 19685 349285 19715 349315
rect 19715 349285 19716 349315
rect 19684 349284 19716 349285
rect 19684 349235 19716 349236
rect 19684 349205 19685 349235
rect 19685 349205 19715 349235
rect 19715 349205 19716 349235
rect 19684 349204 19716 349205
rect 19684 349155 19716 349156
rect 19684 349125 19685 349155
rect 19685 349125 19715 349155
rect 19715 349125 19716 349155
rect 19684 349124 19716 349125
rect 19684 349075 19716 349076
rect 19684 349045 19685 349075
rect 19685 349045 19715 349075
rect 19715 349045 19716 349075
rect 19684 349044 19716 349045
rect 19684 348995 19716 348996
rect 19684 348965 19685 348995
rect 19685 348965 19715 348995
rect 19715 348965 19716 348995
rect 19684 348964 19716 348965
rect 19684 348915 19716 348916
rect 19684 348885 19685 348915
rect 19685 348885 19715 348915
rect 19715 348885 19716 348915
rect 19684 348884 19716 348885
rect 19684 348835 19716 348836
rect 19684 348805 19685 348835
rect 19685 348805 19715 348835
rect 19715 348805 19716 348835
rect 19684 348804 19716 348805
rect 19684 348755 19716 348756
rect 19684 348725 19685 348755
rect 19685 348725 19715 348755
rect 19715 348725 19716 348755
rect 19684 348724 19716 348725
rect 19684 348675 19716 348676
rect 19684 348645 19685 348675
rect 19685 348645 19715 348675
rect 19715 348645 19716 348675
rect 19684 348644 19716 348645
rect 19684 348595 19716 348596
rect 19684 348565 19685 348595
rect 19685 348565 19715 348595
rect 19715 348565 19716 348595
rect 19684 348564 19716 348565
rect 19684 348515 19716 348516
rect 19684 348485 19685 348515
rect 19685 348485 19715 348515
rect 19715 348485 19716 348515
rect 19684 348484 19716 348485
rect 19684 348435 19716 348436
rect 19684 348405 19685 348435
rect 19685 348405 19715 348435
rect 19715 348405 19716 348435
rect 19684 348404 19716 348405
rect 19684 348355 19716 348356
rect 19684 348325 19685 348355
rect 19685 348325 19715 348355
rect 19715 348325 19716 348355
rect 19684 348324 19716 348325
rect 19684 348275 19716 348276
rect 19684 348245 19685 348275
rect 19685 348245 19715 348275
rect 19715 348245 19716 348275
rect 19684 348244 19716 348245
rect 19684 348195 19716 348196
rect 19684 348165 19685 348195
rect 19685 348165 19715 348195
rect 19715 348165 19716 348195
rect 19684 348164 19716 348165
rect 19684 348115 19716 348116
rect 19684 348085 19685 348115
rect 19685 348085 19715 348115
rect 19715 348085 19716 348115
rect 19684 348084 19716 348085
rect 19684 348035 19716 348036
rect 19684 348005 19685 348035
rect 19685 348005 19715 348035
rect 19715 348005 19716 348035
rect 19684 348004 19716 348005
rect 19684 347955 19716 347956
rect 19684 347925 19685 347955
rect 19685 347925 19715 347955
rect 19715 347925 19716 347955
rect 19684 347924 19716 347925
rect 19684 347875 19716 347876
rect 19684 347845 19685 347875
rect 19685 347845 19715 347875
rect 19715 347845 19716 347875
rect 19684 347844 19716 347845
rect 19684 347795 19716 347796
rect 19684 347765 19685 347795
rect 19685 347765 19715 347795
rect 19715 347765 19716 347795
rect 19684 347764 19716 347765
rect 19684 347715 19716 347716
rect 19684 347685 19685 347715
rect 19685 347685 19715 347715
rect 19715 347685 19716 347715
rect 19684 347684 19716 347685
rect 19684 347635 19716 347636
rect 19684 347605 19685 347635
rect 19685 347605 19715 347635
rect 19715 347605 19716 347635
rect 19684 347604 19716 347605
rect 19684 347555 19716 347556
rect 19684 347525 19685 347555
rect 19685 347525 19715 347555
rect 19715 347525 19716 347555
rect 19684 347524 19716 347525
rect 19684 347475 19716 347476
rect 19684 347445 19685 347475
rect 19685 347445 19715 347475
rect 19715 347445 19716 347475
rect 19684 347444 19716 347445
rect 19684 347395 19716 347396
rect 19684 347365 19685 347395
rect 19685 347365 19715 347395
rect 19715 347365 19716 347395
rect 19684 347364 19716 347365
rect 19684 347315 19716 347316
rect 19684 347285 19685 347315
rect 19685 347285 19715 347315
rect 19715 347285 19716 347315
rect 19684 347284 19716 347285
rect 19684 347235 19716 347236
rect 19684 347205 19685 347235
rect 19685 347205 19715 347235
rect 19715 347205 19716 347235
rect 19684 347204 19716 347205
rect 19684 347155 19716 347156
rect 19684 347125 19685 347155
rect 19685 347125 19715 347155
rect 19715 347125 19716 347155
rect 19684 347124 19716 347125
rect 19684 347075 19716 347076
rect 19684 347045 19685 347075
rect 19685 347045 19715 347075
rect 19715 347045 19716 347075
rect 19684 347044 19716 347045
rect 19684 346995 19716 346996
rect 19684 346965 19685 346995
rect 19685 346965 19715 346995
rect 19715 346965 19716 346995
rect 19684 346964 19716 346965
rect 19684 346915 19716 346916
rect 19684 346885 19685 346915
rect 19685 346885 19715 346915
rect 19715 346885 19716 346915
rect 19684 346884 19716 346885
rect 19684 346835 19716 346836
rect 19684 346805 19685 346835
rect 19685 346805 19715 346835
rect 19715 346805 19716 346835
rect 19684 346804 19716 346805
rect 19684 346755 19716 346756
rect 19684 346725 19685 346755
rect 19685 346725 19715 346755
rect 19715 346725 19716 346755
rect 19684 346724 19716 346725
rect 19684 346675 19716 346676
rect 19684 346645 19685 346675
rect 19685 346645 19715 346675
rect 19715 346645 19716 346675
rect 19684 346644 19716 346645
rect 19684 346595 19716 346596
rect 19684 346565 19685 346595
rect 19685 346565 19715 346595
rect 19715 346565 19716 346595
rect 19684 346564 19716 346565
rect 19684 346515 19716 346516
rect 19684 346485 19685 346515
rect 19685 346485 19715 346515
rect 19715 346485 19716 346515
rect 19684 346484 19716 346485
rect 19684 346435 19716 346436
rect 19684 346405 19685 346435
rect 19685 346405 19715 346435
rect 19715 346405 19716 346435
rect 19684 346404 19716 346405
rect 19684 346355 19716 346356
rect 19684 346325 19685 346355
rect 19685 346325 19715 346355
rect 19715 346325 19716 346355
rect 19684 346324 19716 346325
rect 19684 346275 19716 346276
rect 19684 346245 19685 346275
rect 19685 346245 19715 346275
rect 19715 346245 19716 346275
rect 19684 346244 19716 346245
rect 19684 346195 19716 346196
rect 19684 346165 19685 346195
rect 19685 346165 19715 346195
rect 19715 346165 19716 346195
rect 19684 346164 19716 346165
rect 19684 346115 19716 346116
rect 19684 346085 19685 346115
rect 19685 346085 19715 346115
rect 19715 346085 19716 346115
rect 19684 346084 19716 346085
rect 19684 346035 19716 346036
rect 19684 346005 19685 346035
rect 19685 346005 19715 346035
rect 19715 346005 19716 346035
rect 19684 346004 19716 346005
rect 19684 345955 19716 345956
rect 19684 345925 19685 345955
rect 19685 345925 19715 345955
rect 19715 345925 19716 345955
rect 19684 345924 19716 345925
rect 19684 345875 19716 345876
rect 19684 345845 19685 345875
rect 19685 345845 19715 345875
rect 19715 345845 19716 345875
rect 19684 345844 19716 345845
rect 19684 345795 19716 345796
rect 19684 345765 19685 345795
rect 19685 345765 19715 345795
rect 19715 345765 19716 345795
rect 19684 345764 19716 345765
rect 19684 345715 19716 345716
rect 19684 345685 19685 345715
rect 19685 345685 19715 345715
rect 19715 345685 19716 345715
rect 19684 345684 19716 345685
rect 19684 345635 19716 345636
rect 19684 345605 19685 345635
rect 19685 345605 19715 345635
rect 19715 345605 19716 345635
rect 19684 345604 19716 345605
rect 19684 345555 19716 345556
rect 19684 345525 19685 345555
rect 19685 345525 19715 345555
rect 19715 345525 19716 345555
rect 19684 345524 19716 345525
rect 19684 345475 19716 345476
rect 19684 345445 19685 345475
rect 19685 345445 19715 345475
rect 19715 345445 19716 345475
rect 19684 345444 19716 345445
rect 19684 345395 19716 345396
rect 19684 345365 19685 345395
rect 19685 345365 19715 345395
rect 19715 345365 19716 345395
rect 19684 345364 19716 345365
rect 19684 345315 19716 345316
rect 19684 345285 19685 345315
rect 19685 345285 19715 345315
rect 19715 345285 19716 345315
rect 19684 345284 19716 345285
rect 19684 345235 19716 345236
rect 19684 345205 19685 345235
rect 19685 345205 19715 345235
rect 19715 345205 19716 345235
rect 19684 345204 19716 345205
rect 19684 345155 19716 345156
rect 19684 345125 19685 345155
rect 19685 345125 19715 345155
rect 19715 345125 19716 345155
rect 19684 345124 19716 345125
rect 19684 345075 19716 345076
rect 19684 345045 19685 345075
rect 19685 345045 19715 345075
rect 19715 345045 19716 345075
rect 19684 345044 19716 345045
rect 19684 344995 19716 344996
rect 19684 344965 19685 344995
rect 19685 344965 19715 344995
rect 19715 344965 19716 344995
rect 19684 344964 19716 344965
rect 19684 344915 19716 344916
rect 19684 344885 19685 344915
rect 19685 344885 19715 344915
rect 19715 344885 19716 344915
rect 19684 344884 19716 344885
rect 19684 344835 19716 344836
rect 19684 344805 19685 344835
rect 19685 344805 19715 344835
rect 19715 344805 19716 344835
rect 19684 344804 19716 344805
rect 19684 344755 19716 344756
rect 19684 344725 19685 344755
rect 19685 344725 19715 344755
rect 19715 344725 19716 344755
rect 19684 344724 19716 344725
rect 19684 344675 19716 344676
rect 19684 344645 19685 344675
rect 19685 344645 19715 344675
rect 19715 344645 19716 344675
rect 19684 344644 19716 344645
rect 19684 344595 19716 344596
rect 19684 344565 19685 344595
rect 19685 344565 19715 344595
rect 19715 344565 19716 344595
rect 19684 344564 19716 344565
rect 19684 344515 19716 344516
rect 19684 344485 19685 344515
rect 19685 344485 19715 344515
rect 19715 344485 19716 344515
rect 19684 344484 19716 344485
rect 19684 344435 19716 344436
rect 19684 344405 19685 344435
rect 19685 344405 19715 344435
rect 19715 344405 19716 344435
rect 19684 344404 19716 344405
rect 19684 344355 19716 344356
rect 19684 344325 19685 344355
rect 19685 344325 19715 344355
rect 19715 344325 19716 344355
rect 19684 344324 19716 344325
rect 19684 344275 19716 344276
rect 19684 344245 19685 344275
rect 19685 344245 19715 344275
rect 19715 344245 19716 344275
rect 19684 344244 19716 344245
rect 19684 344195 19716 344196
rect 19684 344165 19685 344195
rect 19685 344165 19715 344195
rect 19715 344165 19716 344195
rect 19684 344164 19716 344165
rect 19684 344115 19716 344116
rect 19684 344085 19685 344115
rect 19685 344085 19715 344115
rect 19715 344085 19716 344115
rect 19684 344084 19716 344085
rect 19684 344035 19716 344036
rect 19684 344005 19685 344035
rect 19685 344005 19715 344035
rect 19715 344005 19716 344035
rect 19684 344004 19716 344005
rect 19684 343955 19716 343956
rect 19684 343925 19685 343955
rect 19685 343925 19715 343955
rect 19715 343925 19716 343955
rect 19684 343924 19716 343925
rect 19684 343875 19716 343876
rect 19684 343845 19685 343875
rect 19685 343845 19715 343875
rect 19715 343845 19716 343875
rect 19684 343844 19716 343845
rect 19684 343795 19716 343796
rect 19684 343765 19685 343795
rect 19685 343765 19715 343795
rect 19715 343765 19716 343795
rect 19684 343764 19716 343765
rect 19684 343715 19716 343716
rect 19684 343685 19685 343715
rect 19685 343685 19715 343715
rect 19715 343685 19716 343715
rect 19684 343684 19716 343685
rect 19684 343635 19716 343636
rect 19684 343605 19685 343635
rect 19685 343605 19715 343635
rect 19715 343605 19716 343635
rect 19684 343604 19716 343605
rect 19684 343555 19716 343556
rect 19684 343525 19685 343555
rect 19685 343525 19715 343555
rect 19715 343525 19716 343555
rect 19684 343524 19716 343525
rect 19684 343475 19716 343476
rect 19684 343445 19685 343475
rect 19685 343445 19715 343475
rect 19715 343445 19716 343475
rect 19684 343444 19716 343445
rect 19684 343395 19716 343396
rect 19684 343365 19685 343395
rect 19685 343365 19715 343395
rect 19715 343365 19716 343395
rect 19684 343364 19716 343365
rect 19684 343315 19716 343316
rect 19684 343285 19685 343315
rect 19685 343285 19715 343315
rect 19715 343285 19716 343315
rect 19684 343284 19716 343285
rect 19684 343235 19716 343236
rect 19684 343205 19685 343235
rect 19685 343205 19715 343235
rect 19715 343205 19716 343235
rect 19684 343204 19716 343205
rect 19684 343155 19716 343156
rect 19684 343125 19685 343155
rect 19685 343125 19715 343155
rect 19715 343125 19716 343155
rect 19684 343124 19716 343125
rect 19684 343075 19716 343076
rect 19684 343045 19685 343075
rect 19685 343045 19715 343075
rect 19715 343045 19716 343075
rect 19684 343044 19716 343045
rect 19684 342995 19716 342996
rect 19684 342965 19685 342995
rect 19685 342965 19715 342995
rect 19715 342965 19716 342995
rect 19684 342964 19716 342965
rect 19684 342915 19716 342916
rect 19684 342885 19685 342915
rect 19685 342885 19715 342915
rect 19715 342885 19716 342915
rect 19684 342884 19716 342885
rect 19684 342835 19716 342836
rect 19684 342805 19685 342835
rect 19685 342805 19715 342835
rect 19715 342805 19716 342835
rect 19684 342804 19716 342805
rect 19684 342755 19716 342756
rect 19684 342725 19685 342755
rect 19685 342725 19715 342755
rect 19715 342725 19716 342755
rect 19684 342724 19716 342725
rect 19684 342675 19716 342676
rect 19684 342645 19685 342675
rect 19685 342645 19715 342675
rect 19715 342645 19716 342675
rect 19684 342644 19716 342645
rect 19684 342595 19716 342596
rect 19684 342565 19685 342595
rect 19685 342565 19715 342595
rect 19715 342565 19716 342595
rect 19684 342564 19716 342565
rect 19684 342515 19716 342516
rect 19684 342485 19685 342515
rect 19685 342485 19715 342515
rect 19715 342485 19716 342515
rect 19684 342484 19716 342485
rect 19684 342435 19716 342436
rect 19684 342405 19685 342435
rect 19685 342405 19715 342435
rect 19715 342405 19716 342435
rect 19684 342404 19716 342405
rect 19684 342355 19716 342356
rect 19684 342325 19685 342355
rect 19685 342325 19715 342355
rect 19715 342325 19716 342355
rect 19684 342324 19716 342325
rect 19684 342275 19716 342276
rect 19684 342245 19685 342275
rect 19685 342245 19715 342275
rect 19715 342245 19716 342275
rect 19684 342244 19716 342245
rect 19684 342195 19716 342196
rect 19684 342165 19685 342195
rect 19685 342165 19715 342195
rect 19715 342165 19716 342195
rect 19684 342164 19716 342165
rect 19684 342115 19716 342116
rect 19684 342085 19685 342115
rect 19685 342085 19715 342115
rect 19715 342085 19716 342115
rect 19684 342084 19716 342085
rect 19684 342035 19716 342036
rect 19684 342005 19685 342035
rect 19685 342005 19715 342035
rect 19715 342005 19716 342035
rect 19684 342004 19716 342005
rect 19684 341955 19716 341956
rect 19684 341925 19685 341955
rect 19685 341925 19715 341955
rect 19715 341925 19716 341955
rect 19684 341924 19716 341925
rect 19684 341875 19716 341876
rect 19684 341845 19685 341875
rect 19685 341845 19715 341875
rect 19715 341845 19716 341875
rect 19684 341844 19716 341845
rect 19684 341795 19716 341796
rect 19684 341765 19685 341795
rect 19685 341765 19715 341795
rect 19715 341765 19716 341795
rect 19684 341764 19716 341765
rect 19684 341715 19716 341716
rect 19684 341685 19685 341715
rect 19685 341685 19715 341715
rect 19715 341685 19716 341715
rect 19684 341684 19716 341685
rect 19684 341635 19716 341636
rect 19684 341605 19685 341635
rect 19685 341605 19715 341635
rect 19715 341605 19716 341635
rect 19684 341604 19716 341605
rect 19684 341555 19716 341556
rect 19684 341525 19685 341555
rect 19685 341525 19715 341555
rect 19715 341525 19716 341555
rect 19684 341524 19716 341525
rect 19684 341475 19716 341476
rect 19684 341445 19685 341475
rect 19685 341445 19715 341475
rect 19715 341445 19716 341475
rect 19684 341444 19716 341445
rect 19684 341395 19716 341396
rect 19684 341365 19685 341395
rect 19685 341365 19715 341395
rect 19715 341365 19716 341395
rect 19684 341364 19716 341365
rect 19684 341315 19716 341316
rect 19684 341285 19685 341315
rect 19685 341285 19715 341315
rect 19715 341285 19716 341315
rect 19684 341284 19716 341285
rect 19684 341235 19716 341236
rect 19684 341205 19685 341235
rect 19685 341205 19715 341235
rect 19715 341205 19716 341235
rect 19684 341204 19716 341205
rect 19684 341155 19716 341156
rect 19684 341125 19685 341155
rect 19685 341125 19715 341155
rect 19715 341125 19716 341155
rect 19684 341124 19716 341125
rect 19684 341075 19716 341076
rect 19684 341045 19685 341075
rect 19685 341045 19715 341075
rect 19715 341045 19716 341075
rect 19684 341044 19716 341045
rect 19684 340995 19716 340996
rect 19684 340965 19685 340995
rect 19685 340965 19715 340995
rect 19715 340965 19716 340995
rect 19684 340964 19716 340965
rect 19684 340915 19716 340916
rect 19684 340885 19685 340915
rect 19685 340885 19715 340915
rect 19715 340885 19716 340915
rect 19684 340884 19716 340885
rect 19684 340835 19716 340836
rect 19684 340805 19685 340835
rect 19685 340805 19715 340835
rect 19715 340805 19716 340835
rect 19684 340804 19716 340805
rect 19684 340755 19716 340756
rect 19684 340725 19685 340755
rect 19685 340725 19715 340755
rect 19715 340725 19716 340755
rect 19684 340724 19716 340725
rect 19684 340675 19716 340676
rect 19684 340645 19685 340675
rect 19685 340645 19715 340675
rect 19715 340645 19716 340675
rect 19684 340644 19716 340645
rect 19684 340595 19716 340596
rect 19684 340565 19685 340595
rect 19685 340565 19715 340595
rect 19715 340565 19716 340595
rect 19684 340564 19716 340565
rect 19684 340515 19716 340516
rect 19684 340485 19685 340515
rect 19685 340485 19715 340515
rect 19715 340485 19716 340515
rect 19684 340484 19716 340485
rect 19684 340435 19716 340436
rect 19684 340405 19685 340435
rect 19685 340405 19715 340435
rect 19715 340405 19716 340435
rect 19684 340404 19716 340405
rect 19684 340355 19716 340356
rect 19684 340325 19685 340355
rect 19685 340325 19715 340355
rect 19715 340325 19716 340355
rect 19684 340324 19716 340325
rect 19684 340275 19716 340276
rect 19684 340245 19685 340275
rect 19685 340245 19715 340275
rect 19715 340245 19716 340275
rect 19684 340244 19716 340245
rect 19684 340195 19716 340196
rect 19684 340165 19685 340195
rect 19685 340165 19715 340195
rect 19715 340165 19716 340195
rect 19684 340164 19716 340165
rect 19684 340115 19716 340116
rect 19684 340085 19685 340115
rect 19685 340085 19715 340115
rect 19715 340085 19716 340115
rect 19684 340084 19716 340085
rect 19684 340035 19716 340036
rect 19684 340005 19685 340035
rect 19685 340005 19715 340035
rect 19715 340005 19716 340035
rect 19684 340004 19716 340005
rect 19684 339955 19716 339956
rect 19684 339925 19685 339955
rect 19685 339925 19715 339955
rect 19715 339925 19716 339955
rect 19684 339924 19716 339925
rect 19684 339875 19716 339876
rect 19684 339845 19685 339875
rect 19685 339845 19715 339875
rect 19715 339845 19716 339875
rect 19684 339844 19716 339845
rect 19684 339795 19716 339796
rect 19684 339765 19685 339795
rect 19685 339765 19715 339795
rect 19715 339765 19716 339795
rect 19684 339764 19716 339765
rect 19684 339715 19716 339716
rect 19684 339685 19685 339715
rect 19685 339685 19715 339715
rect 19715 339685 19716 339715
rect 19684 339684 19716 339685
rect 19684 339635 19716 339636
rect 19684 339605 19685 339635
rect 19685 339605 19715 339635
rect 19715 339605 19716 339635
rect 19684 339604 19716 339605
rect 19684 339555 19716 339556
rect 19684 339525 19685 339555
rect 19685 339525 19715 339555
rect 19715 339525 19716 339555
rect 19684 339524 19716 339525
rect 19684 339475 19716 339476
rect 19684 339445 19685 339475
rect 19685 339445 19715 339475
rect 19715 339445 19716 339475
rect 19684 339444 19716 339445
rect 19684 339395 19716 339396
rect 19684 339365 19685 339395
rect 19685 339365 19715 339395
rect 19715 339365 19716 339395
rect 19684 339364 19716 339365
rect 19684 339315 19716 339316
rect 19684 339285 19685 339315
rect 19685 339285 19715 339315
rect 19715 339285 19716 339315
rect 19684 339284 19716 339285
rect 19684 339235 19716 339236
rect 19684 339205 19685 339235
rect 19685 339205 19715 339235
rect 19715 339205 19716 339235
rect 19684 339204 19716 339205
rect 19684 339155 19716 339156
rect 19684 339125 19685 339155
rect 19685 339125 19715 339155
rect 19715 339125 19716 339155
rect 19684 339124 19716 339125
rect 19684 339075 19716 339076
rect 19684 339045 19685 339075
rect 19685 339045 19715 339075
rect 19715 339045 19716 339075
rect 19684 339044 19716 339045
rect 19684 338995 19716 338996
rect 19684 338965 19685 338995
rect 19685 338965 19715 338995
rect 19715 338965 19716 338995
rect 19684 338964 19716 338965
rect 19684 338915 19716 338916
rect 19684 338885 19685 338915
rect 19685 338885 19715 338915
rect 19715 338885 19716 338915
rect 19684 338884 19716 338885
rect 19684 338835 19716 338836
rect 19684 338805 19685 338835
rect 19685 338805 19715 338835
rect 19715 338805 19716 338835
rect 19684 338804 19716 338805
rect 19684 338755 19716 338756
rect 19684 338725 19685 338755
rect 19685 338725 19715 338755
rect 19715 338725 19716 338755
rect 19684 338724 19716 338725
rect 19684 338675 19716 338676
rect 19684 338645 19685 338675
rect 19685 338645 19715 338675
rect 19715 338645 19716 338675
rect 19684 338644 19716 338645
rect 19684 338595 19716 338596
rect 19684 338565 19685 338595
rect 19685 338565 19715 338595
rect 19715 338565 19716 338595
rect 19684 338564 19716 338565
rect 19684 338515 19716 338516
rect 19684 338485 19685 338515
rect 19685 338485 19715 338515
rect 19715 338485 19716 338515
rect 19684 338484 19716 338485
rect 19684 338435 19716 338436
rect 19684 338405 19685 338435
rect 19685 338405 19715 338435
rect 19715 338405 19716 338435
rect 19684 338404 19716 338405
rect 19684 338355 19716 338356
rect 19684 338325 19685 338355
rect 19685 338325 19715 338355
rect 19715 338325 19716 338355
rect 19684 338324 19716 338325
rect 19684 338275 19716 338276
rect 19684 338245 19685 338275
rect 19685 338245 19715 338275
rect 19715 338245 19716 338275
rect 19684 338244 19716 338245
rect 19684 338195 19716 338196
rect 19684 338165 19685 338195
rect 19685 338165 19715 338195
rect 19715 338165 19716 338195
rect 19684 338164 19716 338165
rect 19684 338115 19716 338116
rect 19684 338085 19685 338115
rect 19685 338085 19715 338115
rect 19715 338085 19716 338115
rect 19684 338084 19716 338085
rect 19684 338035 19716 338036
rect 19684 338005 19685 338035
rect 19685 338005 19715 338035
rect 19715 338005 19716 338035
rect 19684 338004 19716 338005
rect 19684 337955 19716 337956
rect 19684 337925 19685 337955
rect 19685 337925 19715 337955
rect 19715 337925 19716 337955
rect 19684 337924 19716 337925
rect 19684 337875 19716 337876
rect 19684 337845 19685 337875
rect 19685 337845 19715 337875
rect 19715 337845 19716 337875
rect 19684 337844 19716 337845
rect 19684 337795 19716 337796
rect 19684 337765 19685 337795
rect 19685 337765 19715 337795
rect 19715 337765 19716 337795
rect 19684 337764 19716 337765
rect 19684 337715 19716 337716
rect 19684 337685 19685 337715
rect 19685 337685 19715 337715
rect 19715 337685 19716 337715
rect 19684 337684 19716 337685
rect 19684 337635 19716 337636
rect 19684 337605 19685 337635
rect 19685 337605 19715 337635
rect 19715 337605 19716 337635
rect 19684 337604 19716 337605
rect 19684 337555 19716 337556
rect 19684 337525 19685 337555
rect 19685 337525 19715 337555
rect 19715 337525 19716 337555
rect 19684 337524 19716 337525
rect 19684 337475 19716 337476
rect 19684 337445 19685 337475
rect 19685 337445 19715 337475
rect 19715 337445 19716 337475
rect 19684 337444 19716 337445
rect 19684 337395 19716 337396
rect 19684 337365 19685 337395
rect 19685 337365 19715 337395
rect 19715 337365 19716 337395
rect 19684 337364 19716 337365
rect 19684 337315 19716 337316
rect 19684 337285 19685 337315
rect 19685 337285 19715 337315
rect 19715 337285 19716 337315
rect 19684 337284 19716 337285
rect 19684 337235 19716 337236
rect 19684 337205 19685 337235
rect 19685 337205 19715 337235
rect 19715 337205 19716 337235
rect 19684 337204 19716 337205
rect 19684 337155 19716 337156
rect 19684 337125 19685 337155
rect 19685 337125 19715 337155
rect 19715 337125 19716 337155
rect 19684 337124 19716 337125
rect 19684 337075 19716 337076
rect 19684 337045 19685 337075
rect 19685 337045 19715 337075
rect 19715 337045 19716 337075
rect 19684 337044 19716 337045
rect 19684 336995 19716 336996
rect 19684 336965 19685 336995
rect 19685 336965 19715 336995
rect 19715 336965 19716 336995
rect 19684 336964 19716 336965
rect 19684 336915 19716 336916
rect 19684 336885 19685 336915
rect 19685 336885 19715 336915
rect 19715 336885 19716 336915
rect 19684 336884 19716 336885
rect 19684 336835 19716 336836
rect 19684 336805 19685 336835
rect 19685 336805 19715 336835
rect 19715 336805 19716 336835
rect 19684 336804 19716 336805
rect 19684 336755 19716 336756
rect 19684 336725 19685 336755
rect 19685 336725 19715 336755
rect 19715 336725 19716 336755
rect 19684 336724 19716 336725
rect 19684 336675 19716 336676
rect 19684 336645 19685 336675
rect 19685 336645 19715 336675
rect 19715 336645 19716 336675
rect 19684 336644 19716 336645
rect 19684 336595 19716 336596
rect 19684 336565 19685 336595
rect 19685 336565 19715 336595
rect 19715 336565 19716 336595
rect 19684 336564 19716 336565
rect 19684 336515 19716 336516
rect 19684 336485 19685 336515
rect 19685 336485 19715 336515
rect 19715 336485 19716 336515
rect 19684 336484 19716 336485
rect 19684 336435 19716 336436
rect 19684 336405 19685 336435
rect 19685 336405 19715 336435
rect 19715 336405 19716 336435
rect 19684 336404 19716 336405
rect 19684 336355 19716 336356
rect 19684 336325 19685 336355
rect 19685 336325 19715 336355
rect 19715 336325 19716 336355
rect 19684 336324 19716 336325
rect 19684 336275 19716 336276
rect 19684 336245 19685 336275
rect 19685 336245 19715 336275
rect 19715 336245 19716 336275
rect 19684 336244 19716 336245
rect 19684 336195 19716 336196
rect 19684 336165 19685 336195
rect 19685 336165 19715 336195
rect 19715 336165 19716 336195
rect 19684 336164 19716 336165
rect 19684 336115 19716 336116
rect 19684 336085 19685 336115
rect 19685 336085 19715 336115
rect 19715 336085 19716 336115
rect 19684 336084 19716 336085
rect 19684 336035 19716 336036
rect 19684 336005 19685 336035
rect 19685 336005 19715 336035
rect 19715 336005 19716 336035
rect 19684 336004 19716 336005
rect 19684 335955 19716 335956
rect 19684 335925 19685 335955
rect 19685 335925 19715 335955
rect 19715 335925 19716 335955
rect 19684 335924 19716 335925
rect 19684 335875 19716 335876
rect 19684 335845 19685 335875
rect 19685 335845 19715 335875
rect 19715 335845 19716 335875
rect 19684 335844 19716 335845
rect 19684 335795 19716 335796
rect 19684 335765 19685 335795
rect 19685 335765 19715 335795
rect 19715 335765 19716 335795
rect 19684 335764 19716 335765
rect 19684 335715 19716 335716
rect 19684 335685 19685 335715
rect 19685 335685 19715 335715
rect 19715 335685 19716 335715
rect 19684 335684 19716 335685
rect 19684 335635 19716 335636
rect 19684 335605 19685 335635
rect 19685 335605 19715 335635
rect 19715 335605 19716 335635
rect 19684 335604 19716 335605
rect 19684 335555 19716 335556
rect 19684 335525 19685 335555
rect 19685 335525 19715 335555
rect 19715 335525 19716 335555
rect 19684 335524 19716 335525
rect 19684 335475 19716 335476
rect 19684 335445 19685 335475
rect 19685 335445 19715 335475
rect 19715 335445 19716 335475
rect 19684 335444 19716 335445
rect 19684 335395 19716 335396
rect 19684 335365 19685 335395
rect 19685 335365 19715 335395
rect 19715 335365 19716 335395
rect 19684 335364 19716 335365
rect 19684 335315 19716 335316
rect 19684 335285 19685 335315
rect 19685 335285 19715 335315
rect 19715 335285 19716 335315
rect 19684 335284 19716 335285
rect 19684 335235 19716 335236
rect 19684 335205 19685 335235
rect 19685 335205 19715 335235
rect 19715 335205 19716 335235
rect 19684 335204 19716 335205
rect 19684 335155 19716 335156
rect 19684 335125 19685 335155
rect 19685 335125 19715 335155
rect 19715 335125 19716 335155
rect 19684 335124 19716 335125
rect 19684 335075 19716 335076
rect 19684 335045 19685 335075
rect 19685 335045 19715 335075
rect 19715 335045 19716 335075
rect 19684 335044 19716 335045
rect 19684 334995 19716 334996
rect 19684 334965 19685 334995
rect 19685 334965 19715 334995
rect 19715 334965 19716 334995
rect 19684 334964 19716 334965
rect 19684 334915 19716 334916
rect 19684 334885 19685 334915
rect 19685 334885 19715 334915
rect 19715 334885 19716 334915
rect 19684 334884 19716 334885
rect 19684 334835 19716 334836
rect 19684 334805 19685 334835
rect 19685 334805 19715 334835
rect 19715 334805 19716 334835
rect 19684 334804 19716 334805
rect 19684 334755 19716 334756
rect 19684 334725 19685 334755
rect 19685 334725 19715 334755
rect 19715 334725 19716 334755
rect 19684 334724 19716 334725
rect 19684 334675 19716 334676
rect 19684 334645 19685 334675
rect 19685 334645 19715 334675
rect 19715 334645 19716 334675
rect 19684 334644 19716 334645
rect 19684 334595 19716 334596
rect 19684 334565 19685 334595
rect 19685 334565 19715 334595
rect 19715 334565 19716 334595
rect 19684 334564 19716 334565
rect 19684 334515 19716 334516
rect 19684 334485 19685 334515
rect 19685 334485 19715 334515
rect 19715 334485 19716 334515
rect 19684 334484 19716 334485
rect 19684 334435 19716 334436
rect 19684 334405 19685 334435
rect 19685 334405 19715 334435
rect 19715 334405 19716 334435
rect 19684 334404 19716 334405
rect 19684 334355 19716 334356
rect 19684 334325 19685 334355
rect 19685 334325 19715 334355
rect 19715 334325 19716 334355
rect 19684 334324 19716 334325
rect 19684 334275 19716 334276
rect 19684 334245 19685 334275
rect 19685 334245 19715 334275
rect 19715 334245 19716 334275
rect 19684 334244 19716 334245
rect 19684 334195 19716 334196
rect 19684 334165 19685 334195
rect 19685 334165 19715 334195
rect 19715 334165 19716 334195
rect 19684 334164 19716 334165
rect 19684 334115 19716 334116
rect 19684 334085 19685 334115
rect 19685 334085 19715 334115
rect 19715 334085 19716 334115
rect 19684 334084 19716 334085
rect 19684 334035 19716 334036
rect 19684 334005 19685 334035
rect 19685 334005 19715 334035
rect 19715 334005 19716 334035
rect 19684 334004 19716 334005
rect 19684 333955 19716 333956
rect 19684 333925 19685 333955
rect 19685 333925 19715 333955
rect 19715 333925 19716 333955
rect 19684 333924 19716 333925
rect 19684 333875 19716 333876
rect 19684 333845 19685 333875
rect 19685 333845 19715 333875
rect 19715 333845 19716 333875
rect 19684 333844 19716 333845
rect 19684 333795 19716 333796
rect 19684 333765 19685 333795
rect 19685 333765 19715 333795
rect 19715 333765 19716 333795
rect 19684 333764 19716 333765
rect 19684 333715 19716 333716
rect 19684 333685 19685 333715
rect 19685 333685 19715 333715
rect 19715 333685 19716 333715
rect 19684 333684 19716 333685
rect 19684 333635 19716 333636
rect 19684 333605 19685 333635
rect 19685 333605 19715 333635
rect 19715 333605 19716 333635
rect 19684 333604 19716 333605
rect 19684 333555 19716 333556
rect 19684 333525 19685 333555
rect 19685 333525 19715 333555
rect 19715 333525 19716 333555
rect 19684 333524 19716 333525
rect 19684 333475 19716 333476
rect 19684 333445 19685 333475
rect 19685 333445 19715 333475
rect 19715 333445 19716 333475
rect 19684 333444 19716 333445
rect 19684 333395 19716 333396
rect 19684 333365 19685 333395
rect 19685 333365 19715 333395
rect 19715 333365 19716 333395
rect 19684 333364 19716 333365
rect 19684 333315 19716 333316
rect 19684 333285 19685 333315
rect 19685 333285 19715 333315
rect 19715 333285 19716 333315
rect 19684 333284 19716 333285
rect 19684 333235 19716 333236
rect 19684 333205 19685 333235
rect 19685 333205 19715 333235
rect 19715 333205 19716 333235
rect 19684 333204 19716 333205
rect 19684 333155 19716 333156
rect 19684 333125 19685 333155
rect 19685 333125 19715 333155
rect 19715 333125 19716 333155
rect 19684 333124 19716 333125
rect 19684 333075 19716 333076
rect 19684 333045 19685 333075
rect 19685 333045 19715 333075
rect 19715 333045 19716 333075
rect 19684 333044 19716 333045
rect 19684 332995 19716 332996
rect 19684 332965 19685 332995
rect 19685 332965 19715 332995
rect 19715 332965 19716 332995
rect 19684 332964 19716 332965
rect 19684 332915 19716 332916
rect 19684 332885 19685 332915
rect 19685 332885 19715 332915
rect 19715 332885 19716 332915
rect 19684 332884 19716 332885
rect 19684 332835 19716 332836
rect 19684 332805 19685 332835
rect 19685 332805 19715 332835
rect 19715 332805 19716 332835
rect 19684 332804 19716 332805
rect 19684 332755 19716 332756
rect 19684 332725 19685 332755
rect 19685 332725 19715 332755
rect 19715 332725 19716 332755
rect 19684 332724 19716 332725
rect 19684 332675 19716 332676
rect 19684 332645 19685 332675
rect 19685 332645 19715 332675
rect 19715 332645 19716 332675
rect 19684 332644 19716 332645
rect 19684 332595 19716 332596
rect 19684 332565 19685 332595
rect 19685 332565 19715 332595
rect 19715 332565 19716 332595
rect 19684 332564 19716 332565
rect 19684 332515 19716 332516
rect 19684 332485 19685 332515
rect 19685 332485 19715 332515
rect 19715 332485 19716 332515
rect 19684 332484 19716 332485
rect 19684 332435 19716 332436
rect 19684 332405 19685 332435
rect 19685 332405 19715 332435
rect 19715 332405 19716 332435
rect 19684 332404 19716 332405
rect 19684 332355 19716 332356
rect 19684 332325 19685 332355
rect 19685 332325 19715 332355
rect 19715 332325 19716 332355
rect 19684 332324 19716 332325
rect 19684 332275 19716 332276
rect 19684 332245 19685 332275
rect 19685 332245 19715 332275
rect 19715 332245 19716 332275
rect 19684 332244 19716 332245
rect 19684 332195 19716 332196
rect 19684 332165 19685 332195
rect 19685 332165 19715 332195
rect 19715 332165 19716 332195
rect 19684 332164 19716 332165
rect 19684 332115 19716 332116
rect 19684 332085 19685 332115
rect 19685 332085 19715 332115
rect 19715 332085 19716 332115
rect 19684 332084 19716 332085
rect 19684 332035 19716 332036
rect 19684 332005 19685 332035
rect 19685 332005 19715 332035
rect 19715 332005 19716 332035
rect 19684 332004 19716 332005
rect 19684 331955 19716 331956
rect 19684 331925 19685 331955
rect 19685 331925 19715 331955
rect 19715 331925 19716 331955
rect 19684 331924 19716 331925
rect 19684 331875 19716 331876
rect 19684 331845 19685 331875
rect 19685 331845 19715 331875
rect 19715 331845 19716 331875
rect 19684 331844 19716 331845
rect 19684 331795 19716 331796
rect 19684 331765 19685 331795
rect 19685 331765 19715 331795
rect 19715 331765 19716 331795
rect 19684 331764 19716 331765
rect 19684 331715 19716 331716
rect 19684 331685 19685 331715
rect 19685 331685 19715 331715
rect 19715 331685 19716 331715
rect 19684 331684 19716 331685
rect 19684 331635 19716 331636
rect 19684 331605 19685 331635
rect 19685 331605 19715 331635
rect 19715 331605 19716 331635
rect 19684 331604 19716 331605
rect 19684 331555 19716 331556
rect 19684 331525 19685 331555
rect 19685 331525 19715 331555
rect 19715 331525 19716 331555
rect 19684 331524 19716 331525
rect 19684 331475 19716 331476
rect 19684 331445 19685 331475
rect 19685 331445 19715 331475
rect 19715 331445 19716 331475
rect 19684 331444 19716 331445
rect 19684 331395 19716 331396
rect 19684 331365 19685 331395
rect 19685 331365 19715 331395
rect 19715 331365 19716 331395
rect 19684 331364 19716 331365
rect 19684 331315 19716 331316
rect 19684 331285 19685 331315
rect 19685 331285 19715 331315
rect 19715 331285 19716 331315
rect 19684 331284 19716 331285
rect 19684 331235 19716 331236
rect 19684 331205 19685 331235
rect 19685 331205 19715 331235
rect 19715 331205 19716 331235
rect 19684 331204 19716 331205
rect 19684 331155 19716 331156
rect 19684 331125 19685 331155
rect 19685 331125 19715 331155
rect 19715 331125 19716 331155
rect 19684 331124 19716 331125
rect 19684 331075 19716 331076
rect 19684 331045 19685 331075
rect 19685 331045 19715 331075
rect 19715 331045 19716 331075
rect 19684 331044 19716 331045
rect 19684 330995 19716 330996
rect 19684 330965 19685 330995
rect 19685 330965 19715 330995
rect 19715 330965 19716 330995
rect 19684 330964 19716 330965
rect 19684 330915 19716 330916
rect 19684 330885 19685 330915
rect 19685 330885 19715 330915
rect 19715 330885 19716 330915
rect 19684 330884 19716 330885
rect 19684 330835 19716 330836
rect 19684 330805 19685 330835
rect 19685 330805 19715 330835
rect 19715 330805 19716 330835
rect 19684 330804 19716 330805
rect 19684 330755 19716 330756
rect 19684 330725 19685 330755
rect 19685 330725 19715 330755
rect 19715 330725 19716 330755
rect 19684 330724 19716 330725
rect 19684 330675 19716 330676
rect 19684 330645 19685 330675
rect 19685 330645 19715 330675
rect 19715 330645 19716 330675
rect 19684 330644 19716 330645
rect 19684 330595 19716 330596
rect 19684 330565 19685 330595
rect 19685 330565 19715 330595
rect 19715 330565 19716 330595
rect 19684 330564 19716 330565
rect 19684 330515 19716 330516
rect 19684 330485 19685 330515
rect 19685 330485 19715 330515
rect 19715 330485 19716 330515
rect 19684 330484 19716 330485
rect 19684 330435 19716 330436
rect 19684 330405 19685 330435
rect 19685 330405 19715 330435
rect 19715 330405 19716 330435
rect 19684 330404 19716 330405
rect 19684 330355 19716 330356
rect 19684 330325 19685 330355
rect 19685 330325 19715 330355
rect 19715 330325 19716 330355
rect 19684 330324 19716 330325
rect 19684 330275 19716 330276
rect 19684 330245 19685 330275
rect 19685 330245 19715 330275
rect 19715 330245 19716 330275
rect 19684 330244 19716 330245
rect 19684 330195 19716 330196
rect 19684 330165 19685 330195
rect 19685 330165 19715 330195
rect 19715 330165 19716 330195
rect 19684 330164 19716 330165
rect 19684 330115 19716 330116
rect 19684 330085 19685 330115
rect 19685 330085 19715 330115
rect 19715 330085 19716 330115
rect 19684 330084 19716 330085
rect 19684 330035 19716 330036
rect 19684 330005 19685 330035
rect 19685 330005 19715 330035
rect 19715 330005 19716 330035
rect 19684 330004 19716 330005
rect 19684 329955 19716 329956
rect 19684 329925 19685 329955
rect 19685 329925 19715 329955
rect 19715 329925 19716 329955
rect 19684 329924 19716 329925
rect 19684 329875 19716 329876
rect 19684 329845 19685 329875
rect 19685 329845 19715 329875
rect 19715 329845 19716 329875
rect 19684 329844 19716 329845
rect 19684 329795 19716 329796
rect 19684 329765 19685 329795
rect 19685 329765 19715 329795
rect 19715 329765 19716 329795
rect 19684 329764 19716 329765
rect 19684 329715 19716 329716
rect 19684 329685 19685 329715
rect 19685 329685 19715 329715
rect 19715 329685 19716 329715
rect 19684 329684 19716 329685
rect 19684 329635 19716 329636
rect 19684 329605 19685 329635
rect 19685 329605 19715 329635
rect 19715 329605 19716 329635
rect 19684 329604 19716 329605
rect 19684 329555 19716 329556
rect 19684 329525 19685 329555
rect 19685 329525 19715 329555
rect 19715 329525 19716 329555
rect 19684 329524 19716 329525
rect 19684 329475 19716 329476
rect 19684 329445 19685 329475
rect 19685 329445 19715 329475
rect 19715 329445 19716 329475
rect 19684 329444 19716 329445
rect 19684 329395 19716 329396
rect 19684 329365 19685 329395
rect 19685 329365 19715 329395
rect 19715 329365 19716 329395
rect 19684 329364 19716 329365
rect 19684 329315 19716 329316
rect 19684 329285 19685 329315
rect 19685 329285 19715 329315
rect 19715 329285 19716 329315
rect 19684 329284 19716 329285
rect 19684 329235 19716 329236
rect 19684 329205 19685 329235
rect 19685 329205 19715 329235
rect 19715 329205 19716 329235
rect 19684 329204 19716 329205
rect 19684 329155 19716 329156
rect 19684 329125 19685 329155
rect 19685 329125 19715 329155
rect 19715 329125 19716 329155
rect 19684 329124 19716 329125
rect 19684 329075 19716 329076
rect 19684 329045 19685 329075
rect 19685 329045 19715 329075
rect 19715 329045 19716 329075
rect 19684 329044 19716 329045
rect 19684 328995 19716 328996
rect 19684 328965 19685 328995
rect 19685 328965 19715 328995
rect 19715 328965 19716 328995
rect 19684 328964 19716 328965
rect 19684 328915 19716 328916
rect 19684 328885 19685 328915
rect 19685 328885 19715 328915
rect 19715 328885 19716 328915
rect 19684 328884 19716 328885
rect 19684 328835 19716 328836
rect 19684 328805 19685 328835
rect 19685 328805 19715 328835
rect 19715 328805 19716 328835
rect 19684 328804 19716 328805
rect 19684 328755 19716 328756
rect 19684 328725 19685 328755
rect 19685 328725 19715 328755
rect 19715 328725 19716 328755
rect 19684 328724 19716 328725
rect 19684 328675 19716 328676
rect 19684 328645 19685 328675
rect 19685 328645 19715 328675
rect 19715 328645 19716 328675
rect 19684 328644 19716 328645
rect 19684 328595 19716 328596
rect 19684 328565 19685 328595
rect 19685 328565 19715 328595
rect 19715 328565 19716 328595
rect 19684 328564 19716 328565
rect 19684 328515 19716 328516
rect 19684 328485 19685 328515
rect 19685 328485 19715 328515
rect 19715 328485 19716 328515
rect 19684 328484 19716 328485
rect 19684 328435 19716 328436
rect 19684 328405 19685 328435
rect 19685 328405 19715 328435
rect 19715 328405 19716 328435
rect 19684 328404 19716 328405
rect 19684 328355 19716 328356
rect 19684 328325 19685 328355
rect 19685 328325 19715 328355
rect 19715 328325 19716 328355
rect 19684 328324 19716 328325
rect 19684 328275 19716 328276
rect 19684 328245 19685 328275
rect 19685 328245 19715 328275
rect 19715 328245 19716 328275
rect 19684 328244 19716 328245
rect 19684 328195 19716 328196
rect 19684 328165 19685 328195
rect 19685 328165 19715 328195
rect 19715 328165 19716 328195
rect 19684 328164 19716 328165
rect 19684 328115 19716 328116
rect 19684 328085 19685 328115
rect 19685 328085 19715 328115
rect 19715 328085 19716 328115
rect 19684 328084 19716 328085
rect 19684 328035 19716 328036
rect 19684 328005 19685 328035
rect 19685 328005 19715 328035
rect 19715 328005 19716 328035
rect 19684 328004 19716 328005
rect 19684 327955 19716 327956
rect 19684 327925 19685 327955
rect 19685 327925 19715 327955
rect 19715 327925 19716 327955
rect 19684 327924 19716 327925
rect 19684 327875 19716 327876
rect 19684 327845 19685 327875
rect 19685 327845 19715 327875
rect 19715 327845 19716 327875
rect 19684 327844 19716 327845
rect 19684 327795 19716 327796
rect 19684 327765 19685 327795
rect 19685 327765 19715 327795
rect 19715 327765 19716 327795
rect 19684 327764 19716 327765
rect 19684 327715 19716 327716
rect 19684 327685 19685 327715
rect 19685 327685 19715 327715
rect 19715 327685 19716 327715
rect 19684 327684 19716 327685
rect 19684 327635 19716 327636
rect 19684 327605 19685 327635
rect 19685 327605 19715 327635
rect 19715 327605 19716 327635
rect 19684 327604 19716 327605
rect 19684 327555 19716 327556
rect 19684 327525 19685 327555
rect 19685 327525 19715 327555
rect 19715 327525 19716 327555
rect 19684 327524 19716 327525
rect 19684 327475 19716 327476
rect 19684 327445 19685 327475
rect 19685 327445 19715 327475
rect 19715 327445 19716 327475
rect 19684 327444 19716 327445
rect 19684 327395 19716 327396
rect 19684 327365 19685 327395
rect 19685 327365 19715 327395
rect 19715 327365 19716 327395
rect 19684 327364 19716 327365
rect 19684 327315 19716 327316
rect 19684 327285 19685 327315
rect 19685 327285 19715 327315
rect 19715 327285 19716 327315
rect 19684 327284 19716 327285
rect 19684 327235 19716 327236
rect 19684 327205 19685 327235
rect 19685 327205 19715 327235
rect 19715 327205 19716 327235
rect 19684 327204 19716 327205
rect 19684 327155 19716 327156
rect 19684 327125 19685 327155
rect 19685 327125 19715 327155
rect 19715 327125 19716 327155
rect 19684 327124 19716 327125
rect 19684 327075 19716 327076
rect 19684 327045 19685 327075
rect 19685 327045 19715 327075
rect 19715 327045 19716 327075
rect 19684 327044 19716 327045
rect 19684 326995 19716 326996
rect 19684 326965 19685 326995
rect 19685 326965 19715 326995
rect 19715 326965 19716 326995
rect 19684 326964 19716 326965
rect 19684 326915 19716 326916
rect 19684 326885 19685 326915
rect 19685 326885 19715 326915
rect 19715 326885 19716 326915
rect 19684 326884 19716 326885
rect 19684 326835 19716 326836
rect 19684 326805 19685 326835
rect 19685 326805 19715 326835
rect 19715 326805 19716 326835
rect 19684 326804 19716 326805
rect 19684 326755 19716 326756
rect 19684 326725 19685 326755
rect 19685 326725 19715 326755
rect 19715 326725 19716 326755
rect 19684 326724 19716 326725
rect 19684 326675 19716 326676
rect 19684 326645 19685 326675
rect 19685 326645 19715 326675
rect 19715 326645 19716 326675
rect 19684 326644 19716 326645
rect 19684 326595 19716 326596
rect 19684 326565 19685 326595
rect 19685 326565 19715 326595
rect 19715 326565 19716 326595
rect 19684 326564 19716 326565
rect 19684 326515 19716 326516
rect 19684 326485 19685 326515
rect 19685 326485 19715 326515
rect 19715 326485 19716 326515
rect 19684 326484 19716 326485
rect 19684 326435 19716 326436
rect 19684 326405 19685 326435
rect 19685 326405 19715 326435
rect 19715 326405 19716 326435
rect 19684 326404 19716 326405
rect 19684 326355 19716 326356
rect 19684 326325 19685 326355
rect 19685 326325 19715 326355
rect 19715 326325 19716 326355
rect 19684 326324 19716 326325
rect 19684 326275 19716 326276
rect 19684 326245 19685 326275
rect 19685 326245 19715 326275
rect 19715 326245 19716 326275
rect 19684 326244 19716 326245
rect 19684 326195 19716 326196
rect 19684 326165 19685 326195
rect 19685 326165 19715 326195
rect 19715 326165 19716 326195
rect 19684 326164 19716 326165
rect 19684 326115 19716 326116
rect 19684 326085 19685 326115
rect 19685 326085 19715 326115
rect 19715 326085 19716 326115
rect 19684 326084 19716 326085
rect 19684 326035 19716 326036
rect 19684 326005 19685 326035
rect 19685 326005 19715 326035
rect 19715 326005 19716 326035
rect 19684 326004 19716 326005
rect 19684 325955 19716 325956
rect 19684 325925 19685 325955
rect 19685 325925 19715 325955
rect 19715 325925 19716 325955
rect 19684 325924 19716 325925
rect 19684 325875 19716 325876
rect 19684 325845 19685 325875
rect 19685 325845 19715 325875
rect 19715 325845 19716 325875
rect 19684 325844 19716 325845
rect 19684 325795 19716 325796
rect 19684 325765 19685 325795
rect 19685 325765 19715 325795
rect 19715 325765 19716 325795
rect 19684 325764 19716 325765
rect 19684 325715 19716 325716
rect 19684 325685 19685 325715
rect 19685 325685 19715 325715
rect 19715 325685 19716 325715
rect 19684 325684 19716 325685
rect 19684 325635 19716 325636
rect 19684 325605 19685 325635
rect 19685 325605 19715 325635
rect 19715 325605 19716 325635
rect 19684 325604 19716 325605
rect 19684 325555 19716 325556
rect 19684 325525 19685 325555
rect 19685 325525 19715 325555
rect 19715 325525 19716 325555
rect 19684 325524 19716 325525
rect 19684 325475 19716 325476
rect 19684 325445 19685 325475
rect 19685 325445 19715 325475
rect 19715 325445 19716 325475
rect 19684 325444 19716 325445
rect 19684 325395 19716 325396
rect 19684 325365 19685 325395
rect 19685 325365 19715 325395
rect 19715 325365 19716 325395
rect 19684 325364 19716 325365
rect 19684 325315 19716 325316
rect 19684 325285 19685 325315
rect 19685 325285 19715 325315
rect 19715 325285 19716 325315
rect 19684 325284 19716 325285
rect 19684 325235 19716 325236
rect 19684 325205 19685 325235
rect 19685 325205 19715 325235
rect 19715 325205 19716 325235
rect 19684 325204 19716 325205
rect 19684 325155 19716 325156
rect 19684 325125 19685 325155
rect 19685 325125 19715 325155
rect 19715 325125 19716 325155
rect 19684 325124 19716 325125
rect 19684 325075 19716 325076
rect 19684 325045 19685 325075
rect 19685 325045 19715 325075
rect 19715 325045 19716 325075
rect 19684 325044 19716 325045
rect 19684 324995 19716 324996
rect 19684 324965 19685 324995
rect 19685 324965 19715 324995
rect 19715 324965 19716 324995
rect 19684 324964 19716 324965
rect 19684 324915 19716 324916
rect 19684 324885 19685 324915
rect 19685 324885 19715 324915
rect 19715 324885 19716 324915
rect 19684 324884 19716 324885
rect 19684 324835 19716 324836
rect 19684 324805 19685 324835
rect 19685 324805 19715 324835
rect 19715 324805 19716 324835
rect 19684 324804 19716 324805
rect 19684 324755 19716 324756
rect 19684 324725 19685 324755
rect 19685 324725 19715 324755
rect 19715 324725 19716 324755
rect 19684 324724 19716 324725
rect 19684 324675 19716 324676
rect 19684 324645 19685 324675
rect 19685 324645 19715 324675
rect 19715 324645 19716 324675
rect 19684 324644 19716 324645
rect 19684 324595 19716 324596
rect 19684 324565 19685 324595
rect 19685 324565 19715 324595
rect 19715 324565 19716 324595
rect 19684 324564 19716 324565
rect 19684 324515 19716 324516
rect 19684 324485 19685 324515
rect 19685 324485 19715 324515
rect 19715 324485 19716 324515
rect 19684 324484 19716 324485
rect 19684 324435 19716 324436
rect 19684 324405 19685 324435
rect 19685 324405 19715 324435
rect 19715 324405 19716 324435
rect 19684 324404 19716 324405
rect 19684 324355 19716 324356
rect 19684 324325 19685 324355
rect 19685 324325 19715 324355
rect 19715 324325 19716 324355
rect 19684 324324 19716 324325
rect 19684 324275 19716 324276
rect 19684 324245 19685 324275
rect 19685 324245 19715 324275
rect 19715 324245 19716 324275
rect 19684 324244 19716 324245
rect 19684 324195 19716 324196
rect 19684 324165 19685 324195
rect 19685 324165 19715 324195
rect 19715 324165 19716 324195
rect 19684 324164 19716 324165
rect 19684 324115 19716 324116
rect 19684 324085 19685 324115
rect 19685 324085 19715 324115
rect 19715 324085 19716 324115
rect 19684 324084 19716 324085
rect 19684 324035 19716 324036
rect 19684 324005 19685 324035
rect 19685 324005 19715 324035
rect 19715 324005 19716 324035
rect 19684 324004 19716 324005
rect 19684 323955 19716 323956
rect 19684 323925 19685 323955
rect 19685 323925 19715 323955
rect 19715 323925 19716 323955
rect 19684 323924 19716 323925
rect 19684 323875 19716 323876
rect 19684 323845 19685 323875
rect 19685 323845 19715 323875
rect 19715 323845 19716 323875
rect 19684 323844 19716 323845
rect 19684 323795 19716 323796
rect 19684 323765 19685 323795
rect 19685 323765 19715 323795
rect 19715 323765 19716 323795
rect 19684 323764 19716 323765
rect 19684 323715 19716 323716
rect 19684 323685 19685 323715
rect 19685 323685 19715 323715
rect 19715 323685 19716 323715
rect 19684 323684 19716 323685
rect 19684 323635 19716 323636
rect 19684 323605 19685 323635
rect 19685 323605 19715 323635
rect 19715 323605 19716 323635
rect 19684 323604 19716 323605
rect 19684 323555 19716 323556
rect 19684 323525 19685 323555
rect 19685 323525 19715 323555
rect 19715 323525 19716 323555
rect 19684 323524 19716 323525
rect 19684 323475 19716 323476
rect 19684 323445 19685 323475
rect 19685 323445 19715 323475
rect 19715 323445 19716 323475
rect 19684 323444 19716 323445
rect 19684 323395 19716 323396
rect 19684 323365 19685 323395
rect 19685 323365 19715 323395
rect 19715 323365 19716 323395
rect 19684 323364 19716 323365
rect 19684 323315 19716 323316
rect 19684 323285 19685 323315
rect 19685 323285 19715 323315
rect 19715 323285 19716 323315
rect 19684 323284 19716 323285
rect 19684 323235 19716 323236
rect 19684 323205 19685 323235
rect 19685 323205 19715 323235
rect 19715 323205 19716 323235
rect 19684 323204 19716 323205
rect 19684 323155 19716 323156
rect 19684 323125 19685 323155
rect 19685 323125 19715 323155
rect 19715 323125 19716 323155
rect 19684 323124 19716 323125
rect 19684 323075 19716 323076
rect 19684 323045 19685 323075
rect 19685 323045 19715 323075
rect 19715 323045 19716 323075
rect 19684 323044 19716 323045
rect 19684 322995 19716 322996
rect 19684 322965 19685 322995
rect 19685 322965 19715 322995
rect 19715 322965 19716 322995
rect 19684 322964 19716 322965
rect 19684 322915 19716 322916
rect 19684 322885 19685 322915
rect 19685 322885 19715 322915
rect 19715 322885 19716 322915
rect 19684 322884 19716 322885
rect 19684 322835 19716 322836
rect 19684 322805 19685 322835
rect 19685 322805 19715 322835
rect 19715 322805 19716 322835
rect 19684 322804 19716 322805
rect 19684 322755 19716 322756
rect 19684 322725 19685 322755
rect 19685 322725 19715 322755
rect 19715 322725 19716 322755
rect 19684 322724 19716 322725
rect 19684 322675 19716 322676
rect 19684 322645 19685 322675
rect 19685 322645 19715 322675
rect 19715 322645 19716 322675
rect 19684 322644 19716 322645
rect 19684 322595 19716 322596
rect 19684 322565 19685 322595
rect 19685 322565 19715 322595
rect 19715 322565 19716 322595
rect 19684 322564 19716 322565
rect 19684 322515 19716 322516
rect 19684 322485 19685 322515
rect 19685 322485 19715 322515
rect 19715 322485 19716 322515
rect 19684 322484 19716 322485
rect 19684 322435 19716 322436
rect 19684 322405 19685 322435
rect 19685 322405 19715 322435
rect 19715 322405 19716 322435
rect 19684 322404 19716 322405
rect 19684 322355 19716 322356
rect 19684 322325 19685 322355
rect 19685 322325 19715 322355
rect 19715 322325 19716 322355
rect 19684 322324 19716 322325
rect 19684 322275 19716 322276
rect 19684 322245 19685 322275
rect 19685 322245 19715 322275
rect 19715 322245 19716 322275
rect 19684 322244 19716 322245
rect 19684 322195 19716 322196
rect 19684 322165 19685 322195
rect 19685 322165 19715 322195
rect 19715 322165 19716 322195
rect 19684 322164 19716 322165
rect 19684 322115 19716 322116
rect 19684 322085 19685 322115
rect 19685 322085 19715 322115
rect 19715 322085 19716 322115
rect 19684 322084 19716 322085
rect 19684 322035 19716 322036
rect 19684 322005 19685 322035
rect 19685 322005 19715 322035
rect 19715 322005 19716 322035
rect 19684 322004 19716 322005
rect 19684 321955 19716 321956
rect 19684 321925 19685 321955
rect 19685 321925 19715 321955
rect 19715 321925 19716 321955
rect 19684 321924 19716 321925
rect 19684 321875 19716 321876
rect 19684 321845 19685 321875
rect 19685 321845 19715 321875
rect 19715 321845 19716 321875
rect 19684 321844 19716 321845
rect 19684 321795 19716 321796
rect 19684 321765 19685 321795
rect 19685 321765 19715 321795
rect 19715 321765 19716 321795
rect 19684 321764 19716 321765
rect 19684 321715 19716 321716
rect 19684 321685 19685 321715
rect 19685 321685 19715 321715
rect 19715 321685 19716 321715
rect 19684 321684 19716 321685
rect 19684 321635 19716 321636
rect 19684 321605 19685 321635
rect 19685 321605 19715 321635
rect 19715 321605 19716 321635
rect 19684 321604 19716 321605
rect 19684 321555 19716 321556
rect 19684 321525 19685 321555
rect 19685 321525 19715 321555
rect 19715 321525 19716 321555
rect 19684 321524 19716 321525
rect 19684 321475 19716 321476
rect 19684 321445 19685 321475
rect 19685 321445 19715 321475
rect 19715 321445 19716 321475
rect 19684 321444 19716 321445
rect 19684 321395 19716 321396
rect 19684 321365 19685 321395
rect 19685 321365 19715 321395
rect 19715 321365 19716 321395
rect 19684 321364 19716 321365
rect 19684 321315 19716 321316
rect 19684 321285 19685 321315
rect 19685 321285 19715 321315
rect 19715 321285 19716 321315
rect 19684 321284 19716 321285
rect 19684 321235 19716 321236
rect 19684 321205 19685 321235
rect 19685 321205 19715 321235
rect 19715 321205 19716 321235
rect 19684 321204 19716 321205
rect 19684 321155 19716 321156
rect 19684 321125 19685 321155
rect 19685 321125 19715 321155
rect 19715 321125 19716 321155
rect 19684 321124 19716 321125
rect 19684 321075 19716 321076
rect 19684 321045 19685 321075
rect 19685 321045 19715 321075
rect 19715 321045 19716 321075
rect 19684 321044 19716 321045
rect 19684 320995 19716 320996
rect 19684 320965 19685 320995
rect 19685 320965 19715 320995
rect 19715 320965 19716 320995
rect 19684 320964 19716 320965
rect 19684 320915 19716 320916
rect 19684 320885 19685 320915
rect 19685 320885 19715 320915
rect 19715 320885 19716 320915
rect 19684 320884 19716 320885
rect 19684 320835 19716 320836
rect 19684 320805 19685 320835
rect 19685 320805 19715 320835
rect 19715 320805 19716 320835
rect 19684 320804 19716 320805
rect 19684 320755 19716 320756
rect 19684 320725 19685 320755
rect 19685 320725 19715 320755
rect 19715 320725 19716 320755
rect 19684 320724 19716 320725
rect 19684 320675 19716 320676
rect 19684 320645 19685 320675
rect 19685 320645 19715 320675
rect 19715 320645 19716 320675
rect 19684 320644 19716 320645
rect 19684 320595 19716 320596
rect 19684 320565 19685 320595
rect 19685 320565 19715 320595
rect 19715 320565 19716 320595
rect 19684 320564 19716 320565
rect 19684 320515 19716 320516
rect 19684 320485 19685 320515
rect 19685 320485 19715 320515
rect 19715 320485 19716 320515
rect 19684 320484 19716 320485
rect 19684 320435 19716 320436
rect 19684 320405 19685 320435
rect 19685 320405 19715 320435
rect 19715 320405 19716 320435
rect 19684 320404 19716 320405
rect 19684 320355 19716 320356
rect 19684 320325 19685 320355
rect 19685 320325 19715 320355
rect 19715 320325 19716 320355
rect 19684 320324 19716 320325
rect 19684 320275 19716 320276
rect 19684 320245 19685 320275
rect 19685 320245 19715 320275
rect 19715 320245 19716 320275
rect 19684 320244 19716 320245
rect 19684 320195 19716 320196
rect 19684 320165 19685 320195
rect 19685 320165 19715 320195
rect 19715 320165 19716 320195
rect 19684 320164 19716 320165
rect 19684 320115 19716 320116
rect 19684 320085 19685 320115
rect 19685 320085 19715 320115
rect 19715 320085 19716 320115
rect 19684 320084 19716 320085
rect 19684 320035 19716 320036
rect 19684 320005 19685 320035
rect 19685 320005 19715 320035
rect 19715 320005 19716 320035
rect 19684 320004 19716 320005
rect 19684 319955 19716 319956
rect 19684 319925 19685 319955
rect 19685 319925 19715 319955
rect 19715 319925 19716 319955
rect 19684 319924 19716 319925
rect 19684 319875 19716 319876
rect 19684 319845 19685 319875
rect 19685 319845 19715 319875
rect 19715 319845 19716 319875
rect 19684 319844 19716 319845
rect 19684 319795 19716 319796
rect 19684 319765 19685 319795
rect 19685 319765 19715 319795
rect 19715 319765 19716 319795
rect 19684 319764 19716 319765
rect 19684 319715 19716 319716
rect 19684 319685 19685 319715
rect 19685 319685 19715 319715
rect 19715 319685 19716 319715
rect 19684 319684 19716 319685
rect 19684 319635 19716 319636
rect 19684 319605 19685 319635
rect 19685 319605 19715 319635
rect 19715 319605 19716 319635
rect 19684 319604 19716 319605
rect 19684 319555 19716 319556
rect 19684 319525 19685 319555
rect 19685 319525 19715 319555
rect 19715 319525 19716 319555
rect 19684 319524 19716 319525
rect 19684 319475 19716 319476
rect 19684 319445 19685 319475
rect 19685 319445 19715 319475
rect 19715 319445 19716 319475
rect 19684 319444 19716 319445
rect 19684 319395 19716 319396
rect 19684 319365 19685 319395
rect 19685 319365 19715 319395
rect 19715 319365 19716 319395
rect 19684 319364 19716 319365
rect 19684 319315 19716 319316
rect 19684 319285 19685 319315
rect 19685 319285 19715 319315
rect 19715 319285 19716 319315
rect 19684 319284 19716 319285
rect 19684 319235 19716 319236
rect 19684 319205 19685 319235
rect 19685 319205 19715 319235
rect 19715 319205 19716 319235
rect 19684 319204 19716 319205
rect 19684 319155 19716 319156
rect 19684 319125 19685 319155
rect 19685 319125 19715 319155
rect 19715 319125 19716 319155
rect 19684 319124 19716 319125
rect 19684 319075 19716 319076
rect 19684 319045 19685 319075
rect 19685 319045 19715 319075
rect 19715 319045 19716 319075
rect 19684 319044 19716 319045
rect 19684 318995 19716 318996
rect 19684 318965 19685 318995
rect 19685 318965 19715 318995
rect 19715 318965 19716 318995
rect 19684 318964 19716 318965
rect 19684 318915 19716 318916
rect 19684 318885 19685 318915
rect 19685 318885 19715 318915
rect 19715 318885 19716 318915
rect 19684 318884 19716 318885
rect 19684 318835 19716 318836
rect 19684 318805 19685 318835
rect 19685 318805 19715 318835
rect 19715 318805 19716 318835
rect 19684 318804 19716 318805
rect 19684 318755 19716 318756
rect 19684 318725 19685 318755
rect 19685 318725 19715 318755
rect 19715 318725 19716 318755
rect 19684 318724 19716 318725
rect 19684 318675 19716 318676
rect 19684 318645 19685 318675
rect 19685 318645 19715 318675
rect 19715 318645 19716 318675
rect 19684 318644 19716 318645
rect 19684 318595 19716 318596
rect 19684 318565 19685 318595
rect 19685 318565 19715 318595
rect 19715 318565 19716 318595
rect 19684 318564 19716 318565
rect 19684 318515 19716 318516
rect 19684 318485 19685 318515
rect 19685 318485 19715 318515
rect 19715 318485 19716 318515
rect 19684 318484 19716 318485
rect 19684 318435 19716 318436
rect 19684 318405 19685 318435
rect 19685 318405 19715 318435
rect 19715 318405 19716 318435
rect 19684 318404 19716 318405
rect 19684 318355 19716 318356
rect 19684 318325 19685 318355
rect 19685 318325 19715 318355
rect 19715 318325 19716 318355
rect 19684 318324 19716 318325
rect 19684 318275 19716 318276
rect 19684 318245 19685 318275
rect 19685 318245 19715 318275
rect 19715 318245 19716 318275
rect 19684 318244 19716 318245
rect 19684 318195 19716 318196
rect 19684 318165 19685 318195
rect 19685 318165 19715 318195
rect 19715 318165 19716 318195
rect 19684 318164 19716 318165
rect 19684 318115 19716 318116
rect 19684 318085 19685 318115
rect 19685 318085 19715 318115
rect 19715 318085 19716 318115
rect 19684 318084 19716 318085
rect 19684 318035 19716 318036
rect 19684 318005 19685 318035
rect 19685 318005 19715 318035
rect 19715 318005 19716 318035
rect 19684 318004 19716 318005
rect 19684 317955 19716 317956
rect 19684 317925 19685 317955
rect 19685 317925 19715 317955
rect 19715 317925 19716 317955
rect 19684 317924 19716 317925
rect 19684 317875 19716 317876
rect 19684 317845 19685 317875
rect 19685 317845 19715 317875
rect 19715 317845 19716 317875
rect 19684 317844 19716 317845
rect 19684 317795 19716 317796
rect 19684 317765 19685 317795
rect 19685 317765 19715 317795
rect 19715 317765 19716 317795
rect 19684 317764 19716 317765
rect 19684 317715 19716 317716
rect 19684 317685 19685 317715
rect 19685 317685 19715 317715
rect 19715 317685 19716 317715
rect 19684 317684 19716 317685
rect 19684 317635 19716 317636
rect 19684 317605 19685 317635
rect 19685 317605 19715 317635
rect 19715 317605 19716 317635
rect 19684 317604 19716 317605
rect 19684 317555 19716 317556
rect 19684 317525 19685 317555
rect 19685 317525 19715 317555
rect 19715 317525 19716 317555
rect 19684 317524 19716 317525
rect 19684 317475 19716 317476
rect 19684 317445 19685 317475
rect 19685 317445 19715 317475
rect 19715 317445 19716 317475
rect 19684 317444 19716 317445
rect 19684 317395 19716 317396
rect 19684 317365 19685 317395
rect 19685 317365 19715 317395
rect 19715 317365 19716 317395
rect 19684 317364 19716 317365
rect 19684 317315 19716 317316
rect 19684 317285 19685 317315
rect 19685 317285 19715 317315
rect 19715 317285 19716 317315
rect 19684 317284 19716 317285
rect 19684 317235 19716 317236
rect 19684 317205 19685 317235
rect 19685 317205 19715 317235
rect 19715 317205 19716 317235
rect 19684 317204 19716 317205
rect 19684 317155 19716 317156
rect 19684 317125 19685 317155
rect 19685 317125 19715 317155
rect 19715 317125 19716 317155
rect 19684 317124 19716 317125
rect 19684 317075 19716 317076
rect 19684 317045 19685 317075
rect 19685 317045 19715 317075
rect 19715 317045 19716 317075
rect 19684 317044 19716 317045
rect 19684 316995 19716 316996
rect 19684 316965 19685 316995
rect 19685 316965 19715 316995
rect 19715 316965 19716 316995
rect 19684 316964 19716 316965
rect 19684 316915 19716 316916
rect 19684 316885 19685 316915
rect 19685 316885 19715 316915
rect 19715 316885 19716 316915
rect 19684 316884 19716 316885
rect 19684 316835 19716 316836
rect 19684 316805 19685 316835
rect 19685 316805 19715 316835
rect 19715 316805 19716 316835
rect 19684 316804 19716 316805
rect 19684 316755 19716 316756
rect 19684 316725 19685 316755
rect 19685 316725 19715 316755
rect 19715 316725 19716 316755
rect 19684 316724 19716 316725
rect 19684 316675 19716 316676
rect 19684 316645 19685 316675
rect 19685 316645 19715 316675
rect 19715 316645 19716 316675
rect 19684 316644 19716 316645
rect 19684 316595 19716 316596
rect 19684 316565 19685 316595
rect 19685 316565 19715 316595
rect 19715 316565 19716 316595
rect 19684 316564 19716 316565
rect 19684 316515 19716 316516
rect 19684 316485 19685 316515
rect 19685 316485 19715 316515
rect 19715 316485 19716 316515
rect 19684 316484 19716 316485
rect 19684 316435 19716 316436
rect 19684 316405 19685 316435
rect 19685 316405 19715 316435
rect 19715 316405 19716 316435
rect 19684 316404 19716 316405
rect 19684 316355 19716 316356
rect 19684 316325 19685 316355
rect 19685 316325 19715 316355
rect 19715 316325 19716 316355
rect 19684 316324 19716 316325
rect 19684 316275 19716 316276
rect 19684 316245 19685 316275
rect 19685 316245 19715 316275
rect 19715 316245 19716 316275
rect 19684 316244 19716 316245
rect 19684 316195 19716 316196
rect 19684 316165 19685 316195
rect 19685 316165 19715 316195
rect 19715 316165 19716 316195
rect 19684 316164 19716 316165
rect 19684 316115 19716 316116
rect 19684 316085 19685 316115
rect 19685 316085 19715 316115
rect 19715 316085 19716 316115
rect 19684 316084 19716 316085
rect 19684 316035 19716 316036
rect 19684 316005 19685 316035
rect 19685 316005 19715 316035
rect 19715 316005 19716 316035
rect 19684 316004 19716 316005
rect 19684 315955 19716 315956
rect 19684 315925 19685 315955
rect 19685 315925 19715 315955
rect 19715 315925 19716 315955
rect 19684 315924 19716 315925
rect 19684 315875 19716 315876
rect 19684 315845 19685 315875
rect 19685 315845 19715 315875
rect 19715 315845 19716 315875
rect 19684 315844 19716 315845
rect 19684 315795 19716 315796
rect 19684 315765 19685 315795
rect 19685 315765 19715 315795
rect 19715 315765 19716 315795
rect 19684 315764 19716 315765
rect 19684 315715 19716 315716
rect 19684 315685 19685 315715
rect 19685 315685 19715 315715
rect 19715 315685 19716 315715
rect 19684 315684 19716 315685
rect 19684 315635 19716 315636
rect 19684 315605 19685 315635
rect 19685 315605 19715 315635
rect 19715 315605 19716 315635
rect 19684 315604 19716 315605
rect 19684 315555 19716 315556
rect 19684 315525 19685 315555
rect 19685 315525 19715 315555
rect 19715 315525 19716 315555
rect 19684 315524 19716 315525
rect 19684 315475 19716 315476
rect 19684 315445 19685 315475
rect 19685 315445 19715 315475
rect 19715 315445 19716 315475
rect 19684 315444 19716 315445
rect 19684 315395 19716 315396
rect 19684 315365 19685 315395
rect 19685 315365 19715 315395
rect 19715 315365 19716 315395
rect 19684 315364 19716 315365
rect 19684 315315 19716 315316
rect 19684 315285 19685 315315
rect 19685 315285 19715 315315
rect 19715 315285 19716 315315
rect 19684 315284 19716 315285
rect 19684 315235 19716 315236
rect 19684 315205 19685 315235
rect 19685 315205 19715 315235
rect 19715 315205 19716 315235
rect 19684 315204 19716 315205
rect 19684 315155 19716 315156
rect 19684 315125 19685 315155
rect 19685 315125 19715 315155
rect 19715 315125 19716 315155
rect 19684 315124 19716 315125
rect 19684 315075 19716 315076
rect 19684 315045 19685 315075
rect 19685 315045 19715 315075
rect 19715 315045 19716 315075
rect 19684 315044 19716 315045
rect 19684 314995 19716 314996
rect 19684 314965 19685 314995
rect 19685 314965 19715 314995
rect 19715 314965 19716 314995
rect 19684 314964 19716 314965
rect 19684 314915 19716 314916
rect 19684 314885 19685 314915
rect 19685 314885 19715 314915
rect 19715 314885 19716 314915
rect 19684 314884 19716 314885
rect 19684 314835 19716 314836
rect 19684 314805 19685 314835
rect 19685 314805 19715 314835
rect 19715 314805 19716 314835
rect 19684 314804 19716 314805
rect 19684 314755 19716 314756
rect 19684 314725 19685 314755
rect 19685 314725 19715 314755
rect 19715 314725 19716 314755
rect 19684 314724 19716 314725
rect 19684 314675 19716 314676
rect 19684 314645 19685 314675
rect 19685 314645 19715 314675
rect 19715 314645 19716 314675
rect 19684 314644 19716 314645
rect 19684 314595 19716 314596
rect 19684 314565 19685 314595
rect 19685 314565 19715 314595
rect 19715 314565 19716 314595
rect 19684 314564 19716 314565
rect 19684 314515 19716 314516
rect 19684 314485 19685 314515
rect 19685 314485 19715 314515
rect 19715 314485 19716 314515
rect 19684 314484 19716 314485
rect 19684 314435 19716 314436
rect 19684 314405 19685 314435
rect 19685 314405 19715 314435
rect 19715 314405 19716 314435
rect 19684 314404 19716 314405
rect 19684 314355 19716 314356
rect 19684 314325 19685 314355
rect 19685 314325 19715 314355
rect 19715 314325 19716 314355
rect 19684 314324 19716 314325
rect 19684 314275 19716 314276
rect 19684 314245 19685 314275
rect 19685 314245 19715 314275
rect 19715 314245 19716 314275
rect 19684 314244 19716 314245
rect 19684 314195 19716 314196
rect 19684 314165 19685 314195
rect 19685 314165 19715 314195
rect 19715 314165 19716 314195
rect 19684 314164 19716 314165
rect 19684 314115 19716 314116
rect 19684 314085 19685 314115
rect 19685 314085 19715 314115
rect 19715 314085 19716 314115
rect 19684 314084 19716 314085
rect 19684 314035 19716 314036
rect 19684 314005 19685 314035
rect 19685 314005 19715 314035
rect 19715 314005 19716 314035
rect 19684 314004 19716 314005
rect 19684 313955 19716 313956
rect 19684 313925 19685 313955
rect 19685 313925 19715 313955
rect 19715 313925 19716 313955
rect 19684 313924 19716 313925
rect 19684 313875 19716 313876
rect 19684 313845 19685 313875
rect 19685 313845 19715 313875
rect 19715 313845 19716 313875
rect 19684 313844 19716 313845
rect 19684 313795 19716 313796
rect 19684 313765 19685 313795
rect 19685 313765 19715 313795
rect 19715 313765 19716 313795
rect 19684 313764 19716 313765
rect 19684 313715 19716 313716
rect 19684 313685 19685 313715
rect 19685 313685 19715 313715
rect 19715 313685 19716 313715
rect 19684 313684 19716 313685
rect 19684 313635 19716 313636
rect 19684 313605 19685 313635
rect 19685 313605 19715 313635
rect 19715 313605 19716 313635
rect 19684 313604 19716 313605
rect 19684 313555 19716 313556
rect 19684 313525 19685 313555
rect 19685 313525 19715 313555
rect 19715 313525 19716 313555
rect 19684 313524 19716 313525
rect 19684 313475 19716 313476
rect 19684 313445 19685 313475
rect 19685 313445 19715 313475
rect 19715 313445 19716 313475
rect 19684 313444 19716 313445
rect 19684 313395 19716 313396
rect 19684 313365 19685 313395
rect 19685 313365 19715 313395
rect 19715 313365 19716 313395
rect 19684 313364 19716 313365
rect 19684 313315 19716 313316
rect 19684 313285 19685 313315
rect 19685 313285 19715 313315
rect 19715 313285 19716 313315
rect 19684 313284 19716 313285
rect 19684 313235 19716 313236
rect 19684 313205 19685 313235
rect 19685 313205 19715 313235
rect 19715 313205 19716 313235
rect 19684 313204 19716 313205
rect 19684 313155 19716 313156
rect 19684 313125 19685 313155
rect 19685 313125 19715 313155
rect 19715 313125 19716 313155
rect 19684 313124 19716 313125
rect 19684 313075 19716 313076
rect 19684 313045 19685 313075
rect 19685 313045 19715 313075
rect 19715 313045 19716 313075
rect 19684 313044 19716 313045
rect 19684 312995 19716 312996
rect 19684 312965 19685 312995
rect 19685 312965 19715 312995
rect 19715 312965 19716 312995
rect 19684 312964 19716 312965
rect 19684 312915 19716 312916
rect 19684 312885 19685 312915
rect 19685 312885 19715 312915
rect 19715 312885 19716 312915
rect 19684 312884 19716 312885
rect 19684 312835 19716 312836
rect 19684 312805 19685 312835
rect 19685 312805 19715 312835
rect 19715 312805 19716 312835
rect 19684 312804 19716 312805
rect 19684 312755 19716 312756
rect 19684 312725 19685 312755
rect 19685 312725 19715 312755
rect 19715 312725 19716 312755
rect 19684 312724 19716 312725
rect 19684 312675 19716 312676
rect 19684 312645 19685 312675
rect 19685 312645 19715 312675
rect 19715 312645 19716 312675
rect 19684 312644 19716 312645
rect 19684 312595 19716 312596
rect 19684 312565 19685 312595
rect 19685 312565 19715 312595
rect 19715 312565 19716 312595
rect 19684 312564 19716 312565
rect 19684 312515 19716 312516
rect 19684 312485 19685 312515
rect 19685 312485 19715 312515
rect 19715 312485 19716 312515
rect 19684 312484 19716 312485
rect 19684 312435 19716 312436
rect 19684 312405 19685 312435
rect 19685 312405 19715 312435
rect 19715 312405 19716 312435
rect 19684 312404 19716 312405
rect 19684 312355 19716 312356
rect 19684 312325 19685 312355
rect 19685 312325 19715 312355
rect 19715 312325 19716 312355
rect 19684 312324 19716 312325
rect 19684 312275 19716 312276
rect 19684 312245 19685 312275
rect 19685 312245 19715 312275
rect 19715 312245 19716 312275
rect 19684 312244 19716 312245
rect 19684 312195 19716 312196
rect 19684 312165 19685 312195
rect 19685 312165 19715 312195
rect 19715 312165 19716 312195
rect 19684 312164 19716 312165
rect 19684 312115 19716 312116
rect 19684 312085 19685 312115
rect 19685 312085 19715 312115
rect 19715 312085 19716 312115
rect 19684 312084 19716 312085
rect 19684 312035 19716 312036
rect 19684 312005 19685 312035
rect 19685 312005 19715 312035
rect 19715 312005 19716 312035
rect 19684 312004 19716 312005
rect 19684 311955 19716 311956
rect 19684 311925 19685 311955
rect 19685 311925 19715 311955
rect 19715 311925 19716 311955
rect 19684 311924 19716 311925
rect 19684 311875 19716 311876
rect 19684 311845 19685 311875
rect 19685 311845 19715 311875
rect 19715 311845 19716 311875
rect 19684 311844 19716 311845
rect 19684 311795 19716 311796
rect 19684 311765 19685 311795
rect 19685 311765 19715 311795
rect 19715 311765 19716 311795
rect 19684 311764 19716 311765
rect 19684 311715 19716 311716
rect 19684 311685 19685 311715
rect 19685 311685 19715 311715
rect 19715 311685 19716 311715
rect 19684 311684 19716 311685
rect 19684 311635 19716 311636
rect 19684 311605 19685 311635
rect 19685 311605 19715 311635
rect 19715 311605 19716 311635
rect 19684 311604 19716 311605
rect 19684 311555 19716 311556
rect 19684 311525 19685 311555
rect 19685 311525 19715 311555
rect 19715 311525 19716 311555
rect 19684 311524 19716 311525
rect 19684 311475 19716 311476
rect 19684 311445 19685 311475
rect 19685 311445 19715 311475
rect 19715 311445 19716 311475
rect 19684 311444 19716 311445
rect 19684 311395 19716 311396
rect 19684 311365 19685 311395
rect 19685 311365 19715 311395
rect 19715 311365 19716 311395
rect 19684 311364 19716 311365
rect 19684 311315 19716 311316
rect 19684 311285 19685 311315
rect 19685 311285 19715 311315
rect 19715 311285 19716 311315
rect 19684 311284 19716 311285
rect 19684 311235 19716 311236
rect 19684 311205 19685 311235
rect 19685 311205 19715 311235
rect 19715 311205 19716 311235
rect 19684 311204 19716 311205
rect 19684 311155 19716 311156
rect 19684 311125 19685 311155
rect 19685 311125 19715 311155
rect 19715 311125 19716 311155
rect 19684 311124 19716 311125
rect 19684 311075 19716 311076
rect 19684 311045 19685 311075
rect 19685 311045 19715 311075
rect 19715 311045 19716 311075
rect 19684 311044 19716 311045
rect 19684 310995 19716 310996
rect 19684 310965 19685 310995
rect 19685 310965 19715 310995
rect 19715 310965 19716 310995
rect 19684 310964 19716 310965
rect 19684 310915 19716 310916
rect 19684 310885 19685 310915
rect 19685 310885 19715 310915
rect 19715 310885 19716 310915
rect 19684 310884 19716 310885
rect 19684 310835 19716 310836
rect 19684 310805 19685 310835
rect 19685 310805 19715 310835
rect 19715 310805 19716 310835
rect 19684 310804 19716 310805
rect 19684 310755 19716 310756
rect 19684 310725 19685 310755
rect 19685 310725 19715 310755
rect 19715 310725 19716 310755
rect 19684 310724 19716 310725
rect 19684 310675 19716 310676
rect 19684 310645 19685 310675
rect 19685 310645 19715 310675
rect 19715 310645 19716 310675
rect 19684 310644 19716 310645
rect 19684 310595 19716 310596
rect 19684 310565 19685 310595
rect 19685 310565 19715 310595
rect 19715 310565 19716 310595
rect 19684 310564 19716 310565
rect 19684 310515 19716 310516
rect 19684 310485 19685 310515
rect 19685 310485 19715 310515
rect 19715 310485 19716 310515
rect 19684 310484 19716 310485
rect 19684 310435 19716 310436
rect 19684 310405 19685 310435
rect 19685 310405 19715 310435
rect 19715 310405 19716 310435
rect 19684 310404 19716 310405
rect 19684 310355 19716 310356
rect 19684 310325 19685 310355
rect 19685 310325 19715 310355
rect 19715 310325 19716 310355
rect 19684 310324 19716 310325
rect 19684 310275 19716 310276
rect 19684 310245 19685 310275
rect 19685 310245 19715 310275
rect 19715 310245 19716 310275
rect 19684 310244 19716 310245
rect 19684 310195 19716 310196
rect 19684 310165 19685 310195
rect 19685 310165 19715 310195
rect 19715 310165 19716 310195
rect 19684 310164 19716 310165
rect 19684 310115 19716 310116
rect 19684 310085 19685 310115
rect 19685 310085 19715 310115
rect 19715 310085 19716 310115
rect 19684 310084 19716 310085
rect 19684 310035 19716 310036
rect 19684 310005 19685 310035
rect 19685 310005 19715 310035
rect 19715 310005 19716 310035
rect 19684 310004 19716 310005
rect 19684 309955 19716 309956
rect 19684 309925 19685 309955
rect 19685 309925 19715 309955
rect 19715 309925 19716 309955
rect 19684 309924 19716 309925
rect 19684 309875 19716 309876
rect 19684 309845 19685 309875
rect 19685 309845 19715 309875
rect 19715 309845 19716 309875
rect 19684 309844 19716 309845
rect 19684 309795 19716 309796
rect 19684 309765 19685 309795
rect 19685 309765 19715 309795
rect 19715 309765 19716 309795
rect 19684 309764 19716 309765
rect 19684 309715 19716 309716
rect 19684 309685 19685 309715
rect 19685 309685 19715 309715
rect 19715 309685 19716 309715
rect 19684 309684 19716 309685
rect 19684 309635 19716 309636
rect 19684 309605 19685 309635
rect 19685 309605 19715 309635
rect 19715 309605 19716 309635
rect 19684 309604 19716 309605
rect 19684 309555 19716 309556
rect 19684 309525 19685 309555
rect 19685 309525 19715 309555
rect 19715 309525 19716 309555
rect 19684 309524 19716 309525
rect 19684 309475 19716 309476
rect 19684 309445 19685 309475
rect 19685 309445 19715 309475
rect 19715 309445 19716 309475
rect 19684 309444 19716 309445
rect 19684 309395 19716 309396
rect 19684 309365 19685 309395
rect 19685 309365 19715 309395
rect 19715 309365 19716 309395
rect 19684 309364 19716 309365
rect 19684 309315 19716 309316
rect 19684 309285 19685 309315
rect 19685 309285 19715 309315
rect 19715 309285 19716 309315
rect 19684 309284 19716 309285
rect 19684 309235 19716 309236
rect 19684 309205 19685 309235
rect 19685 309205 19715 309235
rect 19715 309205 19716 309235
rect 19684 309204 19716 309205
rect 19684 309155 19716 309156
rect 19684 309125 19685 309155
rect 19685 309125 19715 309155
rect 19715 309125 19716 309155
rect 19684 309124 19716 309125
rect 19684 309075 19716 309076
rect 19684 309045 19685 309075
rect 19685 309045 19715 309075
rect 19715 309045 19716 309075
rect 19684 309044 19716 309045
rect 19684 308995 19716 308996
rect 19684 308965 19685 308995
rect 19685 308965 19715 308995
rect 19715 308965 19716 308995
rect 19684 308964 19716 308965
rect 19684 308915 19716 308916
rect 19684 308885 19685 308915
rect 19685 308885 19715 308915
rect 19715 308885 19716 308915
rect 19684 308884 19716 308885
rect 19684 308835 19716 308836
rect 19684 308805 19685 308835
rect 19685 308805 19715 308835
rect 19715 308805 19716 308835
rect 19684 308804 19716 308805
rect 19684 308755 19716 308756
rect 19684 308725 19685 308755
rect 19685 308725 19715 308755
rect 19715 308725 19716 308755
rect 19684 308724 19716 308725
rect 19684 308675 19716 308676
rect 19684 308645 19685 308675
rect 19685 308645 19715 308675
rect 19715 308645 19716 308675
rect 19684 308644 19716 308645
rect 19684 308595 19716 308596
rect 19684 308565 19685 308595
rect 19685 308565 19715 308595
rect 19715 308565 19716 308595
rect 19684 308564 19716 308565
rect 19684 308515 19716 308516
rect 19684 308485 19685 308515
rect 19685 308485 19715 308515
rect 19715 308485 19716 308515
rect 19684 308484 19716 308485
rect 19684 308435 19716 308436
rect 19684 308405 19685 308435
rect 19685 308405 19715 308435
rect 19715 308405 19716 308435
rect 19684 308404 19716 308405
rect 19684 308355 19716 308356
rect 19684 308325 19685 308355
rect 19685 308325 19715 308355
rect 19715 308325 19716 308355
rect 19684 308324 19716 308325
rect 19684 308275 19716 308276
rect 19684 308245 19685 308275
rect 19685 308245 19715 308275
rect 19715 308245 19716 308275
rect 19684 308244 19716 308245
rect 19684 308195 19716 308196
rect 19684 308165 19685 308195
rect 19685 308165 19715 308195
rect 19715 308165 19716 308195
rect 19684 308164 19716 308165
rect 19684 308115 19716 308116
rect 19684 308085 19685 308115
rect 19685 308085 19715 308115
rect 19715 308085 19716 308115
rect 19684 308084 19716 308085
rect 19684 308035 19716 308036
rect 19684 308005 19685 308035
rect 19685 308005 19715 308035
rect 19715 308005 19716 308035
rect 19684 308004 19716 308005
rect 19684 307955 19716 307956
rect 19684 307925 19685 307955
rect 19685 307925 19715 307955
rect 19715 307925 19716 307955
rect 19684 307924 19716 307925
rect 19684 307875 19716 307876
rect 19684 307845 19685 307875
rect 19685 307845 19715 307875
rect 19715 307845 19716 307875
rect 19684 307844 19716 307845
rect 19684 307795 19716 307796
rect 19684 307765 19685 307795
rect 19685 307765 19715 307795
rect 19715 307765 19716 307795
rect 19684 307764 19716 307765
rect 19684 307715 19716 307716
rect 19684 307685 19685 307715
rect 19685 307685 19715 307715
rect 19715 307685 19716 307715
rect 19684 307684 19716 307685
rect 19684 307635 19716 307636
rect 19684 307605 19685 307635
rect 19685 307605 19715 307635
rect 19715 307605 19716 307635
rect 19684 307604 19716 307605
rect 19684 307555 19716 307556
rect 19684 307525 19685 307555
rect 19685 307525 19715 307555
rect 19715 307525 19716 307555
rect 19684 307524 19716 307525
rect 19684 307475 19716 307476
rect 19684 307445 19685 307475
rect 19685 307445 19715 307475
rect 19715 307445 19716 307475
rect 19684 307444 19716 307445
rect 19684 307395 19716 307396
rect 19684 307365 19685 307395
rect 19685 307365 19715 307395
rect 19715 307365 19716 307395
rect 19684 307364 19716 307365
rect 19684 307315 19716 307316
rect 19684 307285 19685 307315
rect 19685 307285 19715 307315
rect 19715 307285 19716 307315
rect 19684 307284 19716 307285
rect 19684 307235 19716 307236
rect 19684 307205 19685 307235
rect 19685 307205 19715 307235
rect 19715 307205 19716 307235
rect 19684 307204 19716 307205
rect 19684 307155 19716 307156
rect 19684 307125 19685 307155
rect 19685 307125 19715 307155
rect 19715 307125 19716 307155
rect 19684 307124 19716 307125
rect 19684 307075 19716 307076
rect 19684 307045 19685 307075
rect 19685 307045 19715 307075
rect 19715 307045 19716 307075
rect 19684 307044 19716 307045
rect 19684 306995 19716 306996
rect 19684 306965 19685 306995
rect 19685 306965 19715 306995
rect 19715 306965 19716 306995
rect 19684 306964 19716 306965
rect 19684 306915 19716 306916
rect 19684 306885 19685 306915
rect 19685 306885 19715 306915
rect 19715 306885 19716 306915
rect 19684 306884 19716 306885
rect 19684 306835 19716 306836
rect 19684 306805 19685 306835
rect 19685 306805 19715 306835
rect 19715 306805 19716 306835
rect 19684 306804 19716 306805
rect 19684 306755 19716 306756
rect 19684 306725 19685 306755
rect 19685 306725 19715 306755
rect 19715 306725 19716 306755
rect 19684 306724 19716 306725
rect 19684 306675 19716 306676
rect 19684 306645 19685 306675
rect 19685 306645 19715 306675
rect 19715 306645 19716 306675
rect 19684 306644 19716 306645
rect 19684 306595 19716 306596
rect 19684 306565 19685 306595
rect 19685 306565 19715 306595
rect 19715 306565 19716 306595
rect 19684 306564 19716 306565
rect 19684 306515 19716 306516
rect 19684 306485 19685 306515
rect 19685 306485 19715 306515
rect 19715 306485 19716 306515
rect 19684 306484 19716 306485
rect 19684 306435 19716 306436
rect 19684 306405 19685 306435
rect 19685 306405 19715 306435
rect 19715 306405 19716 306435
rect 19684 306404 19716 306405
rect 19684 306355 19716 306356
rect 19684 306325 19685 306355
rect 19685 306325 19715 306355
rect 19715 306325 19716 306355
rect 19684 306324 19716 306325
rect 19684 306275 19716 306276
rect 19684 306245 19685 306275
rect 19685 306245 19715 306275
rect 19715 306245 19716 306275
rect 19684 306244 19716 306245
rect 19684 306195 19716 306196
rect 19684 306165 19685 306195
rect 19685 306165 19715 306195
rect 19715 306165 19716 306195
rect 19684 306164 19716 306165
rect 19684 306115 19716 306116
rect 19684 306085 19685 306115
rect 19685 306085 19715 306115
rect 19715 306085 19716 306115
rect 19684 306084 19716 306085
rect 19684 306035 19716 306036
rect 19684 306005 19685 306035
rect 19685 306005 19715 306035
rect 19715 306005 19716 306035
rect 19684 306004 19716 306005
rect 19684 305955 19716 305956
rect 19684 305925 19685 305955
rect 19685 305925 19715 305955
rect 19715 305925 19716 305955
rect 19684 305924 19716 305925
rect 19684 305875 19716 305876
rect 19684 305845 19685 305875
rect 19685 305845 19715 305875
rect 19715 305845 19716 305875
rect 19684 305844 19716 305845
rect 19684 305795 19716 305796
rect 19684 305765 19685 305795
rect 19685 305765 19715 305795
rect 19715 305765 19716 305795
rect 19684 305764 19716 305765
rect 19684 305715 19716 305716
rect 19684 305685 19685 305715
rect 19685 305685 19715 305715
rect 19715 305685 19716 305715
rect 19684 305684 19716 305685
rect 19684 305635 19716 305636
rect 19684 305605 19685 305635
rect 19685 305605 19715 305635
rect 19715 305605 19716 305635
rect 19684 305604 19716 305605
rect 19684 305555 19716 305556
rect 19684 305525 19685 305555
rect 19685 305525 19715 305555
rect 19715 305525 19716 305555
rect 19684 305524 19716 305525
rect 19684 305475 19716 305476
rect 19684 305445 19685 305475
rect 19685 305445 19715 305475
rect 19715 305445 19716 305475
rect 19684 305444 19716 305445
rect 19684 305395 19716 305396
rect 19684 305365 19685 305395
rect 19685 305365 19715 305395
rect 19715 305365 19716 305395
rect 19684 305364 19716 305365
rect 19684 305315 19716 305316
rect 19684 305285 19685 305315
rect 19685 305285 19715 305315
rect 19715 305285 19716 305315
rect 19684 305284 19716 305285
rect 19684 305235 19716 305236
rect 19684 305205 19685 305235
rect 19685 305205 19715 305235
rect 19715 305205 19716 305235
rect 19684 305204 19716 305205
rect 19684 305155 19716 305156
rect 19684 305125 19685 305155
rect 19685 305125 19715 305155
rect 19715 305125 19716 305155
rect 19684 305124 19716 305125
rect 19684 305075 19716 305076
rect 19684 305045 19685 305075
rect 19685 305045 19715 305075
rect 19715 305045 19716 305075
rect 19684 305044 19716 305045
rect 19684 304995 19716 304996
rect 19684 304965 19685 304995
rect 19685 304965 19715 304995
rect 19715 304965 19716 304995
rect 19684 304964 19716 304965
rect 19684 304915 19716 304916
rect 19684 304885 19685 304915
rect 19685 304885 19715 304915
rect 19715 304885 19716 304915
rect 19684 304884 19716 304885
rect 19684 304835 19716 304836
rect 19684 304805 19685 304835
rect 19685 304805 19715 304835
rect 19715 304805 19716 304835
rect 19684 304804 19716 304805
rect 19684 304755 19716 304756
rect 19684 304725 19685 304755
rect 19685 304725 19715 304755
rect 19715 304725 19716 304755
rect 19684 304724 19716 304725
rect 19684 304675 19716 304676
rect 19684 304645 19685 304675
rect 19685 304645 19715 304675
rect 19715 304645 19716 304675
rect 19684 304644 19716 304645
rect 19684 304595 19716 304596
rect 19684 304565 19685 304595
rect 19685 304565 19715 304595
rect 19715 304565 19716 304595
rect 19684 304564 19716 304565
rect 19684 304515 19716 304516
rect 19684 304485 19685 304515
rect 19685 304485 19715 304515
rect 19715 304485 19716 304515
rect 19684 304484 19716 304485
rect 19684 304435 19716 304436
rect 19684 304405 19685 304435
rect 19685 304405 19715 304435
rect 19715 304405 19716 304435
rect 19684 304404 19716 304405
rect 19684 304355 19716 304356
rect 19684 304325 19685 304355
rect 19685 304325 19715 304355
rect 19715 304325 19716 304355
rect 19684 304324 19716 304325
rect 19684 304275 19716 304276
rect 19684 304245 19685 304275
rect 19685 304245 19715 304275
rect 19715 304245 19716 304275
rect 19684 304244 19716 304245
rect 19684 304195 19716 304196
rect 19684 304165 19685 304195
rect 19685 304165 19715 304195
rect 19715 304165 19716 304195
rect 19684 304164 19716 304165
rect 19684 304115 19716 304116
rect 19684 304085 19685 304115
rect 19685 304085 19715 304115
rect 19715 304085 19716 304115
rect 19684 304084 19716 304085
rect 19684 304035 19716 304036
rect 19684 304005 19685 304035
rect 19685 304005 19715 304035
rect 19715 304005 19716 304035
rect 19684 304004 19716 304005
rect 19684 303955 19716 303956
rect 19684 303925 19685 303955
rect 19685 303925 19715 303955
rect 19715 303925 19716 303955
rect 19684 303924 19716 303925
rect 19684 303875 19716 303876
rect 19684 303845 19685 303875
rect 19685 303845 19715 303875
rect 19715 303845 19716 303875
rect 19684 303844 19716 303845
rect 19684 303795 19716 303796
rect 19684 303765 19685 303795
rect 19685 303765 19715 303795
rect 19715 303765 19716 303795
rect 19684 303764 19716 303765
rect 19684 303715 19716 303716
rect 19684 303685 19685 303715
rect 19685 303685 19715 303715
rect 19715 303685 19716 303715
rect 19684 303684 19716 303685
rect 19684 303635 19716 303636
rect 19684 303605 19685 303635
rect 19685 303605 19715 303635
rect 19715 303605 19716 303635
rect 19684 303604 19716 303605
rect 19684 303555 19716 303556
rect 19684 303525 19685 303555
rect 19685 303525 19715 303555
rect 19715 303525 19716 303555
rect 19684 303524 19716 303525
rect 19684 303475 19716 303476
rect 19684 303445 19685 303475
rect 19685 303445 19715 303475
rect 19715 303445 19716 303475
rect 19684 303444 19716 303445
rect 19684 303395 19716 303396
rect 19684 303365 19685 303395
rect 19685 303365 19715 303395
rect 19715 303365 19716 303395
rect 19684 303364 19716 303365
rect 19684 303315 19716 303316
rect 19684 303285 19685 303315
rect 19685 303285 19715 303315
rect 19715 303285 19716 303315
rect 19684 303284 19716 303285
rect 19684 303235 19716 303236
rect 19684 303205 19685 303235
rect 19685 303205 19715 303235
rect 19715 303205 19716 303235
rect 19684 303204 19716 303205
rect 19684 303155 19716 303156
rect 19684 303125 19685 303155
rect 19685 303125 19715 303155
rect 19715 303125 19716 303155
rect 19684 303124 19716 303125
rect 19684 303075 19716 303076
rect 19684 303045 19685 303075
rect 19685 303045 19715 303075
rect 19715 303045 19716 303075
rect 19684 303044 19716 303045
rect 19684 302995 19716 302996
rect 19684 302965 19685 302995
rect 19685 302965 19715 302995
rect 19715 302965 19716 302995
rect 19684 302964 19716 302965
rect 19684 302915 19716 302916
rect 19684 302885 19685 302915
rect 19685 302885 19715 302915
rect 19715 302885 19716 302915
rect 19684 302884 19716 302885
rect 19684 302835 19716 302836
rect 19684 302805 19685 302835
rect 19685 302805 19715 302835
rect 19715 302805 19716 302835
rect 19684 302804 19716 302805
rect 19684 302755 19716 302756
rect 19684 302725 19685 302755
rect 19685 302725 19715 302755
rect 19715 302725 19716 302755
rect 19684 302724 19716 302725
rect 19684 302675 19716 302676
rect 19684 302645 19685 302675
rect 19685 302645 19715 302675
rect 19715 302645 19716 302675
rect 19684 302644 19716 302645
rect 19684 302595 19716 302596
rect 19684 302565 19685 302595
rect 19685 302565 19715 302595
rect 19715 302565 19716 302595
rect 19684 302564 19716 302565
rect 19684 302515 19716 302516
rect 19684 302485 19685 302515
rect 19685 302485 19715 302515
rect 19715 302485 19716 302515
rect 19684 302484 19716 302485
rect 19684 302435 19716 302436
rect 19684 302405 19685 302435
rect 19685 302405 19715 302435
rect 19715 302405 19716 302435
rect 19684 302404 19716 302405
rect 19684 302355 19716 302356
rect 19684 302325 19685 302355
rect 19685 302325 19715 302355
rect 19715 302325 19716 302355
rect 19684 302324 19716 302325
rect 19684 302275 19716 302276
rect 19684 302245 19685 302275
rect 19685 302245 19715 302275
rect 19715 302245 19716 302275
rect 19684 302244 19716 302245
rect 19684 302195 19716 302196
rect 19684 302165 19685 302195
rect 19685 302165 19715 302195
rect 19715 302165 19716 302195
rect 19684 302164 19716 302165
rect 19684 302115 19716 302116
rect 19684 302085 19685 302115
rect 19685 302085 19715 302115
rect 19715 302085 19716 302115
rect 19684 302084 19716 302085
rect 19684 302035 19716 302036
rect 19684 302005 19685 302035
rect 19685 302005 19715 302035
rect 19715 302005 19716 302035
rect 19684 302004 19716 302005
rect 19684 301955 19716 301956
rect 19684 301925 19685 301955
rect 19685 301925 19715 301955
rect 19715 301925 19716 301955
rect 19684 301924 19716 301925
rect 19684 301875 19716 301876
rect 19684 301845 19685 301875
rect 19685 301845 19715 301875
rect 19715 301845 19716 301875
rect 19684 301844 19716 301845
rect 19684 301795 19716 301796
rect 19684 301765 19685 301795
rect 19685 301765 19715 301795
rect 19715 301765 19716 301795
rect 19684 301764 19716 301765
rect 19684 301715 19716 301716
rect 19684 301685 19685 301715
rect 19685 301685 19715 301715
rect 19715 301685 19716 301715
rect 19684 301684 19716 301685
rect 19684 301635 19716 301636
rect 19684 301605 19685 301635
rect 19685 301605 19715 301635
rect 19715 301605 19716 301635
rect 19684 301604 19716 301605
rect 19684 301555 19716 301556
rect 19684 301525 19685 301555
rect 19685 301525 19715 301555
rect 19715 301525 19716 301555
rect 19684 301524 19716 301525
rect 19684 301475 19716 301476
rect 19684 301445 19685 301475
rect 19685 301445 19715 301475
rect 19715 301445 19716 301475
rect 19684 301444 19716 301445
rect 19684 301395 19716 301396
rect 19684 301365 19685 301395
rect 19685 301365 19715 301395
rect 19715 301365 19716 301395
rect 19684 301364 19716 301365
rect 19684 301315 19716 301316
rect 19684 301285 19685 301315
rect 19685 301285 19715 301315
rect 19715 301285 19716 301315
rect 19684 301284 19716 301285
rect 19684 301235 19716 301236
rect 19684 301205 19685 301235
rect 19685 301205 19715 301235
rect 19715 301205 19716 301235
rect 19684 301204 19716 301205
rect 19684 301155 19716 301156
rect 19684 301125 19685 301155
rect 19685 301125 19715 301155
rect 19715 301125 19716 301155
rect 19684 301124 19716 301125
rect 19684 301075 19716 301076
rect 19684 301045 19685 301075
rect 19685 301045 19715 301075
rect 19715 301045 19716 301075
rect 19684 301044 19716 301045
rect 19684 300995 19716 300996
rect 19684 300965 19685 300995
rect 19685 300965 19715 300995
rect 19715 300965 19716 300995
rect 19684 300964 19716 300965
rect 19684 300915 19716 300916
rect 19684 300885 19685 300915
rect 19685 300885 19715 300915
rect 19715 300885 19716 300915
rect 19684 300884 19716 300885
rect 19684 300835 19716 300836
rect 19684 300805 19685 300835
rect 19685 300805 19715 300835
rect 19715 300805 19716 300835
rect 19684 300804 19716 300805
rect 19684 300755 19716 300756
rect 19684 300725 19685 300755
rect 19685 300725 19715 300755
rect 19715 300725 19716 300755
rect 19684 300724 19716 300725
rect 19684 300675 19716 300676
rect 19684 300645 19685 300675
rect 19685 300645 19715 300675
rect 19715 300645 19716 300675
rect 19684 300644 19716 300645
rect 19684 300595 19716 300596
rect 19684 300565 19685 300595
rect 19685 300565 19715 300595
rect 19715 300565 19716 300595
rect 19684 300564 19716 300565
rect 19684 300515 19716 300516
rect 19684 300485 19685 300515
rect 19685 300485 19715 300515
rect 19715 300485 19716 300515
rect 19684 300484 19716 300485
rect 19684 300435 19716 300436
rect 19684 300405 19685 300435
rect 19685 300405 19715 300435
rect 19715 300405 19716 300435
rect 19684 300404 19716 300405
rect 19684 300355 19716 300356
rect 19684 300325 19685 300355
rect 19685 300325 19715 300355
rect 19715 300325 19716 300355
rect 19684 300324 19716 300325
rect 19684 300275 19716 300276
rect 19684 300245 19685 300275
rect 19685 300245 19715 300275
rect 19715 300245 19716 300275
rect 19684 300244 19716 300245
rect 19684 300195 19716 300196
rect 19684 300165 19685 300195
rect 19685 300165 19715 300195
rect 19715 300165 19716 300195
rect 19684 300164 19716 300165
rect 19684 300115 19716 300116
rect 19684 300085 19685 300115
rect 19685 300085 19715 300115
rect 19715 300085 19716 300115
rect 19684 300084 19716 300085
rect 19684 300035 19716 300036
rect 19684 300005 19685 300035
rect 19685 300005 19715 300035
rect 19715 300005 19716 300035
rect 19684 300004 19716 300005
rect 19684 299955 19716 299956
rect 19684 299925 19685 299955
rect 19685 299925 19715 299955
rect 19715 299925 19716 299955
rect 19684 299924 19716 299925
rect 19684 299875 19716 299876
rect 19684 299845 19685 299875
rect 19685 299845 19715 299875
rect 19715 299845 19716 299875
rect 19684 299844 19716 299845
rect 19684 299795 19716 299796
rect 19684 299765 19685 299795
rect 19685 299765 19715 299795
rect 19715 299765 19716 299795
rect 19684 299764 19716 299765
rect 19684 299715 19716 299716
rect 19684 299685 19685 299715
rect 19685 299685 19715 299715
rect 19715 299685 19716 299715
rect 19684 299684 19716 299685
rect 19684 299635 19716 299636
rect 19684 299605 19685 299635
rect 19685 299605 19715 299635
rect 19715 299605 19716 299635
rect 19684 299604 19716 299605
rect 19684 299555 19716 299556
rect 19684 299525 19685 299555
rect 19685 299525 19715 299555
rect 19715 299525 19716 299555
rect 19684 299524 19716 299525
rect 19684 299475 19716 299476
rect 19684 299445 19685 299475
rect 19685 299445 19715 299475
rect 19715 299445 19716 299475
rect 19684 299444 19716 299445
rect 19684 299395 19716 299396
rect 19684 299365 19685 299395
rect 19685 299365 19715 299395
rect 19715 299365 19716 299395
rect 19684 299364 19716 299365
rect 19684 299315 19716 299316
rect 19684 299285 19685 299315
rect 19685 299285 19715 299315
rect 19715 299285 19716 299315
rect 19684 299284 19716 299285
rect 19684 299235 19716 299236
rect 19684 299205 19685 299235
rect 19685 299205 19715 299235
rect 19715 299205 19716 299235
rect 19684 299204 19716 299205
rect 19684 299155 19716 299156
rect 19684 299125 19685 299155
rect 19685 299125 19715 299155
rect 19715 299125 19716 299155
rect 19684 299124 19716 299125
rect 19684 299075 19716 299076
rect 19684 299045 19685 299075
rect 19685 299045 19715 299075
rect 19715 299045 19716 299075
rect 19684 299044 19716 299045
rect 19684 298995 19716 298996
rect 19684 298965 19685 298995
rect 19685 298965 19715 298995
rect 19715 298965 19716 298995
rect 19684 298964 19716 298965
rect 19684 298915 19716 298916
rect 19684 298885 19685 298915
rect 19685 298885 19715 298915
rect 19715 298885 19716 298915
rect 19684 298884 19716 298885
rect 19684 298835 19716 298836
rect 19684 298805 19685 298835
rect 19685 298805 19715 298835
rect 19715 298805 19716 298835
rect 19684 298804 19716 298805
rect 19684 298755 19716 298756
rect 19684 298725 19685 298755
rect 19685 298725 19715 298755
rect 19715 298725 19716 298755
rect 19684 298724 19716 298725
rect 19684 298675 19716 298676
rect 19684 298645 19685 298675
rect 19685 298645 19715 298675
rect 19715 298645 19716 298675
rect 19684 298644 19716 298645
rect 19684 298595 19716 298596
rect 19684 298565 19685 298595
rect 19685 298565 19715 298595
rect 19715 298565 19716 298595
rect 19684 298564 19716 298565
rect 19684 298515 19716 298516
rect 19684 298485 19685 298515
rect 19685 298485 19715 298515
rect 19715 298485 19716 298515
rect 19684 298484 19716 298485
rect 19684 298435 19716 298436
rect 19684 298405 19685 298435
rect 19685 298405 19715 298435
rect 19715 298405 19716 298435
rect 19684 298404 19716 298405
rect 19684 298355 19716 298356
rect 19684 298325 19685 298355
rect 19685 298325 19715 298355
rect 19715 298325 19716 298355
rect 19684 298324 19716 298325
rect 19684 298275 19716 298276
rect 19684 298245 19685 298275
rect 19685 298245 19715 298275
rect 19715 298245 19716 298275
rect 19684 298244 19716 298245
rect 19684 298195 19716 298196
rect 19684 298165 19685 298195
rect 19685 298165 19715 298195
rect 19715 298165 19716 298195
rect 19684 298164 19716 298165
rect 19684 298115 19716 298116
rect 19684 298085 19685 298115
rect 19685 298085 19715 298115
rect 19715 298085 19716 298115
rect 19684 298084 19716 298085
rect 19684 298035 19716 298036
rect 19684 298005 19685 298035
rect 19685 298005 19715 298035
rect 19715 298005 19716 298035
rect 19684 298004 19716 298005
rect 19684 297955 19716 297956
rect 19684 297925 19685 297955
rect 19685 297925 19715 297955
rect 19715 297925 19716 297955
rect 19684 297924 19716 297925
rect 19684 297875 19716 297876
rect 19684 297845 19685 297875
rect 19685 297845 19715 297875
rect 19715 297845 19716 297875
rect 19684 297844 19716 297845
rect 19684 297795 19716 297796
rect 19684 297765 19685 297795
rect 19685 297765 19715 297795
rect 19715 297765 19716 297795
rect 19684 297764 19716 297765
rect 19684 297715 19716 297716
rect 19684 297685 19685 297715
rect 19685 297685 19715 297715
rect 19715 297685 19716 297715
rect 19684 297684 19716 297685
rect 19684 297635 19716 297636
rect 19684 297605 19685 297635
rect 19685 297605 19715 297635
rect 19715 297605 19716 297635
rect 19684 297604 19716 297605
rect 19684 297555 19716 297556
rect 19684 297525 19685 297555
rect 19685 297525 19715 297555
rect 19715 297525 19716 297555
rect 19684 297524 19716 297525
rect 19684 297475 19716 297476
rect 19684 297445 19685 297475
rect 19685 297445 19715 297475
rect 19715 297445 19716 297475
rect 19684 297444 19716 297445
rect 19684 297395 19716 297396
rect 19684 297365 19685 297395
rect 19685 297365 19715 297395
rect 19715 297365 19716 297395
rect 19684 297364 19716 297365
rect 19684 297315 19716 297316
rect 19684 297285 19685 297315
rect 19685 297285 19715 297315
rect 19715 297285 19716 297315
rect 19684 297284 19716 297285
rect 19684 297235 19716 297236
rect 19684 297205 19685 297235
rect 19685 297205 19715 297235
rect 19715 297205 19716 297235
rect 19684 297204 19716 297205
rect 19684 297155 19716 297156
rect 19684 297125 19685 297155
rect 19685 297125 19715 297155
rect 19715 297125 19716 297155
rect 19684 297124 19716 297125
rect 19684 297075 19716 297076
rect 19684 297045 19685 297075
rect 19685 297045 19715 297075
rect 19715 297045 19716 297075
rect 19684 297044 19716 297045
rect 19684 296995 19716 296996
rect 19684 296965 19685 296995
rect 19685 296965 19715 296995
rect 19715 296965 19716 296995
rect 19684 296964 19716 296965
rect 19684 296915 19716 296916
rect 19684 296885 19685 296915
rect 19685 296885 19715 296915
rect 19715 296885 19716 296915
rect 19684 296884 19716 296885
rect 19684 296835 19716 296836
rect 19684 296805 19685 296835
rect 19685 296805 19715 296835
rect 19715 296805 19716 296835
rect 19684 296804 19716 296805
rect 19684 296755 19716 296756
rect 19684 296725 19685 296755
rect 19685 296725 19715 296755
rect 19715 296725 19716 296755
rect 19684 296724 19716 296725
rect 19684 296675 19716 296676
rect 19684 296645 19685 296675
rect 19685 296645 19715 296675
rect 19715 296645 19716 296675
rect 19684 296644 19716 296645
rect 19684 296595 19716 296596
rect 19684 296565 19685 296595
rect 19685 296565 19715 296595
rect 19715 296565 19716 296595
rect 19684 296564 19716 296565
rect 19684 296515 19716 296516
rect 19684 296485 19685 296515
rect 19685 296485 19715 296515
rect 19715 296485 19716 296515
rect 19684 296484 19716 296485
rect 19684 296435 19716 296436
rect 19684 296405 19685 296435
rect 19685 296405 19715 296435
rect 19715 296405 19716 296435
rect 19684 296404 19716 296405
rect 19684 296355 19716 296356
rect 19684 296325 19685 296355
rect 19685 296325 19715 296355
rect 19715 296325 19716 296355
rect 19684 296324 19716 296325
rect 19684 296275 19716 296276
rect 19684 296245 19685 296275
rect 19685 296245 19715 296275
rect 19715 296245 19716 296275
rect 19684 296244 19716 296245
rect 19684 296195 19716 296196
rect 19684 296165 19685 296195
rect 19685 296165 19715 296195
rect 19715 296165 19716 296195
rect 19684 296164 19716 296165
rect 19684 296115 19716 296116
rect 19684 296085 19685 296115
rect 19685 296085 19715 296115
rect 19715 296085 19716 296115
rect 19684 296084 19716 296085
rect 19684 296035 19716 296036
rect 19684 296005 19685 296035
rect 19685 296005 19715 296035
rect 19715 296005 19716 296035
rect 19684 296004 19716 296005
rect 19684 295955 19716 295956
rect 19684 295925 19685 295955
rect 19685 295925 19715 295955
rect 19715 295925 19716 295955
rect 19684 295924 19716 295925
rect 19684 295875 19716 295876
rect 19684 295845 19685 295875
rect 19685 295845 19715 295875
rect 19715 295845 19716 295875
rect 19684 295844 19716 295845
rect 19684 295795 19716 295796
rect 19684 295765 19685 295795
rect 19685 295765 19715 295795
rect 19715 295765 19716 295795
rect 19684 295764 19716 295765
rect 19684 295715 19716 295716
rect 19684 295685 19685 295715
rect 19685 295685 19715 295715
rect 19715 295685 19716 295715
rect 19684 295684 19716 295685
rect 19684 295635 19716 295636
rect 19684 295605 19685 295635
rect 19685 295605 19715 295635
rect 19715 295605 19716 295635
rect 19684 295604 19716 295605
rect 19684 295555 19716 295556
rect 19684 295525 19685 295555
rect 19685 295525 19715 295555
rect 19715 295525 19716 295555
rect 19684 295524 19716 295525
rect 19684 295475 19716 295476
rect 19684 295445 19685 295475
rect 19685 295445 19715 295475
rect 19715 295445 19716 295475
rect 19684 295444 19716 295445
rect 19684 295395 19716 295396
rect 19684 295365 19685 295395
rect 19685 295365 19715 295395
rect 19715 295365 19716 295395
rect 19684 295364 19716 295365
rect 19684 295315 19716 295316
rect 19684 295285 19685 295315
rect 19685 295285 19715 295315
rect 19715 295285 19716 295315
rect 19684 295284 19716 295285
rect 19684 295235 19716 295236
rect 19684 295205 19685 295235
rect 19685 295205 19715 295235
rect 19715 295205 19716 295235
rect 19684 295204 19716 295205
rect 19684 295155 19716 295156
rect 19684 295125 19685 295155
rect 19685 295125 19715 295155
rect 19715 295125 19716 295155
rect 19684 295124 19716 295125
rect 19684 295075 19716 295076
rect 19684 295045 19685 295075
rect 19685 295045 19715 295075
rect 19715 295045 19716 295075
rect 19684 295044 19716 295045
rect 19684 294995 19716 294996
rect 19684 294965 19685 294995
rect 19685 294965 19715 294995
rect 19715 294965 19716 294995
rect 19684 294964 19716 294965
rect 19684 294915 19716 294916
rect 19684 294885 19685 294915
rect 19685 294885 19715 294915
rect 19715 294885 19716 294915
rect 19684 294884 19716 294885
rect 19684 294835 19716 294836
rect 19684 294805 19685 294835
rect 19685 294805 19715 294835
rect 19715 294805 19716 294835
rect 19684 294804 19716 294805
rect 19684 294755 19716 294756
rect 19684 294725 19685 294755
rect 19685 294725 19715 294755
rect 19715 294725 19716 294755
rect 19684 294724 19716 294725
rect 19684 294675 19716 294676
rect 19684 294645 19685 294675
rect 19685 294645 19715 294675
rect 19715 294645 19716 294675
rect 19684 294644 19716 294645
rect 19684 294595 19716 294596
rect 19684 294565 19685 294595
rect 19685 294565 19715 294595
rect 19715 294565 19716 294595
rect 19684 294564 19716 294565
rect 19684 294515 19716 294516
rect 19684 294485 19685 294515
rect 19685 294485 19715 294515
rect 19715 294485 19716 294515
rect 19684 294484 19716 294485
rect 19684 294435 19716 294436
rect 19684 294405 19685 294435
rect 19685 294405 19715 294435
rect 19715 294405 19716 294435
rect 19684 294404 19716 294405
rect 19684 294355 19716 294356
rect 19684 294325 19685 294355
rect 19685 294325 19715 294355
rect 19715 294325 19716 294355
rect 19684 294324 19716 294325
rect 19684 294275 19716 294276
rect 19684 294245 19685 294275
rect 19685 294245 19715 294275
rect 19715 294245 19716 294275
rect 19684 294244 19716 294245
rect 19684 294195 19716 294196
rect 19684 294165 19685 294195
rect 19685 294165 19715 294195
rect 19715 294165 19716 294195
rect 19684 294164 19716 294165
rect 19684 294115 19716 294116
rect 19684 294085 19685 294115
rect 19685 294085 19715 294115
rect 19715 294085 19716 294115
rect 19684 294084 19716 294085
rect 19684 294035 19716 294036
rect 19684 294005 19685 294035
rect 19685 294005 19715 294035
rect 19715 294005 19716 294035
rect 19684 294004 19716 294005
rect 19684 293955 19716 293956
rect 19684 293925 19685 293955
rect 19685 293925 19715 293955
rect 19715 293925 19716 293955
rect 19684 293924 19716 293925
rect 19684 293875 19716 293876
rect 19684 293845 19685 293875
rect 19685 293845 19715 293875
rect 19715 293845 19716 293875
rect 19684 293844 19716 293845
rect 19684 293795 19716 293796
rect 19684 293765 19685 293795
rect 19685 293765 19715 293795
rect 19715 293765 19716 293795
rect 19684 293764 19716 293765
rect 19684 293715 19716 293716
rect 19684 293685 19685 293715
rect 19685 293685 19715 293715
rect 19715 293685 19716 293715
rect 19684 293684 19716 293685
rect 19684 293635 19716 293636
rect 19684 293605 19685 293635
rect 19685 293605 19715 293635
rect 19715 293605 19716 293635
rect 19684 293604 19716 293605
rect 19684 293555 19716 293556
rect 19684 293525 19685 293555
rect 19685 293525 19715 293555
rect 19715 293525 19716 293555
rect 19684 293524 19716 293525
rect 19684 293475 19716 293476
rect 19684 293445 19685 293475
rect 19685 293445 19715 293475
rect 19715 293445 19716 293475
rect 19684 293444 19716 293445
rect 19684 293395 19716 293396
rect 19684 293365 19685 293395
rect 19685 293365 19715 293395
rect 19715 293365 19716 293395
rect 19684 293364 19716 293365
rect 19684 293315 19716 293316
rect 19684 293285 19685 293315
rect 19685 293285 19715 293315
rect 19715 293285 19716 293315
rect 19684 293284 19716 293285
rect 19684 293235 19716 293236
rect 19684 293205 19685 293235
rect 19685 293205 19715 293235
rect 19715 293205 19716 293235
rect 19684 293204 19716 293205
rect 19684 293155 19716 293156
rect 19684 293125 19685 293155
rect 19685 293125 19715 293155
rect 19715 293125 19716 293155
rect 19684 293124 19716 293125
rect 19684 293075 19716 293076
rect 19684 293045 19685 293075
rect 19685 293045 19715 293075
rect 19715 293045 19716 293075
rect 19684 293044 19716 293045
rect 19684 292995 19716 292996
rect 19684 292965 19685 292995
rect 19685 292965 19715 292995
rect 19715 292965 19716 292995
rect 19684 292964 19716 292965
rect 19684 292915 19716 292916
rect 19684 292885 19685 292915
rect 19685 292885 19715 292915
rect 19715 292885 19716 292915
rect 19684 292884 19716 292885
rect 19684 292835 19716 292836
rect 19684 292805 19685 292835
rect 19685 292805 19715 292835
rect 19715 292805 19716 292835
rect 19684 292804 19716 292805
rect 19684 292755 19716 292756
rect 19684 292725 19685 292755
rect 19685 292725 19715 292755
rect 19715 292725 19716 292755
rect 19684 292724 19716 292725
rect 19684 292675 19716 292676
rect 19684 292645 19685 292675
rect 19685 292645 19715 292675
rect 19715 292645 19716 292675
rect 19684 292644 19716 292645
rect 19684 292595 19716 292596
rect 19684 292565 19685 292595
rect 19685 292565 19715 292595
rect 19715 292565 19716 292595
rect 19684 292564 19716 292565
rect 19684 292515 19716 292516
rect 19684 292485 19685 292515
rect 19685 292485 19715 292515
rect 19715 292485 19716 292515
rect 19684 292484 19716 292485
rect 19684 292435 19716 292436
rect 19684 292405 19685 292435
rect 19685 292405 19715 292435
rect 19715 292405 19716 292435
rect 19684 292404 19716 292405
rect 19684 292355 19716 292356
rect 19684 292325 19685 292355
rect 19685 292325 19715 292355
rect 19715 292325 19716 292355
rect 19684 292324 19716 292325
rect 19684 292275 19716 292276
rect 19684 292245 19685 292275
rect 19685 292245 19715 292275
rect 19715 292245 19716 292275
rect 19684 292244 19716 292245
rect 19684 292195 19716 292196
rect 19684 292165 19685 292195
rect 19685 292165 19715 292195
rect 19715 292165 19716 292195
rect 19684 292164 19716 292165
rect 19684 292115 19716 292116
rect 19684 292085 19685 292115
rect 19685 292085 19715 292115
rect 19715 292085 19716 292115
rect 19684 292084 19716 292085
rect 19684 292035 19716 292036
rect 19684 292005 19685 292035
rect 19685 292005 19715 292035
rect 19715 292005 19716 292035
rect 19684 292004 19716 292005
rect 19684 291955 19716 291956
rect 19684 291925 19685 291955
rect 19685 291925 19715 291955
rect 19715 291925 19716 291955
rect 19684 291924 19716 291925
rect 19684 291875 19716 291876
rect 19684 291845 19685 291875
rect 19685 291845 19715 291875
rect 19715 291845 19716 291875
rect 19684 291844 19716 291845
rect 19684 291795 19716 291796
rect 19684 291765 19685 291795
rect 19685 291765 19715 291795
rect 19715 291765 19716 291795
rect 19684 291764 19716 291765
rect 19684 291715 19716 291716
rect 19684 291685 19685 291715
rect 19685 291685 19715 291715
rect 19715 291685 19716 291715
rect 19684 291684 19716 291685
rect 19684 291635 19716 291636
rect 19684 291605 19685 291635
rect 19685 291605 19715 291635
rect 19715 291605 19716 291635
rect 19684 291604 19716 291605
rect 19684 291555 19716 291556
rect 19684 291525 19685 291555
rect 19685 291525 19715 291555
rect 19715 291525 19716 291555
rect 19684 291524 19716 291525
rect 19684 291475 19716 291476
rect 19684 291445 19685 291475
rect 19685 291445 19715 291475
rect 19715 291445 19716 291475
rect 19684 291444 19716 291445
rect 19684 291395 19716 291396
rect 19684 291365 19685 291395
rect 19685 291365 19715 291395
rect 19715 291365 19716 291395
rect 19684 291364 19716 291365
rect 19684 291315 19716 291316
rect 19684 291285 19685 291315
rect 19685 291285 19715 291315
rect 19715 291285 19716 291315
rect 19684 291284 19716 291285
rect 19684 291235 19716 291236
rect 19684 291205 19685 291235
rect 19685 291205 19715 291235
rect 19715 291205 19716 291235
rect 19684 291204 19716 291205
rect 19684 291155 19716 291156
rect 19684 291125 19685 291155
rect 19685 291125 19715 291155
rect 19715 291125 19716 291155
rect 19684 291124 19716 291125
rect 19684 291075 19716 291076
rect 19684 291045 19685 291075
rect 19685 291045 19715 291075
rect 19715 291045 19716 291075
rect 19684 291044 19716 291045
rect 19684 290995 19716 290996
rect 19684 290965 19685 290995
rect 19685 290965 19715 290995
rect 19715 290965 19716 290995
rect 19684 290964 19716 290965
rect 19684 290915 19716 290916
rect 19684 290885 19685 290915
rect 19685 290885 19715 290915
rect 19715 290885 19716 290915
rect 19684 290884 19716 290885
rect 19684 290835 19716 290836
rect 19684 290805 19685 290835
rect 19685 290805 19715 290835
rect 19715 290805 19716 290835
rect 19684 290804 19716 290805
rect 19684 290755 19716 290756
rect 19684 290725 19685 290755
rect 19685 290725 19715 290755
rect 19715 290725 19716 290755
rect 19684 290724 19716 290725
rect 19684 290675 19716 290676
rect 19684 290645 19685 290675
rect 19685 290645 19715 290675
rect 19715 290645 19716 290675
rect 19684 290644 19716 290645
rect 19684 290595 19716 290596
rect 19684 290565 19685 290595
rect 19685 290565 19715 290595
rect 19715 290565 19716 290595
rect 19684 290564 19716 290565
rect 19684 290515 19716 290516
rect 19684 290485 19685 290515
rect 19685 290485 19715 290515
rect 19715 290485 19716 290515
rect 19684 290484 19716 290485
rect 19684 290435 19716 290436
rect 19684 290405 19685 290435
rect 19685 290405 19715 290435
rect 19715 290405 19716 290435
rect 19684 290404 19716 290405
rect 19684 290355 19716 290356
rect 19684 290325 19685 290355
rect 19685 290325 19715 290355
rect 19715 290325 19716 290355
rect 19684 290324 19716 290325
rect 19684 290275 19716 290276
rect 19684 290245 19685 290275
rect 19685 290245 19715 290275
rect 19715 290245 19716 290275
rect 19684 290244 19716 290245
rect 19684 290195 19716 290196
rect 19684 290165 19685 290195
rect 19685 290165 19715 290195
rect 19715 290165 19716 290195
rect 19684 290164 19716 290165
rect 19684 290115 19716 290116
rect 19684 290085 19685 290115
rect 19685 290085 19715 290115
rect 19715 290085 19716 290115
rect 19684 290084 19716 290085
rect 19684 290035 19716 290036
rect 19684 290005 19685 290035
rect 19685 290005 19715 290035
rect 19715 290005 19716 290035
rect 19684 290004 19716 290005
rect 19684 289955 19716 289956
rect 19684 289925 19685 289955
rect 19685 289925 19715 289955
rect 19715 289925 19716 289955
rect 19684 289924 19716 289925
rect 19684 289875 19716 289876
rect 19684 289845 19685 289875
rect 19685 289845 19715 289875
rect 19715 289845 19716 289875
rect 19684 289844 19716 289845
rect 19684 289795 19716 289796
rect 19684 289765 19685 289795
rect 19685 289765 19715 289795
rect 19715 289765 19716 289795
rect 19684 289764 19716 289765
rect 19684 289715 19716 289716
rect 19684 289685 19685 289715
rect 19685 289685 19715 289715
rect 19715 289685 19716 289715
rect 19684 289684 19716 289685
rect 19684 289635 19716 289636
rect 19684 289605 19685 289635
rect 19685 289605 19715 289635
rect 19715 289605 19716 289635
rect 19684 289604 19716 289605
rect 19684 289555 19716 289556
rect 19684 289525 19685 289555
rect 19685 289525 19715 289555
rect 19715 289525 19716 289555
rect 19684 289524 19716 289525
rect 19684 289475 19716 289476
rect 19684 289445 19685 289475
rect 19685 289445 19715 289475
rect 19715 289445 19716 289475
rect 19684 289444 19716 289445
rect 19684 289395 19716 289396
rect 19684 289365 19685 289395
rect 19685 289365 19715 289395
rect 19715 289365 19716 289395
rect 19684 289364 19716 289365
rect 19684 289315 19716 289316
rect 19684 289285 19685 289315
rect 19685 289285 19715 289315
rect 19715 289285 19716 289315
rect 19684 289284 19716 289285
rect 19684 289235 19716 289236
rect 19684 289205 19685 289235
rect 19685 289205 19715 289235
rect 19715 289205 19716 289235
rect 19684 289204 19716 289205
rect 19684 289155 19716 289156
rect 19684 289125 19685 289155
rect 19685 289125 19715 289155
rect 19715 289125 19716 289155
rect 19684 289124 19716 289125
rect 19684 289075 19716 289076
rect 19684 289045 19685 289075
rect 19685 289045 19715 289075
rect 19715 289045 19716 289075
rect 19684 289044 19716 289045
rect 19684 288995 19716 288996
rect 19684 288965 19685 288995
rect 19685 288965 19715 288995
rect 19715 288965 19716 288995
rect 19684 288964 19716 288965
rect 19684 288915 19716 288916
rect 19684 288885 19685 288915
rect 19685 288885 19715 288915
rect 19715 288885 19716 288915
rect 19684 288884 19716 288885
rect 19684 288835 19716 288836
rect 19684 288805 19685 288835
rect 19685 288805 19715 288835
rect 19715 288805 19716 288835
rect 19684 288804 19716 288805
rect 19684 288755 19716 288756
rect 19684 288725 19685 288755
rect 19685 288725 19715 288755
rect 19715 288725 19716 288755
rect 19684 288724 19716 288725
rect 19684 288675 19716 288676
rect 19684 288645 19685 288675
rect 19685 288645 19715 288675
rect 19715 288645 19716 288675
rect 19684 288644 19716 288645
rect 19684 288595 19716 288596
rect 19684 288565 19685 288595
rect 19685 288565 19715 288595
rect 19715 288565 19716 288595
rect 19684 288564 19716 288565
rect 19684 288515 19716 288516
rect 19684 288485 19685 288515
rect 19685 288485 19715 288515
rect 19715 288485 19716 288515
rect 19684 288484 19716 288485
rect 19684 288435 19716 288436
rect 19684 288405 19685 288435
rect 19685 288405 19715 288435
rect 19715 288405 19716 288435
rect 19684 288404 19716 288405
rect 19684 288355 19716 288356
rect 19684 288325 19685 288355
rect 19685 288325 19715 288355
rect 19715 288325 19716 288355
rect 19684 288324 19716 288325
rect 19684 288275 19716 288276
rect 19684 288245 19685 288275
rect 19685 288245 19715 288275
rect 19715 288245 19716 288275
rect 19684 288244 19716 288245
rect 19684 288195 19716 288196
rect 19684 288165 19685 288195
rect 19685 288165 19715 288195
rect 19715 288165 19716 288195
rect 19684 288164 19716 288165
rect 19684 288115 19716 288116
rect 19684 288085 19685 288115
rect 19685 288085 19715 288115
rect 19715 288085 19716 288115
rect 19684 288084 19716 288085
rect 19684 288035 19716 288036
rect 19684 288005 19685 288035
rect 19685 288005 19715 288035
rect 19715 288005 19716 288035
rect 19684 288004 19716 288005
rect 19684 287955 19716 287956
rect 19684 287925 19685 287955
rect 19685 287925 19715 287955
rect 19715 287925 19716 287955
rect 19684 287924 19716 287925
rect 19684 287875 19716 287876
rect 19684 287845 19685 287875
rect 19685 287845 19715 287875
rect 19715 287845 19716 287875
rect 19684 287844 19716 287845
rect 19684 287795 19716 287796
rect 19684 287765 19685 287795
rect 19685 287765 19715 287795
rect 19715 287765 19716 287795
rect 19684 287764 19716 287765
rect 19684 287715 19716 287716
rect 19684 287685 19685 287715
rect 19685 287685 19715 287715
rect 19715 287685 19716 287715
rect 19684 287684 19716 287685
rect 19684 287635 19716 287636
rect 19684 287605 19685 287635
rect 19685 287605 19715 287635
rect 19715 287605 19716 287635
rect 19684 287604 19716 287605
rect 19684 287555 19716 287556
rect 19684 287525 19685 287555
rect 19685 287525 19715 287555
rect 19715 287525 19716 287555
rect 19684 287524 19716 287525
rect 19684 287475 19716 287476
rect 19684 287445 19685 287475
rect 19685 287445 19715 287475
rect 19715 287445 19716 287475
rect 19684 287444 19716 287445
rect 19684 287395 19716 287396
rect 19684 287365 19685 287395
rect 19685 287365 19715 287395
rect 19715 287365 19716 287395
rect 19684 287364 19716 287365
rect 19684 287315 19716 287316
rect 19684 287285 19685 287315
rect 19685 287285 19715 287315
rect 19715 287285 19716 287315
rect 19684 287284 19716 287285
rect 19684 287235 19716 287236
rect 19684 287205 19685 287235
rect 19685 287205 19715 287235
rect 19715 287205 19716 287235
rect 19684 287204 19716 287205
rect 19684 287155 19716 287156
rect 19684 287125 19685 287155
rect 19685 287125 19715 287155
rect 19715 287125 19716 287155
rect 19684 287124 19716 287125
rect 19684 287075 19716 287076
rect 19684 287045 19685 287075
rect 19685 287045 19715 287075
rect 19715 287045 19716 287075
rect 19684 287044 19716 287045
rect 19684 286995 19716 286996
rect 19684 286965 19685 286995
rect 19685 286965 19715 286995
rect 19715 286965 19716 286995
rect 19684 286964 19716 286965
rect 19684 286915 19716 286916
rect 19684 286885 19685 286915
rect 19685 286885 19715 286915
rect 19715 286885 19716 286915
rect 19684 286884 19716 286885
rect 19684 286835 19716 286836
rect 19684 286805 19685 286835
rect 19685 286805 19715 286835
rect 19715 286805 19716 286835
rect 19684 286804 19716 286805
rect 19684 286755 19716 286756
rect 19684 286725 19685 286755
rect 19685 286725 19715 286755
rect 19715 286725 19716 286755
rect 19684 286724 19716 286725
rect 19684 286675 19716 286676
rect 19684 286645 19685 286675
rect 19685 286645 19715 286675
rect 19715 286645 19716 286675
rect 19684 286644 19716 286645
rect 19684 286595 19716 286596
rect 19684 286565 19685 286595
rect 19685 286565 19715 286595
rect 19715 286565 19716 286595
rect 19684 286564 19716 286565
rect 19684 286515 19716 286516
rect 19684 286485 19685 286515
rect 19685 286485 19715 286515
rect 19715 286485 19716 286515
rect 19684 286484 19716 286485
rect 19684 286435 19716 286436
rect 19684 286405 19685 286435
rect 19685 286405 19715 286435
rect 19715 286405 19716 286435
rect 19684 286404 19716 286405
rect 19684 286355 19716 286356
rect 19684 286325 19685 286355
rect 19685 286325 19715 286355
rect 19715 286325 19716 286355
rect 19684 286324 19716 286325
rect 19684 286275 19716 286276
rect 19684 286245 19685 286275
rect 19685 286245 19715 286275
rect 19715 286245 19716 286275
rect 19684 286244 19716 286245
rect 19684 286195 19716 286196
rect 19684 286165 19685 286195
rect 19685 286165 19715 286195
rect 19715 286165 19716 286195
rect 19684 286164 19716 286165
rect 19684 286115 19716 286116
rect 19684 286085 19685 286115
rect 19685 286085 19715 286115
rect 19715 286085 19716 286115
rect 19684 286084 19716 286085
rect 19684 286035 19716 286036
rect 19684 286005 19685 286035
rect 19685 286005 19715 286035
rect 19715 286005 19716 286035
rect 19684 286004 19716 286005
rect 19684 285955 19716 285956
rect 19684 285925 19685 285955
rect 19685 285925 19715 285955
rect 19715 285925 19716 285955
rect 19684 285924 19716 285925
rect 19684 285875 19716 285876
rect 19684 285845 19685 285875
rect 19685 285845 19715 285875
rect 19715 285845 19716 285875
rect 19684 285844 19716 285845
rect 19684 285795 19716 285796
rect 19684 285765 19685 285795
rect 19685 285765 19715 285795
rect 19715 285765 19716 285795
rect 19684 285764 19716 285765
rect 19684 285715 19716 285716
rect 19684 285685 19685 285715
rect 19685 285685 19715 285715
rect 19715 285685 19716 285715
rect 19684 285684 19716 285685
rect 19684 285635 19716 285636
rect 19684 285605 19685 285635
rect 19685 285605 19715 285635
rect 19715 285605 19716 285635
rect 19684 285604 19716 285605
rect 19684 285555 19716 285556
rect 19684 285525 19685 285555
rect 19685 285525 19715 285555
rect 19715 285525 19716 285555
rect 19684 285524 19716 285525
rect 19684 285475 19716 285476
rect 19684 285445 19685 285475
rect 19685 285445 19715 285475
rect 19715 285445 19716 285475
rect 19684 285444 19716 285445
rect 19684 285395 19716 285396
rect 19684 285365 19685 285395
rect 19685 285365 19715 285395
rect 19715 285365 19716 285395
rect 19684 285364 19716 285365
rect 19684 285315 19716 285316
rect 19684 285285 19685 285315
rect 19685 285285 19715 285315
rect 19715 285285 19716 285315
rect 19684 285284 19716 285285
rect 19684 285235 19716 285236
rect 19684 285205 19685 285235
rect 19685 285205 19715 285235
rect 19715 285205 19716 285235
rect 19684 285204 19716 285205
rect 19684 285155 19716 285156
rect 19684 285125 19685 285155
rect 19685 285125 19715 285155
rect 19715 285125 19716 285155
rect 19684 285124 19716 285125
rect 19684 285075 19716 285076
rect 19684 285045 19685 285075
rect 19685 285045 19715 285075
rect 19715 285045 19716 285075
rect 19684 285044 19716 285045
rect 19684 284995 19716 284996
rect 19684 284965 19685 284995
rect 19685 284965 19715 284995
rect 19715 284965 19716 284995
rect 19684 284964 19716 284965
rect 19684 284915 19716 284916
rect 19684 284885 19685 284915
rect 19685 284885 19715 284915
rect 19715 284885 19716 284915
rect 19684 284884 19716 284885
rect 19684 284835 19716 284836
rect 19684 284805 19685 284835
rect 19685 284805 19715 284835
rect 19715 284805 19716 284835
rect 19684 284804 19716 284805
rect 19684 284755 19716 284756
rect 19684 284725 19685 284755
rect 19685 284725 19715 284755
rect 19715 284725 19716 284755
rect 19684 284724 19716 284725
rect 19684 284675 19716 284676
rect 19684 284645 19685 284675
rect 19685 284645 19715 284675
rect 19715 284645 19716 284675
rect 19684 284644 19716 284645
rect 19684 284595 19716 284596
rect 19684 284565 19685 284595
rect 19685 284565 19715 284595
rect 19715 284565 19716 284595
rect 19684 284564 19716 284565
rect 19684 284515 19716 284516
rect 19684 284485 19685 284515
rect 19685 284485 19715 284515
rect 19715 284485 19716 284515
rect 19684 284484 19716 284485
rect 19684 284435 19716 284436
rect 19684 284405 19685 284435
rect 19685 284405 19715 284435
rect 19715 284405 19716 284435
rect 19684 284404 19716 284405
rect 19684 284355 19716 284356
rect 19684 284325 19685 284355
rect 19685 284325 19715 284355
rect 19715 284325 19716 284355
rect 19684 284324 19716 284325
rect 19684 284275 19716 284276
rect 19684 284245 19685 284275
rect 19685 284245 19715 284275
rect 19715 284245 19716 284275
rect 19684 284244 19716 284245
rect 19684 284195 19716 284196
rect 19684 284165 19685 284195
rect 19685 284165 19715 284195
rect 19715 284165 19716 284195
rect 19684 284164 19716 284165
rect 19684 284115 19716 284116
rect 19684 284085 19685 284115
rect 19685 284085 19715 284115
rect 19715 284085 19716 284115
rect 19684 284084 19716 284085
rect 19684 284035 19716 284036
rect 19684 284005 19685 284035
rect 19685 284005 19715 284035
rect 19715 284005 19716 284035
rect 19684 284004 19716 284005
rect 19684 283955 19716 283956
rect 19684 283925 19685 283955
rect 19685 283925 19715 283955
rect 19715 283925 19716 283955
rect 19684 283924 19716 283925
rect 19684 283875 19716 283876
rect 19684 283845 19685 283875
rect 19685 283845 19715 283875
rect 19715 283845 19716 283875
rect 19684 283844 19716 283845
rect 19684 283795 19716 283796
rect 19684 283765 19685 283795
rect 19685 283765 19715 283795
rect 19715 283765 19716 283795
rect 19684 283764 19716 283765
rect 19684 283715 19716 283716
rect 19684 283685 19685 283715
rect 19685 283685 19715 283715
rect 19715 283685 19716 283715
rect 19684 283684 19716 283685
rect 19684 283635 19716 283636
rect 19684 283605 19685 283635
rect 19685 283605 19715 283635
rect 19715 283605 19716 283635
rect 19684 283604 19716 283605
rect 19684 283555 19716 283556
rect 19684 283525 19685 283555
rect 19685 283525 19715 283555
rect 19715 283525 19716 283555
rect 19684 283524 19716 283525
rect 19684 283475 19716 283476
rect 19684 283445 19685 283475
rect 19685 283445 19715 283475
rect 19715 283445 19716 283475
rect 19684 283444 19716 283445
rect 19684 283395 19716 283396
rect 19684 283365 19685 283395
rect 19685 283365 19715 283395
rect 19715 283365 19716 283395
rect 19684 283364 19716 283365
rect 19684 283315 19716 283316
rect 19684 283285 19685 283315
rect 19685 283285 19715 283315
rect 19715 283285 19716 283315
rect 19684 283284 19716 283285
rect 19684 283235 19716 283236
rect 19684 283205 19685 283235
rect 19685 283205 19715 283235
rect 19715 283205 19716 283235
rect 19684 283204 19716 283205
rect 19684 283155 19716 283156
rect 19684 283125 19685 283155
rect 19685 283125 19715 283155
rect 19715 283125 19716 283155
rect 19684 283124 19716 283125
rect 19684 283075 19716 283076
rect 19684 283045 19685 283075
rect 19685 283045 19715 283075
rect 19715 283045 19716 283075
rect 19684 283044 19716 283045
rect 19684 282995 19716 282996
rect 19684 282965 19685 282995
rect 19685 282965 19715 282995
rect 19715 282965 19716 282995
rect 19684 282964 19716 282965
rect 19684 282915 19716 282916
rect 19684 282885 19685 282915
rect 19685 282885 19715 282915
rect 19715 282885 19716 282915
rect 19684 282884 19716 282885
rect 19684 282835 19716 282836
rect 19684 282805 19685 282835
rect 19685 282805 19715 282835
rect 19715 282805 19716 282835
rect 19684 282804 19716 282805
rect 19684 282755 19716 282756
rect 19684 282725 19685 282755
rect 19685 282725 19715 282755
rect 19715 282725 19716 282755
rect 19684 282724 19716 282725
rect 19684 282675 19716 282676
rect 19684 282645 19685 282675
rect 19685 282645 19715 282675
rect 19715 282645 19716 282675
rect 19684 282644 19716 282645
rect 19684 282595 19716 282596
rect 19684 282565 19685 282595
rect 19685 282565 19715 282595
rect 19715 282565 19716 282595
rect 19684 282564 19716 282565
rect 19684 282515 19716 282516
rect 19684 282485 19685 282515
rect 19685 282485 19715 282515
rect 19715 282485 19716 282515
rect 19684 282484 19716 282485
rect 19684 282435 19716 282436
rect 19684 282405 19685 282435
rect 19685 282405 19715 282435
rect 19715 282405 19716 282435
rect 19684 282404 19716 282405
rect 19684 282355 19716 282356
rect 19684 282325 19685 282355
rect 19685 282325 19715 282355
rect 19715 282325 19716 282355
rect 19684 282324 19716 282325
rect 19684 282275 19716 282276
rect 19684 282245 19685 282275
rect 19685 282245 19715 282275
rect 19715 282245 19716 282275
rect 19684 282244 19716 282245
rect 19684 282195 19716 282196
rect 19684 282165 19685 282195
rect 19685 282165 19715 282195
rect 19715 282165 19716 282195
rect 19684 282164 19716 282165
rect 19684 282115 19716 282116
rect 19684 282085 19685 282115
rect 19685 282085 19715 282115
rect 19715 282085 19716 282115
rect 19684 282084 19716 282085
rect 19684 282035 19716 282036
rect 19684 282005 19685 282035
rect 19685 282005 19715 282035
rect 19715 282005 19716 282035
rect 19684 282004 19716 282005
rect 19684 281955 19716 281956
rect 19684 281925 19685 281955
rect 19685 281925 19715 281955
rect 19715 281925 19716 281955
rect 19684 281924 19716 281925
rect 19684 281875 19716 281876
rect 19684 281845 19685 281875
rect 19685 281845 19715 281875
rect 19715 281845 19716 281875
rect 19684 281844 19716 281845
rect 19684 281795 19716 281796
rect 19684 281765 19685 281795
rect 19685 281765 19715 281795
rect 19715 281765 19716 281795
rect 19684 281764 19716 281765
rect 19684 281715 19716 281716
rect 19684 281685 19685 281715
rect 19685 281685 19715 281715
rect 19715 281685 19716 281715
rect 19684 281684 19716 281685
rect 19684 281635 19716 281636
rect 19684 281605 19685 281635
rect 19685 281605 19715 281635
rect 19715 281605 19716 281635
rect 19684 281604 19716 281605
rect 19684 281555 19716 281556
rect 19684 281525 19685 281555
rect 19685 281525 19715 281555
rect 19715 281525 19716 281555
rect 19684 281524 19716 281525
rect 19684 281475 19716 281476
rect 19684 281445 19685 281475
rect 19685 281445 19715 281475
rect 19715 281445 19716 281475
rect 19684 281444 19716 281445
rect 19684 281395 19716 281396
rect 19684 281365 19685 281395
rect 19685 281365 19715 281395
rect 19715 281365 19716 281395
rect 19684 281364 19716 281365
rect 19684 281315 19716 281316
rect 19684 281285 19685 281315
rect 19685 281285 19715 281315
rect 19715 281285 19716 281315
rect 19684 281284 19716 281285
rect 19684 281235 19716 281236
rect 19684 281205 19685 281235
rect 19685 281205 19715 281235
rect 19715 281205 19716 281235
rect 19684 281204 19716 281205
rect 19684 281155 19716 281156
rect 19684 281125 19685 281155
rect 19685 281125 19715 281155
rect 19715 281125 19716 281155
rect 19684 281124 19716 281125
rect 19684 281075 19716 281076
rect 19684 281045 19685 281075
rect 19685 281045 19715 281075
rect 19715 281045 19716 281075
rect 19684 281044 19716 281045
rect 19684 280995 19716 280996
rect 19684 280965 19685 280995
rect 19685 280965 19715 280995
rect 19715 280965 19716 280995
rect 19684 280964 19716 280965
rect 19684 280915 19716 280916
rect 19684 280885 19685 280915
rect 19685 280885 19715 280915
rect 19715 280885 19716 280915
rect 19684 280884 19716 280885
rect 19684 280835 19716 280836
rect 19684 280805 19685 280835
rect 19685 280805 19715 280835
rect 19715 280805 19716 280835
rect 19684 280804 19716 280805
rect 19684 280755 19716 280756
rect 19684 280725 19685 280755
rect 19685 280725 19715 280755
rect 19715 280725 19716 280755
rect 19684 280724 19716 280725
rect 19684 280675 19716 280676
rect 19684 280645 19685 280675
rect 19685 280645 19715 280675
rect 19715 280645 19716 280675
rect 19684 280644 19716 280645
rect 19684 280595 19716 280596
rect 19684 280565 19685 280595
rect 19685 280565 19715 280595
rect 19715 280565 19716 280595
rect 19684 280564 19716 280565
rect 19684 280515 19716 280516
rect 19684 280485 19685 280515
rect 19685 280485 19715 280515
rect 19715 280485 19716 280515
rect 19684 280484 19716 280485
rect 19684 280435 19716 280436
rect 19684 280405 19685 280435
rect 19685 280405 19715 280435
rect 19715 280405 19716 280435
rect 19684 280404 19716 280405
rect 19684 280355 19716 280356
rect 19684 280325 19685 280355
rect 19685 280325 19715 280355
rect 19715 280325 19716 280355
rect 19684 280324 19716 280325
rect 19684 280275 19716 280276
rect 19684 280245 19685 280275
rect 19685 280245 19715 280275
rect 19715 280245 19716 280275
rect 19684 280244 19716 280245
rect 19684 280195 19716 280196
rect 19684 280165 19685 280195
rect 19685 280165 19715 280195
rect 19715 280165 19716 280195
rect 19684 280164 19716 280165
rect 19684 280115 19716 280116
rect 19684 280085 19685 280115
rect 19685 280085 19715 280115
rect 19715 280085 19716 280115
rect 19684 280084 19716 280085
rect 19684 280035 19716 280036
rect 19684 280005 19685 280035
rect 19685 280005 19715 280035
rect 19715 280005 19716 280035
rect 19684 280004 19716 280005
rect 19684 279955 19716 279956
rect 19684 279925 19685 279955
rect 19685 279925 19715 279955
rect 19715 279925 19716 279955
rect 19684 279924 19716 279925
rect 19684 279875 19716 279876
rect 19684 279845 19685 279875
rect 19685 279845 19715 279875
rect 19715 279845 19716 279875
rect 19684 279844 19716 279845
rect 19684 279795 19716 279796
rect 19684 279765 19685 279795
rect 19685 279765 19715 279795
rect 19715 279765 19716 279795
rect 19684 279764 19716 279765
rect 19684 279715 19716 279716
rect 19684 279685 19685 279715
rect 19685 279685 19715 279715
rect 19715 279685 19716 279715
rect 19684 279684 19716 279685
rect 19684 279635 19716 279636
rect 19684 279605 19685 279635
rect 19685 279605 19715 279635
rect 19715 279605 19716 279635
rect 19684 279604 19716 279605
rect 19684 279555 19716 279556
rect 19684 279525 19685 279555
rect 19685 279525 19715 279555
rect 19715 279525 19716 279555
rect 19684 279524 19716 279525
rect 19684 279475 19716 279476
rect 19684 279445 19685 279475
rect 19685 279445 19715 279475
rect 19715 279445 19716 279475
rect 19684 279444 19716 279445
rect 2450 279250 2550 279350
rect 1040 275040 1160 275160
rect 19684 279395 19716 279396
rect 19684 279365 19685 279395
rect 19685 279365 19715 279395
rect 19715 279365 19716 279395
rect 19684 279364 19716 279365
rect 19684 279315 19716 279316
rect 19684 279285 19685 279315
rect 19685 279285 19715 279315
rect 19715 279285 19716 279315
rect 19684 279284 19716 279285
rect 19684 279235 19716 279236
rect 19684 279205 19685 279235
rect 19685 279205 19715 279235
rect 19715 279205 19716 279235
rect 19684 279204 19716 279205
rect 19684 279155 19716 279156
rect 19684 279125 19685 279155
rect 19685 279125 19715 279155
rect 19715 279125 19716 279155
rect 19684 279124 19716 279125
rect 19684 279075 19716 279076
rect 19684 279045 19685 279075
rect 19685 279045 19715 279075
rect 19715 279045 19716 279075
rect 19684 279044 19716 279045
rect 19684 278995 19716 278996
rect 19684 278965 19685 278995
rect 19685 278965 19715 278995
rect 19715 278965 19716 278995
rect 19684 278964 19716 278965
rect 19684 278915 19716 278916
rect 19684 278885 19685 278915
rect 19685 278885 19715 278915
rect 19715 278885 19716 278915
rect 19684 278884 19716 278885
rect 19684 278835 19716 278836
rect 19684 278805 19685 278835
rect 19685 278805 19715 278835
rect 19715 278805 19716 278835
rect 19684 278804 19716 278805
rect 19684 278755 19716 278756
rect 19684 278725 19685 278755
rect 19685 278725 19715 278755
rect 19715 278725 19716 278755
rect 19684 278724 19716 278725
rect 17044 278675 17076 278676
rect 17044 278645 17045 278675
rect 17045 278645 17075 278675
rect 17075 278645 17076 278675
rect 17044 278644 17076 278645
rect 17204 278675 17236 278676
rect 17204 278645 17205 278675
rect 17205 278645 17235 278675
rect 17235 278645 17236 278675
rect 17204 278644 17236 278645
rect 17044 278564 17076 278596
rect 17044 278515 17076 278516
rect 17044 278485 17045 278515
rect 17045 278485 17075 278515
rect 17075 278485 17076 278515
rect 17044 278484 17076 278485
rect 17044 278435 17076 278436
rect 17044 278405 17045 278435
rect 17045 278405 17075 278435
rect 17075 278405 17076 278435
rect 17044 278404 17076 278405
rect 17044 278355 17076 278356
rect 17044 278325 17045 278355
rect 17045 278325 17075 278355
rect 17075 278325 17076 278355
rect 17044 278324 17076 278325
rect 17044 278275 17076 278276
rect 17044 278245 17045 278275
rect 17045 278245 17075 278275
rect 17075 278245 17076 278275
rect 17044 278244 17076 278245
rect 17044 278195 17076 278196
rect 17044 278165 17045 278195
rect 17045 278165 17075 278195
rect 17075 278165 17076 278195
rect 17044 278164 17076 278165
rect 17044 278115 17076 278116
rect 17044 278085 17045 278115
rect 17045 278085 17075 278115
rect 17075 278085 17076 278115
rect 17044 278084 17076 278085
rect 17044 278035 17076 278036
rect 17044 278005 17045 278035
rect 17045 278005 17075 278035
rect 17075 278005 17076 278035
rect 17044 278004 17076 278005
rect 17044 277955 17076 277956
rect 17044 277925 17045 277955
rect 17045 277925 17075 277955
rect 17075 277925 17076 277955
rect 17044 277924 17076 277925
rect 17044 277875 17076 277876
rect 17044 277845 17045 277875
rect 17045 277845 17075 277875
rect 17075 277845 17076 277875
rect 17044 277844 17076 277845
rect 17204 278564 17236 278596
rect 17204 278515 17236 278516
rect 17204 278485 17205 278515
rect 17205 278485 17235 278515
rect 17235 278485 17236 278515
rect 17204 278484 17236 278485
rect 17284 278675 17316 278676
rect 17284 278645 17285 278675
rect 17285 278645 17315 278675
rect 17315 278645 17316 278675
rect 17284 278644 17316 278645
rect 17284 278564 17316 278596
rect 17284 278515 17316 278516
rect 17284 278485 17285 278515
rect 17285 278485 17315 278515
rect 17315 278485 17316 278515
rect 17284 278484 17316 278485
rect 17364 278675 17396 278676
rect 17364 278645 17365 278675
rect 17365 278645 17395 278675
rect 17395 278645 17396 278675
rect 17364 278644 17396 278645
rect 17364 278564 17396 278596
rect 17364 278515 17396 278516
rect 17364 278485 17365 278515
rect 17365 278485 17395 278515
rect 17395 278485 17396 278515
rect 17364 278484 17396 278485
rect 17444 278675 17476 278676
rect 17444 278645 17445 278675
rect 17445 278645 17475 278675
rect 17475 278645 17476 278675
rect 17444 278644 17476 278645
rect 17444 278564 17476 278596
rect 17444 278515 17476 278516
rect 17444 278485 17445 278515
rect 17445 278485 17475 278515
rect 17475 278485 17476 278515
rect 17444 278484 17476 278485
rect 17524 278675 17556 278676
rect 17524 278645 17525 278675
rect 17525 278645 17555 278675
rect 17555 278645 17556 278675
rect 17524 278644 17556 278645
rect 17524 278564 17556 278596
rect 17524 278515 17556 278516
rect 17524 278485 17525 278515
rect 17525 278485 17555 278515
rect 17555 278485 17556 278515
rect 17524 278484 17556 278485
rect 17604 278675 17636 278676
rect 17604 278645 17605 278675
rect 17605 278645 17635 278675
rect 17635 278645 17636 278675
rect 17604 278644 17636 278645
rect 17604 278564 17636 278596
rect 17604 278515 17636 278516
rect 17604 278485 17605 278515
rect 17605 278485 17635 278515
rect 17635 278485 17636 278515
rect 17604 278484 17636 278485
rect 17684 278675 17716 278676
rect 17684 278645 17685 278675
rect 17685 278645 17715 278675
rect 17715 278645 17716 278675
rect 17684 278644 17716 278645
rect 17684 278564 17716 278596
rect 17684 278515 17716 278516
rect 17684 278485 17685 278515
rect 17685 278485 17715 278515
rect 17715 278485 17716 278515
rect 17684 278484 17716 278485
rect 17764 278675 17796 278676
rect 17764 278645 17765 278675
rect 17765 278645 17795 278675
rect 17795 278645 17796 278675
rect 17764 278644 17796 278645
rect 17764 278564 17796 278596
rect 17764 278515 17796 278516
rect 17764 278485 17765 278515
rect 17765 278485 17795 278515
rect 17795 278485 17796 278515
rect 17764 278484 17796 278485
rect 19524 278675 19556 278676
rect 19524 278645 19525 278675
rect 19525 278645 19555 278675
rect 19555 278645 19556 278675
rect 19524 278644 19556 278645
rect 19524 278564 19556 278596
rect 19524 278515 19556 278516
rect 19524 278485 19525 278515
rect 19525 278485 19555 278515
rect 19555 278485 19556 278515
rect 19524 278484 19556 278485
rect 19604 278675 19636 278676
rect 19604 278645 19605 278675
rect 19605 278645 19635 278675
rect 19635 278645 19636 278675
rect 19604 278644 19636 278645
rect 19604 278564 19636 278596
rect 19604 278515 19636 278516
rect 19604 278485 19605 278515
rect 19605 278485 19635 278515
rect 19635 278485 19636 278515
rect 19604 278484 19636 278485
rect 19684 278675 19716 278676
rect 19684 278645 19685 278675
rect 19685 278645 19715 278675
rect 19715 278645 19716 278675
rect 19684 278644 19716 278645
rect 19684 278564 19716 278596
rect 19844 351235 19876 351236
rect 19844 351205 19845 351235
rect 19845 351205 19875 351235
rect 19875 351205 19876 351235
rect 19844 351204 19876 351205
rect 19844 351155 19876 351156
rect 19844 351125 19845 351155
rect 19845 351125 19875 351155
rect 19875 351125 19876 351155
rect 19844 351124 19876 351125
rect 19844 351075 19876 351076
rect 19844 351045 19845 351075
rect 19845 351045 19875 351075
rect 19875 351045 19876 351075
rect 19844 351044 19876 351045
rect 19844 350995 19876 350996
rect 19844 350965 19845 350995
rect 19845 350965 19875 350995
rect 19875 350965 19876 350995
rect 19844 350964 19876 350965
rect 19844 350915 19876 350916
rect 19844 350885 19845 350915
rect 19845 350885 19875 350915
rect 19875 350885 19876 350915
rect 19844 350884 19876 350885
rect 19844 350835 19876 350836
rect 19844 350805 19845 350835
rect 19845 350805 19875 350835
rect 19875 350805 19876 350835
rect 19844 350804 19876 350805
rect 19844 350755 19876 350756
rect 19844 350725 19845 350755
rect 19845 350725 19875 350755
rect 19875 350725 19876 350755
rect 19844 350724 19876 350725
rect 19844 350675 19876 350676
rect 19844 350645 19845 350675
rect 19845 350645 19875 350675
rect 19875 350645 19876 350675
rect 19844 350644 19876 350645
rect 19844 350595 19876 350596
rect 19844 350565 19845 350595
rect 19845 350565 19875 350595
rect 19875 350565 19876 350595
rect 19844 350564 19876 350565
rect 19844 350515 19876 350516
rect 19844 350485 19845 350515
rect 19845 350485 19875 350515
rect 19875 350485 19876 350515
rect 19844 350484 19876 350485
rect 19844 350435 19876 350436
rect 19844 350405 19845 350435
rect 19845 350405 19875 350435
rect 19875 350405 19876 350435
rect 19844 350404 19876 350405
rect 19844 350355 19876 350356
rect 19844 350325 19845 350355
rect 19845 350325 19875 350355
rect 19875 350325 19876 350355
rect 19844 350324 19876 350325
rect 19844 350275 19876 350276
rect 19844 350245 19845 350275
rect 19845 350245 19875 350275
rect 19875 350245 19876 350275
rect 19844 350244 19876 350245
rect 19844 350195 19876 350196
rect 19844 350165 19845 350195
rect 19845 350165 19875 350195
rect 19875 350165 19876 350195
rect 19844 350164 19876 350165
rect 19844 350115 19876 350116
rect 19844 350085 19845 350115
rect 19845 350085 19875 350115
rect 19875 350085 19876 350115
rect 19844 350084 19876 350085
rect 19844 350035 19876 350036
rect 19844 350005 19845 350035
rect 19845 350005 19875 350035
rect 19875 350005 19876 350035
rect 19844 350004 19876 350005
rect 19844 349955 19876 349956
rect 19844 349925 19845 349955
rect 19845 349925 19875 349955
rect 19875 349925 19876 349955
rect 19844 349924 19876 349925
rect 19844 349875 19876 349876
rect 19844 349845 19845 349875
rect 19845 349845 19875 349875
rect 19875 349845 19876 349875
rect 19844 349844 19876 349845
rect 19844 349795 19876 349796
rect 19844 349765 19845 349795
rect 19845 349765 19875 349795
rect 19875 349765 19876 349795
rect 19844 349764 19876 349765
rect 19844 349715 19876 349716
rect 19844 349685 19845 349715
rect 19845 349685 19875 349715
rect 19875 349685 19876 349715
rect 19844 349684 19876 349685
rect 19844 349635 19876 349636
rect 19844 349605 19845 349635
rect 19845 349605 19875 349635
rect 19875 349605 19876 349635
rect 19844 349604 19876 349605
rect 19844 349555 19876 349556
rect 19844 349525 19845 349555
rect 19845 349525 19875 349555
rect 19875 349525 19876 349555
rect 19844 349524 19876 349525
rect 19844 349475 19876 349476
rect 19844 349445 19845 349475
rect 19845 349445 19875 349475
rect 19875 349445 19876 349475
rect 19844 349444 19876 349445
rect 19844 349395 19876 349396
rect 19844 349365 19845 349395
rect 19845 349365 19875 349395
rect 19875 349365 19876 349395
rect 19844 349364 19876 349365
rect 19844 349315 19876 349316
rect 19844 349285 19845 349315
rect 19845 349285 19875 349315
rect 19875 349285 19876 349315
rect 19844 349284 19876 349285
rect 19844 349235 19876 349236
rect 19844 349205 19845 349235
rect 19845 349205 19875 349235
rect 19875 349205 19876 349235
rect 19844 349204 19876 349205
rect 19844 349155 19876 349156
rect 19844 349125 19845 349155
rect 19845 349125 19875 349155
rect 19875 349125 19876 349155
rect 19844 349124 19876 349125
rect 19844 349075 19876 349076
rect 19844 349045 19845 349075
rect 19845 349045 19875 349075
rect 19875 349045 19876 349075
rect 19844 349044 19876 349045
rect 19844 348995 19876 348996
rect 19844 348965 19845 348995
rect 19845 348965 19875 348995
rect 19875 348965 19876 348995
rect 19844 348964 19876 348965
rect 19844 348915 19876 348916
rect 19844 348885 19845 348915
rect 19845 348885 19875 348915
rect 19875 348885 19876 348915
rect 19844 348884 19876 348885
rect 19844 348835 19876 348836
rect 19844 348805 19845 348835
rect 19845 348805 19875 348835
rect 19875 348805 19876 348835
rect 19844 348804 19876 348805
rect 19844 348755 19876 348756
rect 19844 348725 19845 348755
rect 19845 348725 19875 348755
rect 19875 348725 19876 348755
rect 19844 348724 19876 348725
rect 19844 348675 19876 348676
rect 19844 348645 19845 348675
rect 19845 348645 19875 348675
rect 19875 348645 19876 348675
rect 19844 348644 19876 348645
rect 19844 348595 19876 348596
rect 19844 348565 19845 348595
rect 19845 348565 19875 348595
rect 19875 348565 19876 348595
rect 19844 348564 19876 348565
rect 19844 348515 19876 348516
rect 19844 348485 19845 348515
rect 19845 348485 19875 348515
rect 19875 348485 19876 348515
rect 19844 348484 19876 348485
rect 19844 348435 19876 348436
rect 19844 348405 19845 348435
rect 19845 348405 19875 348435
rect 19875 348405 19876 348435
rect 19844 348404 19876 348405
rect 19844 348355 19876 348356
rect 19844 348325 19845 348355
rect 19845 348325 19875 348355
rect 19875 348325 19876 348355
rect 19844 348324 19876 348325
rect 19844 348275 19876 348276
rect 19844 348245 19845 348275
rect 19845 348245 19875 348275
rect 19875 348245 19876 348275
rect 19844 348244 19876 348245
rect 19844 348195 19876 348196
rect 19844 348165 19845 348195
rect 19845 348165 19875 348195
rect 19875 348165 19876 348195
rect 19844 348164 19876 348165
rect 19844 348115 19876 348116
rect 19844 348085 19845 348115
rect 19845 348085 19875 348115
rect 19875 348085 19876 348115
rect 19844 348084 19876 348085
rect 19844 348035 19876 348036
rect 19844 348005 19845 348035
rect 19845 348005 19875 348035
rect 19875 348005 19876 348035
rect 19844 348004 19876 348005
rect 19844 347955 19876 347956
rect 19844 347925 19845 347955
rect 19845 347925 19875 347955
rect 19875 347925 19876 347955
rect 19844 347924 19876 347925
rect 19844 347875 19876 347876
rect 19844 347845 19845 347875
rect 19845 347845 19875 347875
rect 19875 347845 19876 347875
rect 19844 347844 19876 347845
rect 19844 347795 19876 347796
rect 19844 347765 19845 347795
rect 19845 347765 19875 347795
rect 19875 347765 19876 347795
rect 19844 347764 19876 347765
rect 19844 347715 19876 347716
rect 19844 347685 19845 347715
rect 19845 347685 19875 347715
rect 19875 347685 19876 347715
rect 19844 347684 19876 347685
rect 19844 347635 19876 347636
rect 19844 347605 19845 347635
rect 19845 347605 19875 347635
rect 19875 347605 19876 347635
rect 19844 347604 19876 347605
rect 19844 347555 19876 347556
rect 19844 347525 19845 347555
rect 19845 347525 19875 347555
rect 19875 347525 19876 347555
rect 19844 347524 19876 347525
rect 19844 347475 19876 347476
rect 19844 347445 19845 347475
rect 19845 347445 19875 347475
rect 19875 347445 19876 347475
rect 19844 347444 19876 347445
rect 19844 347395 19876 347396
rect 19844 347365 19845 347395
rect 19845 347365 19875 347395
rect 19875 347365 19876 347395
rect 19844 347364 19876 347365
rect 19844 347315 19876 347316
rect 19844 347285 19845 347315
rect 19845 347285 19875 347315
rect 19875 347285 19876 347315
rect 19844 347284 19876 347285
rect 19844 347235 19876 347236
rect 19844 347205 19845 347235
rect 19845 347205 19875 347235
rect 19875 347205 19876 347235
rect 19844 347204 19876 347205
rect 19844 347155 19876 347156
rect 19844 347125 19845 347155
rect 19845 347125 19875 347155
rect 19875 347125 19876 347155
rect 19844 347124 19876 347125
rect 19844 347075 19876 347076
rect 19844 347045 19845 347075
rect 19845 347045 19875 347075
rect 19875 347045 19876 347075
rect 19844 347044 19876 347045
rect 19844 346995 19876 346996
rect 19844 346965 19845 346995
rect 19845 346965 19875 346995
rect 19875 346965 19876 346995
rect 19844 346964 19876 346965
rect 19844 346915 19876 346916
rect 19844 346885 19845 346915
rect 19845 346885 19875 346915
rect 19875 346885 19876 346915
rect 19844 346884 19876 346885
rect 19844 346835 19876 346836
rect 19844 346805 19845 346835
rect 19845 346805 19875 346835
rect 19875 346805 19876 346835
rect 19844 346804 19876 346805
rect 19844 346755 19876 346756
rect 19844 346725 19845 346755
rect 19845 346725 19875 346755
rect 19875 346725 19876 346755
rect 19844 346724 19876 346725
rect 19844 346675 19876 346676
rect 19844 346645 19845 346675
rect 19845 346645 19875 346675
rect 19875 346645 19876 346675
rect 19844 346644 19876 346645
rect 19844 346595 19876 346596
rect 19844 346565 19845 346595
rect 19845 346565 19875 346595
rect 19875 346565 19876 346595
rect 19844 346564 19876 346565
rect 19844 346515 19876 346516
rect 19844 346485 19845 346515
rect 19845 346485 19875 346515
rect 19875 346485 19876 346515
rect 19844 346484 19876 346485
rect 19844 346435 19876 346436
rect 19844 346405 19845 346435
rect 19845 346405 19875 346435
rect 19875 346405 19876 346435
rect 19844 346404 19876 346405
rect 19844 346355 19876 346356
rect 19844 346325 19845 346355
rect 19845 346325 19875 346355
rect 19875 346325 19876 346355
rect 19844 346324 19876 346325
rect 19844 346275 19876 346276
rect 19844 346245 19845 346275
rect 19845 346245 19875 346275
rect 19875 346245 19876 346275
rect 19844 346244 19876 346245
rect 19844 346195 19876 346196
rect 19844 346165 19845 346195
rect 19845 346165 19875 346195
rect 19875 346165 19876 346195
rect 19844 346164 19876 346165
rect 19844 346115 19876 346116
rect 19844 346085 19845 346115
rect 19845 346085 19875 346115
rect 19875 346085 19876 346115
rect 19844 346084 19876 346085
rect 19844 346035 19876 346036
rect 19844 346005 19845 346035
rect 19845 346005 19875 346035
rect 19875 346005 19876 346035
rect 19844 346004 19876 346005
rect 19844 345955 19876 345956
rect 19844 345925 19845 345955
rect 19845 345925 19875 345955
rect 19875 345925 19876 345955
rect 19844 345924 19876 345925
rect 19844 345875 19876 345876
rect 19844 345845 19845 345875
rect 19845 345845 19875 345875
rect 19875 345845 19876 345875
rect 19844 345844 19876 345845
rect 19844 345795 19876 345796
rect 19844 345765 19845 345795
rect 19845 345765 19875 345795
rect 19875 345765 19876 345795
rect 19844 345764 19876 345765
rect 19844 345715 19876 345716
rect 19844 345685 19845 345715
rect 19845 345685 19875 345715
rect 19875 345685 19876 345715
rect 19844 345684 19876 345685
rect 19844 345635 19876 345636
rect 19844 345605 19845 345635
rect 19845 345605 19875 345635
rect 19875 345605 19876 345635
rect 19844 345604 19876 345605
rect 19844 345555 19876 345556
rect 19844 345525 19845 345555
rect 19845 345525 19875 345555
rect 19875 345525 19876 345555
rect 19844 345524 19876 345525
rect 19844 345475 19876 345476
rect 19844 345445 19845 345475
rect 19845 345445 19875 345475
rect 19875 345445 19876 345475
rect 19844 345444 19876 345445
rect 19844 345395 19876 345396
rect 19844 345365 19845 345395
rect 19845 345365 19875 345395
rect 19875 345365 19876 345395
rect 19844 345364 19876 345365
rect 19844 345315 19876 345316
rect 19844 345285 19845 345315
rect 19845 345285 19875 345315
rect 19875 345285 19876 345315
rect 19844 345284 19876 345285
rect 19844 345235 19876 345236
rect 19844 345205 19845 345235
rect 19845 345205 19875 345235
rect 19875 345205 19876 345235
rect 19844 345204 19876 345205
rect 19844 345155 19876 345156
rect 19844 345125 19845 345155
rect 19845 345125 19875 345155
rect 19875 345125 19876 345155
rect 19844 345124 19876 345125
rect 19844 345075 19876 345076
rect 19844 345045 19845 345075
rect 19845 345045 19875 345075
rect 19875 345045 19876 345075
rect 19844 345044 19876 345045
rect 19844 344995 19876 344996
rect 19844 344965 19845 344995
rect 19845 344965 19875 344995
rect 19875 344965 19876 344995
rect 19844 344964 19876 344965
rect 19844 344915 19876 344916
rect 19844 344885 19845 344915
rect 19845 344885 19875 344915
rect 19875 344885 19876 344915
rect 19844 344884 19876 344885
rect 19844 344835 19876 344836
rect 19844 344805 19845 344835
rect 19845 344805 19875 344835
rect 19875 344805 19876 344835
rect 19844 344804 19876 344805
rect 19844 344755 19876 344756
rect 19844 344725 19845 344755
rect 19845 344725 19875 344755
rect 19875 344725 19876 344755
rect 19844 344724 19876 344725
rect 19844 344675 19876 344676
rect 19844 344645 19845 344675
rect 19845 344645 19875 344675
rect 19875 344645 19876 344675
rect 19844 344644 19876 344645
rect 19844 344595 19876 344596
rect 19844 344565 19845 344595
rect 19845 344565 19875 344595
rect 19875 344565 19876 344595
rect 19844 344564 19876 344565
rect 19844 344515 19876 344516
rect 19844 344485 19845 344515
rect 19845 344485 19875 344515
rect 19875 344485 19876 344515
rect 19844 344484 19876 344485
rect 19844 344435 19876 344436
rect 19844 344405 19845 344435
rect 19845 344405 19875 344435
rect 19875 344405 19876 344435
rect 19844 344404 19876 344405
rect 19844 344355 19876 344356
rect 19844 344325 19845 344355
rect 19845 344325 19875 344355
rect 19875 344325 19876 344355
rect 19844 344324 19876 344325
rect 19844 344275 19876 344276
rect 19844 344245 19845 344275
rect 19845 344245 19875 344275
rect 19875 344245 19876 344275
rect 19844 344244 19876 344245
rect 19844 344195 19876 344196
rect 19844 344165 19845 344195
rect 19845 344165 19875 344195
rect 19875 344165 19876 344195
rect 19844 344164 19876 344165
rect 19844 344115 19876 344116
rect 19844 344085 19845 344115
rect 19845 344085 19875 344115
rect 19875 344085 19876 344115
rect 19844 344084 19876 344085
rect 19844 344035 19876 344036
rect 19844 344005 19845 344035
rect 19845 344005 19875 344035
rect 19875 344005 19876 344035
rect 19844 344004 19876 344005
rect 19844 343955 19876 343956
rect 19844 343925 19845 343955
rect 19845 343925 19875 343955
rect 19875 343925 19876 343955
rect 19844 343924 19876 343925
rect 19844 343875 19876 343876
rect 19844 343845 19845 343875
rect 19845 343845 19875 343875
rect 19875 343845 19876 343875
rect 19844 343844 19876 343845
rect 19844 343795 19876 343796
rect 19844 343765 19845 343795
rect 19845 343765 19875 343795
rect 19875 343765 19876 343795
rect 19844 343764 19876 343765
rect 19844 343715 19876 343716
rect 19844 343685 19845 343715
rect 19845 343685 19875 343715
rect 19875 343685 19876 343715
rect 19844 343684 19876 343685
rect 19844 343635 19876 343636
rect 19844 343605 19845 343635
rect 19845 343605 19875 343635
rect 19875 343605 19876 343635
rect 19844 343604 19876 343605
rect 19844 343555 19876 343556
rect 19844 343525 19845 343555
rect 19845 343525 19875 343555
rect 19875 343525 19876 343555
rect 19844 343524 19876 343525
rect 19844 343475 19876 343476
rect 19844 343445 19845 343475
rect 19845 343445 19875 343475
rect 19875 343445 19876 343475
rect 19844 343444 19876 343445
rect 19844 343395 19876 343396
rect 19844 343365 19845 343395
rect 19845 343365 19875 343395
rect 19875 343365 19876 343395
rect 19844 343364 19876 343365
rect 19844 343315 19876 343316
rect 19844 343285 19845 343315
rect 19845 343285 19875 343315
rect 19875 343285 19876 343315
rect 19844 343284 19876 343285
rect 19844 343235 19876 343236
rect 19844 343205 19845 343235
rect 19845 343205 19875 343235
rect 19875 343205 19876 343235
rect 19844 343204 19876 343205
rect 19844 343155 19876 343156
rect 19844 343125 19845 343155
rect 19845 343125 19875 343155
rect 19875 343125 19876 343155
rect 19844 343124 19876 343125
rect 19844 343075 19876 343076
rect 19844 343045 19845 343075
rect 19845 343045 19875 343075
rect 19875 343045 19876 343075
rect 19844 343044 19876 343045
rect 19844 342995 19876 342996
rect 19844 342965 19845 342995
rect 19845 342965 19875 342995
rect 19875 342965 19876 342995
rect 19844 342964 19876 342965
rect 19844 342915 19876 342916
rect 19844 342885 19845 342915
rect 19845 342885 19875 342915
rect 19875 342885 19876 342915
rect 19844 342884 19876 342885
rect 19844 342835 19876 342836
rect 19844 342805 19845 342835
rect 19845 342805 19875 342835
rect 19875 342805 19876 342835
rect 19844 342804 19876 342805
rect 19844 342755 19876 342756
rect 19844 342725 19845 342755
rect 19845 342725 19875 342755
rect 19875 342725 19876 342755
rect 19844 342724 19876 342725
rect 19844 342675 19876 342676
rect 19844 342645 19845 342675
rect 19845 342645 19875 342675
rect 19875 342645 19876 342675
rect 19844 342644 19876 342645
rect 19844 342595 19876 342596
rect 19844 342565 19845 342595
rect 19845 342565 19875 342595
rect 19875 342565 19876 342595
rect 19844 342564 19876 342565
rect 19844 342515 19876 342516
rect 19844 342485 19845 342515
rect 19845 342485 19875 342515
rect 19875 342485 19876 342515
rect 19844 342484 19876 342485
rect 19844 342435 19876 342436
rect 19844 342405 19845 342435
rect 19845 342405 19875 342435
rect 19875 342405 19876 342435
rect 19844 342404 19876 342405
rect 19844 342355 19876 342356
rect 19844 342325 19845 342355
rect 19845 342325 19875 342355
rect 19875 342325 19876 342355
rect 19844 342324 19876 342325
rect 19844 342275 19876 342276
rect 19844 342245 19845 342275
rect 19845 342245 19875 342275
rect 19875 342245 19876 342275
rect 19844 342244 19876 342245
rect 19844 342195 19876 342196
rect 19844 342165 19845 342195
rect 19845 342165 19875 342195
rect 19875 342165 19876 342195
rect 19844 342164 19876 342165
rect 19844 342115 19876 342116
rect 19844 342085 19845 342115
rect 19845 342085 19875 342115
rect 19875 342085 19876 342115
rect 19844 342084 19876 342085
rect 19844 342035 19876 342036
rect 19844 342005 19845 342035
rect 19845 342005 19875 342035
rect 19875 342005 19876 342035
rect 19844 342004 19876 342005
rect 19844 341955 19876 341956
rect 19844 341925 19845 341955
rect 19845 341925 19875 341955
rect 19875 341925 19876 341955
rect 19844 341924 19876 341925
rect 19844 341875 19876 341876
rect 19844 341845 19845 341875
rect 19845 341845 19875 341875
rect 19875 341845 19876 341875
rect 19844 341844 19876 341845
rect 19844 341795 19876 341796
rect 19844 341765 19845 341795
rect 19845 341765 19875 341795
rect 19875 341765 19876 341795
rect 19844 341764 19876 341765
rect 19844 341715 19876 341716
rect 19844 341685 19845 341715
rect 19845 341685 19875 341715
rect 19875 341685 19876 341715
rect 19844 341684 19876 341685
rect 19844 341635 19876 341636
rect 19844 341605 19845 341635
rect 19845 341605 19875 341635
rect 19875 341605 19876 341635
rect 19844 341604 19876 341605
rect 19844 341555 19876 341556
rect 19844 341525 19845 341555
rect 19845 341525 19875 341555
rect 19875 341525 19876 341555
rect 19844 341524 19876 341525
rect 19844 341475 19876 341476
rect 19844 341445 19845 341475
rect 19845 341445 19875 341475
rect 19875 341445 19876 341475
rect 19844 341444 19876 341445
rect 19844 341395 19876 341396
rect 19844 341365 19845 341395
rect 19845 341365 19875 341395
rect 19875 341365 19876 341395
rect 19844 341364 19876 341365
rect 19844 341315 19876 341316
rect 19844 341285 19845 341315
rect 19845 341285 19875 341315
rect 19875 341285 19876 341315
rect 19844 341284 19876 341285
rect 19844 341235 19876 341236
rect 19844 341205 19845 341235
rect 19845 341205 19875 341235
rect 19875 341205 19876 341235
rect 19844 341204 19876 341205
rect 19844 341155 19876 341156
rect 19844 341125 19845 341155
rect 19845 341125 19875 341155
rect 19875 341125 19876 341155
rect 19844 341124 19876 341125
rect 19844 341075 19876 341076
rect 19844 341045 19845 341075
rect 19845 341045 19875 341075
rect 19875 341045 19876 341075
rect 19844 341044 19876 341045
rect 19844 340995 19876 340996
rect 19844 340965 19845 340995
rect 19845 340965 19875 340995
rect 19875 340965 19876 340995
rect 19844 340964 19876 340965
rect 19844 340915 19876 340916
rect 19844 340885 19845 340915
rect 19845 340885 19875 340915
rect 19875 340885 19876 340915
rect 19844 340884 19876 340885
rect 19844 340835 19876 340836
rect 19844 340805 19845 340835
rect 19845 340805 19875 340835
rect 19875 340805 19876 340835
rect 19844 340804 19876 340805
rect 19844 340755 19876 340756
rect 19844 340725 19845 340755
rect 19845 340725 19875 340755
rect 19875 340725 19876 340755
rect 19844 340724 19876 340725
rect 19844 340675 19876 340676
rect 19844 340645 19845 340675
rect 19845 340645 19875 340675
rect 19875 340645 19876 340675
rect 19844 340644 19876 340645
rect 19844 340595 19876 340596
rect 19844 340565 19845 340595
rect 19845 340565 19875 340595
rect 19875 340565 19876 340595
rect 19844 340564 19876 340565
rect 19844 340515 19876 340516
rect 19844 340485 19845 340515
rect 19845 340485 19875 340515
rect 19875 340485 19876 340515
rect 19844 340484 19876 340485
rect 19844 340435 19876 340436
rect 19844 340405 19845 340435
rect 19845 340405 19875 340435
rect 19875 340405 19876 340435
rect 19844 340404 19876 340405
rect 19844 340355 19876 340356
rect 19844 340325 19845 340355
rect 19845 340325 19875 340355
rect 19875 340325 19876 340355
rect 19844 340324 19876 340325
rect 19844 340275 19876 340276
rect 19844 340245 19845 340275
rect 19845 340245 19875 340275
rect 19875 340245 19876 340275
rect 19844 340244 19876 340245
rect 19844 340195 19876 340196
rect 19844 340165 19845 340195
rect 19845 340165 19875 340195
rect 19875 340165 19876 340195
rect 19844 340164 19876 340165
rect 19844 340115 19876 340116
rect 19844 340085 19845 340115
rect 19845 340085 19875 340115
rect 19875 340085 19876 340115
rect 19844 340084 19876 340085
rect 19844 340035 19876 340036
rect 19844 340005 19845 340035
rect 19845 340005 19875 340035
rect 19875 340005 19876 340035
rect 19844 340004 19876 340005
rect 19844 339955 19876 339956
rect 19844 339925 19845 339955
rect 19845 339925 19875 339955
rect 19875 339925 19876 339955
rect 19844 339924 19876 339925
rect 19844 339875 19876 339876
rect 19844 339845 19845 339875
rect 19845 339845 19875 339875
rect 19875 339845 19876 339875
rect 19844 339844 19876 339845
rect 19844 339795 19876 339796
rect 19844 339765 19845 339795
rect 19845 339765 19875 339795
rect 19875 339765 19876 339795
rect 19844 339764 19876 339765
rect 19844 339715 19876 339716
rect 19844 339685 19845 339715
rect 19845 339685 19875 339715
rect 19875 339685 19876 339715
rect 19844 339684 19876 339685
rect 19844 339635 19876 339636
rect 19844 339605 19845 339635
rect 19845 339605 19875 339635
rect 19875 339605 19876 339635
rect 19844 339604 19876 339605
rect 19844 339555 19876 339556
rect 19844 339525 19845 339555
rect 19845 339525 19875 339555
rect 19875 339525 19876 339555
rect 19844 339524 19876 339525
rect 19844 339475 19876 339476
rect 19844 339445 19845 339475
rect 19845 339445 19875 339475
rect 19875 339445 19876 339475
rect 19844 339444 19876 339445
rect 19844 339395 19876 339396
rect 19844 339365 19845 339395
rect 19845 339365 19875 339395
rect 19875 339365 19876 339395
rect 19844 339364 19876 339365
rect 19844 339315 19876 339316
rect 19844 339285 19845 339315
rect 19845 339285 19875 339315
rect 19875 339285 19876 339315
rect 19844 339284 19876 339285
rect 19844 339235 19876 339236
rect 19844 339205 19845 339235
rect 19845 339205 19875 339235
rect 19875 339205 19876 339235
rect 19844 339204 19876 339205
rect 19844 339155 19876 339156
rect 19844 339125 19845 339155
rect 19845 339125 19875 339155
rect 19875 339125 19876 339155
rect 19844 339124 19876 339125
rect 19844 339075 19876 339076
rect 19844 339045 19845 339075
rect 19845 339045 19875 339075
rect 19875 339045 19876 339075
rect 19844 339044 19876 339045
rect 19844 338995 19876 338996
rect 19844 338965 19845 338995
rect 19845 338965 19875 338995
rect 19875 338965 19876 338995
rect 19844 338964 19876 338965
rect 19844 338915 19876 338916
rect 19844 338885 19845 338915
rect 19845 338885 19875 338915
rect 19875 338885 19876 338915
rect 19844 338884 19876 338885
rect 19844 338835 19876 338836
rect 19844 338805 19845 338835
rect 19845 338805 19875 338835
rect 19875 338805 19876 338835
rect 19844 338804 19876 338805
rect 19844 338755 19876 338756
rect 19844 338725 19845 338755
rect 19845 338725 19875 338755
rect 19875 338725 19876 338755
rect 19844 338724 19876 338725
rect 19844 338675 19876 338676
rect 19844 338645 19845 338675
rect 19845 338645 19875 338675
rect 19875 338645 19876 338675
rect 19844 338644 19876 338645
rect 19844 338595 19876 338596
rect 19844 338565 19845 338595
rect 19845 338565 19875 338595
rect 19875 338565 19876 338595
rect 19844 338564 19876 338565
rect 19844 338515 19876 338516
rect 19844 338485 19845 338515
rect 19845 338485 19875 338515
rect 19875 338485 19876 338515
rect 19844 338484 19876 338485
rect 19844 338435 19876 338436
rect 19844 338405 19845 338435
rect 19845 338405 19875 338435
rect 19875 338405 19876 338435
rect 19844 338404 19876 338405
rect 19844 338355 19876 338356
rect 19844 338325 19845 338355
rect 19845 338325 19875 338355
rect 19875 338325 19876 338355
rect 19844 338324 19876 338325
rect 19844 338275 19876 338276
rect 19844 338245 19845 338275
rect 19845 338245 19875 338275
rect 19875 338245 19876 338275
rect 19844 338244 19876 338245
rect 19844 338195 19876 338196
rect 19844 338165 19845 338195
rect 19845 338165 19875 338195
rect 19875 338165 19876 338195
rect 19844 338164 19876 338165
rect 19844 338115 19876 338116
rect 19844 338085 19845 338115
rect 19845 338085 19875 338115
rect 19875 338085 19876 338115
rect 19844 338084 19876 338085
rect 19844 338035 19876 338036
rect 19844 338005 19845 338035
rect 19845 338005 19875 338035
rect 19875 338005 19876 338035
rect 19844 338004 19876 338005
rect 19844 337955 19876 337956
rect 19844 337925 19845 337955
rect 19845 337925 19875 337955
rect 19875 337925 19876 337955
rect 19844 337924 19876 337925
rect 19844 337875 19876 337876
rect 19844 337845 19845 337875
rect 19845 337845 19875 337875
rect 19875 337845 19876 337875
rect 19844 337844 19876 337845
rect 19844 337795 19876 337796
rect 19844 337765 19845 337795
rect 19845 337765 19875 337795
rect 19875 337765 19876 337795
rect 19844 337764 19876 337765
rect 19844 337715 19876 337716
rect 19844 337685 19845 337715
rect 19845 337685 19875 337715
rect 19875 337685 19876 337715
rect 19844 337684 19876 337685
rect 19844 337635 19876 337636
rect 19844 337605 19845 337635
rect 19845 337605 19875 337635
rect 19875 337605 19876 337635
rect 19844 337604 19876 337605
rect 19844 337555 19876 337556
rect 19844 337525 19845 337555
rect 19845 337525 19875 337555
rect 19875 337525 19876 337555
rect 19844 337524 19876 337525
rect 19844 337475 19876 337476
rect 19844 337445 19845 337475
rect 19845 337445 19875 337475
rect 19875 337445 19876 337475
rect 19844 337444 19876 337445
rect 19844 337395 19876 337396
rect 19844 337365 19845 337395
rect 19845 337365 19875 337395
rect 19875 337365 19876 337395
rect 19844 337364 19876 337365
rect 19844 337315 19876 337316
rect 19844 337285 19845 337315
rect 19845 337285 19875 337315
rect 19875 337285 19876 337315
rect 19844 337284 19876 337285
rect 19844 337235 19876 337236
rect 19844 337205 19845 337235
rect 19845 337205 19875 337235
rect 19875 337205 19876 337235
rect 19844 337204 19876 337205
rect 19844 337155 19876 337156
rect 19844 337125 19845 337155
rect 19845 337125 19875 337155
rect 19875 337125 19876 337155
rect 19844 337124 19876 337125
rect 19844 337075 19876 337076
rect 19844 337045 19845 337075
rect 19845 337045 19875 337075
rect 19875 337045 19876 337075
rect 19844 337044 19876 337045
rect 19844 336995 19876 336996
rect 19844 336965 19845 336995
rect 19845 336965 19875 336995
rect 19875 336965 19876 336995
rect 19844 336964 19876 336965
rect 19844 336915 19876 336916
rect 19844 336885 19845 336915
rect 19845 336885 19875 336915
rect 19875 336885 19876 336915
rect 19844 336884 19876 336885
rect 19844 336835 19876 336836
rect 19844 336805 19845 336835
rect 19845 336805 19875 336835
rect 19875 336805 19876 336835
rect 19844 336804 19876 336805
rect 19844 336755 19876 336756
rect 19844 336725 19845 336755
rect 19845 336725 19875 336755
rect 19875 336725 19876 336755
rect 19844 336724 19876 336725
rect 19844 336675 19876 336676
rect 19844 336645 19845 336675
rect 19845 336645 19875 336675
rect 19875 336645 19876 336675
rect 19844 336644 19876 336645
rect 19844 336595 19876 336596
rect 19844 336565 19845 336595
rect 19845 336565 19875 336595
rect 19875 336565 19876 336595
rect 19844 336564 19876 336565
rect 19844 336515 19876 336516
rect 19844 336485 19845 336515
rect 19845 336485 19875 336515
rect 19875 336485 19876 336515
rect 19844 336484 19876 336485
rect 19844 336435 19876 336436
rect 19844 336405 19845 336435
rect 19845 336405 19875 336435
rect 19875 336405 19876 336435
rect 19844 336404 19876 336405
rect 19844 336355 19876 336356
rect 19844 336325 19845 336355
rect 19845 336325 19875 336355
rect 19875 336325 19876 336355
rect 19844 336324 19876 336325
rect 19844 336275 19876 336276
rect 19844 336245 19845 336275
rect 19845 336245 19875 336275
rect 19875 336245 19876 336275
rect 19844 336244 19876 336245
rect 19844 336195 19876 336196
rect 19844 336165 19845 336195
rect 19845 336165 19875 336195
rect 19875 336165 19876 336195
rect 19844 336164 19876 336165
rect 19844 336115 19876 336116
rect 19844 336085 19845 336115
rect 19845 336085 19875 336115
rect 19875 336085 19876 336115
rect 19844 336084 19876 336085
rect 19844 336035 19876 336036
rect 19844 336005 19845 336035
rect 19845 336005 19875 336035
rect 19875 336005 19876 336035
rect 19844 336004 19876 336005
rect 19844 335955 19876 335956
rect 19844 335925 19845 335955
rect 19845 335925 19875 335955
rect 19875 335925 19876 335955
rect 19844 335924 19876 335925
rect 19844 335875 19876 335876
rect 19844 335845 19845 335875
rect 19845 335845 19875 335875
rect 19875 335845 19876 335875
rect 19844 335844 19876 335845
rect 19844 335795 19876 335796
rect 19844 335765 19845 335795
rect 19845 335765 19875 335795
rect 19875 335765 19876 335795
rect 19844 335764 19876 335765
rect 19844 335715 19876 335716
rect 19844 335685 19845 335715
rect 19845 335685 19875 335715
rect 19875 335685 19876 335715
rect 19844 335684 19876 335685
rect 19844 335635 19876 335636
rect 19844 335605 19845 335635
rect 19845 335605 19875 335635
rect 19875 335605 19876 335635
rect 19844 335604 19876 335605
rect 19844 335555 19876 335556
rect 19844 335525 19845 335555
rect 19845 335525 19875 335555
rect 19875 335525 19876 335555
rect 19844 335524 19876 335525
rect 19844 335475 19876 335476
rect 19844 335445 19845 335475
rect 19845 335445 19875 335475
rect 19875 335445 19876 335475
rect 19844 335444 19876 335445
rect 19844 335395 19876 335396
rect 19844 335365 19845 335395
rect 19845 335365 19875 335395
rect 19875 335365 19876 335395
rect 19844 335364 19876 335365
rect 19844 335315 19876 335316
rect 19844 335285 19845 335315
rect 19845 335285 19875 335315
rect 19875 335285 19876 335315
rect 19844 335284 19876 335285
rect 19844 335235 19876 335236
rect 19844 335205 19845 335235
rect 19845 335205 19875 335235
rect 19875 335205 19876 335235
rect 19844 335204 19876 335205
rect 19844 335155 19876 335156
rect 19844 335125 19845 335155
rect 19845 335125 19875 335155
rect 19875 335125 19876 335155
rect 19844 335124 19876 335125
rect 19844 335075 19876 335076
rect 19844 335045 19845 335075
rect 19845 335045 19875 335075
rect 19875 335045 19876 335075
rect 19844 335044 19876 335045
rect 19844 334995 19876 334996
rect 19844 334965 19845 334995
rect 19845 334965 19875 334995
rect 19875 334965 19876 334995
rect 19844 334964 19876 334965
rect 19844 334915 19876 334916
rect 19844 334885 19845 334915
rect 19845 334885 19875 334915
rect 19875 334885 19876 334915
rect 19844 334884 19876 334885
rect 19844 334835 19876 334836
rect 19844 334805 19845 334835
rect 19845 334805 19875 334835
rect 19875 334805 19876 334835
rect 19844 334804 19876 334805
rect 19844 334755 19876 334756
rect 19844 334725 19845 334755
rect 19845 334725 19875 334755
rect 19875 334725 19876 334755
rect 19844 334724 19876 334725
rect 19844 334675 19876 334676
rect 19844 334645 19845 334675
rect 19845 334645 19875 334675
rect 19875 334645 19876 334675
rect 19844 334644 19876 334645
rect 19844 334595 19876 334596
rect 19844 334565 19845 334595
rect 19845 334565 19875 334595
rect 19875 334565 19876 334595
rect 19844 334564 19876 334565
rect 19844 334515 19876 334516
rect 19844 334485 19845 334515
rect 19845 334485 19875 334515
rect 19875 334485 19876 334515
rect 19844 334484 19876 334485
rect 19844 334435 19876 334436
rect 19844 334405 19845 334435
rect 19845 334405 19875 334435
rect 19875 334405 19876 334435
rect 19844 334404 19876 334405
rect 19844 334355 19876 334356
rect 19844 334325 19845 334355
rect 19845 334325 19875 334355
rect 19875 334325 19876 334355
rect 19844 334324 19876 334325
rect 19844 334275 19876 334276
rect 19844 334245 19845 334275
rect 19845 334245 19875 334275
rect 19875 334245 19876 334275
rect 19844 334244 19876 334245
rect 19844 334195 19876 334196
rect 19844 334165 19845 334195
rect 19845 334165 19875 334195
rect 19875 334165 19876 334195
rect 19844 334164 19876 334165
rect 19844 334115 19876 334116
rect 19844 334085 19845 334115
rect 19845 334085 19875 334115
rect 19875 334085 19876 334115
rect 19844 334084 19876 334085
rect 19844 334035 19876 334036
rect 19844 334005 19845 334035
rect 19845 334005 19875 334035
rect 19875 334005 19876 334035
rect 19844 334004 19876 334005
rect 19844 333955 19876 333956
rect 19844 333925 19845 333955
rect 19845 333925 19875 333955
rect 19875 333925 19876 333955
rect 19844 333924 19876 333925
rect 19844 333875 19876 333876
rect 19844 333845 19845 333875
rect 19845 333845 19875 333875
rect 19875 333845 19876 333875
rect 19844 333844 19876 333845
rect 19844 333795 19876 333796
rect 19844 333765 19845 333795
rect 19845 333765 19875 333795
rect 19875 333765 19876 333795
rect 19844 333764 19876 333765
rect 19844 333715 19876 333716
rect 19844 333685 19845 333715
rect 19845 333685 19875 333715
rect 19875 333685 19876 333715
rect 19844 333684 19876 333685
rect 19844 333635 19876 333636
rect 19844 333605 19845 333635
rect 19845 333605 19875 333635
rect 19875 333605 19876 333635
rect 19844 333604 19876 333605
rect 19844 333555 19876 333556
rect 19844 333525 19845 333555
rect 19845 333525 19875 333555
rect 19875 333525 19876 333555
rect 19844 333524 19876 333525
rect 19844 333475 19876 333476
rect 19844 333445 19845 333475
rect 19845 333445 19875 333475
rect 19875 333445 19876 333475
rect 19844 333444 19876 333445
rect 19844 333395 19876 333396
rect 19844 333365 19845 333395
rect 19845 333365 19875 333395
rect 19875 333365 19876 333395
rect 19844 333364 19876 333365
rect 19844 333315 19876 333316
rect 19844 333285 19845 333315
rect 19845 333285 19875 333315
rect 19875 333285 19876 333315
rect 19844 333284 19876 333285
rect 19844 333235 19876 333236
rect 19844 333205 19845 333235
rect 19845 333205 19875 333235
rect 19875 333205 19876 333235
rect 19844 333204 19876 333205
rect 19844 333155 19876 333156
rect 19844 333125 19845 333155
rect 19845 333125 19875 333155
rect 19875 333125 19876 333155
rect 19844 333124 19876 333125
rect 19844 333075 19876 333076
rect 19844 333045 19845 333075
rect 19845 333045 19875 333075
rect 19875 333045 19876 333075
rect 19844 333044 19876 333045
rect 19844 332995 19876 332996
rect 19844 332965 19845 332995
rect 19845 332965 19875 332995
rect 19875 332965 19876 332995
rect 19844 332964 19876 332965
rect 19844 332915 19876 332916
rect 19844 332885 19845 332915
rect 19845 332885 19875 332915
rect 19875 332885 19876 332915
rect 19844 332884 19876 332885
rect 19844 332835 19876 332836
rect 19844 332805 19845 332835
rect 19845 332805 19875 332835
rect 19875 332805 19876 332835
rect 19844 332804 19876 332805
rect 19844 332755 19876 332756
rect 19844 332725 19845 332755
rect 19845 332725 19875 332755
rect 19875 332725 19876 332755
rect 19844 332724 19876 332725
rect 19844 332675 19876 332676
rect 19844 332645 19845 332675
rect 19845 332645 19875 332675
rect 19875 332645 19876 332675
rect 19844 332644 19876 332645
rect 19844 332595 19876 332596
rect 19844 332565 19845 332595
rect 19845 332565 19875 332595
rect 19875 332565 19876 332595
rect 19844 332564 19876 332565
rect 19844 332515 19876 332516
rect 19844 332485 19845 332515
rect 19845 332485 19875 332515
rect 19875 332485 19876 332515
rect 19844 332484 19876 332485
rect 19844 332435 19876 332436
rect 19844 332405 19845 332435
rect 19845 332405 19875 332435
rect 19875 332405 19876 332435
rect 19844 332404 19876 332405
rect 19844 332355 19876 332356
rect 19844 332325 19845 332355
rect 19845 332325 19875 332355
rect 19875 332325 19876 332355
rect 19844 332324 19876 332325
rect 19844 332275 19876 332276
rect 19844 332245 19845 332275
rect 19845 332245 19875 332275
rect 19875 332245 19876 332275
rect 19844 332244 19876 332245
rect 19844 332195 19876 332196
rect 19844 332165 19845 332195
rect 19845 332165 19875 332195
rect 19875 332165 19876 332195
rect 19844 332164 19876 332165
rect 19844 332115 19876 332116
rect 19844 332085 19845 332115
rect 19845 332085 19875 332115
rect 19875 332085 19876 332115
rect 19844 332084 19876 332085
rect 19844 332035 19876 332036
rect 19844 332005 19845 332035
rect 19845 332005 19875 332035
rect 19875 332005 19876 332035
rect 19844 332004 19876 332005
rect 19844 331955 19876 331956
rect 19844 331925 19845 331955
rect 19845 331925 19875 331955
rect 19875 331925 19876 331955
rect 19844 331924 19876 331925
rect 19844 331875 19876 331876
rect 19844 331845 19845 331875
rect 19845 331845 19875 331875
rect 19875 331845 19876 331875
rect 19844 331844 19876 331845
rect 19844 331795 19876 331796
rect 19844 331765 19845 331795
rect 19845 331765 19875 331795
rect 19875 331765 19876 331795
rect 19844 331764 19876 331765
rect 19844 331715 19876 331716
rect 19844 331685 19845 331715
rect 19845 331685 19875 331715
rect 19875 331685 19876 331715
rect 19844 331684 19876 331685
rect 19844 331635 19876 331636
rect 19844 331605 19845 331635
rect 19845 331605 19875 331635
rect 19875 331605 19876 331635
rect 19844 331604 19876 331605
rect 19844 331555 19876 331556
rect 19844 331525 19845 331555
rect 19845 331525 19875 331555
rect 19875 331525 19876 331555
rect 19844 331524 19876 331525
rect 19844 331475 19876 331476
rect 19844 331445 19845 331475
rect 19845 331445 19875 331475
rect 19875 331445 19876 331475
rect 19844 331444 19876 331445
rect 19844 331395 19876 331396
rect 19844 331365 19845 331395
rect 19845 331365 19875 331395
rect 19875 331365 19876 331395
rect 19844 331364 19876 331365
rect 19844 331315 19876 331316
rect 19844 331285 19845 331315
rect 19845 331285 19875 331315
rect 19875 331285 19876 331315
rect 19844 331284 19876 331285
rect 19844 331235 19876 331236
rect 19844 331205 19845 331235
rect 19845 331205 19875 331235
rect 19875 331205 19876 331235
rect 19844 331204 19876 331205
rect 19844 331155 19876 331156
rect 19844 331125 19845 331155
rect 19845 331125 19875 331155
rect 19875 331125 19876 331155
rect 19844 331124 19876 331125
rect 19844 331075 19876 331076
rect 19844 331045 19845 331075
rect 19845 331045 19875 331075
rect 19875 331045 19876 331075
rect 19844 331044 19876 331045
rect 19844 330995 19876 330996
rect 19844 330965 19845 330995
rect 19845 330965 19875 330995
rect 19875 330965 19876 330995
rect 19844 330964 19876 330965
rect 19844 330915 19876 330916
rect 19844 330885 19845 330915
rect 19845 330885 19875 330915
rect 19875 330885 19876 330915
rect 19844 330884 19876 330885
rect 19844 330835 19876 330836
rect 19844 330805 19845 330835
rect 19845 330805 19875 330835
rect 19875 330805 19876 330835
rect 19844 330804 19876 330805
rect 19844 330755 19876 330756
rect 19844 330725 19845 330755
rect 19845 330725 19875 330755
rect 19875 330725 19876 330755
rect 19844 330724 19876 330725
rect 19844 330675 19876 330676
rect 19844 330645 19845 330675
rect 19845 330645 19875 330675
rect 19875 330645 19876 330675
rect 19844 330644 19876 330645
rect 19844 330595 19876 330596
rect 19844 330565 19845 330595
rect 19845 330565 19875 330595
rect 19875 330565 19876 330595
rect 19844 330564 19876 330565
rect 19844 330515 19876 330516
rect 19844 330485 19845 330515
rect 19845 330485 19875 330515
rect 19875 330485 19876 330515
rect 19844 330484 19876 330485
rect 19844 330435 19876 330436
rect 19844 330405 19845 330435
rect 19845 330405 19875 330435
rect 19875 330405 19876 330435
rect 19844 330404 19876 330405
rect 19844 330355 19876 330356
rect 19844 330325 19845 330355
rect 19845 330325 19875 330355
rect 19875 330325 19876 330355
rect 19844 330324 19876 330325
rect 19844 330275 19876 330276
rect 19844 330245 19845 330275
rect 19845 330245 19875 330275
rect 19875 330245 19876 330275
rect 19844 330244 19876 330245
rect 19844 330195 19876 330196
rect 19844 330165 19845 330195
rect 19845 330165 19875 330195
rect 19875 330165 19876 330195
rect 19844 330164 19876 330165
rect 19844 330115 19876 330116
rect 19844 330085 19845 330115
rect 19845 330085 19875 330115
rect 19875 330085 19876 330115
rect 19844 330084 19876 330085
rect 19844 330035 19876 330036
rect 19844 330005 19845 330035
rect 19845 330005 19875 330035
rect 19875 330005 19876 330035
rect 19844 330004 19876 330005
rect 19844 329955 19876 329956
rect 19844 329925 19845 329955
rect 19845 329925 19875 329955
rect 19875 329925 19876 329955
rect 19844 329924 19876 329925
rect 19844 329875 19876 329876
rect 19844 329845 19845 329875
rect 19845 329845 19875 329875
rect 19875 329845 19876 329875
rect 19844 329844 19876 329845
rect 19844 329795 19876 329796
rect 19844 329765 19845 329795
rect 19845 329765 19875 329795
rect 19875 329765 19876 329795
rect 19844 329764 19876 329765
rect 19844 329715 19876 329716
rect 19844 329685 19845 329715
rect 19845 329685 19875 329715
rect 19875 329685 19876 329715
rect 19844 329684 19876 329685
rect 19844 329635 19876 329636
rect 19844 329605 19845 329635
rect 19845 329605 19875 329635
rect 19875 329605 19876 329635
rect 19844 329604 19876 329605
rect 19844 329555 19876 329556
rect 19844 329525 19845 329555
rect 19845 329525 19875 329555
rect 19875 329525 19876 329555
rect 19844 329524 19876 329525
rect 19844 329475 19876 329476
rect 19844 329445 19845 329475
rect 19845 329445 19875 329475
rect 19875 329445 19876 329475
rect 19844 329444 19876 329445
rect 19844 329395 19876 329396
rect 19844 329365 19845 329395
rect 19845 329365 19875 329395
rect 19875 329365 19876 329395
rect 19844 329364 19876 329365
rect 19844 329315 19876 329316
rect 19844 329285 19845 329315
rect 19845 329285 19875 329315
rect 19875 329285 19876 329315
rect 19844 329284 19876 329285
rect 19844 329235 19876 329236
rect 19844 329205 19845 329235
rect 19845 329205 19875 329235
rect 19875 329205 19876 329235
rect 19844 329204 19876 329205
rect 19844 329155 19876 329156
rect 19844 329125 19845 329155
rect 19845 329125 19875 329155
rect 19875 329125 19876 329155
rect 19844 329124 19876 329125
rect 19844 329075 19876 329076
rect 19844 329045 19845 329075
rect 19845 329045 19875 329075
rect 19875 329045 19876 329075
rect 19844 329044 19876 329045
rect 19844 328995 19876 328996
rect 19844 328965 19845 328995
rect 19845 328965 19875 328995
rect 19875 328965 19876 328995
rect 19844 328964 19876 328965
rect 19844 328915 19876 328916
rect 19844 328885 19845 328915
rect 19845 328885 19875 328915
rect 19875 328885 19876 328915
rect 19844 328884 19876 328885
rect 19844 328835 19876 328836
rect 19844 328805 19845 328835
rect 19845 328805 19875 328835
rect 19875 328805 19876 328835
rect 19844 328804 19876 328805
rect 19844 328755 19876 328756
rect 19844 328725 19845 328755
rect 19845 328725 19875 328755
rect 19875 328725 19876 328755
rect 19844 328724 19876 328725
rect 19844 328675 19876 328676
rect 19844 328645 19845 328675
rect 19845 328645 19875 328675
rect 19875 328645 19876 328675
rect 19844 328644 19876 328645
rect 19844 328595 19876 328596
rect 19844 328565 19845 328595
rect 19845 328565 19875 328595
rect 19875 328565 19876 328595
rect 19844 328564 19876 328565
rect 19844 328515 19876 328516
rect 19844 328485 19845 328515
rect 19845 328485 19875 328515
rect 19875 328485 19876 328515
rect 19844 328484 19876 328485
rect 19844 328435 19876 328436
rect 19844 328405 19845 328435
rect 19845 328405 19875 328435
rect 19875 328405 19876 328435
rect 19844 328404 19876 328405
rect 19844 328355 19876 328356
rect 19844 328325 19845 328355
rect 19845 328325 19875 328355
rect 19875 328325 19876 328355
rect 19844 328324 19876 328325
rect 19844 328275 19876 328276
rect 19844 328245 19845 328275
rect 19845 328245 19875 328275
rect 19875 328245 19876 328275
rect 19844 328244 19876 328245
rect 19844 328195 19876 328196
rect 19844 328165 19845 328195
rect 19845 328165 19875 328195
rect 19875 328165 19876 328195
rect 19844 328164 19876 328165
rect 19844 328115 19876 328116
rect 19844 328085 19845 328115
rect 19845 328085 19875 328115
rect 19875 328085 19876 328115
rect 19844 328084 19876 328085
rect 19844 328035 19876 328036
rect 19844 328005 19845 328035
rect 19845 328005 19875 328035
rect 19875 328005 19876 328035
rect 19844 328004 19876 328005
rect 19844 327955 19876 327956
rect 19844 327925 19845 327955
rect 19845 327925 19875 327955
rect 19875 327925 19876 327955
rect 19844 327924 19876 327925
rect 19844 327875 19876 327876
rect 19844 327845 19845 327875
rect 19845 327845 19875 327875
rect 19875 327845 19876 327875
rect 19844 327844 19876 327845
rect 19844 327795 19876 327796
rect 19844 327765 19845 327795
rect 19845 327765 19875 327795
rect 19875 327765 19876 327795
rect 19844 327764 19876 327765
rect 19844 327715 19876 327716
rect 19844 327685 19845 327715
rect 19845 327685 19875 327715
rect 19875 327685 19876 327715
rect 19844 327684 19876 327685
rect 19844 327635 19876 327636
rect 19844 327605 19845 327635
rect 19845 327605 19875 327635
rect 19875 327605 19876 327635
rect 19844 327604 19876 327605
rect 19844 327555 19876 327556
rect 19844 327525 19845 327555
rect 19845 327525 19875 327555
rect 19875 327525 19876 327555
rect 19844 327524 19876 327525
rect 19844 327475 19876 327476
rect 19844 327445 19845 327475
rect 19845 327445 19875 327475
rect 19875 327445 19876 327475
rect 19844 327444 19876 327445
rect 19844 327395 19876 327396
rect 19844 327365 19845 327395
rect 19845 327365 19875 327395
rect 19875 327365 19876 327395
rect 19844 327364 19876 327365
rect 19844 327315 19876 327316
rect 19844 327285 19845 327315
rect 19845 327285 19875 327315
rect 19875 327285 19876 327315
rect 19844 327284 19876 327285
rect 19844 327235 19876 327236
rect 19844 327205 19845 327235
rect 19845 327205 19875 327235
rect 19875 327205 19876 327235
rect 19844 327204 19876 327205
rect 19844 327155 19876 327156
rect 19844 327125 19845 327155
rect 19845 327125 19875 327155
rect 19875 327125 19876 327155
rect 19844 327124 19876 327125
rect 19844 327075 19876 327076
rect 19844 327045 19845 327075
rect 19845 327045 19875 327075
rect 19875 327045 19876 327075
rect 19844 327044 19876 327045
rect 19844 326995 19876 326996
rect 19844 326965 19845 326995
rect 19845 326965 19875 326995
rect 19875 326965 19876 326995
rect 19844 326964 19876 326965
rect 19844 326915 19876 326916
rect 19844 326885 19845 326915
rect 19845 326885 19875 326915
rect 19875 326885 19876 326915
rect 19844 326884 19876 326885
rect 19844 326835 19876 326836
rect 19844 326805 19845 326835
rect 19845 326805 19875 326835
rect 19875 326805 19876 326835
rect 19844 326804 19876 326805
rect 19844 326755 19876 326756
rect 19844 326725 19845 326755
rect 19845 326725 19875 326755
rect 19875 326725 19876 326755
rect 19844 326724 19876 326725
rect 19844 326675 19876 326676
rect 19844 326645 19845 326675
rect 19845 326645 19875 326675
rect 19875 326645 19876 326675
rect 19844 326644 19876 326645
rect 19844 326595 19876 326596
rect 19844 326565 19845 326595
rect 19845 326565 19875 326595
rect 19875 326565 19876 326595
rect 19844 326564 19876 326565
rect 19844 326515 19876 326516
rect 19844 326485 19845 326515
rect 19845 326485 19875 326515
rect 19875 326485 19876 326515
rect 19844 326484 19876 326485
rect 19844 326435 19876 326436
rect 19844 326405 19845 326435
rect 19845 326405 19875 326435
rect 19875 326405 19876 326435
rect 19844 326404 19876 326405
rect 19844 326355 19876 326356
rect 19844 326325 19845 326355
rect 19845 326325 19875 326355
rect 19875 326325 19876 326355
rect 19844 326324 19876 326325
rect 19844 326275 19876 326276
rect 19844 326245 19845 326275
rect 19845 326245 19875 326275
rect 19875 326245 19876 326275
rect 19844 326244 19876 326245
rect 19844 326195 19876 326196
rect 19844 326165 19845 326195
rect 19845 326165 19875 326195
rect 19875 326165 19876 326195
rect 19844 326164 19876 326165
rect 19844 326115 19876 326116
rect 19844 326085 19845 326115
rect 19845 326085 19875 326115
rect 19875 326085 19876 326115
rect 19844 326084 19876 326085
rect 19844 326035 19876 326036
rect 19844 326005 19845 326035
rect 19845 326005 19875 326035
rect 19875 326005 19876 326035
rect 19844 326004 19876 326005
rect 19844 325955 19876 325956
rect 19844 325925 19845 325955
rect 19845 325925 19875 325955
rect 19875 325925 19876 325955
rect 19844 325924 19876 325925
rect 19844 325875 19876 325876
rect 19844 325845 19845 325875
rect 19845 325845 19875 325875
rect 19875 325845 19876 325875
rect 19844 325844 19876 325845
rect 19844 325795 19876 325796
rect 19844 325765 19845 325795
rect 19845 325765 19875 325795
rect 19875 325765 19876 325795
rect 19844 325764 19876 325765
rect 19844 325715 19876 325716
rect 19844 325685 19845 325715
rect 19845 325685 19875 325715
rect 19875 325685 19876 325715
rect 19844 325684 19876 325685
rect 19844 325635 19876 325636
rect 19844 325605 19845 325635
rect 19845 325605 19875 325635
rect 19875 325605 19876 325635
rect 19844 325604 19876 325605
rect 19844 325555 19876 325556
rect 19844 325525 19845 325555
rect 19845 325525 19875 325555
rect 19875 325525 19876 325555
rect 19844 325524 19876 325525
rect 19844 325475 19876 325476
rect 19844 325445 19845 325475
rect 19845 325445 19875 325475
rect 19875 325445 19876 325475
rect 19844 325444 19876 325445
rect 19844 325395 19876 325396
rect 19844 325365 19845 325395
rect 19845 325365 19875 325395
rect 19875 325365 19876 325395
rect 19844 325364 19876 325365
rect 19844 325315 19876 325316
rect 19844 325285 19845 325315
rect 19845 325285 19875 325315
rect 19875 325285 19876 325315
rect 19844 325284 19876 325285
rect 19844 325235 19876 325236
rect 19844 325205 19845 325235
rect 19845 325205 19875 325235
rect 19875 325205 19876 325235
rect 19844 325204 19876 325205
rect 19844 325155 19876 325156
rect 19844 325125 19845 325155
rect 19845 325125 19875 325155
rect 19875 325125 19876 325155
rect 19844 325124 19876 325125
rect 19844 325075 19876 325076
rect 19844 325045 19845 325075
rect 19845 325045 19875 325075
rect 19875 325045 19876 325075
rect 19844 325044 19876 325045
rect 19844 324995 19876 324996
rect 19844 324965 19845 324995
rect 19845 324965 19875 324995
rect 19875 324965 19876 324995
rect 19844 324964 19876 324965
rect 19844 324915 19876 324916
rect 19844 324885 19845 324915
rect 19845 324885 19875 324915
rect 19875 324885 19876 324915
rect 19844 324884 19876 324885
rect 19844 324835 19876 324836
rect 19844 324805 19845 324835
rect 19845 324805 19875 324835
rect 19875 324805 19876 324835
rect 19844 324804 19876 324805
rect 19844 324755 19876 324756
rect 19844 324725 19845 324755
rect 19845 324725 19875 324755
rect 19875 324725 19876 324755
rect 19844 324724 19876 324725
rect 19844 324675 19876 324676
rect 19844 324645 19845 324675
rect 19845 324645 19875 324675
rect 19875 324645 19876 324675
rect 19844 324644 19876 324645
rect 19844 324595 19876 324596
rect 19844 324565 19845 324595
rect 19845 324565 19875 324595
rect 19875 324565 19876 324595
rect 19844 324564 19876 324565
rect 19844 324515 19876 324516
rect 19844 324485 19845 324515
rect 19845 324485 19875 324515
rect 19875 324485 19876 324515
rect 19844 324484 19876 324485
rect 19844 324435 19876 324436
rect 19844 324405 19845 324435
rect 19845 324405 19875 324435
rect 19875 324405 19876 324435
rect 19844 324404 19876 324405
rect 19844 324355 19876 324356
rect 19844 324325 19845 324355
rect 19845 324325 19875 324355
rect 19875 324325 19876 324355
rect 19844 324324 19876 324325
rect 19844 324275 19876 324276
rect 19844 324245 19845 324275
rect 19845 324245 19875 324275
rect 19875 324245 19876 324275
rect 19844 324244 19876 324245
rect 19844 324195 19876 324196
rect 19844 324165 19845 324195
rect 19845 324165 19875 324195
rect 19875 324165 19876 324195
rect 19844 324164 19876 324165
rect 19844 324115 19876 324116
rect 19844 324085 19845 324115
rect 19845 324085 19875 324115
rect 19875 324085 19876 324115
rect 19844 324084 19876 324085
rect 19844 324035 19876 324036
rect 19844 324005 19845 324035
rect 19845 324005 19875 324035
rect 19875 324005 19876 324035
rect 19844 324004 19876 324005
rect 19844 323955 19876 323956
rect 19844 323925 19845 323955
rect 19845 323925 19875 323955
rect 19875 323925 19876 323955
rect 19844 323924 19876 323925
rect 19844 323875 19876 323876
rect 19844 323845 19845 323875
rect 19845 323845 19875 323875
rect 19875 323845 19876 323875
rect 19844 323844 19876 323845
rect 19844 323795 19876 323796
rect 19844 323765 19845 323795
rect 19845 323765 19875 323795
rect 19875 323765 19876 323795
rect 19844 323764 19876 323765
rect 19844 323715 19876 323716
rect 19844 323685 19845 323715
rect 19845 323685 19875 323715
rect 19875 323685 19876 323715
rect 19844 323684 19876 323685
rect 19844 323635 19876 323636
rect 19844 323605 19845 323635
rect 19845 323605 19875 323635
rect 19875 323605 19876 323635
rect 19844 323604 19876 323605
rect 19844 323555 19876 323556
rect 19844 323525 19845 323555
rect 19845 323525 19875 323555
rect 19875 323525 19876 323555
rect 19844 323524 19876 323525
rect 19844 323475 19876 323476
rect 19844 323445 19845 323475
rect 19845 323445 19875 323475
rect 19875 323445 19876 323475
rect 19844 323444 19876 323445
rect 19844 323395 19876 323396
rect 19844 323365 19845 323395
rect 19845 323365 19875 323395
rect 19875 323365 19876 323395
rect 19844 323364 19876 323365
rect 19844 323315 19876 323316
rect 19844 323285 19845 323315
rect 19845 323285 19875 323315
rect 19875 323285 19876 323315
rect 19844 323284 19876 323285
rect 19844 323235 19876 323236
rect 19844 323205 19845 323235
rect 19845 323205 19875 323235
rect 19875 323205 19876 323235
rect 19844 323204 19876 323205
rect 19844 323155 19876 323156
rect 19844 323125 19845 323155
rect 19845 323125 19875 323155
rect 19875 323125 19876 323155
rect 19844 323124 19876 323125
rect 19844 323075 19876 323076
rect 19844 323045 19845 323075
rect 19845 323045 19875 323075
rect 19875 323045 19876 323075
rect 19844 323044 19876 323045
rect 19844 322995 19876 322996
rect 19844 322965 19845 322995
rect 19845 322965 19875 322995
rect 19875 322965 19876 322995
rect 19844 322964 19876 322965
rect 19844 322915 19876 322916
rect 19844 322885 19845 322915
rect 19845 322885 19875 322915
rect 19875 322885 19876 322915
rect 19844 322884 19876 322885
rect 19844 322835 19876 322836
rect 19844 322805 19845 322835
rect 19845 322805 19875 322835
rect 19875 322805 19876 322835
rect 19844 322804 19876 322805
rect 19844 322755 19876 322756
rect 19844 322725 19845 322755
rect 19845 322725 19875 322755
rect 19875 322725 19876 322755
rect 19844 322724 19876 322725
rect 19844 322675 19876 322676
rect 19844 322645 19845 322675
rect 19845 322645 19875 322675
rect 19875 322645 19876 322675
rect 19844 322644 19876 322645
rect 19844 322595 19876 322596
rect 19844 322565 19845 322595
rect 19845 322565 19875 322595
rect 19875 322565 19876 322595
rect 19844 322564 19876 322565
rect 19844 322515 19876 322516
rect 19844 322485 19845 322515
rect 19845 322485 19875 322515
rect 19875 322485 19876 322515
rect 19844 322484 19876 322485
rect 19844 322435 19876 322436
rect 19844 322405 19845 322435
rect 19845 322405 19875 322435
rect 19875 322405 19876 322435
rect 19844 322404 19876 322405
rect 19844 322355 19876 322356
rect 19844 322325 19845 322355
rect 19845 322325 19875 322355
rect 19875 322325 19876 322355
rect 19844 322324 19876 322325
rect 19844 322275 19876 322276
rect 19844 322245 19845 322275
rect 19845 322245 19875 322275
rect 19875 322245 19876 322275
rect 19844 322244 19876 322245
rect 19844 322195 19876 322196
rect 19844 322165 19845 322195
rect 19845 322165 19875 322195
rect 19875 322165 19876 322195
rect 19844 322164 19876 322165
rect 19844 322115 19876 322116
rect 19844 322085 19845 322115
rect 19845 322085 19875 322115
rect 19875 322085 19876 322115
rect 19844 322084 19876 322085
rect 19844 322035 19876 322036
rect 19844 322005 19845 322035
rect 19845 322005 19875 322035
rect 19875 322005 19876 322035
rect 19844 322004 19876 322005
rect 19844 321955 19876 321956
rect 19844 321925 19845 321955
rect 19845 321925 19875 321955
rect 19875 321925 19876 321955
rect 19844 321924 19876 321925
rect 19844 321875 19876 321876
rect 19844 321845 19845 321875
rect 19845 321845 19875 321875
rect 19875 321845 19876 321875
rect 19844 321844 19876 321845
rect 19844 321795 19876 321796
rect 19844 321765 19845 321795
rect 19845 321765 19875 321795
rect 19875 321765 19876 321795
rect 19844 321764 19876 321765
rect 19844 321715 19876 321716
rect 19844 321685 19845 321715
rect 19845 321685 19875 321715
rect 19875 321685 19876 321715
rect 19844 321684 19876 321685
rect 19844 321635 19876 321636
rect 19844 321605 19845 321635
rect 19845 321605 19875 321635
rect 19875 321605 19876 321635
rect 19844 321604 19876 321605
rect 19844 321555 19876 321556
rect 19844 321525 19845 321555
rect 19845 321525 19875 321555
rect 19875 321525 19876 321555
rect 19844 321524 19876 321525
rect 19844 321475 19876 321476
rect 19844 321445 19845 321475
rect 19845 321445 19875 321475
rect 19875 321445 19876 321475
rect 19844 321444 19876 321445
rect 19844 321395 19876 321396
rect 19844 321365 19845 321395
rect 19845 321365 19875 321395
rect 19875 321365 19876 321395
rect 19844 321364 19876 321365
rect 19844 321315 19876 321316
rect 19844 321285 19845 321315
rect 19845 321285 19875 321315
rect 19875 321285 19876 321315
rect 19844 321284 19876 321285
rect 19844 321235 19876 321236
rect 19844 321205 19845 321235
rect 19845 321205 19875 321235
rect 19875 321205 19876 321235
rect 19844 321204 19876 321205
rect 19844 321155 19876 321156
rect 19844 321125 19845 321155
rect 19845 321125 19875 321155
rect 19875 321125 19876 321155
rect 19844 321124 19876 321125
rect 19844 321075 19876 321076
rect 19844 321045 19845 321075
rect 19845 321045 19875 321075
rect 19875 321045 19876 321075
rect 19844 321044 19876 321045
rect 19844 320995 19876 320996
rect 19844 320965 19845 320995
rect 19845 320965 19875 320995
rect 19875 320965 19876 320995
rect 19844 320964 19876 320965
rect 19844 320915 19876 320916
rect 19844 320885 19845 320915
rect 19845 320885 19875 320915
rect 19875 320885 19876 320915
rect 19844 320884 19876 320885
rect 19844 320835 19876 320836
rect 19844 320805 19845 320835
rect 19845 320805 19875 320835
rect 19875 320805 19876 320835
rect 19844 320804 19876 320805
rect 19844 320755 19876 320756
rect 19844 320725 19845 320755
rect 19845 320725 19875 320755
rect 19875 320725 19876 320755
rect 19844 320724 19876 320725
rect 19844 320675 19876 320676
rect 19844 320645 19845 320675
rect 19845 320645 19875 320675
rect 19875 320645 19876 320675
rect 19844 320644 19876 320645
rect 19844 320595 19876 320596
rect 19844 320565 19845 320595
rect 19845 320565 19875 320595
rect 19875 320565 19876 320595
rect 19844 320564 19876 320565
rect 19844 320515 19876 320516
rect 19844 320485 19845 320515
rect 19845 320485 19875 320515
rect 19875 320485 19876 320515
rect 19844 320484 19876 320485
rect 19844 320435 19876 320436
rect 19844 320405 19845 320435
rect 19845 320405 19875 320435
rect 19875 320405 19876 320435
rect 19844 320404 19876 320405
rect 19844 320355 19876 320356
rect 19844 320325 19845 320355
rect 19845 320325 19875 320355
rect 19875 320325 19876 320355
rect 19844 320324 19876 320325
rect 19844 320275 19876 320276
rect 19844 320245 19845 320275
rect 19845 320245 19875 320275
rect 19875 320245 19876 320275
rect 19844 320244 19876 320245
rect 19844 320195 19876 320196
rect 19844 320165 19845 320195
rect 19845 320165 19875 320195
rect 19875 320165 19876 320195
rect 19844 320164 19876 320165
rect 19844 320115 19876 320116
rect 19844 320085 19845 320115
rect 19845 320085 19875 320115
rect 19875 320085 19876 320115
rect 19844 320084 19876 320085
rect 19844 320035 19876 320036
rect 19844 320005 19845 320035
rect 19845 320005 19875 320035
rect 19875 320005 19876 320035
rect 19844 320004 19876 320005
rect 19844 319955 19876 319956
rect 19844 319925 19845 319955
rect 19845 319925 19875 319955
rect 19875 319925 19876 319955
rect 19844 319924 19876 319925
rect 19844 319875 19876 319876
rect 19844 319845 19845 319875
rect 19845 319845 19875 319875
rect 19875 319845 19876 319875
rect 19844 319844 19876 319845
rect 19844 319795 19876 319796
rect 19844 319765 19845 319795
rect 19845 319765 19875 319795
rect 19875 319765 19876 319795
rect 19844 319764 19876 319765
rect 19844 319715 19876 319716
rect 19844 319685 19845 319715
rect 19845 319685 19875 319715
rect 19875 319685 19876 319715
rect 19844 319684 19876 319685
rect 19844 319635 19876 319636
rect 19844 319605 19845 319635
rect 19845 319605 19875 319635
rect 19875 319605 19876 319635
rect 19844 319604 19876 319605
rect 19844 319555 19876 319556
rect 19844 319525 19845 319555
rect 19845 319525 19875 319555
rect 19875 319525 19876 319555
rect 19844 319524 19876 319525
rect 19844 319475 19876 319476
rect 19844 319445 19845 319475
rect 19845 319445 19875 319475
rect 19875 319445 19876 319475
rect 19844 319444 19876 319445
rect 19844 319395 19876 319396
rect 19844 319365 19845 319395
rect 19845 319365 19875 319395
rect 19875 319365 19876 319395
rect 19844 319364 19876 319365
rect 19844 319315 19876 319316
rect 19844 319285 19845 319315
rect 19845 319285 19875 319315
rect 19875 319285 19876 319315
rect 19844 319284 19876 319285
rect 19844 319235 19876 319236
rect 19844 319205 19845 319235
rect 19845 319205 19875 319235
rect 19875 319205 19876 319235
rect 19844 319204 19876 319205
rect 19844 319155 19876 319156
rect 19844 319125 19845 319155
rect 19845 319125 19875 319155
rect 19875 319125 19876 319155
rect 19844 319124 19876 319125
rect 19844 319075 19876 319076
rect 19844 319045 19845 319075
rect 19845 319045 19875 319075
rect 19875 319045 19876 319075
rect 19844 319044 19876 319045
rect 19844 318995 19876 318996
rect 19844 318965 19845 318995
rect 19845 318965 19875 318995
rect 19875 318965 19876 318995
rect 19844 318964 19876 318965
rect 19844 318915 19876 318916
rect 19844 318885 19845 318915
rect 19845 318885 19875 318915
rect 19875 318885 19876 318915
rect 19844 318884 19876 318885
rect 19844 318835 19876 318836
rect 19844 318805 19845 318835
rect 19845 318805 19875 318835
rect 19875 318805 19876 318835
rect 19844 318804 19876 318805
rect 19844 318755 19876 318756
rect 19844 318725 19845 318755
rect 19845 318725 19875 318755
rect 19875 318725 19876 318755
rect 19844 318724 19876 318725
rect 19844 318675 19876 318676
rect 19844 318645 19845 318675
rect 19845 318645 19875 318675
rect 19875 318645 19876 318675
rect 19844 318644 19876 318645
rect 19844 318595 19876 318596
rect 19844 318565 19845 318595
rect 19845 318565 19875 318595
rect 19875 318565 19876 318595
rect 19844 318564 19876 318565
rect 19844 318515 19876 318516
rect 19844 318485 19845 318515
rect 19845 318485 19875 318515
rect 19875 318485 19876 318515
rect 19844 318484 19876 318485
rect 19844 318435 19876 318436
rect 19844 318405 19845 318435
rect 19845 318405 19875 318435
rect 19875 318405 19876 318435
rect 19844 318404 19876 318405
rect 19844 318355 19876 318356
rect 19844 318325 19845 318355
rect 19845 318325 19875 318355
rect 19875 318325 19876 318355
rect 19844 318324 19876 318325
rect 19844 318275 19876 318276
rect 19844 318245 19845 318275
rect 19845 318245 19875 318275
rect 19875 318245 19876 318275
rect 19844 318244 19876 318245
rect 19844 318195 19876 318196
rect 19844 318165 19845 318195
rect 19845 318165 19875 318195
rect 19875 318165 19876 318195
rect 19844 318164 19876 318165
rect 19844 318115 19876 318116
rect 19844 318085 19845 318115
rect 19845 318085 19875 318115
rect 19875 318085 19876 318115
rect 19844 318084 19876 318085
rect 19844 318035 19876 318036
rect 19844 318005 19845 318035
rect 19845 318005 19875 318035
rect 19875 318005 19876 318035
rect 19844 318004 19876 318005
rect 19844 317955 19876 317956
rect 19844 317925 19845 317955
rect 19845 317925 19875 317955
rect 19875 317925 19876 317955
rect 19844 317924 19876 317925
rect 19844 317875 19876 317876
rect 19844 317845 19845 317875
rect 19845 317845 19875 317875
rect 19875 317845 19876 317875
rect 19844 317844 19876 317845
rect 19844 317795 19876 317796
rect 19844 317765 19845 317795
rect 19845 317765 19875 317795
rect 19875 317765 19876 317795
rect 19844 317764 19876 317765
rect 19844 317715 19876 317716
rect 19844 317685 19845 317715
rect 19845 317685 19875 317715
rect 19875 317685 19876 317715
rect 19844 317684 19876 317685
rect 19844 317635 19876 317636
rect 19844 317605 19845 317635
rect 19845 317605 19875 317635
rect 19875 317605 19876 317635
rect 19844 317604 19876 317605
rect 19844 317555 19876 317556
rect 19844 317525 19845 317555
rect 19845 317525 19875 317555
rect 19875 317525 19876 317555
rect 19844 317524 19876 317525
rect 19844 317475 19876 317476
rect 19844 317445 19845 317475
rect 19845 317445 19875 317475
rect 19875 317445 19876 317475
rect 19844 317444 19876 317445
rect 19844 317395 19876 317396
rect 19844 317365 19845 317395
rect 19845 317365 19875 317395
rect 19875 317365 19876 317395
rect 19844 317364 19876 317365
rect 19844 317315 19876 317316
rect 19844 317285 19845 317315
rect 19845 317285 19875 317315
rect 19875 317285 19876 317315
rect 19844 317284 19876 317285
rect 19844 317235 19876 317236
rect 19844 317205 19845 317235
rect 19845 317205 19875 317235
rect 19875 317205 19876 317235
rect 19844 317204 19876 317205
rect 19844 317155 19876 317156
rect 19844 317125 19845 317155
rect 19845 317125 19875 317155
rect 19875 317125 19876 317155
rect 19844 317124 19876 317125
rect 19844 317075 19876 317076
rect 19844 317045 19845 317075
rect 19845 317045 19875 317075
rect 19875 317045 19876 317075
rect 19844 317044 19876 317045
rect 19844 316995 19876 316996
rect 19844 316965 19845 316995
rect 19845 316965 19875 316995
rect 19875 316965 19876 316995
rect 19844 316964 19876 316965
rect 19844 316915 19876 316916
rect 19844 316885 19845 316915
rect 19845 316885 19875 316915
rect 19875 316885 19876 316915
rect 19844 316884 19876 316885
rect 19844 316835 19876 316836
rect 19844 316805 19845 316835
rect 19845 316805 19875 316835
rect 19875 316805 19876 316835
rect 19844 316804 19876 316805
rect 19844 316755 19876 316756
rect 19844 316725 19845 316755
rect 19845 316725 19875 316755
rect 19875 316725 19876 316755
rect 19844 316724 19876 316725
rect 19844 316675 19876 316676
rect 19844 316645 19845 316675
rect 19845 316645 19875 316675
rect 19875 316645 19876 316675
rect 19844 316644 19876 316645
rect 19844 316595 19876 316596
rect 19844 316565 19845 316595
rect 19845 316565 19875 316595
rect 19875 316565 19876 316595
rect 19844 316564 19876 316565
rect 19844 316515 19876 316516
rect 19844 316485 19845 316515
rect 19845 316485 19875 316515
rect 19875 316485 19876 316515
rect 19844 316484 19876 316485
rect 19844 316435 19876 316436
rect 19844 316405 19845 316435
rect 19845 316405 19875 316435
rect 19875 316405 19876 316435
rect 19844 316404 19876 316405
rect 19844 316355 19876 316356
rect 19844 316325 19845 316355
rect 19845 316325 19875 316355
rect 19875 316325 19876 316355
rect 19844 316324 19876 316325
rect 19844 316275 19876 316276
rect 19844 316245 19845 316275
rect 19845 316245 19875 316275
rect 19875 316245 19876 316275
rect 19844 316244 19876 316245
rect 19844 316195 19876 316196
rect 19844 316165 19845 316195
rect 19845 316165 19875 316195
rect 19875 316165 19876 316195
rect 19844 316164 19876 316165
rect 19844 316115 19876 316116
rect 19844 316085 19845 316115
rect 19845 316085 19875 316115
rect 19875 316085 19876 316115
rect 19844 316084 19876 316085
rect 19844 316035 19876 316036
rect 19844 316005 19845 316035
rect 19845 316005 19875 316035
rect 19875 316005 19876 316035
rect 19844 316004 19876 316005
rect 19844 315955 19876 315956
rect 19844 315925 19845 315955
rect 19845 315925 19875 315955
rect 19875 315925 19876 315955
rect 19844 315924 19876 315925
rect 19844 315875 19876 315876
rect 19844 315845 19845 315875
rect 19845 315845 19875 315875
rect 19875 315845 19876 315875
rect 19844 315844 19876 315845
rect 19844 315795 19876 315796
rect 19844 315765 19845 315795
rect 19845 315765 19875 315795
rect 19875 315765 19876 315795
rect 19844 315764 19876 315765
rect 19844 315715 19876 315716
rect 19844 315685 19845 315715
rect 19845 315685 19875 315715
rect 19875 315685 19876 315715
rect 19844 315684 19876 315685
rect 19844 315635 19876 315636
rect 19844 315605 19845 315635
rect 19845 315605 19875 315635
rect 19875 315605 19876 315635
rect 19844 315604 19876 315605
rect 19844 315555 19876 315556
rect 19844 315525 19845 315555
rect 19845 315525 19875 315555
rect 19875 315525 19876 315555
rect 19844 315524 19876 315525
rect 19844 315475 19876 315476
rect 19844 315445 19845 315475
rect 19845 315445 19875 315475
rect 19875 315445 19876 315475
rect 19844 315444 19876 315445
rect 19844 315395 19876 315396
rect 19844 315365 19845 315395
rect 19845 315365 19875 315395
rect 19875 315365 19876 315395
rect 19844 315364 19876 315365
rect 19844 315315 19876 315316
rect 19844 315285 19845 315315
rect 19845 315285 19875 315315
rect 19875 315285 19876 315315
rect 19844 315284 19876 315285
rect 19844 315235 19876 315236
rect 19844 315205 19845 315235
rect 19845 315205 19875 315235
rect 19875 315205 19876 315235
rect 19844 315204 19876 315205
rect 19844 315155 19876 315156
rect 19844 315125 19845 315155
rect 19845 315125 19875 315155
rect 19875 315125 19876 315155
rect 19844 315124 19876 315125
rect 19844 315075 19876 315076
rect 19844 315045 19845 315075
rect 19845 315045 19875 315075
rect 19875 315045 19876 315075
rect 19844 315044 19876 315045
rect 19844 314995 19876 314996
rect 19844 314965 19845 314995
rect 19845 314965 19875 314995
rect 19875 314965 19876 314995
rect 19844 314964 19876 314965
rect 19844 314915 19876 314916
rect 19844 314885 19845 314915
rect 19845 314885 19875 314915
rect 19875 314885 19876 314915
rect 19844 314884 19876 314885
rect 19844 314835 19876 314836
rect 19844 314805 19845 314835
rect 19845 314805 19875 314835
rect 19875 314805 19876 314835
rect 19844 314804 19876 314805
rect 19844 314755 19876 314756
rect 19844 314725 19845 314755
rect 19845 314725 19875 314755
rect 19875 314725 19876 314755
rect 19844 314724 19876 314725
rect 19844 314675 19876 314676
rect 19844 314645 19845 314675
rect 19845 314645 19875 314675
rect 19875 314645 19876 314675
rect 19844 314644 19876 314645
rect 19844 314595 19876 314596
rect 19844 314565 19845 314595
rect 19845 314565 19875 314595
rect 19875 314565 19876 314595
rect 19844 314564 19876 314565
rect 19844 314515 19876 314516
rect 19844 314485 19845 314515
rect 19845 314485 19875 314515
rect 19875 314485 19876 314515
rect 19844 314484 19876 314485
rect 19844 314435 19876 314436
rect 19844 314405 19845 314435
rect 19845 314405 19875 314435
rect 19875 314405 19876 314435
rect 19844 314404 19876 314405
rect 19844 314355 19876 314356
rect 19844 314325 19845 314355
rect 19845 314325 19875 314355
rect 19875 314325 19876 314355
rect 19844 314324 19876 314325
rect 19844 314275 19876 314276
rect 19844 314245 19845 314275
rect 19845 314245 19875 314275
rect 19875 314245 19876 314275
rect 19844 314244 19876 314245
rect 19844 314195 19876 314196
rect 19844 314165 19845 314195
rect 19845 314165 19875 314195
rect 19875 314165 19876 314195
rect 19844 314164 19876 314165
rect 19844 314115 19876 314116
rect 19844 314085 19845 314115
rect 19845 314085 19875 314115
rect 19875 314085 19876 314115
rect 19844 314084 19876 314085
rect 19844 314035 19876 314036
rect 19844 314005 19845 314035
rect 19845 314005 19875 314035
rect 19875 314005 19876 314035
rect 19844 314004 19876 314005
rect 19844 313955 19876 313956
rect 19844 313925 19845 313955
rect 19845 313925 19875 313955
rect 19875 313925 19876 313955
rect 19844 313924 19876 313925
rect 19844 313875 19876 313876
rect 19844 313845 19845 313875
rect 19845 313845 19875 313875
rect 19875 313845 19876 313875
rect 19844 313844 19876 313845
rect 19844 313795 19876 313796
rect 19844 313765 19845 313795
rect 19845 313765 19875 313795
rect 19875 313765 19876 313795
rect 19844 313764 19876 313765
rect 19844 313715 19876 313716
rect 19844 313685 19845 313715
rect 19845 313685 19875 313715
rect 19875 313685 19876 313715
rect 19844 313684 19876 313685
rect 19844 313635 19876 313636
rect 19844 313605 19845 313635
rect 19845 313605 19875 313635
rect 19875 313605 19876 313635
rect 19844 313604 19876 313605
rect 19844 313555 19876 313556
rect 19844 313525 19845 313555
rect 19845 313525 19875 313555
rect 19875 313525 19876 313555
rect 19844 313524 19876 313525
rect 19844 313475 19876 313476
rect 19844 313445 19845 313475
rect 19845 313445 19875 313475
rect 19875 313445 19876 313475
rect 19844 313444 19876 313445
rect 19844 313395 19876 313396
rect 19844 313365 19845 313395
rect 19845 313365 19875 313395
rect 19875 313365 19876 313395
rect 19844 313364 19876 313365
rect 19844 313315 19876 313316
rect 19844 313285 19845 313315
rect 19845 313285 19875 313315
rect 19875 313285 19876 313315
rect 19844 313284 19876 313285
rect 19844 313235 19876 313236
rect 19844 313205 19845 313235
rect 19845 313205 19875 313235
rect 19875 313205 19876 313235
rect 19844 313204 19876 313205
rect 19844 313155 19876 313156
rect 19844 313125 19845 313155
rect 19845 313125 19875 313155
rect 19875 313125 19876 313155
rect 19844 313124 19876 313125
rect 19844 313075 19876 313076
rect 19844 313045 19845 313075
rect 19845 313045 19875 313075
rect 19875 313045 19876 313075
rect 19844 313044 19876 313045
rect 19844 312995 19876 312996
rect 19844 312965 19845 312995
rect 19845 312965 19875 312995
rect 19875 312965 19876 312995
rect 19844 312964 19876 312965
rect 19844 312915 19876 312916
rect 19844 312885 19845 312915
rect 19845 312885 19875 312915
rect 19875 312885 19876 312915
rect 19844 312884 19876 312885
rect 19844 312835 19876 312836
rect 19844 312805 19845 312835
rect 19845 312805 19875 312835
rect 19875 312805 19876 312835
rect 19844 312804 19876 312805
rect 19844 312755 19876 312756
rect 19844 312725 19845 312755
rect 19845 312725 19875 312755
rect 19875 312725 19876 312755
rect 19844 312724 19876 312725
rect 19844 312675 19876 312676
rect 19844 312645 19845 312675
rect 19845 312645 19875 312675
rect 19875 312645 19876 312675
rect 19844 312644 19876 312645
rect 19844 312595 19876 312596
rect 19844 312565 19845 312595
rect 19845 312565 19875 312595
rect 19875 312565 19876 312595
rect 19844 312564 19876 312565
rect 19844 312515 19876 312516
rect 19844 312485 19845 312515
rect 19845 312485 19875 312515
rect 19875 312485 19876 312515
rect 19844 312484 19876 312485
rect 19844 312435 19876 312436
rect 19844 312405 19845 312435
rect 19845 312405 19875 312435
rect 19875 312405 19876 312435
rect 19844 312404 19876 312405
rect 19844 312355 19876 312356
rect 19844 312325 19845 312355
rect 19845 312325 19875 312355
rect 19875 312325 19876 312355
rect 19844 312324 19876 312325
rect 19844 312275 19876 312276
rect 19844 312245 19845 312275
rect 19845 312245 19875 312275
rect 19875 312245 19876 312275
rect 19844 312244 19876 312245
rect 19844 312195 19876 312196
rect 19844 312165 19845 312195
rect 19845 312165 19875 312195
rect 19875 312165 19876 312195
rect 19844 312164 19876 312165
rect 19844 312115 19876 312116
rect 19844 312085 19845 312115
rect 19845 312085 19875 312115
rect 19875 312085 19876 312115
rect 19844 312084 19876 312085
rect 19844 312035 19876 312036
rect 19844 312005 19845 312035
rect 19845 312005 19875 312035
rect 19875 312005 19876 312035
rect 19844 312004 19876 312005
rect 19844 311955 19876 311956
rect 19844 311925 19845 311955
rect 19845 311925 19875 311955
rect 19875 311925 19876 311955
rect 19844 311924 19876 311925
rect 19844 311875 19876 311876
rect 19844 311845 19845 311875
rect 19845 311845 19875 311875
rect 19875 311845 19876 311875
rect 19844 311844 19876 311845
rect 19844 311795 19876 311796
rect 19844 311765 19845 311795
rect 19845 311765 19875 311795
rect 19875 311765 19876 311795
rect 19844 311764 19876 311765
rect 19844 311715 19876 311716
rect 19844 311685 19845 311715
rect 19845 311685 19875 311715
rect 19875 311685 19876 311715
rect 19844 311684 19876 311685
rect 19844 311635 19876 311636
rect 19844 311605 19845 311635
rect 19845 311605 19875 311635
rect 19875 311605 19876 311635
rect 19844 311604 19876 311605
rect 19844 311555 19876 311556
rect 19844 311525 19845 311555
rect 19845 311525 19875 311555
rect 19875 311525 19876 311555
rect 19844 311524 19876 311525
rect 19844 311475 19876 311476
rect 19844 311445 19845 311475
rect 19845 311445 19875 311475
rect 19875 311445 19876 311475
rect 19844 311444 19876 311445
rect 19844 311395 19876 311396
rect 19844 311365 19845 311395
rect 19845 311365 19875 311395
rect 19875 311365 19876 311395
rect 19844 311364 19876 311365
rect 19844 311315 19876 311316
rect 19844 311285 19845 311315
rect 19845 311285 19875 311315
rect 19875 311285 19876 311315
rect 19844 311284 19876 311285
rect 19844 311235 19876 311236
rect 19844 311205 19845 311235
rect 19845 311205 19875 311235
rect 19875 311205 19876 311235
rect 19844 311204 19876 311205
rect 19844 311155 19876 311156
rect 19844 311125 19845 311155
rect 19845 311125 19875 311155
rect 19875 311125 19876 311155
rect 19844 311124 19876 311125
rect 19844 311075 19876 311076
rect 19844 311045 19845 311075
rect 19845 311045 19875 311075
rect 19875 311045 19876 311075
rect 19844 311044 19876 311045
rect 19844 310995 19876 310996
rect 19844 310965 19845 310995
rect 19845 310965 19875 310995
rect 19875 310965 19876 310995
rect 19844 310964 19876 310965
rect 19844 310915 19876 310916
rect 19844 310885 19845 310915
rect 19845 310885 19875 310915
rect 19875 310885 19876 310915
rect 19844 310884 19876 310885
rect 19844 310835 19876 310836
rect 19844 310805 19845 310835
rect 19845 310805 19875 310835
rect 19875 310805 19876 310835
rect 19844 310804 19876 310805
rect 19844 310755 19876 310756
rect 19844 310725 19845 310755
rect 19845 310725 19875 310755
rect 19875 310725 19876 310755
rect 19844 310724 19876 310725
rect 19844 310675 19876 310676
rect 19844 310645 19845 310675
rect 19845 310645 19875 310675
rect 19875 310645 19876 310675
rect 19844 310644 19876 310645
rect 19844 310595 19876 310596
rect 19844 310565 19845 310595
rect 19845 310565 19875 310595
rect 19875 310565 19876 310595
rect 19844 310564 19876 310565
rect 19844 310515 19876 310516
rect 19844 310485 19845 310515
rect 19845 310485 19875 310515
rect 19875 310485 19876 310515
rect 19844 310484 19876 310485
rect 19844 310435 19876 310436
rect 19844 310405 19845 310435
rect 19845 310405 19875 310435
rect 19875 310405 19876 310435
rect 19844 310404 19876 310405
rect 19844 310355 19876 310356
rect 19844 310325 19845 310355
rect 19845 310325 19875 310355
rect 19875 310325 19876 310355
rect 19844 310324 19876 310325
rect 19844 310275 19876 310276
rect 19844 310245 19845 310275
rect 19845 310245 19875 310275
rect 19875 310245 19876 310275
rect 19844 310244 19876 310245
rect 19844 310195 19876 310196
rect 19844 310165 19845 310195
rect 19845 310165 19875 310195
rect 19875 310165 19876 310195
rect 19844 310164 19876 310165
rect 19844 310115 19876 310116
rect 19844 310085 19845 310115
rect 19845 310085 19875 310115
rect 19875 310085 19876 310115
rect 19844 310084 19876 310085
rect 19844 310035 19876 310036
rect 19844 310005 19845 310035
rect 19845 310005 19875 310035
rect 19875 310005 19876 310035
rect 19844 310004 19876 310005
rect 19844 309955 19876 309956
rect 19844 309925 19845 309955
rect 19845 309925 19875 309955
rect 19875 309925 19876 309955
rect 19844 309924 19876 309925
rect 19844 309875 19876 309876
rect 19844 309845 19845 309875
rect 19845 309845 19875 309875
rect 19875 309845 19876 309875
rect 19844 309844 19876 309845
rect 19844 309795 19876 309796
rect 19844 309765 19845 309795
rect 19845 309765 19875 309795
rect 19875 309765 19876 309795
rect 19844 309764 19876 309765
rect 19844 309715 19876 309716
rect 19844 309685 19845 309715
rect 19845 309685 19875 309715
rect 19875 309685 19876 309715
rect 19844 309684 19876 309685
rect 19844 309635 19876 309636
rect 19844 309605 19845 309635
rect 19845 309605 19875 309635
rect 19875 309605 19876 309635
rect 19844 309604 19876 309605
rect 19844 309555 19876 309556
rect 19844 309525 19845 309555
rect 19845 309525 19875 309555
rect 19875 309525 19876 309555
rect 19844 309524 19876 309525
rect 19844 309475 19876 309476
rect 19844 309445 19845 309475
rect 19845 309445 19875 309475
rect 19875 309445 19876 309475
rect 19844 309444 19876 309445
rect 19844 309395 19876 309396
rect 19844 309365 19845 309395
rect 19845 309365 19875 309395
rect 19875 309365 19876 309395
rect 19844 309364 19876 309365
rect 19844 309315 19876 309316
rect 19844 309285 19845 309315
rect 19845 309285 19875 309315
rect 19875 309285 19876 309315
rect 19844 309284 19876 309285
rect 19844 309235 19876 309236
rect 19844 309205 19845 309235
rect 19845 309205 19875 309235
rect 19875 309205 19876 309235
rect 19844 309204 19876 309205
rect 19844 309155 19876 309156
rect 19844 309125 19845 309155
rect 19845 309125 19875 309155
rect 19875 309125 19876 309155
rect 19844 309124 19876 309125
rect 19844 309075 19876 309076
rect 19844 309045 19845 309075
rect 19845 309045 19875 309075
rect 19875 309045 19876 309075
rect 19844 309044 19876 309045
rect 19844 308995 19876 308996
rect 19844 308965 19845 308995
rect 19845 308965 19875 308995
rect 19875 308965 19876 308995
rect 19844 308964 19876 308965
rect 19844 308915 19876 308916
rect 19844 308885 19845 308915
rect 19845 308885 19875 308915
rect 19875 308885 19876 308915
rect 19844 308884 19876 308885
rect 19844 308835 19876 308836
rect 19844 308805 19845 308835
rect 19845 308805 19875 308835
rect 19875 308805 19876 308835
rect 19844 308804 19876 308805
rect 19844 308755 19876 308756
rect 19844 308725 19845 308755
rect 19845 308725 19875 308755
rect 19875 308725 19876 308755
rect 19844 308724 19876 308725
rect 19844 308675 19876 308676
rect 19844 308645 19845 308675
rect 19845 308645 19875 308675
rect 19875 308645 19876 308675
rect 19844 308644 19876 308645
rect 19844 308595 19876 308596
rect 19844 308565 19845 308595
rect 19845 308565 19875 308595
rect 19875 308565 19876 308595
rect 19844 308564 19876 308565
rect 19844 308515 19876 308516
rect 19844 308485 19845 308515
rect 19845 308485 19875 308515
rect 19875 308485 19876 308515
rect 19844 308484 19876 308485
rect 19844 308435 19876 308436
rect 19844 308405 19845 308435
rect 19845 308405 19875 308435
rect 19875 308405 19876 308435
rect 19844 308404 19876 308405
rect 19844 308355 19876 308356
rect 19844 308325 19845 308355
rect 19845 308325 19875 308355
rect 19875 308325 19876 308355
rect 19844 308324 19876 308325
rect 19844 308275 19876 308276
rect 19844 308245 19845 308275
rect 19845 308245 19875 308275
rect 19875 308245 19876 308275
rect 19844 308244 19876 308245
rect 19844 308195 19876 308196
rect 19844 308165 19845 308195
rect 19845 308165 19875 308195
rect 19875 308165 19876 308195
rect 19844 308164 19876 308165
rect 19844 308115 19876 308116
rect 19844 308085 19845 308115
rect 19845 308085 19875 308115
rect 19875 308085 19876 308115
rect 19844 308084 19876 308085
rect 19844 308035 19876 308036
rect 19844 308005 19845 308035
rect 19845 308005 19875 308035
rect 19875 308005 19876 308035
rect 19844 308004 19876 308005
rect 19844 307955 19876 307956
rect 19844 307925 19845 307955
rect 19845 307925 19875 307955
rect 19875 307925 19876 307955
rect 19844 307924 19876 307925
rect 19844 307875 19876 307876
rect 19844 307845 19845 307875
rect 19845 307845 19875 307875
rect 19875 307845 19876 307875
rect 19844 307844 19876 307845
rect 19844 307795 19876 307796
rect 19844 307765 19845 307795
rect 19845 307765 19875 307795
rect 19875 307765 19876 307795
rect 19844 307764 19876 307765
rect 19844 307715 19876 307716
rect 19844 307685 19845 307715
rect 19845 307685 19875 307715
rect 19875 307685 19876 307715
rect 19844 307684 19876 307685
rect 19844 307635 19876 307636
rect 19844 307605 19845 307635
rect 19845 307605 19875 307635
rect 19875 307605 19876 307635
rect 19844 307604 19876 307605
rect 19844 307555 19876 307556
rect 19844 307525 19845 307555
rect 19845 307525 19875 307555
rect 19875 307525 19876 307555
rect 19844 307524 19876 307525
rect 19844 307475 19876 307476
rect 19844 307445 19845 307475
rect 19845 307445 19875 307475
rect 19875 307445 19876 307475
rect 19844 307444 19876 307445
rect 19844 307395 19876 307396
rect 19844 307365 19845 307395
rect 19845 307365 19875 307395
rect 19875 307365 19876 307395
rect 19844 307364 19876 307365
rect 19844 307315 19876 307316
rect 19844 307285 19845 307315
rect 19845 307285 19875 307315
rect 19875 307285 19876 307315
rect 19844 307284 19876 307285
rect 19844 307235 19876 307236
rect 19844 307205 19845 307235
rect 19845 307205 19875 307235
rect 19875 307205 19876 307235
rect 19844 307204 19876 307205
rect 19844 307155 19876 307156
rect 19844 307125 19845 307155
rect 19845 307125 19875 307155
rect 19875 307125 19876 307155
rect 19844 307124 19876 307125
rect 19844 307075 19876 307076
rect 19844 307045 19845 307075
rect 19845 307045 19875 307075
rect 19875 307045 19876 307075
rect 19844 307044 19876 307045
rect 19844 306995 19876 306996
rect 19844 306965 19845 306995
rect 19845 306965 19875 306995
rect 19875 306965 19876 306995
rect 19844 306964 19876 306965
rect 19844 306915 19876 306916
rect 19844 306885 19845 306915
rect 19845 306885 19875 306915
rect 19875 306885 19876 306915
rect 19844 306884 19876 306885
rect 19844 306835 19876 306836
rect 19844 306805 19845 306835
rect 19845 306805 19875 306835
rect 19875 306805 19876 306835
rect 19844 306804 19876 306805
rect 19844 306755 19876 306756
rect 19844 306725 19845 306755
rect 19845 306725 19875 306755
rect 19875 306725 19876 306755
rect 19844 306724 19876 306725
rect 19844 306675 19876 306676
rect 19844 306645 19845 306675
rect 19845 306645 19875 306675
rect 19875 306645 19876 306675
rect 19844 306644 19876 306645
rect 19844 306595 19876 306596
rect 19844 306565 19845 306595
rect 19845 306565 19875 306595
rect 19875 306565 19876 306595
rect 19844 306564 19876 306565
rect 19844 306515 19876 306516
rect 19844 306485 19845 306515
rect 19845 306485 19875 306515
rect 19875 306485 19876 306515
rect 19844 306484 19876 306485
rect 19844 306435 19876 306436
rect 19844 306405 19845 306435
rect 19845 306405 19875 306435
rect 19875 306405 19876 306435
rect 19844 306404 19876 306405
rect 19844 306355 19876 306356
rect 19844 306325 19845 306355
rect 19845 306325 19875 306355
rect 19875 306325 19876 306355
rect 19844 306324 19876 306325
rect 19844 306275 19876 306276
rect 19844 306245 19845 306275
rect 19845 306245 19875 306275
rect 19875 306245 19876 306275
rect 19844 306244 19876 306245
rect 19844 306195 19876 306196
rect 19844 306165 19845 306195
rect 19845 306165 19875 306195
rect 19875 306165 19876 306195
rect 19844 306164 19876 306165
rect 19844 306115 19876 306116
rect 19844 306085 19845 306115
rect 19845 306085 19875 306115
rect 19875 306085 19876 306115
rect 19844 306084 19876 306085
rect 19844 306035 19876 306036
rect 19844 306005 19845 306035
rect 19845 306005 19875 306035
rect 19875 306005 19876 306035
rect 19844 306004 19876 306005
rect 19844 305955 19876 305956
rect 19844 305925 19845 305955
rect 19845 305925 19875 305955
rect 19875 305925 19876 305955
rect 19844 305924 19876 305925
rect 19844 305875 19876 305876
rect 19844 305845 19845 305875
rect 19845 305845 19875 305875
rect 19875 305845 19876 305875
rect 19844 305844 19876 305845
rect 19844 305795 19876 305796
rect 19844 305765 19845 305795
rect 19845 305765 19875 305795
rect 19875 305765 19876 305795
rect 19844 305764 19876 305765
rect 19844 305715 19876 305716
rect 19844 305685 19845 305715
rect 19845 305685 19875 305715
rect 19875 305685 19876 305715
rect 19844 305684 19876 305685
rect 19844 305635 19876 305636
rect 19844 305605 19845 305635
rect 19845 305605 19875 305635
rect 19875 305605 19876 305635
rect 19844 305604 19876 305605
rect 19844 305555 19876 305556
rect 19844 305525 19845 305555
rect 19845 305525 19875 305555
rect 19875 305525 19876 305555
rect 19844 305524 19876 305525
rect 19844 305475 19876 305476
rect 19844 305445 19845 305475
rect 19845 305445 19875 305475
rect 19875 305445 19876 305475
rect 19844 305444 19876 305445
rect 19844 305395 19876 305396
rect 19844 305365 19845 305395
rect 19845 305365 19875 305395
rect 19875 305365 19876 305395
rect 19844 305364 19876 305365
rect 19844 305315 19876 305316
rect 19844 305285 19845 305315
rect 19845 305285 19875 305315
rect 19875 305285 19876 305315
rect 19844 305284 19876 305285
rect 19844 305235 19876 305236
rect 19844 305205 19845 305235
rect 19845 305205 19875 305235
rect 19875 305205 19876 305235
rect 19844 305204 19876 305205
rect 19844 305155 19876 305156
rect 19844 305125 19845 305155
rect 19845 305125 19875 305155
rect 19875 305125 19876 305155
rect 19844 305124 19876 305125
rect 19844 305075 19876 305076
rect 19844 305045 19845 305075
rect 19845 305045 19875 305075
rect 19875 305045 19876 305075
rect 19844 305044 19876 305045
rect 19844 304995 19876 304996
rect 19844 304965 19845 304995
rect 19845 304965 19875 304995
rect 19875 304965 19876 304995
rect 19844 304964 19876 304965
rect 19844 304915 19876 304916
rect 19844 304885 19845 304915
rect 19845 304885 19875 304915
rect 19875 304885 19876 304915
rect 19844 304884 19876 304885
rect 19844 304835 19876 304836
rect 19844 304805 19845 304835
rect 19845 304805 19875 304835
rect 19875 304805 19876 304835
rect 19844 304804 19876 304805
rect 19844 304755 19876 304756
rect 19844 304725 19845 304755
rect 19845 304725 19875 304755
rect 19875 304725 19876 304755
rect 19844 304724 19876 304725
rect 19844 304675 19876 304676
rect 19844 304645 19845 304675
rect 19845 304645 19875 304675
rect 19875 304645 19876 304675
rect 19844 304644 19876 304645
rect 19844 304595 19876 304596
rect 19844 304565 19845 304595
rect 19845 304565 19875 304595
rect 19875 304565 19876 304595
rect 19844 304564 19876 304565
rect 19844 304515 19876 304516
rect 19844 304485 19845 304515
rect 19845 304485 19875 304515
rect 19875 304485 19876 304515
rect 19844 304484 19876 304485
rect 19844 304435 19876 304436
rect 19844 304405 19845 304435
rect 19845 304405 19875 304435
rect 19875 304405 19876 304435
rect 19844 304404 19876 304405
rect 19844 304355 19876 304356
rect 19844 304325 19845 304355
rect 19845 304325 19875 304355
rect 19875 304325 19876 304355
rect 19844 304324 19876 304325
rect 19844 304275 19876 304276
rect 19844 304245 19845 304275
rect 19845 304245 19875 304275
rect 19875 304245 19876 304275
rect 19844 304244 19876 304245
rect 19844 304195 19876 304196
rect 19844 304165 19845 304195
rect 19845 304165 19875 304195
rect 19875 304165 19876 304195
rect 19844 304164 19876 304165
rect 19844 304115 19876 304116
rect 19844 304085 19845 304115
rect 19845 304085 19875 304115
rect 19875 304085 19876 304115
rect 19844 304084 19876 304085
rect 19844 304035 19876 304036
rect 19844 304005 19845 304035
rect 19845 304005 19875 304035
rect 19875 304005 19876 304035
rect 19844 304004 19876 304005
rect 19844 303955 19876 303956
rect 19844 303925 19845 303955
rect 19845 303925 19875 303955
rect 19875 303925 19876 303955
rect 19844 303924 19876 303925
rect 19844 303875 19876 303876
rect 19844 303845 19845 303875
rect 19845 303845 19875 303875
rect 19875 303845 19876 303875
rect 19844 303844 19876 303845
rect 19844 303795 19876 303796
rect 19844 303765 19845 303795
rect 19845 303765 19875 303795
rect 19875 303765 19876 303795
rect 19844 303764 19876 303765
rect 19844 303715 19876 303716
rect 19844 303685 19845 303715
rect 19845 303685 19875 303715
rect 19875 303685 19876 303715
rect 19844 303684 19876 303685
rect 19844 303635 19876 303636
rect 19844 303605 19845 303635
rect 19845 303605 19875 303635
rect 19875 303605 19876 303635
rect 19844 303604 19876 303605
rect 19844 303555 19876 303556
rect 19844 303525 19845 303555
rect 19845 303525 19875 303555
rect 19875 303525 19876 303555
rect 19844 303524 19876 303525
rect 19844 303475 19876 303476
rect 19844 303445 19845 303475
rect 19845 303445 19875 303475
rect 19875 303445 19876 303475
rect 19844 303444 19876 303445
rect 19844 303395 19876 303396
rect 19844 303365 19845 303395
rect 19845 303365 19875 303395
rect 19875 303365 19876 303395
rect 19844 303364 19876 303365
rect 19844 303315 19876 303316
rect 19844 303285 19845 303315
rect 19845 303285 19875 303315
rect 19875 303285 19876 303315
rect 19844 303284 19876 303285
rect 19844 303235 19876 303236
rect 19844 303205 19845 303235
rect 19845 303205 19875 303235
rect 19875 303205 19876 303235
rect 19844 303204 19876 303205
rect 19844 303155 19876 303156
rect 19844 303125 19845 303155
rect 19845 303125 19875 303155
rect 19875 303125 19876 303155
rect 19844 303124 19876 303125
rect 19844 303075 19876 303076
rect 19844 303045 19845 303075
rect 19845 303045 19875 303075
rect 19875 303045 19876 303075
rect 19844 303044 19876 303045
rect 19844 302995 19876 302996
rect 19844 302965 19845 302995
rect 19845 302965 19875 302995
rect 19875 302965 19876 302995
rect 19844 302964 19876 302965
rect 19844 302915 19876 302916
rect 19844 302885 19845 302915
rect 19845 302885 19875 302915
rect 19875 302885 19876 302915
rect 19844 302884 19876 302885
rect 19844 302835 19876 302836
rect 19844 302805 19845 302835
rect 19845 302805 19875 302835
rect 19875 302805 19876 302835
rect 19844 302804 19876 302805
rect 19844 302755 19876 302756
rect 19844 302725 19845 302755
rect 19845 302725 19875 302755
rect 19875 302725 19876 302755
rect 19844 302724 19876 302725
rect 19844 302675 19876 302676
rect 19844 302645 19845 302675
rect 19845 302645 19875 302675
rect 19875 302645 19876 302675
rect 19844 302644 19876 302645
rect 19844 302595 19876 302596
rect 19844 302565 19845 302595
rect 19845 302565 19875 302595
rect 19875 302565 19876 302595
rect 19844 302564 19876 302565
rect 19844 302515 19876 302516
rect 19844 302485 19845 302515
rect 19845 302485 19875 302515
rect 19875 302485 19876 302515
rect 19844 302484 19876 302485
rect 19844 302435 19876 302436
rect 19844 302405 19845 302435
rect 19845 302405 19875 302435
rect 19875 302405 19876 302435
rect 19844 302404 19876 302405
rect 19844 302355 19876 302356
rect 19844 302325 19845 302355
rect 19845 302325 19875 302355
rect 19875 302325 19876 302355
rect 19844 302324 19876 302325
rect 19844 302275 19876 302276
rect 19844 302245 19845 302275
rect 19845 302245 19875 302275
rect 19875 302245 19876 302275
rect 19844 302244 19876 302245
rect 19844 302195 19876 302196
rect 19844 302165 19845 302195
rect 19845 302165 19875 302195
rect 19875 302165 19876 302195
rect 19844 302164 19876 302165
rect 19844 302115 19876 302116
rect 19844 302085 19845 302115
rect 19845 302085 19875 302115
rect 19875 302085 19876 302115
rect 19844 302084 19876 302085
rect 19844 302035 19876 302036
rect 19844 302005 19845 302035
rect 19845 302005 19875 302035
rect 19875 302005 19876 302035
rect 19844 302004 19876 302005
rect 19844 301955 19876 301956
rect 19844 301925 19845 301955
rect 19845 301925 19875 301955
rect 19875 301925 19876 301955
rect 19844 301924 19876 301925
rect 19844 301875 19876 301876
rect 19844 301845 19845 301875
rect 19845 301845 19875 301875
rect 19875 301845 19876 301875
rect 19844 301844 19876 301845
rect 19844 301795 19876 301796
rect 19844 301765 19845 301795
rect 19845 301765 19875 301795
rect 19875 301765 19876 301795
rect 19844 301764 19876 301765
rect 19844 301715 19876 301716
rect 19844 301685 19845 301715
rect 19845 301685 19875 301715
rect 19875 301685 19876 301715
rect 19844 301684 19876 301685
rect 19844 301635 19876 301636
rect 19844 301605 19845 301635
rect 19845 301605 19875 301635
rect 19875 301605 19876 301635
rect 19844 301604 19876 301605
rect 19844 301555 19876 301556
rect 19844 301525 19845 301555
rect 19845 301525 19875 301555
rect 19875 301525 19876 301555
rect 19844 301524 19876 301525
rect 19844 301475 19876 301476
rect 19844 301445 19845 301475
rect 19845 301445 19875 301475
rect 19875 301445 19876 301475
rect 19844 301444 19876 301445
rect 19844 301395 19876 301396
rect 19844 301365 19845 301395
rect 19845 301365 19875 301395
rect 19875 301365 19876 301395
rect 19844 301364 19876 301365
rect 19844 301315 19876 301316
rect 19844 301285 19845 301315
rect 19845 301285 19875 301315
rect 19875 301285 19876 301315
rect 19844 301284 19876 301285
rect 19844 301235 19876 301236
rect 19844 301205 19845 301235
rect 19845 301205 19875 301235
rect 19875 301205 19876 301235
rect 19844 301204 19876 301205
rect 19844 301155 19876 301156
rect 19844 301125 19845 301155
rect 19845 301125 19875 301155
rect 19875 301125 19876 301155
rect 19844 301124 19876 301125
rect 19844 301075 19876 301076
rect 19844 301045 19845 301075
rect 19845 301045 19875 301075
rect 19875 301045 19876 301075
rect 19844 301044 19876 301045
rect 19844 300995 19876 300996
rect 19844 300965 19845 300995
rect 19845 300965 19875 300995
rect 19875 300965 19876 300995
rect 19844 300964 19876 300965
rect 19844 300915 19876 300916
rect 19844 300885 19845 300915
rect 19845 300885 19875 300915
rect 19875 300885 19876 300915
rect 19844 300884 19876 300885
rect 19844 300835 19876 300836
rect 19844 300805 19845 300835
rect 19845 300805 19875 300835
rect 19875 300805 19876 300835
rect 19844 300804 19876 300805
rect 19844 300755 19876 300756
rect 19844 300725 19845 300755
rect 19845 300725 19875 300755
rect 19875 300725 19876 300755
rect 19844 300724 19876 300725
rect 19844 300675 19876 300676
rect 19844 300645 19845 300675
rect 19845 300645 19875 300675
rect 19875 300645 19876 300675
rect 19844 300644 19876 300645
rect 19844 300595 19876 300596
rect 19844 300565 19845 300595
rect 19845 300565 19875 300595
rect 19875 300565 19876 300595
rect 19844 300564 19876 300565
rect 19844 300515 19876 300516
rect 19844 300485 19845 300515
rect 19845 300485 19875 300515
rect 19875 300485 19876 300515
rect 19844 300484 19876 300485
rect 19844 300435 19876 300436
rect 19844 300405 19845 300435
rect 19845 300405 19875 300435
rect 19875 300405 19876 300435
rect 19844 300404 19876 300405
rect 19844 300355 19876 300356
rect 19844 300325 19845 300355
rect 19845 300325 19875 300355
rect 19875 300325 19876 300355
rect 19844 300324 19876 300325
rect 19844 300275 19876 300276
rect 19844 300245 19845 300275
rect 19845 300245 19875 300275
rect 19875 300245 19876 300275
rect 19844 300244 19876 300245
rect 19844 300195 19876 300196
rect 19844 300165 19845 300195
rect 19845 300165 19875 300195
rect 19875 300165 19876 300195
rect 19844 300164 19876 300165
rect 19844 300115 19876 300116
rect 19844 300085 19845 300115
rect 19845 300085 19875 300115
rect 19875 300085 19876 300115
rect 19844 300084 19876 300085
rect 19844 300035 19876 300036
rect 19844 300005 19845 300035
rect 19845 300005 19875 300035
rect 19875 300005 19876 300035
rect 19844 300004 19876 300005
rect 19844 299955 19876 299956
rect 19844 299925 19845 299955
rect 19845 299925 19875 299955
rect 19875 299925 19876 299955
rect 19844 299924 19876 299925
rect 19844 299875 19876 299876
rect 19844 299845 19845 299875
rect 19845 299845 19875 299875
rect 19875 299845 19876 299875
rect 19844 299844 19876 299845
rect 19844 299795 19876 299796
rect 19844 299765 19845 299795
rect 19845 299765 19875 299795
rect 19875 299765 19876 299795
rect 19844 299764 19876 299765
rect 19844 299715 19876 299716
rect 19844 299685 19845 299715
rect 19845 299685 19875 299715
rect 19875 299685 19876 299715
rect 19844 299684 19876 299685
rect 19844 299635 19876 299636
rect 19844 299605 19845 299635
rect 19845 299605 19875 299635
rect 19875 299605 19876 299635
rect 19844 299604 19876 299605
rect 19844 299555 19876 299556
rect 19844 299525 19845 299555
rect 19845 299525 19875 299555
rect 19875 299525 19876 299555
rect 19844 299524 19876 299525
rect 19844 299475 19876 299476
rect 19844 299445 19845 299475
rect 19845 299445 19875 299475
rect 19875 299445 19876 299475
rect 19844 299444 19876 299445
rect 19844 299395 19876 299396
rect 19844 299365 19845 299395
rect 19845 299365 19875 299395
rect 19875 299365 19876 299395
rect 19844 299364 19876 299365
rect 19844 299315 19876 299316
rect 19844 299285 19845 299315
rect 19845 299285 19875 299315
rect 19875 299285 19876 299315
rect 19844 299284 19876 299285
rect 19844 299235 19876 299236
rect 19844 299205 19845 299235
rect 19845 299205 19875 299235
rect 19875 299205 19876 299235
rect 19844 299204 19876 299205
rect 19844 299155 19876 299156
rect 19844 299125 19845 299155
rect 19845 299125 19875 299155
rect 19875 299125 19876 299155
rect 19844 299124 19876 299125
rect 19844 299075 19876 299076
rect 19844 299045 19845 299075
rect 19845 299045 19875 299075
rect 19875 299045 19876 299075
rect 19844 299044 19876 299045
rect 19844 298995 19876 298996
rect 19844 298965 19845 298995
rect 19845 298965 19875 298995
rect 19875 298965 19876 298995
rect 19844 298964 19876 298965
rect 19844 298915 19876 298916
rect 19844 298885 19845 298915
rect 19845 298885 19875 298915
rect 19875 298885 19876 298915
rect 19844 298884 19876 298885
rect 19844 298835 19876 298836
rect 19844 298805 19845 298835
rect 19845 298805 19875 298835
rect 19875 298805 19876 298835
rect 19844 298804 19876 298805
rect 19844 298755 19876 298756
rect 19844 298725 19845 298755
rect 19845 298725 19875 298755
rect 19875 298725 19876 298755
rect 19844 298724 19876 298725
rect 19844 298675 19876 298676
rect 19844 298645 19845 298675
rect 19845 298645 19875 298675
rect 19875 298645 19876 298675
rect 19844 298644 19876 298645
rect 19844 298595 19876 298596
rect 19844 298565 19845 298595
rect 19845 298565 19875 298595
rect 19875 298565 19876 298595
rect 19844 298564 19876 298565
rect 19844 298515 19876 298516
rect 19844 298485 19845 298515
rect 19845 298485 19875 298515
rect 19875 298485 19876 298515
rect 19844 298484 19876 298485
rect 19844 298435 19876 298436
rect 19844 298405 19845 298435
rect 19845 298405 19875 298435
rect 19875 298405 19876 298435
rect 19844 298404 19876 298405
rect 19844 298355 19876 298356
rect 19844 298325 19845 298355
rect 19845 298325 19875 298355
rect 19875 298325 19876 298355
rect 19844 298324 19876 298325
rect 19844 298275 19876 298276
rect 19844 298245 19845 298275
rect 19845 298245 19875 298275
rect 19875 298245 19876 298275
rect 19844 298244 19876 298245
rect 19844 298195 19876 298196
rect 19844 298165 19845 298195
rect 19845 298165 19875 298195
rect 19875 298165 19876 298195
rect 19844 298164 19876 298165
rect 19844 298115 19876 298116
rect 19844 298085 19845 298115
rect 19845 298085 19875 298115
rect 19875 298085 19876 298115
rect 19844 298084 19876 298085
rect 19844 298035 19876 298036
rect 19844 298005 19845 298035
rect 19845 298005 19875 298035
rect 19875 298005 19876 298035
rect 19844 298004 19876 298005
rect 19844 297955 19876 297956
rect 19844 297925 19845 297955
rect 19845 297925 19875 297955
rect 19875 297925 19876 297955
rect 19844 297924 19876 297925
rect 19844 297875 19876 297876
rect 19844 297845 19845 297875
rect 19845 297845 19875 297875
rect 19875 297845 19876 297875
rect 19844 297844 19876 297845
rect 19844 297795 19876 297796
rect 19844 297765 19845 297795
rect 19845 297765 19875 297795
rect 19875 297765 19876 297795
rect 19844 297764 19876 297765
rect 19844 297715 19876 297716
rect 19844 297685 19845 297715
rect 19845 297685 19875 297715
rect 19875 297685 19876 297715
rect 19844 297684 19876 297685
rect 19844 297635 19876 297636
rect 19844 297605 19845 297635
rect 19845 297605 19875 297635
rect 19875 297605 19876 297635
rect 19844 297604 19876 297605
rect 19844 297555 19876 297556
rect 19844 297525 19845 297555
rect 19845 297525 19875 297555
rect 19875 297525 19876 297555
rect 19844 297524 19876 297525
rect 19844 297475 19876 297476
rect 19844 297445 19845 297475
rect 19845 297445 19875 297475
rect 19875 297445 19876 297475
rect 19844 297444 19876 297445
rect 19844 297395 19876 297396
rect 19844 297365 19845 297395
rect 19845 297365 19875 297395
rect 19875 297365 19876 297395
rect 19844 297364 19876 297365
rect 19844 297315 19876 297316
rect 19844 297285 19845 297315
rect 19845 297285 19875 297315
rect 19875 297285 19876 297315
rect 19844 297284 19876 297285
rect 19844 297235 19876 297236
rect 19844 297205 19845 297235
rect 19845 297205 19875 297235
rect 19875 297205 19876 297235
rect 19844 297204 19876 297205
rect 19844 297155 19876 297156
rect 19844 297125 19845 297155
rect 19845 297125 19875 297155
rect 19875 297125 19876 297155
rect 19844 297124 19876 297125
rect 19844 297075 19876 297076
rect 19844 297045 19845 297075
rect 19845 297045 19875 297075
rect 19875 297045 19876 297075
rect 19844 297044 19876 297045
rect 19844 296995 19876 296996
rect 19844 296965 19845 296995
rect 19845 296965 19875 296995
rect 19875 296965 19876 296995
rect 19844 296964 19876 296965
rect 19844 296915 19876 296916
rect 19844 296885 19845 296915
rect 19845 296885 19875 296915
rect 19875 296885 19876 296915
rect 19844 296884 19876 296885
rect 19844 296835 19876 296836
rect 19844 296805 19845 296835
rect 19845 296805 19875 296835
rect 19875 296805 19876 296835
rect 19844 296804 19876 296805
rect 19844 296755 19876 296756
rect 19844 296725 19845 296755
rect 19845 296725 19875 296755
rect 19875 296725 19876 296755
rect 19844 296724 19876 296725
rect 19844 296675 19876 296676
rect 19844 296645 19845 296675
rect 19845 296645 19875 296675
rect 19875 296645 19876 296675
rect 19844 296644 19876 296645
rect 19844 296595 19876 296596
rect 19844 296565 19845 296595
rect 19845 296565 19875 296595
rect 19875 296565 19876 296595
rect 19844 296564 19876 296565
rect 19844 296515 19876 296516
rect 19844 296485 19845 296515
rect 19845 296485 19875 296515
rect 19875 296485 19876 296515
rect 19844 296484 19876 296485
rect 19844 296435 19876 296436
rect 19844 296405 19845 296435
rect 19845 296405 19875 296435
rect 19875 296405 19876 296435
rect 19844 296404 19876 296405
rect 19844 296355 19876 296356
rect 19844 296325 19845 296355
rect 19845 296325 19875 296355
rect 19875 296325 19876 296355
rect 19844 296324 19876 296325
rect 19844 296275 19876 296276
rect 19844 296245 19845 296275
rect 19845 296245 19875 296275
rect 19875 296245 19876 296275
rect 19844 296244 19876 296245
rect 19844 296195 19876 296196
rect 19844 296165 19845 296195
rect 19845 296165 19875 296195
rect 19875 296165 19876 296195
rect 19844 296164 19876 296165
rect 19844 296115 19876 296116
rect 19844 296085 19845 296115
rect 19845 296085 19875 296115
rect 19875 296085 19876 296115
rect 19844 296084 19876 296085
rect 19844 296035 19876 296036
rect 19844 296005 19845 296035
rect 19845 296005 19875 296035
rect 19875 296005 19876 296035
rect 19844 296004 19876 296005
rect 19844 295955 19876 295956
rect 19844 295925 19845 295955
rect 19845 295925 19875 295955
rect 19875 295925 19876 295955
rect 19844 295924 19876 295925
rect 19844 295875 19876 295876
rect 19844 295845 19845 295875
rect 19845 295845 19875 295875
rect 19875 295845 19876 295875
rect 19844 295844 19876 295845
rect 19844 295795 19876 295796
rect 19844 295765 19845 295795
rect 19845 295765 19875 295795
rect 19875 295765 19876 295795
rect 19844 295764 19876 295765
rect 19844 295715 19876 295716
rect 19844 295685 19845 295715
rect 19845 295685 19875 295715
rect 19875 295685 19876 295715
rect 19844 295684 19876 295685
rect 19844 295635 19876 295636
rect 19844 295605 19845 295635
rect 19845 295605 19875 295635
rect 19875 295605 19876 295635
rect 19844 295604 19876 295605
rect 19844 295555 19876 295556
rect 19844 295525 19845 295555
rect 19845 295525 19875 295555
rect 19875 295525 19876 295555
rect 19844 295524 19876 295525
rect 19844 295475 19876 295476
rect 19844 295445 19845 295475
rect 19845 295445 19875 295475
rect 19875 295445 19876 295475
rect 19844 295444 19876 295445
rect 19844 295395 19876 295396
rect 19844 295365 19845 295395
rect 19845 295365 19875 295395
rect 19875 295365 19876 295395
rect 19844 295364 19876 295365
rect 19844 295315 19876 295316
rect 19844 295285 19845 295315
rect 19845 295285 19875 295315
rect 19875 295285 19876 295315
rect 19844 295284 19876 295285
rect 19844 295235 19876 295236
rect 19844 295205 19845 295235
rect 19845 295205 19875 295235
rect 19875 295205 19876 295235
rect 19844 295204 19876 295205
rect 19844 295155 19876 295156
rect 19844 295125 19845 295155
rect 19845 295125 19875 295155
rect 19875 295125 19876 295155
rect 19844 295124 19876 295125
rect 19844 295075 19876 295076
rect 19844 295045 19845 295075
rect 19845 295045 19875 295075
rect 19875 295045 19876 295075
rect 19844 295044 19876 295045
rect 19844 294995 19876 294996
rect 19844 294965 19845 294995
rect 19845 294965 19875 294995
rect 19875 294965 19876 294995
rect 19844 294964 19876 294965
rect 19844 294915 19876 294916
rect 19844 294885 19845 294915
rect 19845 294885 19875 294915
rect 19875 294885 19876 294915
rect 19844 294884 19876 294885
rect 19844 294835 19876 294836
rect 19844 294805 19845 294835
rect 19845 294805 19875 294835
rect 19875 294805 19876 294835
rect 19844 294804 19876 294805
rect 19844 294755 19876 294756
rect 19844 294725 19845 294755
rect 19845 294725 19875 294755
rect 19875 294725 19876 294755
rect 19844 294724 19876 294725
rect 19844 294675 19876 294676
rect 19844 294645 19845 294675
rect 19845 294645 19875 294675
rect 19875 294645 19876 294675
rect 19844 294644 19876 294645
rect 19844 294595 19876 294596
rect 19844 294565 19845 294595
rect 19845 294565 19875 294595
rect 19875 294565 19876 294595
rect 19844 294564 19876 294565
rect 19844 294515 19876 294516
rect 19844 294485 19845 294515
rect 19845 294485 19875 294515
rect 19875 294485 19876 294515
rect 19844 294484 19876 294485
rect 19844 294435 19876 294436
rect 19844 294405 19845 294435
rect 19845 294405 19875 294435
rect 19875 294405 19876 294435
rect 19844 294404 19876 294405
rect 19844 294355 19876 294356
rect 19844 294325 19845 294355
rect 19845 294325 19875 294355
rect 19875 294325 19876 294355
rect 19844 294324 19876 294325
rect 19844 294275 19876 294276
rect 19844 294245 19845 294275
rect 19845 294245 19875 294275
rect 19875 294245 19876 294275
rect 19844 294244 19876 294245
rect 19844 294195 19876 294196
rect 19844 294165 19845 294195
rect 19845 294165 19875 294195
rect 19875 294165 19876 294195
rect 19844 294164 19876 294165
rect 19844 294115 19876 294116
rect 19844 294085 19845 294115
rect 19845 294085 19875 294115
rect 19875 294085 19876 294115
rect 19844 294084 19876 294085
rect 19844 294035 19876 294036
rect 19844 294005 19845 294035
rect 19845 294005 19875 294035
rect 19875 294005 19876 294035
rect 19844 294004 19876 294005
rect 19844 293955 19876 293956
rect 19844 293925 19845 293955
rect 19845 293925 19875 293955
rect 19875 293925 19876 293955
rect 19844 293924 19876 293925
rect 19844 293875 19876 293876
rect 19844 293845 19845 293875
rect 19845 293845 19875 293875
rect 19875 293845 19876 293875
rect 19844 293844 19876 293845
rect 19844 293795 19876 293796
rect 19844 293765 19845 293795
rect 19845 293765 19875 293795
rect 19875 293765 19876 293795
rect 19844 293764 19876 293765
rect 19844 293715 19876 293716
rect 19844 293685 19845 293715
rect 19845 293685 19875 293715
rect 19875 293685 19876 293715
rect 19844 293684 19876 293685
rect 19844 293635 19876 293636
rect 19844 293605 19845 293635
rect 19845 293605 19875 293635
rect 19875 293605 19876 293635
rect 19844 293604 19876 293605
rect 19844 293555 19876 293556
rect 19844 293525 19845 293555
rect 19845 293525 19875 293555
rect 19875 293525 19876 293555
rect 19844 293524 19876 293525
rect 19844 293475 19876 293476
rect 19844 293445 19845 293475
rect 19845 293445 19875 293475
rect 19875 293445 19876 293475
rect 19844 293444 19876 293445
rect 19844 293395 19876 293396
rect 19844 293365 19845 293395
rect 19845 293365 19875 293395
rect 19875 293365 19876 293395
rect 19844 293364 19876 293365
rect 19844 293315 19876 293316
rect 19844 293285 19845 293315
rect 19845 293285 19875 293315
rect 19875 293285 19876 293315
rect 19844 293284 19876 293285
rect 19844 293235 19876 293236
rect 19844 293205 19845 293235
rect 19845 293205 19875 293235
rect 19875 293205 19876 293235
rect 19844 293204 19876 293205
rect 19844 293155 19876 293156
rect 19844 293125 19845 293155
rect 19845 293125 19875 293155
rect 19875 293125 19876 293155
rect 19844 293124 19876 293125
rect 19844 293075 19876 293076
rect 19844 293045 19845 293075
rect 19845 293045 19875 293075
rect 19875 293045 19876 293075
rect 19844 293044 19876 293045
rect 19844 292995 19876 292996
rect 19844 292965 19845 292995
rect 19845 292965 19875 292995
rect 19875 292965 19876 292995
rect 19844 292964 19876 292965
rect 19844 292915 19876 292916
rect 19844 292885 19845 292915
rect 19845 292885 19875 292915
rect 19875 292885 19876 292915
rect 19844 292884 19876 292885
rect 19844 292835 19876 292836
rect 19844 292805 19845 292835
rect 19845 292805 19875 292835
rect 19875 292805 19876 292835
rect 19844 292804 19876 292805
rect 19844 292755 19876 292756
rect 19844 292725 19845 292755
rect 19845 292725 19875 292755
rect 19875 292725 19876 292755
rect 19844 292724 19876 292725
rect 19844 292675 19876 292676
rect 19844 292645 19845 292675
rect 19845 292645 19875 292675
rect 19875 292645 19876 292675
rect 19844 292644 19876 292645
rect 19844 292595 19876 292596
rect 19844 292565 19845 292595
rect 19845 292565 19875 292595
rect 19875 292565 19876 292595
rect 19844 292564 19876 292565
rect 19844 292515 19876 292516
rect 19844 292485 19845 292515
rect 19845 292485 19875 292515
rect 19875 292485 19876 292515
rect 19844 292484 19876 292485
rect 19844 292435 19876 292436
rect 19844 292405 19845 292435
rect 19845 292405 19875 292435
rect 19875 292405 19876 292435
rect 19844 292404 19876 292405
rect 19844 292355 19876 292356
rect 19844 292325 19845 292355
rect 19845 292325 19875 292355
rect 19875 292325 19876 292355
rect 19844 292324 19876 292325
rect 19844 292275 19876 292276
rect 19844 292245 19845 292275
rect 19845 292245 19875 292275
rect 19875 292245 19876 292275
rect 19844 292244 19876 292245
rect 19844 292195 19876 292196
rect 19844 292165 19845 292195
rect 19845 292165 19875 292195
rect 19875 292165 19876 292195
rect 19844 292164 19876 292165
rect 19844 292115 19876 292116
rect 19844 292085 19845 292115
rect 19845 292085 19875 292115
rect 19875 292085 19876 292115
rect 19844 292084 19876 292085
rect 19844 292035 19876 292036
rect 19844 292005 19845 292035
rect 19845 292005 19875 292035
rect 19875 292005 19876 292035
rect 19844 292004 19876 292005
rect 19844 291955 19876 291956
rect 19844 291925 19845 291955
rect 19845 291925 19875 291955
rect 19875 291925 19876 291955
rect 19844 291924 19876 291925
rect 19844 291875 19876 291876
rect 19844 291845 19845 291875
rect 19845 291845 19875 291875
rect 19875 291845 19876 291875
rect 19844 291844 19876 291845
rect 19844 291795 19876 291796
rect 19844 291765 19845 291795
rect 19845 291765 19875 291795
rect 19875 291765 19876 291795
rect 19844 291764 19876 291765
rect 19844 291715 19876 291716
rect 19844 291685 19845 291715
rect 19845 291685 19875 291715
rect 19875 291685 19876 291715
rect 19844 291684 19876 291685
rect 19844 291635 19876 291636
rect 19844 291605 19845 291635
rect 19845 291605 19875 291635
rect 19875 291605 19876 291635
rect 19844 291604 19876 291605
rect 19844 291555 19876 291556
rect 19844 291525 19845 291555
rect 19845 291525 19875 291555
rect 19875 291525 19876 291555
rect 19844 291524 19876 291525
rect 19844 291475 19876 291476
rect 19844 291445 19845 291475
rect 19845 291445 19875 291475
rect 19875 291445 19876 291475
rect 19844 291444 19876 291445
rect 19844 291395 19876 291396
rect 19844 291365 19845 291395
rect 19845 291365 19875 291395
rect 19875 291365 19876 291395
rect 19844 291364 19876 291365
rect 19844 291315 19876 291316
rect 19844 291285 19845 291315
rect 19845 291285 19875 291315
rect 19875 291285 19876 291315
rect 19844 291284 19876 291285
rect 19844 291235 19876 291236
rect 19844 291205 19845 291235
rect 19845 291205 19875 291235
rect 19875 291205 19876 291235
rect 19844 291204 19876 291205
rect 19844 291155 19876 291156
rect 19844 291125 19845 291155
rect 19845 291125 19875 291155
rect 19875 291125 19876 291155
rect 19844 291124 19876 291125
rect 19844 291075 19876 291076
rect 19844 291045 19845 291075
rect 19845 291045 19875 291075
rect 19875 291045 19876 291075
rect 19844 291044 19876 291045
rect 19844 290995 19876 290996
rect 19844 290965 19845 290995
rect 19845 290965 19875 290995
rect 19875 290965 19876 290995
rect 19844 290964 19876 290965
rect 19844 290915 19876 290916
rect 19844 290885 19845 290915
rect 19845 290885 19875 290915
rect 19875 290885 19876 290915
rect 19844 290884 19876 290885
rect 19844 290835 19876 290836
rect 19844 290805 19845 290835
rect 19845 290805 19875 290835
rect 19875 290805 19876 290835
rect 19844 290804 19876 290805
rect 19844 290755 19876 290756
rect 19844 290725 19845 290755
rect 19845 290725 19875 290755
rect 19875 290725 19876 290755
rect 19844 290724 19876 290725
rect 19844 290675 19876 290676
rect 19844 290645 19845 290675
rect 19845 290645 19875 290675
rect 19875 290645 19876 290675
rect 19844 290644 19876 290645
rect 19844 290595 19876 290596
rect 19844 290565 19845 290595
rect 19845 290565 19875 290595
rect 19875 290565 19876 290595
rect 19844 290564 19876 290565
rect 19844 290515 19876 290516
rect 19844 290485 19845 290515
rect 19845 290485 19875 290515
rect 19875 290485 19876 290515
rect 19844 290484 19876 290485
rect 19844 290435 19876 290436
rect 19844 290405 19845 290435
rect 19845 290405 19875 290435
rect 19875 290405 19876 290435
rect 19844 290404 19876 290405
rect 19844 290355 19876 290356
rect 19844 290325 19845 290355
rect 19845 290325 19875 290355
rect 19875 290325 19876 290355
rect 19844 290324 19876 290325
rect 19844 290275 19876 290276
rect 19844 290245 19845 290275
rect 19845 290245 19875 290275
rect 19875 290245 19876 290275
rect 19844 290244 19876 290245
rect 19844 290195 19876 290196
rect 19844 290165 19845 290195
rect 19845 290165 19875 290195
rect 19875 290165 19876 290195
rect 19844 290164 19876 290165
rect 19844 290115 19876 290116
rect 19844 290085 19845 290115
rect 19845 290085 19875 290115
rect 19875 290085 19876 290115
rect 19844 290084 19876 290085
rect 19844 290035 19876 290036
rect 19844 290005 19845 290035
rect 19845 290005 19875 290035
rect 19875 290005 19876 290035
rect 19844 290004 19876 290005
rect 19844 289955 19876 289956
rect 19844 289925 19845 289955
rect 19845 289925 19875 289955
rect 19875 289925 19876 289955
rect 19844 289924 19876 289925
rect 19844 289875 19876 289876
rect 19844 289845 19845 289875
rect 19845 289845 19875 289875
rect 19875 289845 19876 289875
rect 19844 289844 19876 289845
rect 19844 289795 19876 289796
rect 19844 289765 19845 289795
rect 19845 289765 19875 289795
rect 19875 289765 19876 289795
rect 19844 289764 19876 289765
rect 19844 289715 19876 289716
rect 19844 289685 19845 289715
rect 19845 289685 19875 289715
rect 19875 289685 19876 289715
rect 19844 289684 19876 289685
rect 19844 289635 19876 289636
rect 19844 289605 19845 289635
rect 19845 289605 19875 289635
rect 19875 289605 19876 289635
rect 19844 289604 19876 289605
rect 19844 289555 19876 289556
rect 19844 289525 19845 289555
rect 19845 289525 19875 289555
rect 19875 289525 19876 289555
rect 19844 289524 19876 289525
rect 19844 289475 19876 289476
rect 19844 289445 19845 289475
rect 19845 289445 19875 289475
rect 19875 289445 19876 289475
rect 19844 289444 19876 289445
rect 19844 289395 19876 289396
rect 19844 289365 19845 289395
rect 19845 289365 19875 289395
rect 19875 289365 19876 289395
rect 19844 289364 19876 289365
rect 19844 289315 19876 289316
rect 19844 289285 19845 289315
rect 19845 289285 19875 289315
rect 19875 289285 19876 289315
rect 19844 289284 19876 289285
rect 19844 289235 19876 289236
rect 19844 289205 19845 289235
rect 19845 289205 19875 289235
rect 19875 289205 19876 289235
rect 19844 289204 19876 289205
rect 19844 289155 19876 289156
rect 19844 289125 19845 289155
rect 19845 289125 19875 289155
rect 19875 289125 19876 289155
rect 19844 289124 19876 289125
rect 19844 289075 19876 289076
rect 19844 289045 19845 289075
rect 19845 289045 19875 289075
rect 19875 289045 19876 289075
rect 19844 289044 19876 289045
rect 19844 288995 19876 288996
rect 19844 288965 19845 288995
rect 19845 288965 19875 288995
rect 19875 288965 19876 288995
rect 19844 288964 19876 288965
rect 19844 288915 19876 288916
rect 19844 288885 19845 288915
rect 19845 288885 19875 288915
rect 19875 288885 19876 288915
rect 19844 288884 19876 288885
rect 19844 288835 19876 288836
rect 19844 288805 19845 288835
rect 19845 288805 19875 288835
rect 19875 288805 19876 288835
rect 19844 288804 19876 288805
rect 19844 288755 19876 288756
rect 19844 288725 19845 288755
rect 19845 288725 19875 288755
rect 19875 288725 19876 288755
rect 19844 288724 19876 288725
rect 19844 288675 19876 288676
rect 19844 288645 19845 288675
rect 19845 288645 19875 288675
rect 19875 288645 19876 288675
rect 19844 288644 19876 288645
rect 19844 288595 19876 288596
rect 19844 288565 19845 288595
rect 19845 288565 19875 288595
rect 19875 288565 19876 288595
rect 19844 288564 19876 288565
rect 19844 288515 19876 288516
rect 19844 288485 19845 288515
rect 19845 288485 19875 288515
rect 19875 288485 19876 288515
rect 19844 288484 19876 288485
rect 19844 288435 19876 288436
rect 19844 288405 19845 288435
rect 19845 288405 19875 288435
rect 19875 288405 19876 288435
rect 19844 288404 19876 288405
rect 19844 288355 19876 288356
rect 19844 288325 19845 288355
rect 19845 288325 19875 288355
rect 19875 288325 19876 288355
rect 19844 288324 19876 288325
rect 19844 288275 19876 288276
rect 19844 288245 19845 288275
rect 19845 288245 19875 288275
rect 19875 288245 19876 288275
rect 19844 288244 19876 288245
rect 19844 288195 19876 288196
rect 19844 288165 19845 288195
rect 19845 288165 19875 288195
rect 19875 288165 19876 288195
rect 19844 288164 19876 288165
rect 19844 288115 19876 288116
rect 19844 288085 19845 288115
rect 19845 288085 19875 288115
rect 19875 288085 19876 288115
rect 19844 288084 19876 288085
rect 19844 288035 19876 288036
rect 19844 288005 19845 288035
rect 19845 288005 19875 288035
rect 19875 288005 19876 288035
rect 19844 288004 19876 288005
rect 19844 287955 19876 287956
rect 19844 287925 19845 287955
rect 19845 287925 19875 287955
rect 19875 287925 19876 287955
rect 19844 287924 19876 287925
rect 19844 287875 19876 287876
rect 19844 287845 19845 287875
rect 19845 287845 19875 287875
rect 19875 287845 19876 287875
rect 19844 287844 19876 287845
rect 19844 287795 19876 287796
rect 19844 287765 19845 287795
rect 19845 287765 19875 287795
rect 19875 287765 19876 287795
rect 19844 287764 19876 287765
rect 19844 287715 19876 287716
rect 19844 287685 19845 287715
rect 19845 287685 19875 287715
rect 19875 287685 19876 287715
rect 19844 287684 19876 287685
rect 19844 287635 19876 287636
rect 19844 287605 19845 287635
rect 19845 287605 19875 287635
rect 19875 287605 19876 287635
rect 19844 287604 19876 287605
rect 19844 287555 19876 287556
rect 19844 287525 19845 287555
rect 19845 287525 19875 287555
rect 19875 287525 19876 287555
rect 19844 287524 19876 287525
rect 19844 287475 19876 287476
rect 19844 287445 19845 287475
rect 19845 287445 19875 287475
rect 19875 287445 19876 287475
rect 19844 287444 19876 287445
rect 19844 287395 19876 287396
rect 19844 287365 19845 287395
rect 19845 287365 19875 287395
rect 19875 287365 19876 287395
rect 19844 287364 19876 287365
rect 19844 287315 19876 287316
rect 19844 287285 19845 287315
rect 19845 287285 19875 287315
rect 19875 287285 19876 287315
rect 19844 287284 19876 287285
rect 19844 287235 19876 287236
rect 19844 287205 19845 287235
rect 19845 287205 19875 287235
rect 19875 287205 19876 287235
rect 19844 287204 19876 287205
rect 19844 287155 19876 287156
rect 19844 287125 19845 287155
rect 19845 287125 19875 287155
rect 19875 287125 19876 287155
rect 19844 287124 19876 287125
rect 19844 287075 19876 287076
rect 19844 287045 19845 287075
rect 19845 287045 19875 287075
rect 19875 287045 19876 287075
rect 19844 287044 19876 287045
rect 19844 286995 19876 286996
rect 19844 286965 19845 286995
rect 19845 286965 19875 286995
rect 19875 286965 19876 286995
rect 19844 286964 19876 286965
rect 19844 286915 19876 286916
rect 19844 286885 19845 286915
rect 19845 286885 19875 286915
rect 19875 286885 19876 286915
rect 19844 286884 19876 286885
rect 19844 286835 19876 286836
rect 19844 286805 19845 286835
rect 19845 286805 19875 286835
rect 19875 286805 19876 286835
rect 19844 286804 19876 286805
rect 19844 286755 19876 286756
rect 19844 286725 19845 286755
rect 19845 286725 19875 286755
rect 19875 286725 19876 286755
rect 19844 286724 19876 286725
rect 19844 286675 19876 286676
rect 19844 286645 19845 286675
rect 19845 286645 19875 286675
rect 19875 286645 19876 286675
rect 19844 286644 19876 286645
rect 19844 286595 19876 286596
rect 19844 286565 19845 286595
rect 19845 286565 19875 286595
rect 19875 286565 19876 286595
rect 19844 286564 19876 286565
rect 19844 286515 19876 286516
rect 19844 286485 19845 286515
rect 19845 286485 19875 286515
rect 19875 286485 19876 286515
rect 19844 286484 19876 286485
rect 19844 286435 19876 286436
rect 19844 286405 19845 286435
rect 19845 286405 19875 286435
rect 19875 286405 19876 286435
rect 19844 286404 19876 286405
rect 19844 286355 19876 286356
rect 19844 286325 19845 286355
rect 19845 286325 19875 286355
rect 19875 286325 19876 286355
rect 19844 286324 19876 286325
rect 19844 286275 19876 286276
rect 19844 286245 19845 286275
rect 19845 286245 19875 286275
rect 19875 286245 19876 286275
rect 19844 286244 19876 286245
rect 19844 286195 19876 286196
rect 19844 286165 19845 286195
rect 19845 286165 19875 286195
rect 19875 286165 19876 286195
rect 19844 286164 19876 286165
rect 19844 286115 19876 286116
rect 19844 286085 19845 286115
rect 19845 286085 19875 286115
rect 19875 286085 19876 286115
rect 19844 286084 19876 286085
rect 19844 286035 19876 286036
rect 19844 286005 19845 286035
rect 19845 286005 19875 286035
rect 19875 286005 19876 286035
rect 19844 286004 19876 286005
rect 19844 285955 19876 285956
rect 19844 285925 19845 285955
rect 19845 285925 19875 285955
rect 19875 285925 19876 285955
rect 19844 285924 19876 285925
rect 19844 285875 19876 285876
rect 19844 285845 19845 285875
rect 19845 285845 19875 285875
rect 19875 285845 19876 285875
rect 19844 285844 19876 285845
rect 19844 285795 19876 285796
rect 19844 285765 19845 285795
rect 19845 285765 19875 285795
rect 19875 285765 19876 285795
rect 19844 285764 19876 285765
rect 19844 285715 19876 285716
rect 19844 285685 19845 285715
rect 19845 285685 19875 285715
rect 19875 285685 19876 285715
rect 19844 285684 19876 285685
rect 19844 285635 19876 285636
rect 19844 285605 19845 285635
rect 19845 285605 19875 285635
rect 19875 285605 19876 285635
rect 19844 285604 19876 285605
rect 19844 285555 19876 285556
rect 19844 285525 19845 285555
rect 19845 285525 19875 285555
rect 19875 285525 19876 285555
rect 19844 285524 19876 285525
rect 19844 285475 19876 285476
rect 19844 285445 19845 285475
rect 19845 285445 19875 285475
rect 19875 285445 19876 285475
rect 19844 285444 19876 285445
rect 19844 285395 19876 285396
rect 19844 285365 19845 285395
rect 19845 285365 19875 285395
rect 19875 285365 19876 285395
rect 19844 285364 19876 285365
rect 19844 285315 19876 285316
rect 19844 285285 19845 285315
rect 19845 285285 19875 285315
rect 19875 285285 19876 285315
rect 19844 285284 19876 285285
rect 19844 285235 19876 285236
rect 19844 285205 19845 285235
rect 19845 285205 19875 285235
rect 19875 285205 19876 285235
rect 19844 285204 19876 285205
rect 19844 285155 19876 285156
rect 19844 285125 19845 285155
rect 19845 285125 19875 285155
rect 19875 285125 19876 285155
rect 19844 285124 19876 285125
rect 19844 285075 19876 285076
rect 19844 285045 19845 285075
rect 19845 285045 19875 285075
rect 19875 285045 19876 285075
rect 19844 285044 19876 285045
rect 19844 284995 19876 284996
rect 19844 284965 19845 284995
rect 19845 284965 19875 284995
rect 19875 284965 19876 284995
rect 19844 284964 19876 284965
rect 19844 284915 19876 284916
rect 19844 284885 19845 284915
rect 19845 284885 19875 284915
rect 19875 284885 19876 284915
rect 19844 284884 19876 284885
rect 19844 284835 19876 284836
rect 19844 284805 19845 284835
rect 19845 284805 19875 284835
rect 19875 284805 19876 284835
rect 19844 284804 19876 284805
rect 19844 284755 19876 284756
rect 19844 284725 19845 284755
rect 19845 284725 19875 284755
rect 19875 284725 19876 284755
rect 19844 284724 19876 284725
rect 19844 284675 19876 284676
rect 19844 284645 19845 284675
rect 19845 284645 19875 284675
rect 19875 284645 19876 284675
rect 19844 284644 19876 284645
rect 19844 284595 19876 284596
rect 19844 284565 19845 284595
rect 19845 284565 19875 284595
rect 19875 284565 19876 284595
rect 19844 284564 19876 284565
rect 19844 284515 19876 284516
rect 19844 284485 19845 284515
rect 19845 284485 19875 284515
rect 19875 284485 19876 284515
rect 19844 284484 19876 284485
rect 19844 284435 19876 284436
rect 19844 284405 19845 284435
rect 19845 284405 19875 284435
rect 19875 284405 19876 284435
rect 19844 284404 19876 284405
rect 19844 284355 19876 284356
rect 19844 284325 19845 284355
rect 19845 284325 19875 284355
rect 19875 284325 19876 284355
rect 19844 284324 19876 284325
rect 19844 284275 19876 284276
rect 19844 284245 19845 284275
rect 19845 284245 19875 284275
rect 19875 284245 19876 284275
rect 19844 284244 19876 284245
rect 19844 284195 19876 284196
rect 19844 284165 19845 284195
rect 19845 284165 19875 284195
rect 19875 284165 19876 284195
rect 19844 284164 19876 284165
rect 19844 284115 19876 284116
rect 19844 284085 19845 284115
rect 19845 284085 19875 284115
rect 19875 284085 19876 284115
rect 19844 284084 19876 284085
rect 19844 284035 19876 284036
rect 19844 284005 19845 284035
rect 19845 284005 19875 284035
rect 19875 284005 19876 284035
rect 19844 284004 19876 284005
rect 19844 283955 19876 283956
rect 19844 283925 19845 283955
rect 19845 283925 19875 283955
rect 19875 283925 19876 283955
rect 19844 283924 19876 283925
rect 19844 283875 19876 283876
rect 19844 283845 19845 283875
rect 19845 283845 19875 283875
rect 19875 283845 19876 283875
rect 19844 283844 19876 283845
rect 19844 283795 19876 283796
rect 19844 283765 19845 283795
rect 19845 283765 19875 283795
rect 19875 283765 19876 283795
rect 19844 283764 19876 283765
rect 19844 283715 19876 283716
rect 19844 283685 19845 283715
rect 19845 283685 19875 283715
rect 19875 283685 19876 283715
rect 19844 283684 19876 283685
rect 19844 283635 19876 283636
rect 19844 283605 19845 283635
rect 19845 283605 19875 283635
rect 19875 283605 19876 283635
rect 19844 283604 19876 283605
rect 19844 283555 19876 283556
rect 19844 283525 19845 283555
rect 19845 283525 19875 283555
rect 19875 283525 19876 283555
rect 19844 283524 19876 283525
rect 19844 283475 19876 283476
rect 19844 283445 19845 283475
rect 19845 283445 19875 283475
rect 19875 283445 19876 283475
rect 19844 283444 19876 283445
rect 19844 283395 19876 283396
rect 19844 283365 19845 283395
rect 19845 283365 19875 283395
rect 19875 283365 19876 283395
rect 19844 283364 19876 283365
rect 19844 283315 19876 283316
rect 19844 283285 19845 283315
rect 19845 283285 19875 283315
rect 19875 283285 19876 283315
rect 19844 283284 19876 283285
rect 19844 283235 19876 283236
rect 19844 283205 19845 283235
rect 19845 283205 19875 283235
rect 19875 283205 19876 283235
rect 19844 283204 19876 283205
rect 19844 283155 19876 283156
rect 19844 283125 19845 283155
rect 19845 283125 19875 283155
rect 19875 283125 19876 283155
rect 19844 283124 19876 283125
rect 19844 283075 19876 283076
rect 19844 283045 19845 283075
rect 19845 283045 19875 283075
rect 19875 283045 19876 283075
rect 19844 283044 19876 283045
rect 19844 282995 19876 282996
rect 19844 282965 19845 282995
rect 19845 282965 19875 282995
rect 19875 282965 19876 282995
rect 19844 282964 19876 282965
rect 19844 282915 19876 282916
rect 19844 282885 19845 282915
rect 19845 282885 19875 282915
rect 19875 282885 19876 282915
rect 19844 282884 19876 282885
rect 19844 282835 19876 282836
rect 19844 282805 19845 282835
rect 19845 282805 19875 282835
rect 19875 282805 19876 282835
rect 19844 282804 19876 282805
rect 19844 282755 19876 282756
rect 19844 282725 19845 282755
rect 19845 282725 19875 282755
rect 19875 282725 19876 282755
rect 19844 282724 19876 282725
rect 19844 282675 19876 282676
rect 19844 282645 19845 282675
rect 19845 282645 19875 282675
rect 19875 282645 19876 282675
rect 19844 282644 19876 282645
rect 19844 282595 19876 282596
rect 19844 282565 19845 282595
rect 19845 282565 19875 282595
rect 19875 282565 19876 282595
rect 19844 282564 19876 282565
rect 19844 282515 19876 282516
rect 19844 282485 19845 282515
rect 19845 282485 19875 282515
rect 19875 282485 19876 282515
rect 19844 282484 19876 282485
rect 19844 282435 19876 282436
rect 19844 282405 19845 282435
rect 19845 282405 19875 282435
rect 19875 282405 19876 282435
rect 19844 282404 19876 282405
rect 19844 282355 19876 282356
rect 19844 282325 19845 282355
rect 19845 282325 19875 282355
rect 19875 282325 19876 282355
rect 19844 282324 19876 282325
rect 19844 282275 19876 282276
rect 19844 282245 19845 282275
rect 19845 282245 19875 282275
rect 19875 282245 19876 282275
rect 19844 282244 19876 282245
rect 19844 282195 19876 282196
rect 19844 282165 19845 282195
rect 19845 282165 19875 282195
rect 19875 282165 19876 282195
rect 19844 282164 19876 282165
rect 19844 282115 19876 282116
rect 19844 282085 19845 282115
rect 19845 282085 19875 282115
rect 19875 282085 19876 282115
rect 19844 282084 19876 282085
rect 19844 282035 19876 282036
rect 19844 282005 19845 282035
rect 19845 282005 19875 282035
rect 19875 282005 19876 282035
rect 19844 282004 19876 282005
rect 19844 281955 19876 281956
rect 19844 281925 19845 281955
rect 19845 281925 19875 281955
rect 19875 281925 19876 281955
rect 19844 281924 19876 281925
rect 19844 281875 19876 281876
rect 19844 281845 19845 281875
rect 19845 281845 19875 281875
rect 19875 281845 19876 281875
rect 19844 281844 19876 281845
rect 19844 281795 19876 281796
rect 19844 281765 19845 281795
rect 19845 281765 19875 281795
rect 19875 281765 19876 281795
rect 19844 281764 19876 281765
rect 19844 281715 19876 281716
rect 19844 281685 19845 281715
rect 19845 281685 19875 281715
rect 19875 281685 19876 281715
rect 19844 281684 19876 281685
rect 19844 281635 19876 281636
rect 19844 281605 19845 281635
rect 19845 281605 19875 281635
rect 19875 281605 19876 281635
rect 19844 281604 19876 281605
rect 19844 281555 19876 281556
rect 19844 281525 19845 281555
rect 19845 281525 19875 281555
rect 19875 281525 19876 281555
rect 19844 281524 19876 281525
rect 19844 281475 19876 281476
rect 19844 281445 19845 281475
rect 19845 281445 19875 281475
rect 19875 281445 19876 281475
rect 19844 281444 19876 281445
rect 19844 281395 19876 281396
rect 19844 281365 19845 281395
rect 19845 281365 19875 281395
rect 19875 281365 19876 281395
rect 19844 281364 19876 281365
rect 19844 281315 19876 281316
rect 19844 281285 19845 281315
rect 19845 281285 19875 281315
rect 19875 281285 19876 281315
rect 19844 281284 19876 281285
rect 19844 281235 19876 281236
rect 19844 281205 19845 281235
rect 19845 281205 19875 281235
rect 19875 281205 19876 281235
rect 19844 281204 19876 281205
rect 19844 281155 19876 281156
rect 19844 281125 19845 281155
rect 19845 281125 19875 281155
rect 19875 281125 19876 281155
rect 19844 281124 19876 281125
rect 19844 281075 19876 281076
rect 19844 281045 19845 281075
rect 19845 281045 19875 281075
rect 19875 281045 19876 281075
rect 19844 281044 19876 281045
rect 19844 280995 19876 280996
rect 19844 280965 19845 280995
rect 19845 280965 19875 280995
rect 19875 280965 19876 280995
rect 19844 280964 19876 280965
rect 19844 280915 19876 280916
rect 19844 280885 19845 280915
rect 19845 280885 19875 280915
rect 19875 280885 19876 280915
rect 19844 280884 19876 280885
rect 19844 280835 19876 280836
rect 19844 280805 19845 280835
rect 19845 280805 19875 280835
rect 19875 280805 19876 280835
rect 19844 280804 19876 280805
rect 19844 280755 19876 280756
rect 19844 280725 19845 280755
rect 19845 280725 19875 280755
rect 19875 280725 19876 280755
rect 19844 280724 19876 280725
rect 19844 280675 19876 280676
rect 19844 280645 19845 280675
rect 19845 280645 19875 280675
rect 19875 280645 19876 280675
rect 19844 280644 19876 280645
rect 19844 280595 19876 280596
rect 19844 280565 19845 280595
rect 19845 280565 19875 280595
rect 19875 280565 19876 280595
rect 19844 280564 19876 280565
rect 19844 280515 19876 280516
rect 19844 280485 19845 280515
rect 19845 280485 19875 280515
rect 19875 280485 19876 280515
rect 19844 280484 19876 280485
rect 19844 280435 19876 280436
rect 19844 280405 19845 280435
rect 19845 280405 19875 280435
rect 19875 280405 19876 280435
rect 19844 280404 19876 280405
rect 19844 280355 19876 280356
rect 19844 280325 19845 280355
rect 19845 280325 19875 280355
rect 19875 280325 19876 280355
rect 19844 280324 19876 280325
rect 19844 280275 19876 280276
rect 19844 280245 19845 280275
rect 19845 280245 19875 280275
rect 19875 280245 19876 280275
rect 19844 280244 19876 280245
rect 19844 280195 19876 280196
rect 19844 280165 19845 280195
rect 19845 280165 19875 280195
rect 19875 280165 19876 280195
rect 19844 280164 19876 280165
rect 19844 280115 19876 280116
rect 19844 280085 19845 280115
rect 19845 280085 19875 280115
rect 19875 280085 19876 280115
rect 19844 280084 19876 280085
rect 19844 280035 19876 280036
rect 19844 280005 19845 280035
rect 19845 280005 19875 280035
rect 19875 280005 19876 280035
rect 19844 280004 19876 280005
rect 19844 279955 19876 279956
rect 19844 279925 19845 279955
rect 19845 279925 19875 279955
rect 19875 279925 19876 279955
rect 19844 279924 19876 279925
rect 19844 279875 19876 279876
rect 19844 279845 19845 279875
rect 19845 279845 19875 279875
rect 19875 279845 19876 279875
rect 19844 279844 19876 279845
rect 19844 279795 19876 279796
rect 19844 279765 19845 279795
rect 19845 279765 19875 279795
rect 19875 279765 19876 279795
rect 19844 279764 19876 279765
rect 19844 279715 19876 279716
rect 19844 279685 19845 279715
rect 19845 279685 19875 279715
rect 19875 279685 19876 279715
rect 19844 279684 19876 279685
rect 19844 279635 19876 279636
rect 19844 279605 19845 279635
rect 19845 279605 19875 279635
rect 19875 279605 19876 279635
rect 19844 279604 19876 279605
rect 19844 279555 19876 279556
rect 19844 279525 19845 279555
rect 19845 279525 19875 279555
rect 19875 279525 19876 279555
rect 19844 279524 19876 279525
rect 19844 279475 19876 279476
rect 19844 279445 19845 279475
rect 19845 279445 19875 279475
rect 19875 279445 19876 279475
rect 19844 279444 19876 279445
rect 19844 279395 19876 279396
rect 19844 279365 19845 279395
rect 19845 279365 19875 279395
rect 19875 279365 19876 279395
rect 19844 279364 19876 279365
rect 19844 279315 19876 279316
rect 19844 279285 19845 279315
rect 19845 279285 19875 279315
rect 19875 279285 19876 279315
rect 19844 279284 19876 279285
rect 19844 279235 19876 279236
rect 19844 279205 19845 279235
rect 19845 279205 19875 279235
rect 19875 279205 19876 279235
rect 19844 279204 19876 279205
rect 19844 279155 19876 279156
rect 19844 279125 19845 279155
rect 19845 279125 19875 279155
rect 19875 279125 19876 279155
rect 19844 279124 19876 279125
rect 19844 279075 19876 279076
rect 19844 279045 19845 279075
rect 19845 279045 19875 279075
rect 19875 279045 19876 279075
rect 19844 279044 19876 279045
rect 19844 278995 19876 278996
rect 19844 278965 19845 278995
rect 19845 278965 19875 278995
rect 19875 278965 19876 278995
rect 19844 278964 19876 278965
rect 19844 278915 19876 278916
rect 19844 278885 19845 278915
rect 19845 278885 19875 278915
rect 19875 278885 19876 278915
rect 19844 278884 19876 278885
rect 19844 278835 19876 278836
rect 19844 278805 19845 278835
rect 19845 278805 19875 278835
rect 19875 278805 19876 278835
rect 19844 278804 19876 278805
rect 19844 278755 19876 278756
rect 19844 278725 19845 278755
rect 19845 278725 19875 278755
rect 19875 278725 19876 278755
rect 19844 278724 19876 278725
rect 19844 278675 19876 278676
rect 19844 278645 19845 278675
rect 19845 278645 19875 278675
rect 19875 278645 19876 278675
rect 19844 278644 19876 278645
rect 19684 278515 19716 278516
rect 19684 278485 19685 278515
rect 19685 278485 19715 278515
rect 19715 278485 19716 278515
rect 19684 278484 19716 278485
rect 19844 278515 19876 278516
rect 19844 278485 19845 278515
rect 19845 278485 19875 278515
rect 19875 278485 19876 278515
rect 19844 278484 19876 278485
rect 17204 278435 17236 278436
rect 17204 278405 17205 278435
rect 17205 278405 17235 278435
rect 17235 278405 17236 278435
rect 17204 278404 17236 278405
rect 17204 278355 17236 278356
rect 17204 278325 17205 278355
rect 17205 278325 17235 278355
rect 17235 278325 17236 278355
rect 17204 278324 17236 278325
rect 17204 278275 17236 278276
rect 17204 278245 17205 278275
rect 17205 278245 17235 278275
rect 17235 278245 17236 278275
rect 17204 278244 17236 278245
rect 17204 278195 17236 278196
rect 17204 278165 17205 278195
rect 17205 278165 17235 278195
rect 17235 278165 17236 278195
rect 17204 278164 17236 278165
rect 17204 278115 17236 278116
rect 17204 278085 17205 278115
rect 17205 278085 17235 278115
rect 17235 278085 17236 278115
rect 17204 278084 17236 278085
rect 17204 278035 17236 278036
rect 17204 278005 17205 278035
rect 17205 278005 17235 278035
rect 17235 278005 17236 278035
rect 17204 278004 17236 278005
rect 17204 277955 17236 277956
rect 17204 277925 17205 277955
rect 17205 277925 17235 277955
rect 17235 277925 17236 277955
rect 17204 277924 17236 277925
rect 17204 277875 17236 277876
rect 17204 277845 17205 277875
rect 17205 277845 17235 277875
rect 17235 277845 17236 277875
rect 17204 277844 17236 277845
rect 28404 275355 28436 275356
rect 28404 275325 28405 275355
rect 28405 275325 28435 275355
rect 28435 275325 28436 275355
rect 28404 275324 28436 275325
rect 28404 275275 28436 275276
rect 28404 275245 28405 275275
rect 28405 275245 28435 275275
rect 28435 275245 28436 275275
rect 28404 275244 28436 275245
rect 28564 275355 28596 275356
rect 28564 275325 28565 275355
rect 28565 275325 28595 275355
rect 28595 275325 28596 275355
rect 28564 275324 28596 275325
rect 28564 275275 28596 275276
rect 28564 275245 28565 275275
rect 28565 275245 28595 275275
rect 28595 275245 28596 275275
rect 28564 275244 28596 275245
rect 28724 275355 28756 275356
rect 28724 275325 28725 275355
rect 28725 275325 28755 275355
rect 28755 275325 28756 275355
rect 28724 275324 28756 275325
rect 28724 275275 28756 275276
rect 28724 275245 28725 275275
rect 28725 275245 28755 275275
rect 28755 275245 28756 275275
rect 28724 275244 28756 275245
<< metal4 >>
rect 10720 351396 19880 351400
rect 10720 351364 10724 351396
rect 10756 351364 10804 351396
rect 10836 351364 10884 351396
rect 10916 351364 10964 351396
rect 10996 351364 11044 351396
rect 11076 351364 11124 351396
rect 11156 351364 11204 351396
rect 11236 351364 11284 351396
rect 11316 351364 11364 351396
rect 11396 351364 11444 351396
rect 11476 351364 11524 351396
rect 11556 351364 11604 351396
rect 11636 351364 11684 351396
rect 11716 351364 11764 351396
rect 11796 351364 11844 351396
rect 11876 351364 11924 351396
rect 11956 351364 12004 351396
rect 12036 351364 12084 351396
rect 12116 351364 12164 351396
rect 12196 351364 12244 351396
rect 12276 351364 12324 351396
rect 12356 351364 12404 351396
rect 12436 351364 12484 351396
rect 12516 351364 12564 351396
rect 12596 351364 12644 351396
rect 12676 351364 12724 351396
rect 12756 351364 12804 351396
rect 12836 351364 12884 351396
rect 12916 351364 12964 351396
rect 12996 351364 13044 351396
rect 13076 351364 13124 351396
rect 13156 351364 13204 351396
rect 13236 351364 13284 351396
rect 13316 351364 13364 351396
rect 13396 351364 13444 351396
rect 13476 351364 13524 351396
rect 13556 351364 13604 351396
rect 13636 351364 13684 351396
rect 13716 351364 13764 351396
rect 13796 351364 13844 351396
rect 13876 351364 13924 351396
rect 13956 351364 14004 351396
rect 14036 351364 14084 351396
rect 14116 351364 14164 351396
rect 14196 351364 14244 351396
rect 14276 351364 14324 351396
rect 14356 351364 14404 351396
rect 14436 351364 14484 351396
rect 14516 351364 14564 351396
rect 14596 351364 14644 351396
rect 14676 351364 14724 351396
rect 14756 351364 14804 351396
rect 14836 351364 14884 351396
rect 14916 351364 14964 351396
rect 14996 351364 15044 351396
rect 15076 351364 15124 351396
rect 15156 351364 15204 351396
rect 15236 351364 15284 351396
rect 15316 351364 15364 351396
rect 15396 351364 15444 351396
rect 15476 351364 15524 351396
rect 15556 351364 15604 351396
rect 15636 351364 15684 351396
rect 15716 351364 15764 351396
rect 15796 351364 15844 351396
rect 15876 351364 15924 351396
rect 15956 351364 16004 351396
rect 16036 351364 16084 351396
rect 16116 351364 16164 351396
rect 16196 351364 16244 351396
rect 16276 351364 16324 351396
rect 16356 351364 16404 351396
rect 16436 351364 16484 351396
rect 16516 351364 16564 351396
rect 16596 351364 16644 351396
rect 16676 351364 16724 351396
rect 16756 351364 16804 351396
rect 16836 351364 16884 351396
rect 16916 351364 16964 351396
rect 16996 351364 17044 351396
rect 17076 351364 17124 351396
rect 17156 351364 17204 351396
rect 17236 351364 17284 351396
rect 17316 351364 17364 351396
rect 17396 351364 17444 351396
rect 17476 351364 17524 351396
rect 17556 351364 17604 351396
rect 17636 351364 17684 351396
rect 17716 351364 17764 351396
rect 17796 351364 17844 351396
rect 17876 351364 17924 351396
rect 17956 351364 18004 351396
rect 18036 351364 18084 351396
rect 18116 351364 18164 351396
rect 18196 351364 18244 351396
rect 18276 351364 18324 351396
rect 18356 351364 18404 351396
rect 18436 351364 18484 351396
rect 18516 351364 18564 351396
rect 18596 351364 18644 351396
rect 18676 351364 18724 351396
rect 18756 351364 18804 351396
rect 18836 351364 18884 351396
rect 18916 351364 18964 351396
rect 18996 351364 19044 351396
rect 19076 351364 19124 351396
rect 19156 351364 19204 351396
rect 19236 351364 19284 351396
rect 19316 351364 19364 351396
rect 19396 351364 19444 351396
rect 19476 351364 19524 351396
rect 19556 351364 19604 351396
rect 19636 351364 19684 351396
rect 19716 351364 19844 351396
rect 19876 351364 19880 351396
rect 10720 351360 19880 351364
rect 10640 351316 19800 351320
rect 10640 351284 10724 351316
rect 10756 351284 10804 351316
rect 10836 351284 10884 351316
rect 10916 351284 10964 351316
rect 10996 351284 11044 351316
rect 11076 351284 11124 351316
rect 11156 351284 11204 351316
rect 11236 351284 11284 351316
rect 11316 351284 11364 351316
rect 11396 351284 11444 351316
rect 11476 351284 11524 351316
rect 11556 351284 11604 351316
rect 11636 351284 11684 351316
rect 11716 351284 11764 351316
rect 11796 351284 11844 351316
rect 11876 351284 11924 351316
rect 11956 351284 12004 351316
rect 12036 351284 12084 351316
rect 12116 351284 12164 351316
rect 12196 351284 12244 351316
rect 12276 351284 12324 351316
rect 12356 351284 12404 351316
rect 12436 351284 12484 351316
rect 12516 351284 12564 351316
rect 12596 351284 12644 351316
rect 12676 351284 12724 351316
rect 12756 351284 12804 351316
rect 12836 351284 12884 351316
rect 12916 351284 12964 351316
rect 12996 351284 13044 351316
rect 13076 351284 13124 351316
rect 13156 351284 13204 351316
rect 13236 351284 13284 351316
rect 13316 351284 13364 351316
rect 13396 351284 13444 351316
rect 13476 351284 13524 351316
rect 13556 351284 13604 351316
rect 13636 351284 13684 351316
rect 13716 351284 13764 351316
rect 13796 351284 13844 351316
rect 13876 351284 13924 351316
rect 13956 351284 14004 351316
rect 14036 351284 14084 351316
rect 14116 351284 14164 351316
rect 14196 351284 14244 351316
rect 14276 351284 14324 351316
rect 14356 351284 14404 351316
rect 14436 351284 14484 351316
rect 14516 351284 14564 351316
rect 14596 351284 14644 351316
rect 14676 351284 14724 351316
rect 14756 351284 14804 351316
rect 14836 351284 14884 351316
rect 14916 351284 14964 351316
rect 14996 351284 15044 351316
rect 15076 351284 15124 351316
rect 15156 351284 15204 351316
rect 15236 351284 15284 351316
rect 15316 351284 15364 351316
rect 15396 351284 15444 351316
rect 15476 351284 15524 351316
rect 15556 351284 15604 351316
rect 15636 351284 15684 351316
rect 15716 351284 15764 351316
rect 15796 351284 15844 351316
rect 15876 351284 15924 351316
rect 15956 351284 16004 351316
rect 16036 351284 16084 351316
rect 16116 351284 16164 351316
rect 16196 351284 16244 351316
rect 16276 351284 16324 351316
rect 16356 351284 16404 351316
rect 16436 351284 16484 351316
rect 16516 351284 16564 351316
rect 16596 351284 16644 351316
rect 16676 351284 16724 351316
rect 16756 351284 16804 351316
rect 16836 351284 16884 351316
rect 16916 351284 16964 351316
rect 16996 351284 17044 351316
rect 17076 351284 17124 351316
rect 17156 351284 17204 351316
rect 17236 351284 17284 351316
rect 17316 351284 17364 351316
rect 17396 351284 17444 351316
rect 17476 351284 17524 351316
rect 17556 351284 17604 351316
rect 17636 351284 17684 351316
rect 17716 351284 17764 351316
rect 17796 351284 17844 351316
rect 17876 351284 17924 351316
rect 17956 351284 18004 351316
rect 18036 351284 18084 351316
rect 18116 351284 18164 351316
rect 18196 351284 18244 351316
rect 18276 351284 18324 351316
rect 18356 351284 18404 351316
rect 18436 351284 18484 351316
rect 18516 351284 18564 351316
rect 18596 351284 18644 351316
rect 18676 351284 18724 351316
rect 18756 351284 18804 351316
rect 18836 351284 18884 351316
rect 18916 351284 18964 351316
rect 18996 351284 19044 351316
rect 19076 351284 19124 351316
rect 19156 351284 19204 351316
rect 19236 351284 19284 351316
rect 19316 351284 19364 351316
rect 19396 351284 19444 351316
rect 19476 351284 19524 351316
rect 19556 351284 19604 351316
rect 19636 351284 19684 351316
rect 19716 351284 19800 351316
rect 10640 351280 19800 351284
rect 10720 351236 19880 351240
rect 10720 351204 10724 351236
rect 10756 351204 10804 351236
rect 10836 351204 10884 351236
rect 10916 351204 10964 351236
rect 10996 351204 11044 351236
rect 11076 351204 11124 351236
rect 11156 351204 11204 351236
rect 11236 351204 11284 351236
rect 11316 351204 11364 351236
rect 11396 351204 11444 351236
rect 11476 351204 11524 351236
rect 11556 351204 11604 351236
rect 11636 351204 11684 351236
rect 11716 351204 11764 351236
rect 11796 351204 11844 351236
rect 11876 351204 11924 351236
rect 11956 351204 12004 351236
rect 12036 351204 12084 351236
rect 12116 351204 12164 351236
rect 12196 351204 12244 351236
rect 12276 351204 12324 351236
rect 12356 351204 12404 351236
rect 12436 351204 12484 351236
rect 12516 351204 12564 351236
rect 12596 351204 12644 351236
rect 12676 351204 12724 351236
rect 12756 351204 12804 351236
rect 12836 351204 12884 351236
rect 12916 351204 12964 351236
rect 12996 351204 13044 351236
rect 13076 351204 13124 351236
rect 13156 351204 13204 351236
rect 13236 351204 13284 351236
rect 13316 351204 13364 351236
rect 13396 351204 13444 351236
rect 13476 351204 13524 351236
rect 13556 351204 13604 351236
rect 13636 351204 13684 351236
rect 13716 351204 13764 351236
rect 13796 351204 13844 351236
rect 13876 351204 13924 351236
rect 13956 351204 14004 351236
rect 14036 351204 14084 351236
rect 14116 351204 14164 351236
rect 14196 351204 14244 351236
rect 14276 351204 14324 351236
rect 14356 351204 14404 351236
rect 14436 351204 14484 351236
rect 14516 351204 14564 351236
rect 14596 351204 14644 351236
rect 14676 351204 14724 351236
rect 14756 351204 14804 351236
rect 14836 351204 14884 351236
rect 14916 351204 14964 351236
rect 14996 351204 15044 351236
rect 15076 351204 15124 351236
rect 15156 351204 15204 351236
rect 15236 351204 15284 351236
rect 15316 351204 15364 351236
rect 15396 351204 15444 351236
rect 15476 351204 15524 351236
rect 15556 351204 15604 351236
rect 15636 351204 15684 351236
rect 15716 351204 15764 351236
rect 15796 351204 15844 351236
rect 15876 351204 15924 351236
rect 15956 351204 16004 351236
rect 16036 351204 16084 351236
rect 16116 351204 16164 351236
rect 16196 351204 16244 351236
rect 16276 351204 16324 351236
rect 16356 351204 16404 351236
rect 16436 351204 16484 351236
rect 16516 351204 16564 351236
rect 16596 351204 16644 351236
rect 16676 351204 16724 351236
rect 16756 351204 16804 351236
rect 16836 351204 16884 351236
rect 16916 351204 16964 351236
rect 16996 351204 17044 351236
rect 17076 351204 17124 351236
rect 17156 351204 17204 351236
rect 17236 351204 17284 351236
rect 17316 351204 17364 351236
rect 17396 351204 17444 351236
rect 17476 351204 17524 351236
rect 17556 351204 17604 351236
rect 17636 351204 17684 351236
rect 17716 351204 17764 351236
rect 17796 351204 17844 351236
rect 17876 351204 17924 351236
rect 17956 351204 18004 351236
rect 18036 351204 18084 351236
rect 18116 351204 18164 351236
rect 18196 351204 18244 351236
rect 18276 351204 18324 351236
rect 18356 351204 18404 351236
rect 18436 351204 18484 351236
rect 18516 351204 18564 351236
rect 18596 351204 18644 351236
rect 18676 351204 18724 351236
rect 18756 351204 18804 351236
rect 18836 351204 18884 351236
rect 18916 351204 18964 351236
rect 18996 351204 19044 351236
rect 19076 351204 19124 351236
rect 19156 351204 19204 351236
rect 19236 351204 19284 351236
rect 19316 351204 19364 351236
rect 19396 351204 19444 351236
rect 19476 351204 19524 351236
rect 19556 351204 19604 351236
rect 19636 351204 19684 351236
rect 19716 351204 19844 351236
rect 19876 351204 19880 351236
rect 10720 351200 19880 351204
rect 19680 351156 19880 351160
rect 19680 351124 19684 351156
rect 19716 351124 19844 351156
rect 19876 351124 19880 351156
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
rect 19680 351120 19880 351124
rect 19680 351076 19880 351080
rect 19680 351044 19684 351076
rect 19716 351044 19844 351076
rect 19876 351044 19880 351076
rect 19680 351040 19880 351044
rect 19680 350996 19880 351000
rect 19680 350964 19684 350996
rect 19716 350964 19844 350996
rect 19876 350964 19880 350996
rect 19680 350960 19880 350964
rect 19680 350916 19880 350920
rect 19680 350884 19684 350916
rect 19716 350884 19844 350916
rect 19876 350884 19880 350916
rect 19680 350880 19880 350884
rect 19680 350836 19880 350840
rect 19680 350804 19684 350836
rect 19716 350804 19844 350836
rect 19876 350804 19880 350836
rect 19680 350800 19880 350804
rect 19680 350756 19880 350760
rect 19680 350724 19684 350756
rect 19716 350724 19844 350756
rect 19876 350724 19880 350756
rect 19680 350720 19880 350724
rect 19680 350676 19880 350680
rect 19680 350644 19684 350676
rect 19716 350644 19844 350676
rect 19876 350644 19880 350676
rect 19680 350640 19880 350644
rect 19680 350596 19880 350600
rect 19680 350564 19684 350596
rect 19716 350564 19844 350596
rect 19876 350564 19880 350596
rect 19680 350560 19880 350564
rect 19680 350516 19880 350520
rect 19680 350484 19684 350516
rect 19716 350484 19844 350516
rect 19876 350484 19880 350516
rect 19680 350480 19880 350484
rect 19680 350436 19880 350440
rect 19680 350404 19684 350436
rect 19716 350404 19844 350436
rect 19876 350404 19880 350436
rect 19680 350400 19880 350404
rect 19680 350356 19880 350360
rect 19680 350324 19684 350356
rect 19716 350324 19844 350356
rect 19876 350324 19880 350356
rect 19680 350320 19880 350324
rect 19680 350276 19880 350280
rect 19680 350244 19684 350276
rect 19716 350244 19844 350276
rect 19876 350244 19880 350276
rect 19680 350240 19880 350244
rect 19680 350196 19880 350200
rect 19680 350164 19684 350196
rect 19716 350164 19844 350196
rect 19876 350164 19880 350196
rect 19680 350160 19880 350164
rect 19680 350116 19880 350120
rect 19680 350084 19684 350116
rect 19716 350084 19844 350116
rect 19876 350084 19880 350116
rect 19680 350080 19880 350084
rect 19680 350036 19880 350040
rect 19680 350004 19684 350036
rect 19716 350004 19844 350036
rect 19876 350004 19880 350036
rect 19680 350000 19880 350004
rect 19680 349956 19880 349960
rect 19680 349924 19684 349956
rect 19716 349924 19844 349956
rect 19876 349924 19880 349956
rect 19680 349920 19880 349924
rect 19680 349876 19880 349880
rect 19680 349844 19684 349876
rect 19716 349844 19844 349876
rect 19876 349844 19880 349876
rect 19680 349840 19880 349844
rect 19680 349796 19880 349800
rect 19680 349764 19684 349796
rect 19716 349764 19844 349796
rect 19876 349764 19880 349796
rect 19680 349760 19880 349764
rect 19680 349716 19880 349720
rect 19680 349684 19684 349716
rect 19716 349684 19844 349716
rect 19876 349684 19880 349716
rect 19680 349680 19880 349684
rect 19680 349636 19880 349640
rect 19680 349604 19684 349636
rect 19716 349604 19844 349636
rect 19876 349604 19880 349636
rect 19680 349600 19880 349604
rect 19680 349556 19880 349560
rect 19680 349524 19684 349556
rect 19716 349524 19844 349556
rect 19876 349524 19880 349556
rect 19680 349520 19880 349524
rect 19680 349476 19880 349480
rect 19680 349444 19684 349476
rect 19716 349444 19844 349476
rect 19876 349444 19880 349476
rect 19680 349440 19880 349444
rect 19680 349396 19880 349400
rect 19680 349364 19684 349396
rect 19716 349364 19844 349396
rect 19876 349364 19880 349396
rect 19680 349360 19880 349364
rect 19680 349316 19880 349320
rect 19680 349284 19684 349316
rect 19716 349284 19844 349316
rect 19876 349284 19880 349316
rect 19680 349280 19880 349284
rect 19680 349236 19880 349240
rect 19680 349204 19684 349236
rect 19716 349204 19844 349236
rect 19876 349204 19880 349236
rect 19680 349200 19880 349204
rect 19680 349156 19880 349160
rect 19680 349124 19684 349156
rect 19716 349124 19844 349156
rect 19876 349124 19880 349156
rect 19680 349120 19880 349124
rect 19680 349076 19880 349080
rect 19680 349044 19684 349076
rect 19716 349044 19844 349076
rect 19876 349044 19880 349076
rect 19680 349040 19880 349044
rect 19680 348996 19880 349000
rect 19680 348964 19684 348996
rect 19716 348964 19844 348996
rect 19876 348964 19880 348996
rect 19680 348960 19880 348964
rect 19680 348916 19880 348920
rect 19680 348884 19684 348916
rect 19716 348884 19844 348916
rect 19876 348884 19880 348916
rect 19680 348880 19880 348884
rect 19680 348836 19880 348840
rect 19680 348804 19684 348836
rect 19716 348804 19844 348836
rect 19876 348804 19880 348836
rect 19680 348800 19880 348804
rect 19680 348756 19880 348760
rect 19680 348724 19684 348756
rect 19716 348724 19844 348756
rect 19876 348724 19880 348756
rect 19680 348720 19880 348724
rect 19680 348676 19880 348680
rect 19680 348644 19684 348676
rect 19716 348644 19844 348676
rect 19876 348644 19880 348676
rect 19680 348640 19880 348644
rect 19680 348596 19880 348600
rect 19680 348564 19684 348596
rect 19716 348564 19844 348596
rect 19876 348564 19880 348596
rect 19680 348560 19880 348564
rect 19680 348516 19880 348520
rect 19680 348484 19684 348516
rect 19716 348484 19844 348516
rect 19876 348484 19880 348516
rect 19680 348480 19880 348484
rect 19680 348436 19880 348440
rect 19680 348404 19684 348436
rect 19716 348404 19844 348436
rect 19876 348404 19880 348436
rect 19680 348400 19880 348404
rect 19680 348356 19880 348360
rect 19680 348324 19684 348356
rect 19716 348324 19844 348356
rect 19876 348324 19880 348356
rect 19680 348320 19880 348324
rect 19680 348276 19880 348280
rect 19680 348244 19684 348276
rect 19716 348244 19844 348276
rect 19876 348244 19880 348276
rect 19680 348240 19880 348244
rect 19680 348196 19880 348200
rect 19680 348164 19684 348196
rect 19716 348164 19844 348196
rect 19876 348164 19880 348196
rect 19680 348160 19880 348164
rect 19680 348116 19880 348120
rect 19680 348084 19684 348116
rect 19716 348084 19844 348116
rect 19876 348084 19880 348116
rect 19680 348080 19880 348084
rect 19680 348036 19880 348040
rect 19680 348004 19684 348036
rect 19716 348004 19844 348036
rect 19876 348004 19880 348036
rect 19680 348000 19880 348004
rect 19680 347956 19880 347960
rect 19680 347924 19684 347956
rect 19716 347924 19844 347956
rect 19876 347924 19880 347956
rect 19680 347920 19880 347924
rect 19680 347876 19880 347880
rect 19680 347844 19684 347876
rect 19716 347844 19844 347876
rect 19876 347844 19880 347876
rect 19680 347840 19880 347844
rect 19680 347796 19880 347800
rect 19680 347764 19684 347796
rect 19716 347764 19844 347796
rect 19876 347764 19880 347796
rect 19680 347760 19880 347764
rect 19680 347716 19880 347720
rect 19680 347684 19684 347716
rect 19716 347684 19844 347716
rect 19876 347684 19880 347716
rect 19680 347680 19880 347684
rect 19680 347636 19880 347640
rect 19680 347604 19684 347636
rect 19716 347604 19844 347636
rect 19876 347604 19880 347636
rect 19680 347600 19880 347604
rect 19680 347556 19880 347560
rect 19680 347524 19684 347556
rect 19716 347524 19844 347556
rect 19876 347524 19880 347556
rect 19680 347520 19880 347524
rect 19680 347476 19880 347480
rect 19680 347444 19684 347476
rect 19716 347444 19844 347476
rect 19876 347444 19880 347476
rect 19680 347440 19880 347444
rect 19680 347396 19880 347400
rect 19680 347364 19684 347396
rect 19716 347364 19844 347396
rect 19876 347364 19880 347396
rect 19680 347360 19880 347364
rect 19680 347316 19880 347320
rect 19680 347284 19684 347316
rect 19716 347284 19844 347316
rect 19876 347284 19880 347316
rect 19680 347280 19880 347284
rect 19680 347236 19880 347240
rect 19680 347204 19684 347236
rect 19716 347204 19844 347236
rect 19876 347204 19880 347236
rect 19680 347200 19880 347204
rect 19680 347156 19880 347160
rect 19680 347124 19684 347156
rect 19716 347124 19844 347156
rect 19876 347124 19880 347156
rect 19680 347120 19880 347124
rect 19680 347076 19880 347080
rect 19680 347044 19684 347076
rect 19716 347044 19844 347076
rect 19876 347044 19880 347076
rect 19680 347040 19880 347044
rect 19680 346996 19880 347000
rect 19680 346964 19684 346996
rect 19716 346964 19844 346996
rect 19876 346964 19880 346996
rect 19680 346960 19880 346964
rect 19680 346916 19880 346920
rect 19680 346884 19684 346916
rect 19716 346884 19844 346916
rect 19876 346884 19880 346916
rect 19680 346880 19880 346884
rect 19680 346836 19880 346840
rect 19680 346804 19684 346836
rect 19716 346804 19844 346836
rect 19876 346804 19880 346836
rect 19680 346800 19880 346804
rect 19680 346756 19880 346760
rect 19680 346724 19684 346756
rect 19716 346724 19844 346756
rect 19876 346724 19880 346756
rect 19680 346720 19880 346724
rect 19680 346676 19880 346680
rect 19680 346644 19684 346676
rect 19716 346644 19844 346676
rect 19876 346644 19880 346676
rect 19680 346640 19880 346644
rect 19680 346596 19880 346600
rect 19680 346564 19684 346596
rect 19716 346564 19844 346596
rect 19876 346564 19880 346596
rect 19680 346560 19880 346564
rect 19680 346516 19880 346520
rect 19680 346484 19684 346516
rect 19716 346484 19844 346516
rect 19876 346484 19880 346516
rect 19680 346480 19880 346484
rect 19680 346436 19880 346440
rect 19680 346404 19684 346436
rect 19716 346404 19844 346436
rect 19876 346404 19880 346436
rect 19680 346400 19880 346404
rect 19680 346356 19880 346360
rect 19680 346324 19684 346356
rect 19716 346324 19844 346356
rect 19876 346324 19880 346356
rect 19680 346320 19880 346324
rect 19680 346276 19880 346280
rect 19680 346244 19684 346276
rect 19716 346244 19844 346276
rect 19876 346244 19880 346276
rect 19680 346240 19880 346244
rect 19680 346196 19880 346200
rect 19680 346164 19684 346196
rect 19716 346164 19844 346196
rect 19876 346164 19880 346196
rect 19680 346160 19880 346164
rect 19680 346116 19880 346120
rect 19680 346084 19684 346116
rect 19716 346084 19844 346116
rect 19876 346084 19880 346116
rect 19680 346080 19880 346084
rect 19680 346036 19880 346040
rect 19680 346004 19684 346036
rect 19716 346004 19844 346036
rect 19876 346004 19880 346036
rect 19680 346000 19880 346004
rect 19680 345956 19880 345960
rect 19680 345924 19684 345956
rect 19716 345924 19844 345956
rect 19876 345924 19880 345956
rect 19680 345920 19880 345924
rect 19680 345876 19880 345880
rect 19680 345844 19684 345876
rect 19716 345844 19844 345876
rect 19876 345844 19880 345876
rect 19680 345840 19880 345844
rect 19680 345796 19880 345800
rect 19680 345764 19684 345796
rect 19716 345764 19844 345796
rect 19876 345764 19880 345796
rect 19680 345760 19880 345764
rect 19680 345716 19880 345720
rect 19680 345684 19684 345716
rect 19716 345684 19844 345716
rect 19876 345684 19880 345716
rect 19680 345680 19880 345684
rect 19680 345636 19880 345640
rect 19680 345604 19684 345636
rect 19716 345604 19844 345636
rect 19876 345604 19880 345636
rect 19680 345600 19880 345604
rect 19680 345556 19880 345560
rect 19680 345524 19684 345556
rect 19716 345524 19844 345556
rect 19876 345524 19880 345556
rect 19680 345520 19880 345524
rect 19680 345476 19880 345480
rect 19680 345444 19684 345476
rect 19716 345444 19844 345476
rect 19876 345444 19880 345476
rect 19680 345440 19880 345444
rect 19680 345396 19880 345400
rect 19680 345364 19684 345396
rect 19716 345364 19844 345396
rect 19876 345364 19880 345396
rect 19680 345360 19880 345364
rect 19680 345316 19880 345320
rect 19680 345284 19684 345316
rect 19716 345284 19844 345316
rect 19876 345284 19880 345316
rect 19680 345280 19880 345284
rect 19680 345236 19880 345240
rect 19680 345204 19684 345236
rect 19716 345204 19844 345236
rect 19876 345204 19880 345236
rect 19680 345200 19880 345204
rect 19680 345156 19880 345160
rect 19680 345124 19684 345156
rect 19716 345124 19844 345156
rect 19876 345124 19880 345156
rect 19680 345120 19880 345124
rect 19680 345076 19880 345080
rect 19680 345044 19684 345076
rect 19716 345044 19844 345076
rect 19876 345044 19880 345076
rect 19680 345040 19880 345044
rect 19680 344996 19880 345000
rect 19680 344964 19684 344996
rect 19716 344964 19844 344996
rect 19876 344964 19880 344996
rect 19680 344960 19880 344964
rect 19680 344916 19880 344920
rect 19680 344884 19684 344916
rect 19716 344884 19844 344916
rect 19876 344884 19880 344916
rect 19680 344880 19880 344884
rect 19680 344836 19880 344840
rect 19680 344804 19684 344836
rect 19716 344804 19844 344836
rect 19876 344804 19880 344836
rect 19680 344800 19880 344804
rect 19680 344756 19880 344760
rect 19680 344724 19684 344756
rect 19716 344724 19844 344756
rect 19876 344724 19880 344756
rect 19680 344720 19880 344724
rect 19680 344676 19880 344680
rect 19680 344644 19684 344676
rect 19716 344644 19844 344676
rect 19876 344644 19880 344676
rect 19680 344640 19880 344644
rect 19680 344596 19880 344600
rect 19680 344564 19684 344596
rect 19716 344564 19844 344596
rect 19876 344564 19880 344596
rect 19680 344560 19880 344564
rect 19680 344516 19880 344520
rect 19680 344484 19684 344516
rect 19716 344484 19844 344516
rect 19876 344484 19880 344516
rect 19680 344480 19880 344484
rect 19680 344436 19880 344440
rect 19680 344404 19684 344436
rect 19716 344404 19844 344436
rect 19876 344404 19880 344436
rect 19680 344400 19880 344404
rect 19680 344356 19880 344360
rect 19680 344324 19684 344356
rect 19716 344324 19844 344356
rect 19876 344324 19880 344356
rect 19680 344320 19880 344324
rect 19680 344276 19880 344280
rect 19680 344244 19684 344276
rect 19716 344244 19844 344276
rect 19876 344244 19880 344276
rect 19680 344240 19880 344244
rect 19680 344196 19880 344200
rect 19680 344164 19684 344196
rect 19716 344164 19844 344196
rect 19876 344164 19880 344196
rect 19680 344160 19880 344164
rect 19680 344116 19880 344120
rect 19680 344084 19684 344116
rect 19716 344084 19844 344116
rect 19876 344084 19880 344116
rect 19680 344080 19880 344084
rect 19680 344036 19880 344040
rect 19680 344004 19684 344036
rect 19716 344004 19844 344036
rect 19876 344004 19880 344036
rect 19680 344000 19880 344004
rect 19680 343956 19880 343960
rect 19680 343924 19684 343956
rect 19716 343924 19844 343956
rect 19876 343924 19880 343956
rect 19680 343920 19880 343924
rect 19680 343876 19880 343880
rect 19680 343844 19684 343876
rect 19716 343844 19844 343876
rect 19876 343844 19880 343876
rect 19680 343840 19880 343844
rect 19680 343796 19880 343800
rect 19680 343764 19684 343796
rect 19716 343764 19844 343796
rect 19876 343764 19880 343796
rect 19680 343760 19880 343764
rect 19680 343716 19880 343720
rect 19680 343684 19684 343716
rect 19716 343684 19844 343716
rect 19876 343684 19880 343716
rect 19680 343680 19880 343684
rect 19680 343636 19880 343640
rect 19680 343604 19684 343636
rect 19716 343604 19844 343636
rect 19876 343604 19880 343636
rect 19680 343600 19880 343604
rect 19680 343556 19880 343560
rect 19680 343524 19684 343556
rect 19716 343524 19844 343556
rect 19876 343524 19880 343556
rect 19680 343520 19880 343524
rect 19680 343476 19880 343480
rect 19680 343444 19684 343476
rect 19716 343444 19844 343476
rect 19876 343444 19880 343476
rect 19680 343440 19880 343444
rect 19680 343396 19880 343400
rect 19680 343364 19684 343396
rect 19716 343364 19844 343396
rect 19876 343364 19880 343396
rect 19680 343360 19880 343364
rect 19680 343316 19880 343320
rect 19680 343284 19684 343316
rect 19716 343284 19844 343316
rect 19876 343284 19880 343316
rect 19680 343280 19880 343284
rect 19680 343236 19880 343240
rect 19680 343204 19684 343236
rect 19716 343204 19844 343236
rect 19876 343204 19880 343236
rect 19680 343200 19880 343204
rect 19680 343156 19880 343160
rect 19680 343124 19684 343156
rect 19716 343124 19844 343156
rect 19876 343124 19880 343156
rect 19680 343120 19880 343124
rect 19680 343076 19880 343080
rect 19680 343044 19684 343076
rect 19716 343044 19844 343076
rect 19876 343044 19880 343076
rect 19680 343040 19880 343044
rect 19680 342996 19880 343000
rect 19680 342964 19684 342996
rect 19716 342964 19844 342996
rect 19876 342964 19880 342996
rect 19680 342960 19880 342964
rect 19680 342916 19880 342920
rect 19680 342884 19684 342916
rect 19716 342884 19844 342916
rect 19876 342884 19880 342916
rect 19680 342880 19880 342884
rect 19680 342836 19880 342840
rect 19680 342804 19684 342836
rect 19716 342804 19844 342836
rect 19876 342804 19880 342836
rect 19680 342800 19880 342804
rect 19680 342756 19880 342760
rect 19680 342724 19684 342756
rect 19716 342724 19844 342756
rect 19876 342724 19880 342756
rect 19680 342720 19880 342724
rect 19680 342676 19880 342680
rect 19680 342644 19684 342676
rect 19716 342644 19844 342676
rect 19876 342644 19880 342676
rect 19680 342640 19880 342644
rect 19680 342596 19880 342600
rect 19680 342564 19684 342596
rect 19716 342564 19844 342596
rect 19876 342564 19880 342596
rect 19680 342560 19880 342564
rect 19680 342516 19880 342520
rect 19680 342484 19684 342516
rect 19716 342484 19844 342516
rect 19876 342484 19880 342516
rect 19680 342480 19880 342484
rect 19680 342436 19880 342440
rect 19680 342404 19684 342436
rect 19716 342404 19844 342436
rect 19876 342404 19880 342436
rect 19680 342400 19880 342404
rect 19680 342356 19880 342360
rect 19680 342324 19684 342356
rect 19716 342324 19844 342356
rect 19876 342324 19880 342356
rect 19680 342320 19880 342324
rect 19680 342276 19880 342280
rect 19680 342244 19684 342276
rect 19716 342244 19844 342276
rect 19876 342244 19880 342276
rect 19680 342240 19880 342244
rect 19680 342196 19880 342200
rect 19680 342164 19684 342196
rect 19716 342164 19844 342196
rect 19876 342164 19880 342196
rect 19680 342160 19880 342164
rect 19680 342116 19880 342120
rect 19680 342084 19684 342116
rect 19716 342084 19844 342116
rect 19876 342084 19880 342116
rect 19680 342080 19880 342084
rect 19680 342036 19880 342040
rect 19680 342004 19684 342036
rect 19716 342004 19844 342036
rect 19876 342004 19880 342036
rect 19680 342000 19880 342004
rect 19680 341956 19880 341960
rect 19680 341924 19684 341956
rect 19716 341924 19844 341956
rect 19876 341924 19880 341956
rect 19680 341920 19880 341924
rect 19680 341876 19880 341880
rect 19680 341844 19684 341876
rect 19716 341844 19844 341876
rect 19876 341844 19880 341876
rect 19680 341840 19880 341844
rect 19680 341796 19880 341800
rect 19680 341764 19684 341796
rect 19716 341764 19844 341796
rect 19876 341764 19880 341796
rect 19680 341760 19880 341764
rect 19680 341716 19880 341720
rect 19680 341684 19684 341716
rect 19716 341684 19844 341716
rect 19876 341684 19880 341716
rect 19680 341680 19880 341684
rect 19680 341636 19880 341640
rect 19680 341604 19684 341636
rect 19716 341604 19844 341636
rect 19876 341604 19880 341636
rect 19680 341600 19880 341604
rect 19680 341556 19880 341560
rect 19680 341524 19684 341556
rect 19716 341524 19844 341556
rect 19876 341524 19880 341556
rect 19680 341520 19880 341524
rect 19680 341476 19880 341480
rect 19680 341444 19684 341476
rect 19716 341444 19844 341476
rect 19876 341444 19880 341476
rect 19680 341440 19880 341444
rect 19680 341396 19880 341400
rect 19680 341364 19684 341396
rect 19716 341364 19844 341396
rect 19876 341364 19880 341396
rect 19680 341360 19880 341364
rect 19680 341316 19880 341320
rect 19680 341284 19684 341316
rect 19716 341284 19844 341316
rect 19876 341284 19880 341316
rect 19680 341280 19880 341284
rect 19680 341236 19880 341240
rect 19680 341204 19684 341236
rect 19716 341204 19844 341236
rect 19876 341204 19880 341236
rect 19680 341200 19880 341204
rect 19680 341156 19880 341160
rect 19680 341124 19684 341156
rect 19716 341124 19844 341156
rect 19876 341124 19880 341156
rect 19680 341120 19880 341124
rect 19680 341076 19880 341080
rect 19680 341044 19684 341076
rect 19716 341044 19844 341076
rect 19876 341044 19880 341076
rect 19680 341040 19880 341044
rect 19680 340996 19880 341000
rect 19680 340964 19684 340996
rect 19716 340964 19844 340996
rect 19876 340964 19880 340996
rect 19680 340960 19880 340964
rect 19680 340916 19880 340920
rect 19680 340884 19684 340916
rect 19716 340884 19844 340916
rect 19876 340884 19880 340916
rect 19680 340880 19880 340884
rect 19680 340836 19880 340840
rect 19680 340804 19684 340836
rect 19716 340804 19844 340836
rect 19876 340804 19880 340836
rect 19680 340800 19880 340804
rect 19680 340756 19880 340760
rect 19680 340724 19684 340756
rect 19716 340724 19844 340756
rect 19876 340724 19880 340756
rect 19680 340720 19880 340724
rect 19680 340676 19880 340680
rect 19680 340644 19684 340676
rect 19716 340644 19844 340676
rect 19876 340644 19880 340676
rect 19680 340640 19880 340644
rect 19680 340596 19880 340600
rect 19680 340564 19684 340596
rect 19716 340564 19844 340596
rect 19876 340564 19880 340596
rect 19680 340560 19880 340564
rect 19680 340516 19880 340520
rect 19680 340484 19684 340516
rect 19716 340484 19844 340516
rect 19876 340484 19880 340516
rect 19680 340480 19880 340484
rect 19680 340436 19880 340440
rect 19680 340404 19684 340436
rect 19716 340404 19844 340436
rect 19876 340404 19880 340436
rect 19680 340400 19880 340404
rect 19680 340356 19880 340360
rect 19680 340324 19684 340356
rect 19716 340324 19844 340356
rect 19876 340324 19880 340356
rect 19680 340320 19880 340324
rect 19680 340276 19880 340280
rect 19680 340244 19684 340276
rect 19716 340244 19844 340276
rect 19876 340244 19880 340276
rect 19680 340240 19880 340244
rect 19680 340196 19880 340200
rect 19680 340164 19684 340196
rect 19716 340164 19844 340196
rect 19876 340164 19880 340196
rect 19680 340160 19880 340164
rect 19680 340116 19880 340120
rect 19680 340084 19684 340116
rect 19716 340084 19844 340116
rect 19876 340084 19880 340116
rect 19680 340080 19880 340084
rect 19680 340036 19880 340040
rect 19680 340004 19684 340036
rect 19716 340004 19844 340036
rect 19876 340004 19880 340036
rect 19680 340000 19880 340004
rect 19680 339956 19880 339960
rect 19680 339924 19684 339956
rect 19716 339924 19844 339956
rect 19876 339924 19880 339956
rect 19680 339920 19880 339924
rect 19680 339876 19880 339880
rect 19680 339844 19684 339876
rect 19716 339844 19844 339876
rect 19876 339844 19880 339876
rect 19680 339840 19880 339844
rect 19680 339796 19880 339800
rect 19680 339764 19684 339796
rect 19716 339764 19844 339796
rect 19876 339764 19880 339796
rect 19680 339760 19880 339764
rect 19680 339716 19880 339720
rect 19680 339684 19684 339716
rect 19716 339684 19844 339716
rect 19876 339684 19880 339716
rect 19680 339680 19880 339684
rect 19680 339636 19880 339640
rect 19680 339604 19684 339636
rect 19716 339604 19844 339636
rect 19876 339604 19880 339636
rect 19680 339600 19880 339604
rect 19680 339556 19880 339560
rect 19680 339524 19684 339556
rect 19716 339524 19844 339556
rect 19876 339524 19880 339556
rect 19680 339520 19880 339524
rect 19680 339476 19880 339480
rect 19680 339444 19684 339476
rect 19716 339444 19844 339476
rect 19876 339444 19880 339476
rect 19680 339440 19880 339444
rect 19680 339396 19880 339400
rect 19680 339364 19684 339396
rect 19716 339364 19844 339396
rect 19876 339364 19880 339396
rect 19680 339360 19880 339364
rect 19680 339316 19880 339320
rect 19680 339284 19684 339316
rect 19716 339284 19844 339316
rect 19876 339284 19880 339316
rect 19680 339280 19880 339284
rect 19680 339236 19880 339240
rect 19680 339204 19684 339236
rect 19716 339204 19844 339236
rect 19876 339204 19880 339236
rect 19680 339200 19880 339204
rect 19680 339156 19880 339160
rect 19680 339124 19684 339156
rect 19716 339124 19844 339156
rect 19876 339124 19880 339156
rect 19680 339120 19880 339124
rect 19680 339076 19880 339080
rect 19680 339044 19684 339076
rect 19716 339044 19844 339076
rect 19876 339044 19880 339076
rect 19680 339040 19880 339044
rect 19680 338996 19880 339000
rect 19680 338964 19684 338996
rect 19716 338964 19844 338996
rect 19876 338964 19880 338996
rect 19680 338960 19880 338964
rect 19680 338916 19880 338920
rect 19680 338884 19684 338916
rect 19716 338884 19844 338916
rect 19876 338884 19880 338916
rect 19680 338880 19880 338884
rect 19680 338836 19880 338840
rect 19680 338804 19684 338836
rect 19716 338804 19844 338836
rect 19876 338804 19880 338836
rect 19680 338800 19880 338804
rect 19680 338756 19880 338760
rect 19680 338724 19684 338756
rect 19716 338724 19844 338756
rect 19876 338724 19880 338756
rect 19680 338720 19880 338724
rect 19680 338676 19880 338680
rect 19680 338644 19684 338676
rect 19716 338644 19844 338676
rect 19876 338644 19880 338676
rect 19680 338640 19880 338644
rect 19680 338596 19880 338600
rect 19680 338564 19684 338596
rect 19716 338564 19844 338596
rect 19876 338564 19880 338596
rect 19680 338560 19880 338564
rect 19680 338516 19880 338520
rect 19680 338484 19684 338516
rect 19716 338484 19844 338516
rect 19876 338484 19880 338516
rect 19680 338480 19880 338484
rect 19680 338436 19880 338440
rect 19680 338404 19684 338436
rect 19716 338404 19844 338436
rect 19876 338404 19880 338436
rect 19680 338400 19880 338404
rect 19680 338356 19880 338360
rect 19680 338324 19684 338356
rect 19716 338324 19844 338356
rect 19876 338324 19880 338356
rect 19680 338320 19880 338324
rect 19680 338276 19880 338280
rect 19680 338244 19684 338276
rect 19716 338244 19844 338276
rect 19876 338244 19880 338276
rect 19680 338240 19880 338244
rect 19680 338196 19880 338200
rect 19680 338164 19684 338196
rect 19716 338164 19844 338196
rect 19876 338164 19880 338196
rect 19680 338160 19880 338164
rect 19680 338116 19880 338120
rect 19680 338084 19684 338116
rect 19716 338084 19844 338116
rect 19876 338084 19880 338116
rect 19680 338080 19880 338084
rect 19680 338036 19880 338040
rect 19680 338004 19684 338036
rect 19716 338004 19844 338036
rect 19876 338004 19880 338036
rect 19680 338000 19880 338004
rect 19680 337956 19880 337960
rect 19680 337924 19684 337956
rect 19716 337924 19844 337956
rect 19876 337924 19880 337956
rect 19680 337920 19880 337924
rect 19680 337876 19880 337880
rect 19680 337844 19684 337876
rect 19716 337844 19844 337876
rect 19876 337844 19880 337876
rect 19680 337840 19880 337844
rect 19680 337796 19880 337800
rect 19680 337764 19684 337796
rect 19716 337764 19844 337796
rect 19876 337764 19880 337796
rect 19680 337760 19880 337764
rect 19680 337716 19880 337720
rect 19680 337684 19684 337716
rect 19716 337684 19844 337716
rect 19876 337684 19880 337716
rect 19680 337680 19880 337684
rect 19680 337636 19880 337640
rect 19680 337604 19684 337636
rect 19716 337604 19844 337636
rect 19876 337604 19880 337636
rect 19680 337600 19880 337604
rect 19680 337556 19880 337560
rect 19680 337524 19684 337556
rect 19716 337524 19844 337556
rect 19876 337524 19880 337556
rect 19680 337520 19880 337524
rect 19680 337476 19880 337480
rect 19680 337444 19684 337476
rect 19716 337444 19844 337476
rect 19876 337444 19880 337476
rect 19680 337440 19880 337444
rect 19680 337396 19880 337400
rect 19680 337364 19684 337396
rect 19716 337364 19844 337396
rect 19876 337364 19880 337396
rect 19680 337360 19880 337364
rect 19680 337316 19880 337320
rect 19680 337284 19684 337316
rect 19716 337284 19844 337316
rect 19876 337284 19880 337316
rect 19680 337280 19880 337284
rect 19680 337236 19880 337240
rect 19680 337204 19684 337236
rect 19716 337204 19844 337236
rect 19876 337204 19880 337236
rect 19680 337200 19880 337204
rect 19680 337156 19880 337160
rect 19680 337124 19684 337156
rect 19716 337124 19844 337156
rect 19876 337124 19880 337156
rect 19680 337120 19880 337124
rect 19680 337076 19880 337080
rect 19680 337044 19684 337076
rect 19716 337044 19844 337076
rect 19876 337044 19880 337076
rect 19680 337040 19880 337044
rect 19680 336996 19880 337000
rect 19680 336964 19684 336996
rect 19716 336964 19844 336996
rect 19876 336964 19880 336996
rect 19680 336960 19880 336964
rect 19680 336916 19880 336920
rect 19680 336884 19684 336916
rect 19716 336884 19844 336916
rect 19876 336884 19880 336916
rect 19680 336880 19880 336884
rect 19680 336836 19880 336840
rect 19680 336804 19684 336836
rect 19716 336804 19844 336836
rect 19876 336804 19880 336836
rect 19680 336800 19880 336804
rect 19680 336756 19880 336760
rect 19680 336724 19684 336756
rect 19716 336724 19844 336756
rect 19876 336724 19880 336756
rect 19680 336720 19880 336724
rect 19680 336676 19880 336680
rect 19680 336644 19684 336676
rect 19716 336644 19844 336676
rect 19876 336644 19880 336676
rect 19680 336640 19880 336644
rect 19680 336596 19880 336600
rect 19680 336564 19684 336596
rect 19716 336564 19844 336596
rect 19876 336564 19880 336596
rect 19680 336560 19880 336564
rect 19680 336516 19880 336520
rect 19680 336484 19684 336516
rect 19716 336484 19844 336516
rect 19876 336484 19880 336516
rect 19680 336480 19880 336484
rect 19680 336436 19880 336440
rect 19680 336404 19684 336436
rect 19716 336404 19844 336436
rect 19876 336404 19880 336436
rect 19680 336400 19880 336404
rect 19680 336356 19880 336360
rect 19680 336324 19684 336356
rect 19716 336324 19844 336356
rect 19876 336324 19880 336356
rect 19680 336320 19880 336324
rect 19680 336276 19880 336280
rect 19680 336244 19684 336276
rect 19716 336244 19844 336276
rect 19876 336244 19880 336276
rect 19680 336240 19880 336244
rect 19680 336196 19880 336200
rect 19680 336164 19684 336196
rect 19716 336164 19844 336196
rect 19876 336164 19880 336196
rect 19680 336160 19880 336164
rect 19680 336116 19880 336120
rect 19680 336084 19684 336116
rect 19716 336084 19844 336116
rect 19876 336084 19880 336116
rect 19680 336080 19880 336084
rect 19680 336036 19880 336040
rect 19680 336004 19684 336036
rect 19716 336004 19844 336036
rect 19876 336004 19880 336036
rect 19680 336000 19880 336004
rect 19680 335956 19880 335960
rect 19680 335924 19684 335956
rect 19716 335924 19844 335956
rect 19876 335924 19880 335956
rect 19680 335920 19880 335924
rect 19680 335876 19880 335880
rect 19680 335844 19684 335876
rect 19716 335844 19844 335876
rect 19876 335844 19880 335876
rect 19680 335840 19880 335844
rect 19680 335796 19880 335800
rect 19680 335764 19684 335796
rect 19716 335764 19844 335796
rect 19876 335764 19880 335796
rect 19680 335760 19880 335764
rect 19680 335716 19880 335720
rect 19680 335684 19684 335716
rect 19716 335684 19844 335716
rect 19876 335684 19880 335716
rect 19680 335680 19880 335684
rect 19680 335636 19880 335640
rect 19680 335604 19684 335636
rect 19716 335604 19844 335636
rect 19876 335604 19880 335636
rect 19680 335600 19880 335604
rect 19680 335556 19880 335560
rect 19680 335524 19684 335556
rect 19716 335524 19844 335556
rect 19876 335524 19880 335556
rect 19680 335520 19880 335524
rect 19680 335476 19880 335480
rect 19680 335444 19684 335476
rect 19716 335444 19844 335476
rect 19876 335444 19880 335476
rect 19680 335440 19880 335444
rect 19680 335396 19880 335400
rect 19680 335364 19684 335396
rect 19716 335364 19844 335396
rect 19876 335364 19880 335396
rect 19680 335360 19880 335364
rect 19680 335316 19880 335320
rect 19680 335284 19684 335316
rect 19716 335284 19844 335316
rect 19876 335284 19880 335316
rect 19680 335280 19880 335284
rect 19680 335236 19880 335240
rect 19680 335204 19684 335236
rect 19716 335204 19844 335236
rect 19876 335204 19880 335236
rect 19680 335200 19880 335204
rect 19680 335156 19880 335160
rect 19680 335124 19684 335156
rect 19716 335124 19844 335156
rect 19876 335124 19880 335156
rect 19680 335120 19880 335124
rect 19680 335076 19880 335080
rect 19680 335044 19684 335076
rect 19716 335044 19844 335076
rect 19876 335044 19880 335076
rect 19680 335040 19880 335044
rect 19680 334996 19880 335000
rect 19680 334964 19684 334996
rect 19716 334964 19844 334996
rect 19876 334964 19880 334996
rect 19680 334960 19880 334964
rect 19680 334916 19880 334920
rect 19680 334884 19684 334916
rect 19716 334884 19844 334916
rect 19876 334884 19880 334916
rect 19680 334880 19880 334884
rect 19680 334836 19880 334840
rect 19680 334804 19684 334836
rect 19716 334804 19844 334836
rect 19876 334804 19880 334836
rect 19680 334800 19880 334804
rect 19680 334756 19880 334760
rect 19680 334724 19684 334756
rect 19716 334724 19844 334756
rect 19876 334724 19880 334756
rect 19680 334720 19880 334724
rect 19680 334676 19880 334680
rect 19680 334644 19684 334676
rect 19716 334644 19844 334676
rect 19876 334644 19880 334676
rect 19680 334640 19880 334644
rect 19680 334596 19880 334600
rect 19680 334564 19684 334596
rect 19716 334564 19844 334596
rect 19876 334564 19880 334596
rect 19680 334560 19880 334564
rect 19680 334516 19880 334520
rect 19680 334484 19684 334516
rect 19716 334484 19844 334516
rect 19876 334484 19880 334516
rect 19680 334480 19880 334484
rect 19680 334436 19880 334440
rect 19680 334404 19684 334436
rect 19716 334404 19844 334436
rect 19876 334404 19880 334436
rect 19680 334400 19880 334404
rect 19680 334356 19880 334360
rect 19680 334324 19684 334356
rect 19716 334324 19844 334356
rect 19876 334324 19880 334356
rect 19680 334320 19880 334324
rect 19680 334276 19880 334280
rect 19680 334244 19684 334276
rect 19716 334244 19844 334276
rect 19876 334244 19880 334276
rect 19680 334240 19880 334244
rect 19680 334196 19880 334200
rect 19680 334164 19684 334196
rect 19716 334164 19844 334196
rect 19876 334164 19880 334196
rect 19680 334160 19880 334164
rect 19680 334116 19880 334120
rect 19680 334084 19684 334116
rect 19716 334084 19844 334116
rect 19876 334084 19880 334116
rect 19680 334080 19880 334084
rect 19680 334036 19880 334040
rect 19680 334004 19684 334036
rect 19716 334004 19844 334036
rect 19876 334004 19880 334036
rect 19680 334000 19880 334004
rect 19680 333956 19880 333960
rect 19680 333924 19684 333956
rect 19716 333924 19844 333956
rect 19876 333924 19880 333956
rect 19680 333920 19880 333924
rect 19680 333876 19880 333880
rect 19680 333844 19684 333876
rect 19716 333844 19844 333876
rect 19876 333844 19880 333876
rect 19680 333840 19880 333844
rect 19680 333796 19880 333800
rect 19680 333764 19684 333796
rect 19716 333764 19844 333796
rect 19876 333764 19880 333796
rect 19680 333760 19880 333764
rect 19680 333716 19880 333720
rect 19680 333684 19684 333716
rect 19716 333684 19844 333716
rect 19876 333684 19880 333716
rect 19680 333680 19880 333684
rect 19680 333636 19880 333640
rect 19680 333604 19684 333636
rect 19716 333604 19844 333636
rect 19876 333604 19880 333636
rect 19680 333600 19880 333604
rect 19680 333556 19880 333560
rect 19680 333524 19684 333556
rect 19716 333524 19844 333556
rect 19876 333524 19880 333556
rect 19680 333520 19880 333524
rect 19680 333476 19880 333480
rect 19680 333444 19684 333476
rect 19716 333444 19844 333476
rect 19876 333444 19880 333476
rect 19680 333440 19880 333444
rect 19680 333396 19880 333400
rect 19680 333364 19684 333396
rect 19716 333364 19844 333396
rect 19876 333364 19880 333396
rect 19680 333360 19880 333364
rect 19680 333316 19880 333320
rect 19680 333284 19684 333316
rect 19716 333284 19844 333316
rect 19876 333284 19880 333316
rect 19680 333280 19880 333284
rect 19680 333236 19880 333240
rect 19680 333204 19684 333236
rect 19716 333204 19844 333236
rect 19876 333204 19880 333236
rect 19680 333200 19880 333204
rect 19680 333156 19880 333160
rect 19680 333124 19684 333156
rect 19716 333124 19844 333156
rect 19876 333124 19880 333156
rect 19680 333120 19880 333124
rect 19680 333076 19880 333080
rect 19680 333044 19684 333076
rect 19716 333044 19844 333076
rect 19876 333044 19880 333076
rect 19680 333040 19880 333044
rect 19680 332996 19880 333000
rect 19680 332964 19684 332996
rect 19716 332964 19844 332996
rect 19876 332964 19880 332996
rect 19680 332960 19880 332964
rect 19680 332916 19880 332920
rect 19680 332884 19684 332916
rect 19716 332884 19844 332916
rect 19876 332884 19880 332916
rect 19680 332880 19880 332884
rect 19680 332836 19880 332840
rect 19680 332804 19684 332836
rect 19716 332804 19844 332836
rect 19876 332804 19880 332836
rect 19680 332800 19880 332804
rect 19680 332756 19880 332760
rect 19680 332724 19684 332756
rect 19716 332724 19844 332756
rect 19876 332724 19880 332756
rect 19680 332720 19880 332724
rect 19680 332676 19880 332680
rect 19680 332644 19684 332676
rect 19716 332644 19844 332676
rect 19876 332644 19880 332676
rect 19680 332640 19880 332644
rect 19680 332596 19880 332600
rect 19680 332564 19684 332596
rect 19716 332564 19844 332596
rect 19876 332564 19880 332596
rect 19680 332560 19880 332564
rect 19680 332516 19880 332520
rect 19680 332484 19684 332516
rect 19716 332484 19844 332516
rect 19876 332484 19880 332516
rect 19680 332480 19880 332484
rect 19680 332436 19880 332440
rect 19680 332404 19684 332436
rect 19716 332404 19844 332436
rect 19876 332404 19880 332436
rect 19680 332400 19880 332404
rect 19680 332356 19880 332360
rect 19680 332324 19684 332356
rect 19716 332324 19844 332356
rect 19876 332324 19880 332356
rect 19680 332320 19880 332324
rect 19680 332276 19880 332280
rect 19680 332244 19684 332276
rect 19716 332244 19844 332276
rect 19876 332244 19880 332276
rect 19680 332240 19880 332244
rect 19680 332196 19880 332200
rect 19680 332164 19684 332196
rect 19716 332164 19844 332196
rect 19876 332164 19880 332196
rect 19680 332160 19880 332164
rect 19680 332116 19880 332120
rect 19680 332084 19684 332116
rect 19716 332084 19844 332116
rect 19876 332084 19880 332116
rect 19680 332080 19880 332084
rect 19680 332036 19880 332040
rect 19680 332004 19684 332036
rect 19716 332004 19844 332036
rect 19876 332004 19880 332036
rect 19680 332000 19880 332004
rect 19680 331956 19880 331960
rect 19680 331924 19684 331956
rect 19716 331924 19844 331956
rect 19876 331924 19880 331956
rect 19680 331920 19880 331924
rect 19680 331876 19880 331880
rect 19680 331844 19684 331876
rect 19716 331844 19844 331876
rect 19876 331844 19880 331876
rect 19680 331840 19880 331844
rect 19680 331796 19880 331800
rect 19680 331764 19684 331796
rect 19716 331764 19844 331796
rect 19876 331764 19880 331796
rect 19680 331760 19880 331764
rect 19680 331716 19880 331720
rect 19680 331684 19684 331716
rect 19716 331684 19844 331716
rect 19876 331684 19880 331716
rect 19680 331680 19880 331684
rect 19680 331636 19880 331640
rect 19680 331604 19684 331636
rect 19716 331604 19844 331636
rect 19876 331604 19880 331636
rect 19680 331600 19880 331604
rect 19680 331556 19880 331560
rect 19680 331524 19684 331556
rect 19716 331524 19844 331556
rect 19876 331524 19880 331556
rect 19680 331520 19880 331524
rect 19680 331476 19880 331480
rect 19680 331444 19684 331476
rect 19716 331444 19844 331476
rect 19876 331444 19880 331476
rect 19680 331440 19880 331444
rect 19680 331396 19880 331400
rect 19680 331364 19684 331396
rect 19716 331364 19844 331396
rect 19876 331364 19880 331396
rect 19680 331360 19880 331364
rect 19680 331316 19880 331320
rect 19680 331284 19684 331316
rect 19716 331284 19844 331316
rect 19876 331284 19880 331316
rect 19680 331280 19880 331284
rect 19680 331236 19880 331240
rect 19680 331204 19684 331236
rect 19716 331204 19844 331236
rect 19876 331204 19880 331236
rect 19680 331200 19880 331204
rect 19680 331156 19880 331160
rect 19680 331124 19684 331156
rect 19716 331124 19844 331156
rect 19876 331124 19880 331156
rect 19680 331120 19880 331124
rect 19680 331076 19880 331080
rect 19680 331044 19684 331076
rect 19716 331044 19844 331076
rect 19876 331044 19880 331076
rect 19680 331040 19880 331044
rect 19680 330996 19880 331000
rect 19680 330964 19684 330996
rect 19716 330964 19844 330996
rect 19876 330964 19880 330996
rect 19680 330960 19880 330964
rect 19680 330916 19880 330920
rect 19680 330884 19684 330916
rect 19716 330884 19844 330916
rect 19876 330884 19880 330916
rect 19680 330880 19880 330884
rect 19680 330836 19880 330840
rect 19680 330804 19684 330836
rect 19716 330804 19844 330836
rect 19876 330804 19880 330836
rect 19680 330800 19880 330804
rect 19680 330756 19880 330760
rect 19680 330724 19684 330756
rect 19716 330724 19844 330756
rect 19876 330724 19880 330756
rect 19680 330720 19880 330724
rect 19680 330676 19880 330680
rect 19680 330644 19684 330676
rect 19716 330644 19844 330676
rect 19876 330644 19880 330676
rect 19680 330640 19880 330644
rect 19680 330596 19880 330600
rect 19680 330564 19684 330596
rect 19716 330564 19844 330596
rect 19876 330564 19880 330596
rect 19680 330560 19880 330564
rect 19680 330516 19880 330520
rect 19680 330484 19684 330516
rect 19716 330484 19844 330516
rect 19876 330484 19880 330516
rect 19680 330480 19880 330484
rect 19680 330436 19880 330440
rect 19680 330404 19684 330436
rect 19716 330404 19844 330436
rect 19876 330404 19880 330436
rect 19680 330400 19880 330404
rect 19680 330356 19880 330360
rect 19680 330324 19684 330356
rect 19716 330324 19844 330356
rect 19876 330324 19880 330356
rect 19680 330320 19880 330324
rect 19680 330276 19880 330280
rect 19680 330244 19684 330276
rect 19716 330244 19844 330276
rect 19876 330244 19880 330276
rect 19680 330240 19880 330244
rect 19680 330196 19880 330200
rect 19680 330164 19684 330196
rect 19716 330164 19844 330196
rect 19876 330164 19880 330196
rect 19680 330160 19880 330164
rect 19680 330116 19880 330120
rect 19680 330084 19684 330116
rect 19716 330084 19844 330116
rect 19876 330084 19880 330116
rect 19680 330080 19880 330084
rect 19680 330036 19880 330040
rect 19680 330004 19684 330036
rect 19716 330004 19844 330036
rect 19876 330004 19880 330036
rect 19680 330000 19880 330004
rect 19680 329956 19880 329960
rect 19680 329924 19684 329956
rect 19716 329924 19844 329956
rect 19876 329924 19880 329956
rect 19680 329920 19880 329924
rect 19680 329876 19880 329880
rect 19680 329844 19684 329876
rect 19716 329844 19844 329876
rect 19876 329844 19880 329876
rect 19680 329840 19880 329844
rect 19680 329796 19880 329800
rect 19680 329764 19684 329796
rect 19716 329764 19844 329796
rect 19876 329764 19880 329796
rect 19680 329760 19880 329764
rect 19680 329716 19880 329720
rect 19680 329684 19684 329716
rect 19716 329684 19844 329716
rect 19876 329684 19880 329716
rect 19680 329680 19880 329684
rect 19680 329636 19880 329640
rect 19680 329604 19684 329636
rect 19716 329604 19844 329636
rect 19876 329604 19880 329636
rect 19680 329600 19880 329604
rect 19680 329556 19880 329560
rect 19680 329524 19684 329556
rect 19716 329524 19844 329556
rect 19876 329524 19880 329556
rect 19680 329520 19880 329524
rect 19680 329476 19880 329480
rect 19680 329444 19684 329476
rect 19716 329444 19844 329476
rect 19876 329444 19880 329476
rect 19680 329440 19880 329444
rect 19680 329396 19880 329400
rect 19680 329364 19684 329396
rect 19716 329364 19844 329396
rect 19876 329364 19880 329396
rect 19680 329360 19880 329364
rect 19680 329316 19880 329320
rect 19680 329284 19684 329316
rect 19716 329284 19844 329316
rect 19876 329284 19880 329316
rect 19680 329280 19880 329284
rect 19680 329236 19880 329240
rect 19680 329204 19684 329236
rect 19716 329204 19844 329236
rect 19876 329204 19880 329236
rect 19680 329200 19880 329204
rect 19680 329156 19880 329160
rect 19680 329124 19684 329156
rect 19716 329124 19844 329156
rect 19876 329124 19880 329156
rect 19680 329120 19880 329124
rect 19680 329076 19880 329080
rect 19680 329044 19684 329076
rect 19716 329044 19844 329076
rect 19876 329044 19880 329076
rect 19680 329040 19880 329044
rect 19680 328996 19880 329000
rect 19680 328964 19684 328996
rect 19716 328964 19844 328996
rect 19876 328964 19880 328996
rect 19680 328960 19880 328964
rect 19680 328916 19880 328920
rect 19680 328884 19684 328916
rect 19716 328884 19844 328916
rect 19876 328884 19880 328916
rect 19680 328880 19880 328884
rect 19680 328836 19880 328840
rect 19680 328804 19684 328836
rect 19716 328804 19844 328836
rect 19876 328804 19880 328836
rect 19680 328800 19880 328804
rect 19680 328756 19880 328760
rect 19680 328724 19684 328756
rect 19716 328724 19844 328756
rect 19876 328724 19880 328756
rect 19680 328720 19880 328724
rect 19680 328676 19880 328680
rect 19680 328644 19684 328676
rect 19716 328644 19844 328676
rect 19876 328644 19880 328676
rect 19680 328640 19880 328644
rect 19680 328596 19880 328600
rect 19680 328564 19684 328596
rect 19716 328564 19844 328596
rect 19876 328564 19880 328596
rect 19680 328560 19880 328564
rect 19680 328516 19880 328520
rect 19680 328484 19684 328516
rect 19716 328484 19844 328516
rect 19876 328484 19880 328516
rect 19680 328480 19880 328484
rect 19680 328436 19880 328440
rect 19680 328404 19684 328436
rect 19716 328404 19844 328436
rect 19876 328404 19880 328436
rect 19680 328400 19880 328404
rect 19680 328356 19880 328360
rect 19680 328324 19684 328356
rect 19716 328324 19844 328356
rect 19876 328324 19880 328356
rect 19680 328320 19880 328324
rect 19680 328276 19880 328280
rect 19680 328244 19684 328276
rect 19716 328244 19844 328276
rect 19876 328244 19880 328276
rect 19680 328240 19880 328244
rect 19680 328196 19880 328200
rect 19680 328164 19684 328196
rect 19716 328164 19844 328196
rect 19876 328164 19880 328196
rect 19680 328160 19880 328164
rect 19680 328116 19880 328120
rect 19680 328084 19684 328116
rect 19716 328084 19844 328116
rect 19876 328084 19880 328116
rect 19680 328080 19880 328084
rect 19680 328036 19880 328040
rect 19680 328004 19684 328036
rect 19716 328004 19844 328036
rect 19876 328004 19880 328036
rect 19680 328000 19880 328004
rect 19680 327956 19880 327960
rect 19680 327924 19684 327956
rect 19716 327924 19844 327956
rect 19876 327924 19880 327956
rect 19680 327920 19880 327924
rect 19680 327876 19880 327880
rect 19680 327844 19684 327876
rect 19716 327844 19844 327876
rect 19876 327844 19880 327876
rect 19680 327840 19880 327844
rect 19680 327796 19880 327800
rect 19680 327764 19684 327796
rect 19716 327764 19844 327796
rect 19876 327764 19880 327796
rect 19680 327760 19880 327764
rect 19680 327716 19880 327720
rect 19680 327684 19684 327716
rect 19716 327684 19844 327716
rect 19876 327684 19880 327716
rect 19680 327680 19880 327684
rect 19680 327636 19880 327640
rect 19680 327604 19684 327636
rect 19716 327604 19844 327636
rect 19876 327604 19880 327636
rect 19680 327600 19880 327604
rect 19680 327556 19880 327560
rect 19680 327524 19684 327556
rect 19716 327524 19844 327556
rect 19876 327524 19880 327556
rect 19680 327520 19880 327524
rect 19680 327476 19880 327480
rect 19680 327444 19684 327476
rect 19716 327444 19844 327476
rect 19876 327444 19880 327476
rect 19680 327440 19880 327444
rect 19680 327396 19880 327400
rect 19680 327364 19684 327396
rect 19716 327364 19844 327396
rect 19876 327364 19880 327396
rect 19680 327360 19880 327364
rect 19680 327316 19880 327320
rect 19680 327284 19684 327316
rect 19716 327284 19844 327316
rect 19876 327284 19880 327316
rect 19680 327280 19880 327284
rect 19680 327236 19880 327240
rect 19680 327204 19684 327236
rect 19716 327204 19844 327236
rect 19876 327204 19880 327236
rect 19680 327200 19880 327204
rect 19680 327156 19880 327160
rect 19680 327124 19684 327156
rect 19716 327124 19844 327156
rect 19876 327124 19880 327156
rect 19680 327120 19880 327124
rect 19680 327076 19880 327080
rect 19680 327044 19684 327076
rect 19716 327044 19844 327076
rect 19876 327044 19880 327076
rect 19680 327040 19880 327044
rect 19680 326996 19880 327000
rect 19680 326964 19684 326996
rect 19716 326964 19844 326996
rect 19876 326964 19880 326996
rect 19680 326960 19880 326964
rect 19680 326916 19880 326920
rect 19680 326884 19684 326916
rect 19716 326884 19844 326916
rect 19876 326884 19880 326916
rect 19680 326880 19880 326884
rect 19680 326836 19880 326840
rect 19680 326804 19684 326836
rect 19716 326804 19844 326836
rect 19876 326804 19880 326836
rect 19680 326800 19880 326804
rect 19680 326756 19880 326760
rect 19680 326724 19684 326756
rect 19716 326724 19844 326756
rect 19876 326724 19880 326756
rect 19680 326720 19880 326724
rect 19680 326676 19880 326680
rect 19680 326644 19684 326676
rect 19716 326644 19844 326676
rect 19876 326644 19880 326676
rect 19680 326640 19880 326644
rect 19680 326596 19880 326600
rect 19680 326564 19684 326596
rect 19716 326564 19844 326596
rect 19876 326564 19880 326596
rect 19680 326560 19880 326564
rect 19680 326516 19880 326520
rect 19680 326484 19684 326516
rect 19716 326484 19844 326516
rect 19876 326484 19880 326516
rect 19680 326480 19880 326484
rect 19680 326436 19880 326440
rect 19680 326404 19684 326436
rect 19716 326404 19844 326436
rect 19876 326404 19880 326436
rect 19680 326400 19880 326404
rect 19680 326356 19880 326360
rect 19680 326324 19684 326356
rect 19716 326324 19844 326356
rect 19876 326324 19880 326356
rect 19680 326320 19880 326324
rect 19680 326276 19880 326280
rect 19680 326244 19684 326276
rect 19716 326244 19844 326276
rect 19876 326244 19880 326276
rect 19680 326240 19880 326244
rect 19680 326196 19880 326200
rect 19680 326164 19684 326196
rect 19716 326164 19844 326196
rect 19876 326164 19880 326196
rect 19680 326160 19880 326164
rect 19680 326116 19880 326120
rect 19680 326084 19684 326116
rect 19716 326084 19844 326116
rect 19876 326084 19880 326116
rect 19680 326080 19880 326084
rect 19680 326036 19880 326040
rect 19680 326004 19684 326036
rect 19716 326004 19844 326036
rect 19876 326004 19880 326036
rect 19680 326000 19880 326004
rect 19680 325956 19880 325960
rect 19680 325924 19684 325956
rect 19716 325924 19844 325956
rect 19876 325924 19880 325956
rect 19680 325920 19880 325924
rect 19680 325876 19880 325880
rect 19680 325844 19684 325876
rect 19716 325844 19844 325876
rect 19876 325844 19880 325876
rect 19680 325840 19880 325844
rect 19680 325796 19880 325800
rect 19680 325764 19684 325796
rect 19716 325764 19844 325796
rect 19876 325764 19880 325796
rect 19680 325760 19880 325764
rect 19680 325716 19880 325720
rect 19680 325684 19684 325716
rect 19716 325684 19844 325716
rect 19876 325684 19880 325716
rect 19680 325680 19880 325684
rect 19680 325636 19880 325640
rect 19680 325604 19684 325636
rect 19716 325604 19844 325636
rect 19876 325604 19880 325636
rect 19680 325600 19880 325604
rect 19680 325556 19880 325560
rect 19680 325524 19684 325556
rect 19716 325524 19844 325556
rect 19876 325524 19880 325556
rect 19680 325520 19880 325524
rect 19680 325476 19880 325480
rect 19680 325444 19684 325476
rect 19716 325444 19844 325476
rect 19876 325444 19880 325476
rect 19680 325440 19880 325444
rect 19680 325396 19880 325400
rect 19680 325364 19684 325396
rect 19716 325364 19844 325396
rect 19876 325364 19880 325396
rect 19680 325360 19880 325364
rect 19680 325316 19880 325320
rect 19680 325284 19684 325316
rect 19716 325284 19844 325316
rect 19876 325284 19880 325316
rect 19680 325280 19880 325284
rect 19680 325236 19880 325240
rect 19680 325204 19684 325236
rect 19716 325204 19844 325236
rect 19876 325204 19880 325236
rect 19680 325200 19880 325204
rect 19680 325156 19880 325160
rect 19680 325124 19684 325156
rect 19716 325124 19844 325156
rect 19876 325124 19880 325156
rect 19680 325120 19880 325124
rect 19680 325076 19880 325080
rect 19680 325044 19684 325076
rect 19716 325044 19844 325076
rect 19876 325044 19880 325076
rect 19680 325040 19880 325044
rect 19680 324996 19880 325000
rect 19680 324964 19684 324996
rect 19716 324964 19844 324996
rect 19876 324964 19880 324996
rect 19680 324960 19880 324964
rect 19680 324916 19880 324920
rect 19680 324884 19684 324916
rect 19716 324884 19844 324916
rect 19876 324884 19880 324916
rect 19680 324880 19880 324884
rect 19680 324836 19880 324840
rect 19680 324804 19684 324836
rect 19716 324804 19844 324836
rect 19876 324804 19880 324836
rect 19680 324800 19880 324804
rect 19680 324756 19880 324760
rect 19680 324724 19684 324756
rect 19716 324724 19844 324756
rect 19876 324724 19880 324756
rect 19680 324720 19880 324724
rect 19680 324676 19880 324680
rect 19680 324644 19684 324676
rect 19716 324644 19844 324676
rect 19876 324644 19880 324676
rect 19680 324640 19880 324644
rect 19680 324596 19880 324600
rect 19680 324564 19684 324596
rect 19716 324564 19844 324596
rect 19876 324564 19880 324596
rect 19680 324560 19880 324564
rect 19680 324516 19880 324520
rect 19680 324484 19684 324516
rect 19716 324484 19844 324516
rect 19876 324484 19880 324516
rect 19680 324480 19880 324484
rect 19680 324436 19880 324440
rect 19680 324404 19684 324436
rect 19716 324404 19844 324436
rect 19876 324404 19880 324436
rect 19680 324400 19880 324404
rect 19680 324356 19880 324360
rect 19680 324324 19684 324356
rect 19716 324324 19844 324356
rect 19876 324324 19880 324356
rect 19680 324320 19880 324324
rect 19680 324276 19880 324280
rect 19680 324244 19684 324276
rect 19716 324244 19844 324276
rect 19876 324244 19880 324276
rect 19680 324240 19880 324244
rect 19680 324196 19880 324200
rect 19680 324164 19684 324196
rect 19716 324164 19844 324196
rect 19876 324164 19880 324196
rect 19680 324160 19880 324164
rect 19680 324116 19880 324120
rect 19680 324084 19684 324116
rect 19716 324084 19844 324116
rect 19876 324084 19880 324116
rect 19680 324080 19880 324084
rect 19680 324036 19880 324040
rect 19680 324004 19684 324036
rect 19716 324004 19844 324036
rect 19876 324004 19880 324036
rect 19680 324000 19880 324004
rect 19680 323956 19880 323960
rect 19680 323924 19684 323956
rect 19716 323924 19844 323956
rect 19876 323924 19880 323956
rect 19680 323920 19880 323924
rect 19680 323876 19880 323880
rect 19680 323844 19684 323876
rect 19716 323844 19844 323876
rect 19876 323844 19880 323876
rect 19680 323840 19880 323844
rect 19680 323796 19880 323800
rect 19680 323764 19684 323796
rect 19716 323764 19844 323796
rect 19876 323764 19880 323796
rect 19680 323760 19880 323764
rect 19680 323716 19880 323720
rect 19680 323684 19684 323716
rect 19716 323684 19844 323716
rect 19876 323684 19880 323716
rect 19680 323680 19880 323684
rect 19680 323636 19880 323640
rect 19680 323604 19684 323636
rect 19716 323604 19844 323636
rect 19876 323604 19880 323636
rect 19680 323600 19880 323604
rect 19680 323556 19880 323560
rect 19680 323524 19684 323556
rect 19716 323524 19844 323556
rect 19876 323524 19880 323556
rect 19680 323520 19880 323524
rect 19680 323476 19880 323480
rect 19680 323444 19684 323476
rect 19716 323444 19844 323476
rect 19876 323444 19880 323476
rect 19680 323440 19880 323444
rect 19680 323396 19880 323400
rect 19680 323364 19684 323396
rect 19716 323364 19844 323396
rect 19876 323364 19880 323396
rect 19680 323360 19880 323364
rect 19680 323316 19880 323320
rect 19680 323284 19684 323316
rect 19716 323284 19844 323316
rect 19876 323284 19880 323316
rect 19680 323280 19880 323284
rect 19680 323236 19880 323240
rect 19680 323204 19684 323236
rect 19716 323204 19844 323236
rect 19876 323204 19880 323236
rect 19680 323200 19880 323204
rect 19680 323156 19880 323160
rect 19680 323124 19684 323156
rect 19716 323124 19844 323156
rect 19876 323124 19880 323156
rect 19680 323120 19880 323124
rect 19680 323076 19880 323080
rect 19680 323044 19684 323076
rect 19716 323044 19844 323076
rect 19876 323044 19880 323076
rect 19680 323040 19880 323044
rect 19680 322996 19880 323000
rect 19680 322964 19684 322996
rect 19716 322964 19844 322996
rect 19876 322964 19880 322996
rect 19680 322960 19880 322964
rect 19680 322916 19880 322920
rect 19680 322884 19684 322916
rect 19716 322884 19844 322916
rect 19876 322884 19880 322916
rect 19680 322880 19880 322884
rect 19680 322836 19880 322840
rect 19680 322804 19684 322836
rect 19716 322804 19844 322836
rect 19876 322804 19880 322836
rect 19680 322800 19880 322804
rect 19680 322756 19880 322760
rect 19680 322724 19684 322756
rect 19716 322724 19844 322756
rect 19876 322724 19880 322756
rect 19680 322720 19880 322724
rect 19680 322676 19880 322680
rect 19680 322644 19684 322676
rect 19716 322644 19844 322676
rect 19876 322644 19880 322676
rect 19680 322640 19880 322644
rect 19680 322596 19880 322600
rect 19680 322564 19684 322596
rect 19716 322564 19844 322596
rect 19876 322564 19880 322596
rect 19680 322560 19880 322564
rect 19680 322516 19880 322520
rect 19680 322484 19684 322516
rect 19716 322484 19844 322516
rect 19876 322484 19880 322516
rect 19680 322480 19880 322484
rect 19680 322436 19880 322440
rect 19680 322404 19684 322436
rect 19716 322404 19844 322436
rect 19876 322404 19880 322436
rect 19680 322400 19880 322404
rect 19680 322356 19880 322360
rect 19680 322324 19684 322356
rect 19716 322324 19844 322356
rect 19876 322324 19880 322356
rect 19680 322320 19880 322324
rect 19680 322276 19880 322280
rect 19680 322244 19684 322276
rect 19716 322244 19844 322276
rect 19876 322244 19880 322276
rect 19680 322240 19880 322244
rect 19680 322196 19880 322200
rect 19680 322164 19684 322196
rect 19716 322164 19844 322196
rect 19876 322164 19880 322196
rect 19680 322160 19880 322164
rect 19680 322116 19880 322120
rect 19680 322084 19684 322116
rect 19716 322084 19844 322116
rect 19876 322084 19880 322116
rect 19680 322080 19880 322084
rect 19680 322036 19880 322040
rect 19680 322004 19684 322036
rect 19716 322004 19844 322036
rect 19876 322004 19880 322036
rect 19680 322000 19880 322004
rect 19680 321956 19880 321960
rect 19680 321924 19684 321956
rect 19716 321924 19844 321956
rect 19876 321924 19880 321956
rect 19680 321920 19880 321924
rect 19680 321876 19880 321880
rect 19680 321844 19684 321876
rect 19716 321844 19844 321876
rect 19876 321844 19880 321876
rect 19680 321840 19880 321844
rect 19680 321796 19880 321800
rect 19680 321764 19684 321796
rect 19716 321764 19844 321796
rect 19876 321764 19880 321796
rect 19680 321760 19880 321764
rect 19680 321716 19880 321720
rect 19680 321684 19684 321716
rect 19716 321684 19844 321716
rect 19876 321684 19880 321716
rect 19680 321680 19880 321684
rect 19680 321636 19880 321640
rect 19680 321604 19684 321636
rect 19716 321604 19844 321636
rect 19876 321604 19880 321636
rect 19680 321600 19880 321604
rect 19680 321556 19880 321560
rect 19680 321524 19684 321556
rect 19716 321524 19844 321556
rect 19876 321524 19880 321556
rect 19680 321520 19880 321524
rect 19680 321476 19880 321480
rect 19680 321444 19684 321476
rect 19716 321444 19844 321476
rect 19876 321444 19880 321476
rect 19680 321440 19880 321444
rect 19680 321396 19880 321400
rect 19680 321364 19684 321396
rect 19716 321364 19844 321396
rect 19876 321364 19880 321396
rect 19680 321360 19880 321364
rect 19680 321316 19880 321320
rect 19680 321284 19684 321316
rect 19716 321284 19844 321316
rect 19876 321284 19880 321316
rect 19680 321280 19880 321284
rect 19680 321236 19880 321240
rect 19680 321204 19684 321236
rect 19716 321204 19844 321236
rect 19876 321204 19880 321236
rect 19680 321200 19880 321204
rect 19680 321156 19880 321160
rect 19680 321124 19684 321156
rect 19716 321124 19844 321156
rect 19876 321124 19880 321156
rect 19680 321120 19880 321124
rect 19680 321076 19880 321080
rect 19680 321044 19684 321076
rect 19716 321044 19844 321076
rect 19876 321044 19880 321076
rect 19680 321040 19880 321044
rect 19680 320996 19880 321000
rect 19680 320964 19684 320996
rect 19716 320964 19844 320996
rect 19876 320964 19880 320996
rect 19680 320960 19880 320964
rect 19680 320916 19880 320920
rect 19680 320884 19684 320916
rect 19716 320884 19844 320916
rect 19876 320884 19880 320916
rect 19680 320880 19880 320884
rect 19680 320836 19880 320840
rect 19680 320804 19684 320836
rect 19716 320804 19844 320836
rect 19876 320804 19880 320836
rect 19680 320800 19880 320804
rect 19680 320756 19880 320760
rect 19680 320724 19684 320756
rect 19716 320724 19844 320756
rect 19876 320724 19880 320756
rect 19680 320720 19880 320724
rect 19680 320676 19880 320680
rect 19680 320644 19684 320676
rect 19716 320644 19844 320676
rect 19876 320644 19880 320676
rect 19680 320640 19880 320644
rect 19680 320596 19880 320600
rect 19680 320564 19684 320596
rect 19716 320564 19844 320596
rect 19876 320564 19880 320596
rect 19680 320560 19880 320564
rect 19680 320516 19880 320520
rect 19680 320484 19684 320516
rect 19716 320484 19844 320516
rect 19876 320484 19880 320516
rect 19680 320480 19880 320484
rect 19680 320436 19880 320440
rect 19680 320404 19684 320436
rect 19716 320404 19844 320436
rect 19876 320404 19880 320436
rect 19680 320400 19880 320404
rect 19680 320356 19880 320360
rect 19680 320324 19684 320356
rect 19716 320324 19844 320356
rect 19876 320324 19880 320356
rect 19680 320320 19880 320324
rect 19680 320276 19880 320280
rect 19680 320244 19684 320276
rect 19716 320244 19844 320276
rect 19876 320244 19880 320276
rect 19680 320240 19880 320244
rect 19680 320196 19880 320200
rect 19680 320164 19684 320196
rect 19716 320164 19844 320196
rect 19876 320164 19880 320196
rect 19680 320160 19880 320164
rect 19680 320116 19880 320120
rect 19680 320084 19684 320116
rect 19716 320084 19844 320116
rect 19876 320084 19880 320116
rect 19680 320080 19880 320084
rect 19680 320036 19880 320040
rect 19680 320004 19684 320036
rect 19716 320004 19844 320036
rect 19876 320004 19880 320036
rect 19680 320000 19880 320004
rect 19680 319956 19880 319960
rect 19680 319924 19684 319956
rect 19716 319924 19844 319956
rect 19876 319924 19880 319956
rect 19680 319920 19880 319924
rect 19680 319876 19880 319880
rect 19680 319844 19684 319876
rect 19716 319844 19844 319876
rect 19876 319844 19880 319876
rect 19680 319840 19880 319844
rect 19680 319796 19880 319800
rect 19680 319764 19684 319796
rect 19716 319764 19844 319796
rect 19876 319764 19880 319796
rect 19680 319760 19880 319764
rect 19680 319716 19880 319720
rect 19680 319684 19684 319716
rect 19716 319684 19844 319716
rect 19876 319684 19880 319716
rect 19680 319680 19880 319684
rect 19680 319636 19880 319640
rect 19680 319604 19684 319636
rect 19716 319604 19844 319636
rect 19876 319604 19880 319636
rect 19680 319600 19880 319604
rect 19680 319556 19880 319560
rect 19680 319524 19684 319556
rect 19716 319524 19844 319556
rect 19876 319524 19880 319556
rect 19680 319520 19880 319524
rect 19680 319476 19880 319480
rect 19680 319444 19684 319476
rect 19716 319444 19844 319476
rect 19876 319444 19880 319476
rect 19680 319440 19880 319444
rect 19680 319396 19880 319400
rect 19680 319364 19684 319396
rect 19716 319364 19844 319396
rect 19876 319364 19880 319396
rect 19680 319360 19880 319364
rect 19680 319316 19880 319320
rect 19680 319284 19684 319316
rect 19716 319284 19844 319316
rect 19876 319284 19880 319316
rect 19680 319280 19880 319284
rect 19680 319236 19880 319240
rect 19680 319204 19684 319236
rect 19716 319204 19844 319236
rect 19876 319204 19880 319236
rect 19680 319200 19880 319204
rect 19680 319156 19880 319160
rect 19680 319124 19684 319156
rect 19716 319124 19844 319156
rect 19876 319124 19880 319156
rect 19680 319120 19880 319124
rect 19680 319076 19880 319080
rect 19680 319044 19684 319076
rect 19716 319044 19844 319076
rect 19876 319044 19880 319076
rect 19680 319040 19880 319044
rect 19680 318996 19880 319000
rect 19680 318964 19684 318996
rect 19716 318964 19844 318996
rect 19876 318964 19880 318996
rect 19680 318960 19880 318964
rect 19680 318916 19880 318920
rect 19680 318884 19684 318916
rect 19716 318884 19844 318916
rect 19876 318884 19880 318916
rect 19680 318880 19880 318884
rect 19680 318836 19880 318840
rect 19680 318804 19684 318836
rect 19716 318804 19844 318836
rect 19876 318804 19880 318836
rect 19680 318800 19880 318804
rect 19680 318756 19880 318760
rect 19680 318724 19684 318756
rect 19716 318724 19844 318756
rect 19876 318724 19880 318756
rect 19680 318720 19880 318724
rect 19680 318676 19880 318680
rect 19680 318644 19684 318676
rect 19716 318644 19844 318676
rect 19876 318644 19880 318676
rect 19680 318640 19880 318644
rect 19680 318596 19880 318600
rect 19680 318564 19684 318596
rect 19716 318564 19844 318596
rect 19876 318564 19880 318596
rect 19680 318560 19880 318564
rect 19680 318516 19880 318520
rect 19680 318484 19684 318516
rect 19716 318484 19844 318516
rect 19876 318484 19880 318516
rect 19680 318480 19880 318484
rect 19680 318436 19880 318440
rect 19680 318404 19684 318436
rect 19716 318404 19844 318436
rect 19876 318404 19880 318436
rect 19680 318400 19880 318404
rect 19680 318356 19880 318360
rect 19680 318324 19684 318356
rect 19716 318324 19844 318356
rect 19876 318324 19880 318356
rect 19680 318320 19880 318324
rect 19680 318276 19880 318280
rect 19680 318244 19684 318276
rect 19716 318244 19844 318276
rect 19876 318244 19880 318276
rect 19680 318240 19880 318244
rect 19680 318196 19880 318200
rect 19680 318164 19684 318196
rect 19716 318164 19844 318196
rect 19876 318164 19880 318196
rect 19680 318160 19880 318164
rect 19680 318116 19880 318120
rect 19680 318084 19684 318116
rect 19716 318084 19844 318116
rect 19876 318084 19880 318116
rect 19680 318080 19880 318084
rect 19680 318036 19880 318040
rect 19680 318004 19684 318036
rect 19716 318004 19844 318036
rect 19876 318004 19880 318036
rect 19680 318000 19880 318004
rect 19680 317956 19880 317960
rect 19680 317924 19684 317956
rect 19716 317924 19844 317956
rect 19876 317924 19880 317956
rect 19680 317920 19880 317924
rect 19680 317876 19880 317880
rect 19680 317844 19684 317876
rect 19716 317844 19844 317876
rect 19876 317844 19880 317876
rect 19680 317840 19880 317844
rect 19680 317796 19880 317800
rect 19680 317764 19684 317796
rect 19716 317764 19844 317796
rect 19876 317764 19880 317796
rect 19680 317760 19880 317764
rect 19680 317716 19880 317720
rect 19680 317684 19684 317716
rect 19716 317684 19844 317716
rect 19876 317684 19880 317716
rect 19680 317680 19880 317684
rect 19680 317636 19880 317640
rect 19680 317604 19684 317636
rect 19716 317604 19844 317636
rect 19876 317604 19880 317636
rect 19680 317600 19880 317604
rect 19680 317556 19880 317560
rect 19680 317524 19684 317556
rect 19716 317524 19844 317556
rect 19876 317524 19880 317556
rect 19680 317520 19880 317524
rect 19680 317476 19880 317480
rect 19680 317444 19684 317476
rect 19716 317444 19844 317476
rect 19876 317444 19880 317476
rect 19680 317440 19880 317444
rect 19680 317396 19880 317400
rect 19680 317364 19684 317396
rect 19716 317364 19844 317396
rect 19876 317364 19880 317396
rect 19680 317360 19880 317364
rect 19680 317316 19880 317320
rect 19680 317284 19684 317316
rect 19716 317284 19844 317316
rect 19876 317284 19880 317316
rect 19680 317280 19880 317284
rect 19680 317236 19880 317240
rect 19680 317204 19684 317236
rect 19716 317204 19844 317236
rect 19876 317204 19880 317236
rect 19680 317200 19880 317204
rect 19680 317156 19880 317160
rect 19680 317124 19684 317156
rect 19716 317124 19844 317156
rect 19876 317124 19880 317156
rect 19680 317120 19880 317124
rect 19680 317076 19880 317080
rect 19680 317044 19684 317076
rect 19716 317044 19844 317076
rect 19876 317044 19880 317076
rect 19680 317040 19880 317044
rect 19680 316996 19880 317000
rect 19680 316964 19684 316996
rect 19716 316964 19844 316996
rect 19876 316964 19880 316996
rect 19680 316960 19880 316964
rect 19680 316916 19880 316920
rect 19680 316884 19684 316916
rect 19716 316884 19844 316916
rect 19876 316884 19880 316916
rect 19680 316880 19880 316884
rect 19680 316836 19880 316840
rect 19680 316804 19684 316836
rect 19716 316804 19844 316836
rect 19876 316804 19880 316836
rect 19680 316800 19880 316804
rect 19680 316756 19880 316760
rect 19680 316724 19684 316756
rect 19716 316724 19844 316756
rect 19876 316724 19880 316756
rect 19680 316720 19880 316724
rect 19680 316676 19880 316680
rect 19680 316644 19684 316676
rect 19716 316644 19844 316676
rect 19876 316644 19880 316676
rect 19680 316640 19880 316644
rect 19680 316596 19880 316600
rect 19680 316564 19684 316596
rect 19716 316564 19844 316596
rect 19876 316564 19880 316596
rect 19680 316560 19880 316564
rect 19680 316516 19880 316520
rect 19680 316484 19684 316516
rect 19716 316484 19844 316516
rect 19876 316484 19880 316516
rect 19680 316480 19880 316484
rect 19680 316436 19880 316440
rect 19680 316404 19684 316436
rect 19716 316404 19844 316436
rect 19876 316404 19880 316436
rect 19680 316400 19880 316404
rect 19680 316356 19880 316360
rect 19680 316324 19684 316356
rect 19716 316324 19844 316356
rect 19876 316324 19880 316356
rect 19680 316320 19880 316324
rect 19680 316276 19880 316280
rect 19680 316244 19684 316276
rect 19716 316244 19844 316276
rect 19876 316244 19880 316276
rect 19680 316240 19880 316244
rect 19680 316196 19880 316200
rect 19680 316164 19684 316196
rect 19716 316164 19844 316196
rect 19876 316164 19880 316196
rect 19680 316160 19880 316164
rect 19680 316116 19880 316120
rect 19680 316084 19684 316116
rect 19716 316084 19844 316116
rect 19876 316084 19880 316116
rect 19680 316080 19880 316084
rect 19680 316036 19880 316040
rect 19680 316004 19684 316036
rect 19716 316004 19844 316036
rect 19876 316004 19880 316036
rect 19680 316000 19880 316004
rect 19680 315956 19880 315960
rect 19680 315924 19684 315956
rect 19716 315924 19844 315956
rect 19876 315924 19880 315956
rect 19680 315920 19880 315924
rect 19680 315876 19880 315880
rect 19680 315844 19684 315876
rect 19716 315844 19844 315876
rect 19876 315844 19880 315876
rect 19680 315840 19880 315844
rect 19680 315796 19880 315800
rect 19680 315764 19684 315796
rect 19716 315764 19844 315796
rect 19876 315764 19880 315796
rect 19680 315760 19880 315764
rect 19680 315716 19880 315720
rect 19680 315684 19684 315716
rect 19716 315684 19844 315716
rect 19876 315684 19880 315716
rect 19680 315680 19880 315684
rect 19680 315636 19880 315640
rect 19680 315604 19684 315636
rect 19716 315604 19844 315636
rect 19876 315604 19880 315636
rect 19680 315600 19880 315604
rect 19680 315556 19880 315560
rect 19680 315524 19684 315556
rect 19716 315524 19844 315556
rect 19876 315524 19880 315556
rect 19680 315520 19880 315524
rect 19680 315476 19880 315480
rect 19680 315444 19684 315476
rect 19716 315444 19844 315476
rect 19876 315444 19880 315476
rect 19680 315440 19880 315444
rect 19680 315396 19880 315400
rect 19680 315364 19684 315396
rect 19716 315364 19844 315396
rect 19876 315364 19880 315396
rect 19680 315360 19880 315364
rect 19680 315316 19880 315320
rect 19680 315284 19684 315316
rect 19716 315284 19844 315316
rect 19876 315284 19880 315316
rect 19680 315280 19880 315284
rect 19680 315236 19880 315240
rect 19680 315204 19684 315236
rect 19716 315204 19844 315236
rect 19876 315204 19880 315236
rect 19680 315200 19880 315204
rect 19680 315156 19880 315160
rect 19680 315124 19684 315156
rect 19716 315124 19844 315156
rect 19876 315124 19880 315156
rect 19680 315120 19880 315124
rect 19680 315076 19880 315080
rect 19680 315044 19684 315076
rect 19716 315044 19844 315076
rect 19876 315044 19880 315076
rect 19680 315040 19880 315044
rect 19680 314996 19880 315000
rect 19680 314964 19684 314996
rect 19716 314964 19844 314996
rect 19876 314964 19880 314996
rect 19680 314960 19880 314964
rect 19680 314916 19880 314920
rect 19680 314884 19684 314916
rect 19716 314884 19844 314916
rect 19876 314884 19880 314916
rect 19680 314880 19880 314884
rect 19680 314836 19880 314840
rect 19680 314804 19684 314836
rect 19716 314804 19844 314836
rect 19876 314804 19880 314836
rect 19680 314800 19880 314804
rect 19680 314756 19880 314760
rect 19680 314724 19684 314756
rect 19716 314724 19844 314756
rect 19876 314724 19880 314756
rect 19680 314720 19880 314724
rect 19680 314676 19880 314680
rect 19680 314644 19684 314676
rect 19716 314644 19844 314676
rect 19876 314644 19880 314676
rect 19680 314640 19880 314644
rect 19680 314596 19880 314600
rect 19680 314564 19684 314596
rect 19716 314564 19844 314596
rect 19876 314564 19880 314596
rect 19680 314560 19880 314564
rect 19680 314516 19880 314520
rect 19680 314484 19684 314516
rect 19716 314484 19844 314516
rect 19876 314484 19880 314516
rect 19680 314480 19880 314484
rect 19680 314436 19880 314440
rect 19680 314404 19684 314436
rect 19716 314404 19844 314436
rect 19876 314404 19880 314436
rect 19680 314400 19880 314404
rect 19680 314356 19880 314360
rect 19680 314324 19684 314356
rect 19716 314324 19844 314356
rect 19876 314324 19880 314356
rect 19680 314320 19880 314324
rect 19680 314276 19880 314280
rect 19680 314244 19684 314276
rect 19716 314244 19844 314276
rect 19876 314244 19880 314276
rect 19680 314240 19880 314244
rect 19680 314196 19880 314200
rect 19680 314164 19684 314196
rect 19716 314164 19844 314196
rect 19876 314164 19880 314196
rect 19680 314160 19880 314164
rect 19680 314116 19880 314120
rect 19680 314084 19684 314116
rect 19716 314084 19844 314116
rect 19876 314084 19880 314116
rect 19680 314080 19880 314084
rect 19680 314036 19880 314040
rect 19680 314004 19684 314036
rect 19716 314004 19844 314036
rect 19876 314004 19880 314036
rect 19680 314000 19880 314004
rect 19680 313956 19880 313960
rect 19680 313924 19684 313956
rect 19716 313924 19844 313956
rect 19876 313924 19880 313956
rect 19680 313920 19880 313924
rect 19680 313876 19880 313880
rect 19680 313844 19684 313876
rect 19716 313844 19844 313876
rect 19876 313844 19880 313876
rect 19680 313840 19880 313844
rect 19680 313796 19880 313800
rect 19680 313764 19684 313796
rect 19716 313764 19844 313796
rect 19876 313764 19880 313796
rect 19680 313760 19880 313764
rect 19680 313716 19880 313720
rect 19680 313684 19684 313716
rect 19716 313684 19844 313716
rect 19876 313684 19880 313716
rect 19680 313680 19880 313684
rect 19680 313636 19880 313640
rect 19680 313604 19684 313636
rect 19716 313604 19844 313636
rect 19876 313604 19880 313636
rect 19680 313600 19880 313604
rect 19680 313556 19880 313560
rect 19680 313524 19684 313556
rect 19716 313524 19844 313556
rect 19876 313524 19880 313556
rect 19680 313520 19880 313524
rect 19680 313476 19880 313480
rect 19680 313444 19684 313476
rect 19716 313444 19844 313476
rect 19876 313444 19880 313476
rect 19680 313440 19880 313444
rect 19680 313396 19880 313400
rect 19680 313364 19684 313396
rect 19716 313364 19844 313396
rect 19876 313364 19880 313396
rect 19680 313360 19880 313364
rect 19680 313316 19880 313320
rect 19680 313284 19684 313316
rect 19716 313284 19844 313316
rect 19876 313284 19880 313316
rect 19680 313280 19880 313284
rect 19680 313236 19880 313240
rect 19680 313204 19684 313236
rect 19716 313204 19844 313236
rect 19876 313204 19880 313236
rect 19680 313200 19880 313204
rect 19680 313156 19880 313160
rect 19680 313124 19684 313156
rect 19716 313124 19844 313156
rect 19876 313124 19880 313156
rect 19680 313120 19880 313124
rect 19680 313076 19880 313080
rect 19680 313044 19684 313076
rect 19716 313044 19844 313076
rect 19876 313044 19880 313076
rect 19680 313040 19880 313044
rect 19680 312996 19880 313000
rect 19680 312964 19684 312996
rect 19716 312964 19844 312996
rect 19876 312964 19880 312996
rect 19680 312960 19880 312964
rect 19680 312916 19880 312920
rect 19680 312884 19684 312916
rect 19716 312884 19844 312916
rect 19876 312884 19880 312916
rect 19680 312880 19880 312884
rect 19680 312836 19880 312840
rect 19680 312804 19684 312836
rect 19716 312804 19844 312836
rect 19876 312804 19880 312836
rect 19680 312800 19880 312804
rect 19680 312756 19880 312760
rect 19680 312724 19684 312756
rect 19716 312724 19844 312756
rect 19876 312724 19880 312756
rect 19680 312720 19880 312724
rect 19680 312676 19880 312680
rect 19680 312644 19684 312676
rect 19716 312644 19844 312676
rect 19876 312644 19880 312676
rect 19680 312640 19880 312644
rect 19680 312596 19880 312600
rect 19680 312564 19684 312596
rect 19716 312564 19844 312596
rect 19876 312564 19880 312596
rect 19680 312560 19880 312564
rect 19680 312516 19880 312520
rect 19680 312484 19684 312516
rect 19716 312484 19844 312516
rect 19876 312484 19880 312516
rect 19680 312480 19880 312484
rect 19680 312436 19880 312440
rect 19680 312404 19684 312436
rect 19716 312404 19844 312436
rect 19876 312404 19880 312436
rect 19680 312400 19880 312404
rect 19680 312356 19880 312360
rect 19680 312324 19684 312356
rect 19716 312324 19844 312356
rect 19876 312324 19880 312356
rect 19680 312320 19880 312324
rect 19680 312276 19880 312280
rect 19680 312244 19684 312276
rect 19716 312244 19844 312276
rect 19876 312244 19880 312276
rect 19680 312240 19880 312244
rect 19680 312196 19880 312200
rect 19680 312164 19684 312196
rect 19716 312164 19844 312196
rect 19876 312164 19880 312196
rect 19680 312160 19880 312164
rect 19680 312116 19880 312120
rect 19680 312084 19684 312116
rect 19716 312084 19844 312116
rect 19876 312084 19880 312116
rect 19680 312080 19880 312084
rect 19680 312036 19880 312040
rect 19680 312004 19684 312036
rect 19716 312004 19844 312036
rect 19876 312004 19880 312036
rect 19680 312000 19880 312004
rect 19680 311956 19880 311960
rect 19680 311924 19684 311956
rect 19716 311924 19844 311956
rect 19876 311924 19880 311956
rect 19680 311920 19880 311924
rect 19680 311876 19880 311880
rect 19680 311844 19684 311876
rect 19716 311844 19844 311876
rect 19876 311844 19880 311876
rect 19680 311840 19880 311844
rect 19680 311796 19880 311800
rect 19680 311764 19684 311796
rect 19716 311764 19844 311796
rect 19876 311764 19880 311796
rect 19680 311760 19880 311764
rect 19680 311716 19880 311720
rect 19680 311684 19684 311716
rect 19716 311684 19844 311716
rect 19876 311684 19880 311716
rect 19680 311680 19880 311684
rect 19680 311636 19880 311640
rect 19680 311604 19684 311636
rect 19716 311604 19844 311636
rect 19876 311604 19880 311636
rect 19680 311600 19880 311604
rect 19680 311556 19880 311560
rect 19680 311524 19684 311556
rect 19716 311524 19844 311556
rect 19876 311524 19880 311556
rect 19680 311520 19880 311524
rect 19680 311476 19880 311480
rect 19680 311444 19684 311476
rect 19716 311444 19844 311476
rect 19876 311444 19880 311476
rect 19680 311440 19880 311444
rect 19680 311396 19880 311400
rect 19680 311364 19684 311396
rect 19716 311364 19844 311396
rect 19876 311364 19880 311396
rect 19680 311360 19880 311364
rect 19680 311316 19880 311320
rect 19680 311284 19684 311316
rect 19716 311284 19844 311316
rect 19876 311284 19880 311316
rect 19680 311280 19880 311284
rect 19680 311236 19880 311240
rect 19680 311204 19684 311236
rect 19716 311204 19844 311236
rect 19876 311204 19880 311236
rect 19680 311200 19880 311204
rect 19680 311156 19880 311160
rect 19680 311124 19684 311156
rect 19716 311124 19844 311156
rect 19876 311124 19880 311156
rect 19680 311120 19880 311124
rect 19680 311076 19880 311080
rect 19680 311044 19684 311076
rect 19716 311044 19844 311076
rect 19876 311044 19880 311076
rect 19680 311040 19880 311044
rect 19680 310996 19880 311000
rect 19680 310964 19684 310996
rect 19716 310964 19844 310996
rect 19876 310964 19880 310996
rect 19680 310960 19880 310964
rect 19680 310916 19880 310920
rect 19680 310884 19684 310916
rect 19716 310884 19844 310916
rect 19876 310884 19880 310916
rect 19680 310880 19880 310884
rect 19680 310836 19880 310840
rect 19680 310804 19684 310836
rect 19716 310804 19844 310836
rect 19876 310804 19880 310836
rect 19680 310800 19880 310804
rect 19680 310756 19880 310760
rect 19680 310724 19684 310756
rect 19716 310724 19844 310756
rect 19876 310724 19880 310756
rect 19680 310720 19880 310724
rect 19680 310676 19880 310680
rect 19680 310644 19684 310676
rect 19716 310644 19844 310676
rect 19876 310644 19880 310676
rect 19680 310640 19880 310644
rect 19680 310596 19880 310600
rect 19680 310564 19684 310596
rect 19716 310564 19844 310596
rect 19876 310564 19880 310596
rect 19680 310560 19880 310564
rect 19680 310516 19880 310520
rect 19680 310484 19684 310516
rect 19716 310484 19844 310516
rect 19876 310484 19880 310516
rect 19680 310480 19880 310484
rect 19680 310436 19880 310440
rect 19680 310404 19684 310436
rect 19716 310404 19844 310436
rect 19876 310404 19880 310436
rect 19680 310400 19880 310404
rect 19680 310356 19880 310360
rect 19680 310324 19684 310356
rect 19716 310324 19844 310356
rect 19876 310324 19880 310356
rect 19680 310320 19880 310324
rect 19680 310276 19880 310280
rect 19680 310244 19684 310276
rect 19716 310244 19844 310276
rect 19876 310244 19880 310276
rect 19680 310240 19880 310244
rect 19680 310196 19880 310200
rect 19680 310164 19684 310196
rect 19716 310164 19844 310196
rect 19876 310164 19880 310196
rect 19680 310160 19880 310164
rect 19680 310116 19880 310120
rect 19680 310084 19684 310116
rect 19716 310084 19844 310116
rect 19876 310084 19880 310116
rect 19680 310080 19880 310084
rect 19680 310036 19880 310040
rect 19680 310004 19684 310036
rect 19716 310004 19844 310036
rect 19876 310004 19880 310036
rect 19680 310000 19880 310004
rect 19680 309956 19880 309960
rect 19680 309924 19684 309956
rect 19716 309924 19844 309956
rect 19876 309924 19880 309956
rect 19680 309920 19880 309924
rect 19680 309876 19880 309880
rect 19680 309844 19684 309876
rect 19716 309844 19844 309876
rect 19876 309844 19880 309876
rect 19680 309840 19880 309844
rect 19680 309796 19880 309800
rect 19680 309764 19684 309796
rect 19716 309764 19844 309796
rect 19876 309764 19880 309796
rect 19680 309760 19880 309764
rect 19680 309716 19880 309720
rect 19680 309684 19684 309716
rect 19716 309684 19844 309716
rect 19876 309684 19880 309716
rect 19680 309680 19880 309684
rect 19680 309636 19880 309640
rect 19680 309604 19684 309636
rect 19716 309604 19844 309636
rect 19876 309604 19880 309636
rect 19680 309600 19880 309604
rect 19680 309556 19880 309560
rect 19680 309524 19684 309556
rect 19716 309524 19844 309556
rect 19876 309524 19880 309556
rect 19680 309520 19880 309524
rect 19680 309476 19880 309480
rect 19680 309444 19684 309476
rect 19716 309444 19844 309476
rect 19876 309444 19880 309476
rect 19680 309440 19880 309444
rect 19680 309396 19880 309400
rect 19680 309364 19684 309396
rect 19716 309364 19844 309396
rect 19876 309364 19880 309396
rect 19680 309360 19880 309364
rect 19680 309316 19880 309320
rect 19680 309284 19684 309316
rect 19716 309284 19844 309316
rect 19876 309284 19880 309316
rect 19680 309280 19880 309284
rect 19680 309236 19880 309240
rect 19680 309204 19684 309236
rect 19716 309204 19844 309236
rect 19876 309204 19880 309236
rect 19680 309200 19880 309204
rect 19680 309156 19880 309160
rect 19680 309124 19684 309156
rect 19716 309124 19844 309156
rect 19876 309124 19880 309156
rect 19680 309120 19880 309124
rect 19680 309076 19880 309080
rect 19680 309044 19684 309076
rect 19716 309044 19844 309076
rect 19876 309044 19880 309076
rect 19680 309040 19880 309044
rect 19680 308996 19880 309000
rect 19680 308964 19684 308996
rect 19716 308964 19844 308996
rect 19876 308964 19880 308996
rect 19680 308960 19880 308964
rect 19680 308916 19880 308920
rect 19680 308884 19684 308916
rect 19716 308884 19844 308916
rect 19876 308884 19880 308916
rect 19680 308880 19880 308884
rect 19680 308836 19880 308840
rect 19680 308804 19684 308836
rect 19716 308804 19844 308836
rect 19876 308804 19880 308836
rect 19680 308800 19880 308804
rect 19680 308756 19880 308760
rect 19680 308724 19684 308756
rect 19716 308724 19844 308756
rect 19876 308724 19880 308756
rect 19680 308720 19880 308724
rect 19680 308676 19880 308680
rect 19680 308644 19684 308676
rect 19716 308644 19844 308676
rect 19876 308644 19880 308676
rect 19680 308640 19880 308644
rect 19680 308596 19880 308600
rect 19680 308564 19684 308596
rect 19716 308564 19844 308596
rect 19876 308564 19880 308596
rect 19680 308560 19880 308564
rect 19680 308516 19880 308520
rect 19680 308484 19684 308516
rect 19716 308484 19844 308516
rect 19876 308484 19880 308516
rect 19680 308480 19880 308484
rect 19680 308436 19880 308440
rect 19680 308404 19684 308436
rect 19716 308404 19844 308436
rect 19876 308404 19880 308436
rect 19680 308400 19880 308404
rect 19680 308356 19880 308360
rect 19680 308324 19684 308356
rect 19716 308324 19844 308356
rect 19876 308324 19880 308356
rect 19680 308320 19880 308324
rect 19680 308276 19880 308280
rect 19680 308244 19684 308276
rect 19716 308244 19844 308276
rect 19876 308244 19880 308276
rect 19680 308240 19880 308244
rect 19680 308196 19880 308200
rect 19680 308164 19684 308196
rect 19716 308164 19844 308196
rect 19876 308164 19880 308196
rect 19680 308160 19880 308164
rect 19680 308116 19880 308120
rect 19680 308084 19684 308116
rect 19716 308084 19844 308116
rect 19876 308084 19880 308116
rect 19680 308080 19880 308084
rect 19680 308036 19880 308040
rect 19680 308004 19684 308036
rect 19716 308004 19844 308036
rect 19876 308004 19880 308036
rect 19680 308000 19880 308004
rect 19680 307956 19880 307960
rect 19680 307924 19684 307956
rect 19716 307924 19844 307956
rect 19876 307924 19880 307956
rect 19680 307920 19880 307924
rect 19680 307876 19880 307880
rect 19680 307844 19684 307876
rect 19716 307844 19844 307876
rect 19876 307844 19880 307876
rect 19680 307840 19880 307844
rect 19680 307796 19880 307800
rect 19680 307764 19684 307796
rect 19716 307764 19844 307796
rect 19876 307764 19880 307796
rect 19680 307760 19880 307764
rect 19680 307716 19880 307720
rect 19680 307684 19684 307716
rect 19716 307684 19844 307716
rect 19876 307684 19880 307716
rect 19680 307680 19880 307684
rect 19680 307636 19880 307640
rect 19680 307604 19684 307636
rect 19716 307604 19844 307636
rect 19876 307604 19880 307636
rect 19680 307600 19880 307604
rect 19680 307556 19880 307560
rect 19680 307524 19684 307556
rect 19716 307524 19844 307556
rect 19876 307524 19880 307556
rect 19680 307520 19880 307524
rect 19680 307476 19880 307480
rect 19680 307444 19684 307476
rect 19716 307444 19844 307476
rect 19876 307444 19880 307476
rect 19680 307440 19880 307444
rect 19680 307396 19880 307400
rect 19680 307364 19684 307396
rect 19716 307364 19844 307396
rect 19876 307364 19880 307396
rect 19680 307360 19880 307364
rect 19680 307316 19880 307320
rect 19680 307284 19684 307316
rect 19716 307284 19844 307316
rect 19876 307284 19880 307316
rect 19680 307280 19880 307284
rect 19680 307236 19880 307240
rect 19680 307204 19684 307236
rect 19716 307204 19844 307236
rect 19876 307204 19880 307236
rect 19680 307200 19880 307204
rect 19680 307156 19880 307160
rect 19680 307124 19684 307156
rect 19716 307124 19844 307156
rect 19876 307124 19880 307156
rect 19680 307120 19880 307124
rect 19680 307076 19880 307080
rect 19680 307044 19684 307076
rect 19716 307044 19844 307076
rect 19876 307044 19880 307076
rect 19680 307040 19880 307044
rect 19680 306996 19880 307000
rect 19680 306964 19684 306996
rect 19716 306964 19844 306996
rect 19876 306964 19880 306996
rect 19680 306960 19880 306964
rect 19680 306916 19880 306920
rect 19680 306884 19684 306916
rect 19716 306884 19844 306916
rect 19876 306884 19880 306916
rect 19680 306880 19880 306884
rect 19680 306836 19880 306840
rect 19680 306804 19684 306836
rect 19716 306804 19844 306836
rect 19876 306804 19880 306836
rect 19680 306800 19880 306804
rect 19680 306756 19880 306760
rect 19680 306724 19684 306756
rect 19716 306724 19844 306756
rect 19876 306724 19880 306756
rect 19680 306720 19880 306724
rect 19680 306676 19880 306680
rect 19680 306644 19684 306676
rect 19716 306644 19844 306676
rect 19876 306644 19880 306676
rect 19680 306640 19880 306644
rect 19680 306596 19880 306600
rect 19680 306564 19684 306596
rect 19716 306564 19844 306596
rect 19876 306564 19880 306596
rect 19680 306560 19880 306564
rect 19680 306516 19880 306520
rect 19680 306484 19684 306516
rect 19716 306484 19844 306516
rect 19876 306484 19880 306516
rect 19680 306480 19880 306484
rect 19680 306436 19880 306440
rect 19680 306404 19684 306436
rect 19716 306404 19844 306436
rect 19876 306404 19880 306436
rect 19680 306400 19880 306404
rect 19680 306356 19880 306360
rect 19680 306324 19684 306356
rect 19716 306324 19844 306356
rect 19876 306324 19880 306356
rect 19680 306320 19880 306324
rect 19680 306276 19880 306280
rect 19680 306244 19684 306276
rect 19716 306244 19844 306276
rect 19876 306244 19880 306276
rect 19680 306240 19880 306244
rect 19680 306196 19880 306200
rect 19680 306164 19684 306196
rect 19716 306164 19844 306196
rect 19876 306164 19880 306196
rect 19680 306160 19880 306164
rect 19680 306116 19880 306120
rect 19680 306084 19684 306116
rect 19716 306084 19844 306116
rect 19876 306084 19880 306116
rect 19680 306080 19880 306084
rect 19680 306036 19880 306040
rect 19680 306004 19684 306036
rect 19716 306004 19844 306036
rect 19876 306004 19880 306036
rect 19680 306000 19880 306004
rect 19680 305956 19880 305960
rect 19680 305924 19684 305956
rect 19716 305924 19844 305956
rect 19876 305924 19880 305956
rect 19680 305920 19880 305924
rect 19680 305876 19880 305880
rect 19680 305844 19684 305876
rect 19716 305844 19844 305876
rect 19876 305844 19880 305876
rect 19680 305840 19880 305844
rect 19680 305796 19880 305800
rect 19680 305764 19684 305796
rect 19716 305764 19844 305796
rect 19876 305764 19880 305796
rect 19680 305760 19880 305764
rect 19680 305716 19880 305720
rect 19680 305684 19684 305716
rect 19716 305684 19844 305716
rect 19876 305684 19880 305716
rect 19680 305680 19880 305684
rect 19680 305636 19880 305640
rect 19680 305604 19684 305636
rect 19716 305604 19844 305636
rect 19876 305604 19880 305636
rect 19680 305600 19880 305604
rect 19680 305556 19880 305560
rect 19680 305524 19684 305556
rect 19716 305524 19844 305556
rect 19876 305524 19880 305556
rect 19680 305520 19880 305524
rect 19680 305476 19880 305480
rect 19680 305444 19684 305476
rect 19716 305444 19844 305476
rect 19876 305444 19880 305476
rect 19680 305440 19880 305444
rect 19680 305396 19880 305400
rect 19680 305364 19684 305396
rect 19716 305364 19844 305396
rect 19876 305364 19880 305396
rect 19680 305360 19880 305364
rect 19680 305316 19880 305320
rect 19680 305284 19684 305316
rect 19716 305284 19844 305316
rect 19876 305284 19880 305316
rect 19680 305280 19880 305284
rect 19680 305236 19880 305240
rect 19680 305204 19684 305236
rect 19716 305204 19844 305236
rect 19876 305204 19880 305236
rect 19680 305200 19880 305204
rect 19680 305156 19880 305160
rect 19680 305124 19684 305156
rect 19716 305124 19844 305156
rect 19876 305124 19880 305156
rect 19680 305120 19880 305124
rect 19680 305076 19880 305080
rect 19680 305044 19684 305076
rect 19716 305044 19844 305076
rect 19876 305044 19880 305076
rect 19680 305040 19880 305044
rect 19680 304996 19880 305000
rect 19680 304964 19684 304996
rect 19716 304964 19844 304996
rect 19876 304964 19880 304996
rect 19680 304960 19880 304964
rect 19680 304916 19880 304920
rect 19680 304884 19684 304916
rect 19716 304884 19844 304916
rect 19876 304884 19880 304916
rect 19680 304880 19880 304884
rect 19680 304836 19880 304840
rect 19680 304804 19684 304836
rect 19716 304804 19844 304836
rect 19876 304804 19880 304836
rect 19680 304800 19880 304804
rect 19680 304756 19880 304760
rect 19680 304724 19684 304756
rect 19716 304724 19844 304756
rect 19876 304724 19880 304756
rect 19680 304720 19880 304724
rect 19680 304676 19880 304680
rect 19680 304644 19684 304676
rect 19716 304644 19844 304676
rect 19876 304644 19880 304676
rect 19680 304640 19880 304644
rect 19680 304596 19880 304600
rect 19680 304564 19684 304596
rect 19716 304564 19844 304596
rect 19876 304564 19880 304596
rect 19680 304560 19880 304564
rect 19680 304516 19880 304520
rect 19680 304484 19684 304516
rect 19716 304484 19844 304516
rect 19876 304484 19880 304516
rect 19680 304480 19880 304484
rect 19680 304436 19880 304440
rect 19680 304404 19684 304436
rect 19716 304404 19844 304436
rect 19876 304404 19880 304436
rect 19680 304400 19880 304404
rect 19680 304356 19880 304360
rect 19680 304324 19684 304356
rect 19716 304324 19844 304356
rect 19876 304324 19880 304356
rect 19680 304320 19880 304324
rect 19680 304276 19880 304280
rect 19680 304244 19684 304276
rect 19716 304244 19844 304276
rect 19876 304244 19880 304276
rect 19680 304240 19880 304244
rect 19680 304196 19880 304200
rect 19680 304164 19684 304196
rect 19716 304164 19844 304196
rect 19876 304164 19880 304196
rect 19680 304160 19880 304164
rect 19680 304116 19880 304120
rect 19680 304084 19684 304116
rect 19716 304084 19844 304116
rect 19876 304084 19880 304116
rect 19680 304080 19880 304084
rect 19680 304036 19880 304040
rect 19680 304004 19684 304036
rect 19716 304004 19844 304036
rect 19876 304004 19880 304036
rect 19680 304000 19880 304004
rect 19680 303956 19880 303960
rect 19680 303924 19684 303956
rect 19716 303924 19844 303956
rect 19876 303924 19880 303956
rect 19680 303920 19880 303924
rect 19680 303876 19880 303880
rect 19680 303844 19684 303876
rect 19716 303844 19844 303876
rect 19876 303844 19880 303876
rect 19680 303840 19880 303844
rect 19680 303796 19880 303800
rect 19680 303764 19684 303796
rect 19716 303764 19844 303796
rect 19876 303764 19880 303796
rect 19680 303760 19880 303764
rect 19680 303716 19880 303720
rect 19680 303684 19684 303716
rect 19716 303684 19844 303716
rect 19876 303684 19880 303716
rect 19680 303680 19880 303684
rect 19680 303636 19880 303640
rect 19680 303604 19684 303636
rect 19716 303604 19844 303636
rect 19876 303604 19880 303636
rect 19680 303600 19880 303604
rect 19680 303556 19880 303560
rect 19680 303524 19684 303556
rect 19716 303524 19844 303556
rect 19876 303524 19880 303556
rect 19680 303520 19880 303524
rect 19680 303476 19880 303480
rect 19680 303444 19684 303476
rect 19716 303444 19844 303476
rect 19876 303444 19880 303476
rect 19680 303440 19880 303444
rect 19680 303396 19880 303400
rect 19680 303364 19684 303396
rect 19716 303364 19844 303396
rect 19876 303364 19880 303396
rect 19680 303360 19880 303364
rect 19680 303316 19880 303320
rect 19680 303284 19684 303316
rect 19716 303284 19844 303316
rect 19876 303284 19880 303316
rect 19680 303280 19880 303284
rect 19680 303236 19880 303240
rect 19680 303204 19684 303236
rect 19716 303204 19844 303236
rect 19876 303204 19880 303236
rect 19680 303200 19880 303204
rect 19680 303156 19880 303160
rect 19680 303124 19684 303156
rect 19716 303124 19844 303156
rect 19876 303124 19880 303156
rect 19680 303120 19880 303124
rect 19680 303076 19880 303080
rect 19680 303044 19684 303076
rect 19716 303044 19844 303076
rect 19876 303044 19880 303076
rect 19680 303040 19880 303044
rect 19680 302996 19880 303000
rect 19680 302964 19684 302996
rect 19716 302964 19844 302996
rect 19876 302964 19880 302996
rect 19680 302960 19880 302964
rect 19680 302916 19880 302920
rect 19680 302884 19684 302916
rect 19716 302884 19844 302916
rect 19876 302884 19880 302916
rect 19680 302880 19880 302884
rect 19680 302836 19880 302840
rect 19680 302804 19684 302836
rect 19716 302804 19844 302836
rect 19876 302804 19880 302836
rect 19680 302800 19880 302804
rect 19680 302756 19880 302760
rect 19680 302724 19684 302756
rect 19716 302724 19844 302756
rect 19876 302724 19880 302756
rect 19680 302720 19880 302724
rect 19680 302676 19880 302680
rect 19680 302644 19684 302676
rect 19716 302644 19844 302676
rect 19876 302644 19880 302676
rect 19680 302640 19880 302644
rect 19680 302596 19880 302600
rect 19680 302564 19684 302596
rect 19716 302564 19844 302596
rect 19876 302564 19880 302596
rect 19680 302560 19880 302564
rect 19680 302516 19880 302520
rect 19680 302484 19684 302516
rect 19716 302484 19844 302516
rect 19876 302484 19880 302516
rect 19680 302480 19880 302484
rect 19680 302436 19880 302440
rect 19680 302404 19684 302436
rect 19716 302404 19844 302436
rect 19876 302404 19880 302436
rect 19680 302400 19880 302404
rect 19680 302356 19880 302360
rect 19680 302324 19684 302356
rect 19716 302324 19844 302356
rect 19876 302324 19880 302356
rect 19680 302320 19880 302324
rect 19680 302276 19880 302280
rect 19680 302244 19684 302276
rect 19716 302244 19844 302276
rect 19876 302244 19880 302276
rect 19680 302240 19880 302244
rect 19680 302196 19880 302200
rect 19680 302164 19684 302196
rect 19716 302164 19844 302196
rect 19876 302164 19880 302196
rect 19680 302160 19880 302164
rect 19680 302116 19880 302120
rect 19680 302084 19684 302116
rect 19716 302084 19844 302116
rect 19876 302084 19880 302116
rect 19680 302080 19880 302084
rect 19680 302036 19880 302040
rect 19680 302004 19684 302036
rect 19716 302004 19844 302036
rect 19876 302004 19880 302036
rect 19680 302000 19880 302004
rect 19680 301956 19880 301960
rect 19680 301924 19684 301956
rect 19716 301924 19844 301956
rect 19876 301924 19880 301956
rect 19680 301920 19880 301924
rect 19680 301876 19880 301880
rect 19680 301844 19684 301876
rect 19716 301844 19844 301876
rect 19876 301844 19880 301876
rect 19680 301840 19880 301844
rect 19680 301796 19880 301800
rect 19680 301764 19684 301796
rect 19716 301764 19844 301796
rect 19876 301764 19880 301796
rect 19680 301760 19880 301764
rect 19680 301716 19880 301720
rect 19680 301684 19684 301716
rect 19716 301684 19844 301716
rect 19876 301684 19880 301716
rect 19680 301680 19880 301684
rect 19680 301636 19880 301640
rect 19680 301604 19684 301636
rect 19716 301604 19844 301636
rect 19876 301604 19880 301636
rect 19680 301600 19880 301604
rect 19680 301556 19880 301560
rect 19680 301524 19684 301556
rect 19716 301524 19844 301556
rect 19876 301524 19880 301556
rect 19680 301520 19880 301524
rect 19680 301476 19880 301480
rect 19680 301444 19684 301476
rect 19716 301444 19844 301476
rect 19876 301444 19880 301476
rect 19680 301440 19880 301444
rect 19680 301396 19880 301400
rect 19680 301364 19684 301396
rect 19716 301364 19844 301396
rect 19876 301364 19880 301396
rect 19680 301360 19880 301364
rect 19680 301316 19880 301320
rect 19680 301284 19684 301316
rect 19716 301284 19844 301316
rect 19876 301284 19880 301316
rect 19680 301280 19880 301284
rect 19680 301236 19880 301240
rect 19680 301204 19684 301236
rect 19716 301204 19844 301236
rect 19876 301204 19880 301236
rect 19680 301200 19880 301204
rect 19680 301156 19880 301160
rect 19680 301124 19684 301156
rect 19716 301124 19844 301156
rect 19876 301124 19880 301156
rect 19680 301120 19880 301124
rect 19680 301076 19880 301080
rect 19680 301044 19684 301076
rect 19716 301044 19844 301076
rect 19876 301044 19880 301076
rect 19680 301040 19880 301044
rect 19680 300996 19880 301000
rect 19680 300964 19684 300996
rect 19716 300964 19844 300996
rect 19876 300964 19880 300996
rect 19680 300960 19880 300964
rect 19680 300916 19880 300920
rect 19680 300884 19684 300916
rect 19716 300884 19844 300916
rect 19876 300884 19880 300916
rect 19680 300880 19880 300884
rect 19680 300836 19880 300840
rect 19680 300804 19684 300836
rect 19716 300804 19844 300836
rect 19876 300804 19880 300836
rect 19680 300800 19880 300804
rect 19680 300756 19880 300760
rect 19680 300724 19684 300756
rect 19716 300724 19844 300756
rect 19876 300724 19880 300756
rect 19680 300720 19880 300724
rect 19680 300676 19880 300680
rect 19680 300644 19684 300676
rect 19716 300644 19844 300676
rect 19876 300644 19880 300676
rect 19680 300640 19880 300644
rect 19680 300596 19880 300600
rect 19680 300564 19684 300596
rect 19716 300564 19844 300596
rect 19876 300564 19880 300596
rect 19680 300560 19880 300564
rect 19680 300516 19880 300520
rect 19680 300484 19684 300516
rect 19716 300484 19844 300516
rect 19876 300484 19880 300516
rect 19680 300480 19880 300484
rect 19680 300436 19880 300440
rect 19680 300404 19684 300436
rect 19716 300404 19844 300436
rect 19876 300404 19880 300436
rect 19680 300400 19880 300404
rect 19680 300356 19880 300360
rect 19680 300324 19684 300356
rect 19716 300324 19844 300356
rect 19876 300324 19880 300356
rect 19680 300320 19880 300324
rect 19680 300276 19880 300280
rect 19680 300244 19684 300276
rect 19716 300244 19844 300276
rect 19876 300244 19880 300276
rect 19680 300240 19880 300244
rect 19680 300196 19880 300200
rect 19680 300164 19684 300196
rect 19716 300164 19844 300196
rect 19876 300164 19880 300196
rect 19680 300160 19880 300164
rect 19680 300116 19880 300120
rect 19680 300084 19684 300116
rect 19716 300084 19844 300116
rect 19876 300084 19880 300116
rect 19680 300080 19880 300084
rect 19680 300036 19880 300040
rect 19680 300004 19684 300036
rect 19716 300004 19844 300036
rect 19876 300004 19880 300036
rect 19680 300000 19880 300004
rect 19680 299956 19880 299960
rect 19680 299924 19684 299956
rect 19716 299924 19844 299956
rect 19876 299924 19880 299956
rect 19680 299920 19880 299924
rect 19680 299876 19880 299880
rect 19680 299844 19684 299876
rect 19716 299844 19844 299876
rect 19876 299844 19880 299876
rect 19680 299840 19880 299844
rect 19680 299796 19880 299800
rect 19680 299764 19684 299796
rect 19716 299764 19844 299796
rect 19876 299764 19880 299796
rect 19680 299760 19880 299764
rect 19680 299716 19880 299720
rect 19680 299684 19684 299716
rect 19716 299684 19844 299716
rect 19876 299684 19880 299716
rect 19680 299680 19880 299684
rect 19680 299636 19880 299640
rect 19680 299604 19684 299636
rect 19716 299604 19844 299636
rect 19876 299604 19880 299636
rect 19680 299600 19880 299604
rect 19680 299556 19880 299560
rect 19680 299524 19684 299556
rect 19716 299524 19844 299556
rect 19876 299524 19880 299556
rect 19680 299520 19880 299524
rect 19680 299476 19880 299480
rect 19680 299444 19684 299476
rect 19716 299444 19844 299476
rect 19876 299444 19880 299476
rect 19680 299440 19880 299444
rect 19680 299396 19880 299400
rect 19680 299364 19684 299396
rect 19716 299364 19844 299396
rect 19876 299364 19880 299396
rect 19680 299360 19880 299364
rect 19680 299316 19880 299320
rect 19680 299284 19684 299316
rect 19716 299284 19844 299316
rect 19876 299284 19880 299316
rect 19680 299280 19880 299284
rect 19680 299236 19880 299240
rect 19680 299204 19684 299236
rect 19716 299204 19844 299236
rect 19876 299204 19880 299236
rect 19680 299200 19880 299204
rect 19680 299156 19880 299160
rect 19680 299124 19684 299156
rect 19716 299124 19844 299156
rect 19876 299124 19880 299156
rect 19680 299120 19880 299124
rect 19680 299076 19880 299080
rect 19680 299044 19684 299076
rect 19716 299044 19844 299076
rect 19876 299044 19880 299076
rect 19680 299040 19880 299044
rect 19680 298996 19880 299000
rect 19680 298964 19684 298996
rect 19716 298964 19844 298996
rect 19876 298964 19880 298996
rect 19680 298960 19880 298964
rect 19680 298916 19880 298920
rect 19680 298884 19684 298916
rect 19716 298884 19844 298916
rect 19876 298884 19880 298916
rect 19680 298880 19880 298884
rect 19680 298836 19880 298840
rect 19680 298804 19684 298836
rect 19716 298804 19844 298836
rect 19876 298804 19880 298836
rect 19680 298800 19880 298804
rect 19680 298756 19880 298760
rect 19680 298724 19684 298756
rect 19716 298724 19844 298756
rect 19876 298724 19880 298756
rect 19680 298720 19880 298724
rect 19680 298676 19880 298680
rect 19680 298644 19684 298676
rect 19716 298644 19844 298676
rect 19876 298644 19880 298676
rect 19680 298640 19880 298644
rect 19680 298596 19880 298600
rect 19680 298564 19684 298596
rect 19716 298564 19844 298596
rect 19876 298564 19880 298596
rect 19680 298560 19880 298564
rect 19680 298516 19880 298520
rect 19680 298484 19684 298516
rect 19716 298484 19844 298516
rect 19876 298484 19880 298516
rect 19680 298480 19880 298484
rect 19680 298436 19880 298440
rect 19680 298404 19684 298436
rect 19716 298404 19844 298436
rect 19876 298404 19880 298436
rect 19680 298400 19880 298404
rect 19680 298356 19880 298360
rect 19680 298324 19684 298356
rect 19716 298324 19844 298356
rect 19876 298324 19880 298356
rect 19680 298320 19880 298324
rect 19680 298276 19880 298280
rect 19680 298244 19684 298276
rect 19716 298244 19844 298276
rect 19876 298244 19880 298276
rect 19680 298240 19880 298244
rect 19680 298196 19880 298200
rect 19680 298164 19684 298196
rect 19716 298164 19844 298196
rect 19876 298164 19880 298196
rect 19680 298160 19880 298164
rect 19680 298116 19880 298120
rect 19680 298084 19684 298116
rect 19716 298084 19844 298116
rect 19876 298084 19880 298116
rect 19680 298080 19880 298084
rect 19680 298036 19880 298040
rect 19680 298004 19684 298036
rect 19716 298004 19844 298036
rect 19876 298004 19880 298036
rect 19680 298000 19880 298004
rect 19680 297956 19880 297960
rect 19680 297924 19684 297956
rect 19716 297924 19844 297956
rect 19876 297924 19880 297956
rect 19680 297920 19880 297924
rect 19680 297876 19880 297880
rect 19680 297844 19684 297876
rect 19716 297844 19844 297876
rect 19876 297844 19880 297876
rect 19680 297840 19880 297844
rect 19680 297796 19880 297800
rect 19680 297764 19684 297796
rect 19716 297764 19844 297796
rect 19876 297764 19880 297796
rect 19680 297760 19880 297764
rect 19680 297716 19880 297720
rect 19680 297684 19684 297716
rect 19716 297684 19844 297716
rect 19876 297684 19880 297716
rect 19680 297680 19880 297684
rect 19680 297636 19880 297640
rect 19680 297604 19684 297636
rect 19716 297604 19844 297636
rect 19876 297604 19880 297636
rect 19680 297600 19880 297604
rect 19680 297556 19880 297560
rect 19680 297524 19684 297556
rect 19716 297524 19844 297556
rect 19876 297524 19880 297556
rect 19680 297520 19880 297524
rect 19680 297476 19880 297480
rect 19680 297444 19684 297476
rect 19716 297444 19844 297476
rect 19876 297444 19880 297476
rect 19680 297440 19880 297444
rect 19680 297396 19880 297400
rect 19680 297364 19684 297396
rect 19716 297364 19844 297396
rect 19876 297364 19880 297396
rect 19680 297360 19880 297364
rect 19680 297316 19880 297320
rect 19680 297284 19684 297316
rect 19716 297284 19844 297316
rect 19876 297284 19880 297316
rect 19680 297280 19880 297284
rect 19680 297236 19880 297240
rect 19680 297204 19684 297236
rect 19716 297204 19844 297236
rect 19876 297204 19880 297236
rect 19680 297200 19880 297204
rect 19680 297156 19880 297160
rect 19680 297124 19684 297156
rect 19716 297124 19844 297156
rect 19876 297124 19880 297156
rect 19680 297120 19880 297124
rect 19680 297076 19880 297080
rect 19680 297044 19684 297076
rect 19716 297044 19844 297076
rect 19876 297044 19880 297076
rect 19680 297040 19880 297044
rect 19680 296996 19880 297000
rect 19680 296964 19684 296996
rect 19716 296964 19844 296996
rect 19876 296964 19880 296996
rect 19680 296960 19880 296964
rect 19680 296916 19880 296920
rect 19680 296884 19684 296916
rect 19716 296884 19844 296916
rect 19876 296884 19880 296916
rect 19680 296880 19880 296884
rect 19680 296836 19880 296840
rect 19680 296804 19684 296836
rect 19716 296804 19844 296836
rect 19876 296804 19880 296836
rect 19680 296800 19880 296804
rect 19680 296756 19880 296760
rect 19680 296724 19684 296756
rect 19716 296724 19844 296756
rect 19876 296724 19880 296756
rect 19680 296720 19880 296724
rect 19680 296676 19880 296680
rect 19680 296644 19684 296676
rect 19716 296644 19844 296676
rect 19876 296644 19880 296676
rect 19680 296640 19880 296644
rect 19680 296596 19880 296600
rect 19680 296564 19684 296596
rect 19716 296564 19844 296596
rect 19876 296564 19880 296596
rect 19680 296560 19880 296564
rect 19680 296516 19880 296520
rect 19680 296484 19684 296516
rect 19716 296484 19844 296516
rect 19876 296484 19880 296516
rect 19680 296480 19880 296484
rect 19680 296436 19880 296440
rect 19680 296404 19684 296436
rect 19716 296404 19844 296436
rect 19876 296404 19880 296436
rect 19680 296400 19880 296404
rect 19680 296356 19880 296360
rect 19680 296324 19684 296356
rect 19716 296324 19844 296356
rect 19876 296324 19880 296356
rect 19680 296320 19880 296324
rect 19680 296276 19880 296280
rect 19680 296244 19684 296276
rect 19716 296244 19844 296276
rect 19876 296244 19880 296276
rect 19680 296240 19880 296244
rect 19680 296196 19880 296200
rect 19680 296164 19684 296196
rect 19716 296164 19844 296196
rect 19876 296164 19880 296196
rect 19680 296160 19880 296164
rect 19680 296116 19880 296120
rect 19680 296084 19684 296116
rect 19716 296084 19844 296116
rect 19876 296084 19880 296116
rect 19680 296080 19880 296084
rect 19680 296036 19880 296040
rect 19680 296004 19684 296036
rect 19716 296004 19844 296036
rect 19876 296004 19880 296036
rect 19680 296000 19880 296004
rect 19680 295956 19880 295960
rect 19680 295924 19684 295956
rect 19716 295924 19844 295956
rect 19876 295924 19880 295956
rect 19680 295920 19880 295924
rect 19680 295876 19880 295880
rect 19680 295844 19684 295876
rect 19716 295844 19844 295876
rect 19876 295844 19880 295876
rect 19680 295840 19880 295844
rect 19680 295796 19880 295800
rect 19680 295764 19684 295796
rect 19716 295764 19844 295796
rect 19876 295764 19880 295796
rect 19680 295760 19880 295764
rect 19680 295716 19880 295720
rect 19680 295684 19684 295716
rect 19716 295684 19844 295716
rect 19876 295684 19880 295716
rect 19680 295680 19880 295684
rect 19680 295636 19880 295640
rect 19680 295604 19684 295636
rect 19716 295604 19844 295636
rect 19876 295604 19880 295636
rect 19680 295600 19880 295604
rect 19680 295556 19880 295560
rect 19680 295524 19684 295556
rect 19716 295524 19844 295556
rect 19876 295524 19880 295556
rect 19680 295520 19880 295524
rect 19680 295476 19880 295480
rect 19680 295444 19684 295476
rect 19716 295444 19844 295476
rect 19876 295444 19880 295476
rect 19680 295440 19880 295444
rect 19680 295396 19880 295400
rect 19680 295364 19684 295396
rect 19716 295364 19844 295396
rect 19876 295364 19880 295396
rect 19680 295360 19880 295364
rect 19680 295316 19880 295320
rect 19680 295284 19684 295316
rect 19716 295284 19844 295316
rect 19876 295284 19880 295316
rect 19680 295280 19880 295284
rect 19680 295236 19880 295240
rect 19680 295204 19684 295236
rect 19716 295204 19844 295236
rect 19876 295204 19880 295236
rect 19680 295200 19880 295204
rect 19680 295156 19880 295160
rect 19680 295124 19684 295156
rect 19716 295124 19844 295156
rect 19876 295124 19880 295156
rect 19680 295120 19880 295124
rect 19680 295076 19880 295080
rect 19680 295044 19684 295076
rect 19716 295044 19844 295076
rect 19876 295044 19880 295076
rect 19680 295040 19880 295044
rect 19680 294996 19880 295000
rect 19680 294964 19684 294996
rect 19716 294964 19844 294996
rect 19876 294964 19880 294996
rect 19680 294960 19880 294964
rect 19680 294916 19880 294920
rect 19680 294884 19684 294916
rect 19716 294884 19844 294916
rect 19876 294884 19880 294916
rect 19680 294880 19880 294884
rect 19680 294836 19880 294840
rect 19680 294804 19684 294836
rect 19716 294804 19844 294836
rect 19876 294804 19880 294836
rect 19680 294800 19880 294804
rect 19680 294756 19880 294760
rect 19680 294724 19684 294756
rect 19716 294724 19844 294756
rect 19876 294724 19880 294756
rect 19680 294720 19880 294724
rect 19680 294676 19880 294680
rect 19680 294644 19684 294676
rect 19716 294644 19844 294676
rect 19876 294644 19880 294676
rect 19680 294640 19880 294644
rect 19680 294596 19880 294600
rect 19680 294564 19684 294596
rect 19716 294564 19844 294596
rect 19876 294564 19880 294596
rect 19680 294560 19880 294564
rect 19680 294516 19880 294520
rect 19680 294484 19684 294516
rect 19716 294484 19844 294516
rect 19876 294484 19880 294516
rect 19680 294480 19880 294484
rect 19680 294436 19880 294440
rect 19680 294404 19684 294436
rect 19716 294404 19844 294436
rect 19876 294404 19880 294436
rect 19680 294400 19880 294404
rect 19680 294356 19880 294360
rect 19680 294324 19684 294356
rect 19716 294324 19844 294356
rect 19876 294324 19880 294356
rect 19680 294320 19880 294324
rect 19680 294276 19880 294280
rect 19680 294244 19684 294276
rect 19716 294244 19844 294276
rect 19876 294244 19880 294276
rect 19680 294240 19880 294244
rect 19680 294196 19880 294200
rect 19680 294164 19684 294196
rect 19716 294164 19844 294196
rect 19876 294164 19880 294196
rect 19680 294160 19880 294164
rect 19680 294116 19880 294120
rect 19680 294084 19684 294116
rect 19716 294084 19844 294116
rect 19876 294084 19880 294116
rect 19680 294080 19880 294084
rect 19680 294036 19880 294040
rect 19680 294004 19684 294036
rect 19716 294004 19844 294036
rect 19876 294004 19880 294036
rect 19680 294000 19880 294004
rect 19680 293956 19880 293960
rect 19680 293924 19684 293956
rect 19716 293924 19844 293956
rect 19876 293924 19880 293956
rect 19680 293920 19880 293924
rect 19680 293876 19880 293880
rect 19680 293844 19684 293876
rect 19716 293844 19844 293876
rect 19876 293844 19880 293876
rect 19680 293840 19880 293844
rect 19680 293796 19880 293800
rect 19680 293764 19684 293796
rect 19716 293764 19844 293796
rect 19876 293764 19880 293796
rect 19680 293760 19880 293764
rect 19680 293716 19880 293720
rect 19680 293684 19684 293716
rect 19716 293684 19844 293716
rect 19876 293684 19880 293716
rect 19680 293680 19880 293684
rect 19680 293636 19880 293640
rect 19680 293604 19684 293636
rect 19716 293604 19844 293636
rect 19876 293604 19880 293636
rect 19680 293600 19880 293604
rect 19680 293556 19880 293560
rect 19680 293524 19684 293556
rect 19716 293524 19844 293556
rect 19876 293524 19880 293556
rect 19680 293520 19880 293524
rect 19680 293476 19880 293480
rect 19680 293444 19684 293476
rect 19716 293444 19844 293476
rect 19876 293444 19880 293476
rect 19680 293440 19880 293444
rect 19680 293396 19880 293400
rect 19680 293364 19684 293396
rect 19716 293364 19844 293396
rect 19876 293364 19880 293396
rect 19680 293360 19880 293364
rect 19680 293316 19880 293320
rect 19680 293284 19684 293316
rect 19716 293284 19844 293316
rect 19876 293284 19880 293316
rect 19680 293280 19880 293284
rect 19680 293236 19880 293240
rect 19680 293204 19684 293236
rect 19716 293204 19844 293236
rect 19876 293204 19880 293236
rect 19680 293200 19880 293204
rect 19680 293156 19880 293160
rect 19680 293124 19684 293156
rect 19716 293124 19844 293156
rect 19876 293124 19880 293156
rect 19680 293120 19880 293124
rect 19680 293076 19880 293080
rect 19680 293044 19684 293076
rect 19716 293044 19844 293076
rect 19876 293044 19880 293076
rect 19680 293040 19880 293044
rect 19680 292996 19880 293000
rect 19680 292964 19684 292996
rect 19716 292964 19844 292996
rect 19876 292964 19880 292996
rect 19680 292960 19880 292964
rect 19680 292916 19880 292920
rect 19680 292884 19684 292916
rect 19716 292884 19844 292916
rect 19876 292884 19880 292916
rect 19680 292880 19880 292884
rect 19680 292836 19880 292840
rect 19680 292804 19684 292836
rect 19716 292804 19844 292836
rect 19876 292804 19880 292836
rect 19680 292800 19880 292804
rect 19680 292756 19880 292760
rect 19680 292724 19684 292756
rect 19716 292724 19844 292756
rect 19876 292724 19880 292756
rect 19680 292720 19880 292724
rect 19680 292676 19880 292680
rect 19680 292644 19684 292676
rect 19716 292644 19844 292676
rect 19876 292644 19880 292676
rect 19680 292640 19880 292644
rect 19680 292596 19880 292600
rect 19680 292564 19684 292596
rect 19716 292564 19844 292596
rect 19876 292564 19880 292596
rect 19680 292560 19880 292564
rect 19680 292516 19880 292520
rect 19680 292484 19684 292516
rect 19716 292484 19844 292516
rect 19876 292484 19880 292516
rect 19680 292480 19880 292484
rect 19680 292436 19880 292440
rect 19680 292404 19684 292436
rect 19716 292404 19844 292436
rect 19876 292404 19880 292436
rect 19680 292400 19880 292404
rect 19680 292356 19880 292360
rect 19680 292324 19684 292356
rect 19716 292324 19844 292356
rect 19876 292324 19880 292356
rect 19680 292320 19880 292324
rect 19680 292276 19880 292280
rect 19680 292244 19684 292276
rect 19716 292244 19844 292276
rect 19876 292244 19880 292276
rect 19680 292240 19880 292244
rect 19680 292196 19880 292200
rect 19680 292164 19684 292196
rect 19716 292164 19844 292196
rect 19876 292164 19880 292196
rect 19680 292160 19880 292164
rect 19680 292116 19880 292120
rect 19680 292084 19684 292116
rect 19716 292084 19844 292116
rect 19876 292084 19880 292116
rect 19680 292080 19880 292084
rect 19680 292036 19880 292040
rect 19680 292004 19684 292036
rect 19716 292004 19844 292036
rect 19876 292004 19880 292036
rect 19680 292000 19880 292004
rect 19680 291956 19880 291960
rect 19680 291924 19684 291956
rect 19716 291924 19844 291956
rect 19876 291924 19880 291956
rect 19680 291920 19880 291924
rect 19680 291876 19880 291880
rect 19680 291844 19684 291876
rect 19716 291844 19844 291876
rect 19876 291844 19880 291876
rect 19680 291840 19880 291844
rect 19680 291796 19880 291800
rect 19680 291764 19684 291796
rect 19716 291764 19844 291796
rect 19876 291764 19880 291796
rect 19680 291760 19880 291764
rect 19680 291716 19880 291720
rect 19680 291684 19684 291716
rect 19716 291684 19844 291716
rect 19876 291684 19880 291716
rect 19680 291680 19880 291684
rect 19680 291636 19880 291640
rect 19680 291604 19684 291636
rect 19716 291604 19844 291636
rect 19876 291604 19880 291636
rect 19680 291600 19880 291604
rect 19680 291556 19880 291560
rect 19680 291524 19684 291556
rect 19716 291524 19844 291556
rect 19876 291524 19880 291556
rect 19680 291520 19880 291524
rect 19680 291476 19880 291480
rect 19680 291444 19684 291476
rect 19716 291444 19844 291476
rect 19876 291444 19880 291476
rect 19680 291440 19880 291444
rect 19680 291396 19880 291400
rect 19680 291364 19684 291396
rect 19716 291364 19844 291396
rect 19876 291364 19880 291396
rect 19680 291360 19880 291364
rect 19680 291316 19880 291320
rect 19680 291284 19684 291316
rect 19716 291284 19844 291316
rect 19876 291284 19880 291316
rect 19680 291280 19880 291284
rect 19680 291236 19880 291240
rect 19680 291204 19684 291236
rect 19716 291204 19844 291236
rect 19876 291204 19880 291236
rect 19680 291200 19880 291204
rect 19680 291156 19880 291160
rect 19680 291124 19684 291156
rect 19716 291124 19844 291156
rect 19876 291124 19880 291156
rect 19680 291120 19880 291124
rect 19680 291076 19880 291080
rect 19680 291044 19684 291076
rect 19716 291044 19844 291076
rect 19876 291044 19880 291076
rect 19680 291040 19880 291044
rect 19680 290996 19880 291000
rect 19680 290964 19684 290996
rect 19716 290964 19844 290996
rect 19876 290964 19880 290996
rect 19680 290960 19880 290964
rect 19680 290916 19880 290920
rect 19680 290884 19684 290916
rect 19716 290884 19844 290916
rect 19876 290884 19880 290916
rect 19680 290880 19880 290884
rect 19680 290836 19880 290840
rect 19680 290804 19684 290836
rect 19716 290804 19844 290836
rect 19876 290804 19880 290836
rect 19680 290800 19880 290804
rect 19680 290756 19880 290760
rect 19680 290724 19684 290756
rect 19716 290724 19844 290756
rect 19876 290724 19880 290756
rect 19680 290720 19880 290724
rect 19680 290676 19880 290680
rect 19680 290644 19684 290676
rect 19716 290644 19844 290676
rect 19876 290644 19880 290676
rect 19680 290640 19880 290644
rect 19680 290596 19880 290600
rect 19680 290564 19684 290596
rect 19716 290564 19844 290596
rect 19876 290564 19880 290596
rect 19680 290560 19880 290564
rect 19680 290516 19880 290520
rect 19680 290484 19684 290516
rect 19716 290484 19844 290516
rect 19876 290484 19880 290516
rect 19680 290480 19880 290484
rect 19680 290436 19880 290440
rect 19680 290404 19684 290436
rect 19716 290404 19844 290436
rect 19876 290404 19880 290436
rect 19680 290400 19880 290404
rect 19680 290356 19880 290360
rect 19680 290324 19684 290356
rect 19716 290324 19844 290356
rect 19876 290324 19880 290356
rect 19680 290320 19880 290324
rect 19680 290276 19880 290280
rect 19680 290244 19684 290276
rect 19716 290244 19844 290276
rect 19876 290244 19880 290276
rect 19680 290240 19880 290244
rect 19680 290196 19880 290200
rect 19680 290164 19684 290196
rect 19716 290164 19844 290196
rect 19876 290164 19880 290196
rect 19680 290160 19880 290164
rect 19680 290116 19880 290120
rect 19680 290084 19684 290116
rect 19716 290084 19844 290116
rect 19876 290084 19880 290116
rect 19680 290080 19880 290084
rect 19680 290036 19880 290040
rect 19680 290004 19684 290036
rect 19716 290004 19844 290036
rect 19876 290004 19880 290036
rect 19680 290000 19880 290004
rect 19680 289956 19880 289960
rect 19680 289924 19684 289956
rect 19716 289924 19844 289956
rect 19876 289924 19880 289956
rect 19680 289920 19880 289924
rect 19680 289876 19880 289880
rect 19680 289844 19684 289876
rect 19716 289844 19844 289876
rect 19876 289844 19880 289876
rect 19680 289840 19880 289844
rect 19680 289796 19880 289800
rect 19680 289764 19684 289796
rect 19716 289764 19844 289796
rect 19876 289764 19880 289796
rect 19680 289760 19880 289764
rect 19680 289716 19880 289720
rect 19680 289684 19684 289716
rect 19716 289684 19844 289716
rect 19876 289684 19880 289716
rect 19680 289680 19880 289684
rect 19680 289636 19880 289640
rect 19680 289604 19684 289636
rect 19716 289604 19844 289636
rect 19876 289604 19880 289636
rect 19680 289600 19880 289604
rect 19680 289556 19880 289560
rect 19680 289524 19684 289556
rect 19716 289524 19844 289556
rect 19876 289524 19880 289556
rect 19680 289520 19880 289524
rect 19680 289476 19880 289480
rect 19680 289444 19684 289476
rect 19716 289444 19844 289476
rect 19876 289444 19880 289476
rect 19680 289440 19880 289444
rect 19680 289396 19880 289400
rect 19680 289364 19684 289396
rect 19716 289364 19844 289396
rect 19876 289364 19880 289396
rect 19680 289360 19880 289364
rect 19680 289316 19880 289320
rect 19680 289284 19684 289316
rect 19716 289284 19844 289316
rect 19876 289284 19880 289316
rect 19680 289280 19880 289284
rect 19680 289236 19880 289240
rect 19680 289204 19684 289236
rect 19716 289204 19844 289236
rect 19876 289204 19880 289236
rect 19680 289200 19880 289204
rect 19680 289156 19880 289160
rect 19680 289124 19684 289156
rect 19716 289124 19844 289156
rect 19876 289124 19880 289156
rect 19680 289120 19880 289124
rect 19680 289076 19880 289080
rect 19680 289044 19684 289076
rect 19716 289044 19844 289076
rect 19876 289044 19880 289076
rect 19680 289040 19880 289044
rect 19680 288996 19880 289000
rect 19680 288964 19684 288996
rect 19716 288964 19844 288996
rect 19876 288964 19880 288996
rect 19680 288960 19880 288964
rect 19680 288916 19880 288920
rect 19680 288884 19684 288916
rect 19716 288884 19844 288916
rect 19876 288884 19880 288916
rect 19680 288880 19880 288884
rect 19680 288836 19880 288840
rect 19680 288804 19684 288836
rect 19716 288804 19844 288836
rect 19876 288804 19880 288836
rect 19680 288800 19880 288804
rect 19680 288756 19880 288760
rect 19680 288724 19684 288756
rect 19716 288724 19844 288756
rect 19876 288724 19880 288756
rect 19680 288720 19880 288724
rect 19680 288676 19880 288680
rect 19680 288644 19684 288676
rect 19716 288644 19844 288676
rect 19876 288644 19880 288676
rect 19680 288640 19880 288644
rect 19680 288596 19880 288600
rect 19680 288564 19684 288596
rect 19716 288564 19844 288596
rect 19876 288564 19880 288596
rect 19680 288560 19880 288564
rect 19680 288516 19880 288520
rect 19680 288484 19684 288516
rect 19716 288484 19844 288516
rect 19876 288484 19880 288516
rect 19680 288480 19880 288484
rect 19680 288436 19880 288440
rect 19680 288404 19684 288436
rect 19716 288404 19844 288436
rect 19876 288404 19880 288436
rect 19680 288400 19880 288404
rect 19680 288356 19880 288360
rect 19680 288324 19684 288356
rect 19716 288324 19844 288356
rect 19876 288324 19880 288356
rect 19680 288320 19880 288324
rect 19680 288276 19880 288280
rect 19680 288244 19684 288276
rect 19716 288244 19844 288276
rect 19876 288244 19880 288276
rect 19680 288240 19880 288244
rect 19680 288196 19880 288200
rect 19680 288164 19684 288196
rect 19716 288164 19844 288196
rect 19876 288164 19880 288196
rect 19680 288160 19880 288164
rect 19680 288116 19880 288120
rect 19680 288084 19684 288116
rect 19716 288084 19844 288116
rect 19876 288084 19880 288116
rect 19680 288080 19880 288084
rect 19680 288036 19880 288040
rect 19680 288004 19684 288036
rect 19716 288004 19844 288036
rect 19876 288004 19880 288036
rect 19680 288000 19880 288004
rect 19680 287956 19880 287960
rect 19680 287924 19684 287956
rect 19716 287924 19844 287956
rect 19876 287924 19880 287956
rect 19680 287920 19880 287924
rect 19680 287876 19880 287880
rect 19680 287844 19684 287876
rect 19716 287844 19844 287876
rect 19876 287844 19880 287876
rect 19680 287840 19880 287844
rect 19680 287796 19880 287800
rect 19680 287764 19684 287796
rect 19716 287764 19844 287796
rect 19876 287764 19880 287796
rect 19680 287760 19880 287764
rect 19680 287716 19880 287720
rect 19680 287684 19684 287716
rect 19716 287684 19844 287716
rect 19876 287684 19880 287716
rect 19680 287680 19880 287684
rect 19680 287636 19880 287640
rect 19680 287604 19684 287636
rect 19716 287604 19844 287636
rect 19876 287604 19880 287636
rect 19680 287600 19880 287604
rect 19680 287556 19880 287560
rect 19680 287524 19684 287556
rect 19716 287524 19844 287556
rect 19876 287524 19880 287556
rect 19680 287520 19880 287524
rect 19680 287476 19880 287480
rect 19680 287444 19684 287476
rect 19716 287444 19844 287476
rect 19876 287444 19880 287476
rect 19680 287440 19880 287444
rect 19680 287396 19880 287400
rect 19680 287364 19684 287396
rect 19716 287364 19844 287396
rect 19876 287364 19880 287396
rect 19680 287360 19880 287364
rect 19680 287316 19880 287320
rect 19680 287284 19684 287316
rect 19716 287284 19844 287316
rect 19876 287284 19880 287316
rect 19680 287280 19880 287284
rect 19680 287236 19880 287240
rect 19680 287204 19684 287236
rect 19716 287204 19844 287236
rect 19876 287204 19880 287236
rect 19680 287200 19880 287204
rect 19680 287156 19880 287160
rect 19680 287124 19684 287156
rect 19716 287124 19844 287156
rect 19876 287124 19880 287156
rect 19680 287120 19880 287124
rect 19680 287076 19880 287080
rect 19680 287044 19684 287076
rect 19716 287044 19844 287076
rect 19876 287044 19880 287076
rect 19680 287040 19880 287044
rect 19680 286996 19880 287000
rect 19680 286964 19684 286996
rect 19716 286964 19844 286996
rect 19876 286964 19880 286996
rect 19680 286960 19880 286964
rect 19680 286916 19880 286920
rect 19680 286884 19684 286916
rect 19716 286884 19844 286916
rect 19876 286884 19880 286916
rect 19680 286880 19880 286884
rect 19680 286836 19880 286840
rect 19680 286804 19684 286836
rect 19716 286804 19844 286836
rect 19876 286804 19880 286836
rect 19680 286800 19880 286804
rect 19680 286756 19880 286760
rect 19680 286724 19684 286756
rect 19716 286724 19844 286756
rect 19876 286724 19880 286756
rect 19680 286720 19880 286724
rect 19680 286676 19880 286680
rect 19680 286644 19684 286676
rect 19716 286644 19844 286676
rect 19876 286644 19880 286676
rect 19680 286640 19880 286644
rect 19680 286596 19880 286600
rect 19680 286564 19684 286596
rect 19716 286564 19844 286596
rect 19876 286564 19880 286596
rect 19680 286560 19880 286564
rect 19680 286516 19880 286520
rect 19680 286484 19684 286516
rect 19716 286484 19844 286516
rect 19876 286484 19880 286516
rect 19680 286480 19880 286484
rect 19680 286436 19880 286440
rect 19680 286404 19684 286436
rect 19716 286404 19844 286436
rect 19876 286404 19880 286436
rect 19680 286400 19880 286404
rect 19680 286356 19880 286360
rect 19680 286324 19684 286356
rect 19716 286324 19844 286356
rect 19876 286324 19880 286356
rect 19680 286320 19880 286324
rect 19680 286276 19880 286280
rect 19680 286244 19684 286276
rect 19716 286244 19844 286276
rect 19876 286244 19880 286276
rect 19680 286240 19880 286244
rect 19680 286196 19880 286200
rect 19680 286164 19684 286196
rect 19716 286164 19844 286196
rect 19876 286164 19880 286196
rect 19680 286160 19880 286164
rect 19680 286116 19880 286120
rect 19680 286084 19684 286116
rect 19716 286084 19844 286116
rect 19876 286084 19880 286116
rect 19680 286080 19880 286084
rect 19680 286036 19880 286040
rect 19680 286004 19684 286036
rect 19716 286004 19844 286036
rect 19876 286004 19880 286036
rect 19680 286000 19880 286004
rect 19680 285956 19880 285960
rect 19680 285924 19684 285956
rect 19716 285924 19844 285956
rect 19876 285924 19880 285956
rect 19680 285920 19880 285924
rect 19680 285876 19880 285880
rect 19680 285844 19684 285876
rect 19716 285844 19844 285876
rect 19876 285844 19880 285876
rect 19680 285840 19880 285844
rect 19680 285796 19880 285800
rect 19680 285764 19684 285796
rect 19716 285764 19844 285796
rect 19876 285764 19880 285796
rect 19680 285760 19880 285764
rect 19680 285716 19880 285720
rect 19680 285684 19684 285716
rect 19716 285684 19844 285716
rect 19876 285684 19880 285716
rect 19680 285680 19880 285684
rect 19680 285636 19880 285640
rect 19680 285604 19684 285636
rect 19716 285604 19844 285636
rect 19876 285604 19880 285636
rect 19680 285600 19880 285604
rect 19680 285556 19880 285560
rect 19680 285524 19684 285556
rect 19716 285524 19844 285556
rect 19876 285524 19880 285556
rect 19680 285520 19880 285524
rect 19680 285476 19880 285480
rect 19680 285444 19684 285476
rect 19716 285444 19844 285476
rect 19876 285444 19880 285476
rect 19680 285440 19880 285444
rect 19680 285396 19880 285400
rect 19680 285364 19684 285396
rect 19716 285364 19844 285396
rect 19876 285364 19880 285396
rect 19680 285360 19880 285364
rect 19680 285316 19880 285320
rect 19680 285284 19684 285316
rect 19716 285284 19844 285316
rect 19876 285284 19880 285316
rect 19680 285280 19880 285284
rect 19680 285236 19880 285240
rect 19680 285204 19684 285236
rect 19716 285204 19844 285236
rect 19876 285204 19880 285236
rect 19680 285200 19880 285204
rect 19680 285156 19880 285160
rect 19680 285124 19684 285156
rect 19716 285124 19844 285156
rect 19876 285124 19880 285156
rect 19680 285120 19880 285124
rect 19680 285076 19880 285080
rect 19680 285044 19684 285076
rect 19716 285044 19844 285076
rect 19876 285044 19880 285076
rect 19680 285040 19880 285044
rect 19680 284996 19880 285000
rect 19680 284964 19684 284996
rect 19716 284964 19844 284996
rect 19876 284964 19880 284996
rect 19680 284960 19880 284964
rect 19680 284916 19880 284920
rect 19680 284884 19684 284916
rect 19716 284884 19844 284916
rect 19876 284884 19880 284916
rect 19680 284880 19880 284884
rect 19680 284836 19880 284840
rect 19680 284804 19684 284836
rect 19716 284804 19844 284836
rect 19876 284804 19880 284836
rect 19680 284800 19880 284804
rect 19680 284756 19880 284760
rect 19680 284724 19684 284756
rect 19716 284724 19844 284756
rect 19876 284724 19880 284756
rect 19680 284720 19880 284724
rect 19680 284676 19880 284680
rect 19680 284644 19684 284676
rect 19716 284644 19844 284676
rect 19876 284644 19880 284676
rect 19680 284640 19880 284644
rect 19680 284596 19880 284600
rect 19680 284564 19684 284596
rect 19716 284564 19844 284596
rect 19876 284564 19880 284596
rect 19680 284560 19880 284564
rect 19680 284516 19880 284520
rect 19680 284484 19684 284516
rect 19716 284484 19844 284516
rect 19876 284484 19880 284516
rect 19680 284480 19880 284484
rect 19680 284436 19880 284440
rect 19680 284404 19684 284436
rect 19716 284404 19844 284436
rect 19876 284404 19880 284436
rect 19680 284400 19880 284404
rect 19680 284356 19880 284360
rect 19680 284324 19684 284356
rect 19716 284324 19844 284356
rect 19876 284324 19880 284356
rect 19680 284320 19880 284324
rect 19680 284276 19880 284280
rect 19680 284244 19684 284276
rect 19716 284244 19844 284276
rect 19876 284244 19880 284276
rect 19680 284240 19880 284244
rect 19680 284196 19880 284200
rect 19680 284164 19684 284196
rect 19716 284164 19844 284196
rect 19876 284164 19880 284196
rect 19680 284160 19880 284164
rect 19680 284116 19880 284120
rect 19680 284084 19684 284116
rect 19716 284084 19844 284116
rect 19876 284084 19880 284116
rect 19680 284080 19880 284084
rect 19680 284036 19880 284040
rect 19680 284004 19684 284036
rect 19716 284004 19844 284036
rect 19876 284004 19880 284036
rect 19680 284000 19880 284004
rect 19680 283956 19880 283960
rect 19680 283924 19684 283956
rect 19716 283924 19844 283956
rect 19876 283924 19880 283956
rect 19680 283920 19880 283924
rect 19680 283876 19880 283880
rect 19680 283844 19684 283876
rect 19716 283844 19844 283876
rect 19876 283844 19880 283876
rect 19680 283840 19880 283844
rect 19680 283796 19880 283800
rect 19680 283764 19684 283796
rect 19716 283764 19844 283796
rect 19876 283764 19880 283796
rect 19680 283760 19880 283764
rect 19680 283716 19880 283720
rect 19680 283684 19684 283716
rect 19716 283684 19844 283716
rect 19876 283684 19880 283716
rect 19680 283680 19880 283684
rect 19680 283636 19880 283640
rect 19680 283604 19684 283636
rect 19716 283604 19844 283636
rect 19876 283604 19880 283636
rect 19680 283600 19880 283604
rect 19680 283556 19880 283560
rect 19680 283524 19684 283556
rect 19716 283524 19844 283556
rect 19876 283524 19880 283556
rect 19680 283520 19880 283524
rect 19680 283476 19880 283480
rect 19680 283444 19684 283476
rect 19716 283444 19844 283476
rect 19876 283444 19880 283476
rect 19680 283440 19880 283444
rect 19680 283396 19880 283400
rect 19680 283364 19684 283396
rect 19716 283364 19844 283396
rect 19876 283364 19880 283396
rect 19680 283360 19880 283364
rect 19680 283316 19880 283320
rect 19680 283284 19684 283316
rect 19716 283284 19844 283316
rect 19876 283284 19880 283316
rect 19680 283280 19880 283284
rect 19680 283236 19880 283240
rect 19680 283204 19684 283236
rect 19716 283204 19844 283236
rect 19876 283204 19880 283236
rect 19680 283200 19880 283204
rect 19680 283156 19880 283160
rect 19680 283124 19684 283156
rect 19716 283124 19844 283156
rect 19876 283124 19880 283156
rect 19680 283120 19880 283124
rect 19680 283076 19880 283080
rect 19680 283044 19684 283076
rect 19716 283044 19844 283076
rect 19876 283044 19880 283076
rect 19680 283040 19880 283044
rect 19680 282996 19880 283000
rect 19680 282964 19684 282996
rect 19716 282964 19844 282996
rect 19876 282964 19880 282996
rect 19680 282960 19880 282964
rect 19680 282916 19880 282920
rect 19680 282884 19684 282916
rect 19716 282884 19844 282916
rect 19876 282884 19880 282916
rect 19680 282880 19880 282884
rect 19680 282836 19880 282840
rect 19680 282804 19684 282836
rect 19716 282804 19844 282836
rect 19876 282804 19880 282836
rect 19680 282800 19880 282804
rect 19680 282756 19880 282760
rect 19680 282724 19684 282756
rect 19716 282724 19844 282756
rect 19876 282724 19880 282756
rect 19680 282720 19880 282724
rect 19680 282676 19880 282680
rect 19680 282644 19684 282676
rect 19716 282644 19844 282676
rect 19876 282644 19880 282676
rect 19680 282640 19880 282644
rect 19680 282596 19880 282600
rect 19680 282564 19684 282596
rect 19716 282564 19844 282596
rect 19876 282564 19880 282596
rect 19680 282560 19880 282564
rect 19680 282516 19880 282520
rect 19680 282484 19684 282516
rect 19716 282484 19844 282516
rect 19876 282484 19880 282516
rect 19680 282480 19880 282484
rect 19680 282436 19880 282440
rect 19680 282404 19684 282436
rect 19716 282404 19844 282436
rect 19876 282404 19880 282436
rect 19680 282400 19880 282404
rect 19680 282356 19880 282360
rect 19680 282324 19684 282356
rect 19716 282324 19844 282356
rect 19876 282324 19880 282356
rect 19680 282320 19880 282324
rect 19680 282276 19880 282280
rect 19680 282244 19684 282276
rect 19716 282244 19844 282276
rect 19876 282244 19880 282276
rect 19680 282240 19880 282244
rect 19680 282196 19880 282200
rect 19680 282164 19684 282196
rect 19716 282164 19844 282196
rect 19876 282164 19880 282196
rect 19680 282160 19880 282164
rect 19680 282116 19880 282120
rect 19680 282084 19684 282116
rect 19716 282084 19844 282116
rect 19876 282084 19880 282116
rect 19680 282080 19880 282084
rect 19680 282036 19880 282040
rect 19680 282004 19684 282036
rect 19716 282004 19844 282036
rect 19876 282004 19880 282036
rect 19680 282000 19880 282004
rect 19680 281956 19880 281960
rect 19680 281924 19684 281956
rect 19716 281924 19844 281956
rect 19876 281924 19880 281956
rect 19680 281920 19880 281924
rect 19680 281876 19880 281880
rect 19680 281844 19684 281876
rect 19716 281844 19844 281876
rect 19876 281844 19880 281876
rect 19680 281840 19880 281844
rect 19680 281796 19880 281800
rect 19680 281764 19684 281796
rect 19716 281764 19844 281796
rect 19876 281764 19880 281796
rect 19680 281760 19880 281764
rect 19680 281716 19880 281720
rect 19680 281684 19684 281716
rect 19716 281684 19844 281716
rect 19876 281684 19880 281716
rect 19680 281680 19880 281684
rect 19680 281636 19880 281640
rect 19680 281604 19684 281636
rect 19716 281604 19844 281636
rect 19876 281604 19880 281636
rect 19680 281600 19880 281604
rect 19680 281556 19880 281560
rect 19680 281524 19684 281556
rect 19716 281524 19844 281556
rect 19876 281524 19880 281556
rect 19680 281520 19880 281524
rect 19680 281476 19880 281480
rect 19680 281444 19684 281476
rect 19716 281444 19844 281476
rect 19876 281444 19880 281476
rect 19680 281440 19880 281444
rect 19680 281396 19880 281400
rect 19680 281364 19684 281396
rect 19716 281364 19844 281396
rect 19876 281364 19880 281396
rect 19680 281360 19880 281364
rect 19680 281316 19880 281320
rect 19680 281284 19684 281316
rect 19716 281284 19844 281316
rect 19876 281284 19880 281316
rect 19680 281280 19880 281284
rect 19680 281236 19880 281240
rect 19680 281204 19684 281236
rect 19716 281204 19844 281236
rect 19876 281204 19880 281236
rect 19680 281200 19880 281204
rect 19680 281156 19880 281160
rect 19680 281124 19684 281156
rect 19716 281124 19844 281156
rect 19876 281124 19880 281156
rect 19680 281120 19880 281124
rect 19680 281076 19880 281080
rect 19680 281044 19684 281076
rect 19716 281044 19844 281076
rect 19876 281044 19880 281076
rect 19680 281040 19880 281044
rect 19680 280996 19880 281000
rect 19680 280964 19684 280996
rect 19716 280964 19844 280996
rect 19876 280964 19880 280996
rect 19680 280960 19880 280964
rect 19680 280916 19880 280920
rect 19680 280884 19684 280916
rect 19716 280884 19844 280916
rect 19876 280884 19880 280916
rect 19680 280880 19880 280884
rect 19680 280836 19880 280840
rect 19680 280804 19684 280836
rect 19716 280804 19844 280836
rect 19876 280804 19880 280836
rect 19680 280800 19880 280804
rect 19680 280756 19880 280760
rect 19680 280724 19684 280756
rect 19716 280724 19844 280756
rect 19876 280724 19880 280756
rect 19680 280720 19880 280724
rect 19680 280676 19880 280680
rect 19680 280644 19684 280676
rect 19716 280644 19844 280676
rect 19876 280644 19880 280676
rect 19680 280640 19880 280644
rect 19680 280596 19880 280600
rect 19680 280564 19684 280596
rect 19716 280564 19844 280596
rect 19876 280564 19880 280596
rect 19680 280560 19880 280564
rect 19680 280516 19880 280520
rect 19680 280484 19684 280516
rect 19716 280484 19844 280516
rect 19876 280484 19880 280516
rect 19680 280480 19880 280484
rect 19680 280436 19880 280440
rect 19680 280404 19684 280436
rect 19716 280404 19844 280436
rect 19876 280404 19880 280436
rect 19680 280400 19880 280404
rect 19680 280356 19880 280360
rect 19680 280324 19684 280356
rect 19716 280324 19844 280356
rect 19876 280324 19880 280356
rect 19680 280320 19880 280324
rect 19680 280276 19880 280280
rect 19680 280244 19684 280276
rect 19716 280244 19844 280276
rect 19876 280244 19880 280276
rect 19680 280240 19880 280244
rect 19680 280196 19880 280200
rect 19680 280164 19684 280196
rect 19716 280164 19844 280196
rect 19876 280164 19880 280196
rect 19680 280160 19880 280164
rect 19680 280116 19880 280120
rect 19680 280084 19684 280116
rect 19716 280084 19844 280116
rect 19876 280084 19880 280116
rect 19680 280080 19880 280084
rect 19680 280036 19880 280040
rect 19680 280004 19684 280036
rect 19716 280004 19844 280036
rect 19876 280004 19880 280036
rect 19680 280000 19880 280004
rect 19680 279956 19880 279960
rect 19680 279924 19684 279956
rect 19716 279924 19844 279956
rect 19876 279924 19880 279956
rect 19680 279920 19880 279924
rect 19680 279876 19880 279880
rect 19680 279844 19684 279876
rect 19716 279844 19844 279876
rect 19876 279844 19880 279876
rect 19680 279840 19880 279844
rect 19680 279796 19880 279800
rect 19680 279764 19684 279796
rect 19716 279764 19844 279796
rect 19876 279764 19880 279796
rect 19680 279760 19880 279764
rect 19680 279716 19880 279720
rect 19680 279684 19684 279716
rect 19716 279684 19844 279716
rect 19876 279684 19880 279716
rect 19680 279680 19880 279684
rect 19680 279636 19880 279640
rect 19680 279604 19684 279636
rect 19716 279604 19844 279636
rect 19876 279604 19880 279636
rect 19680 279600 19880 279604
rect 19680 279556 19880 279560
rect 19680 279524 19684 279556
rect 19716 279524 19844 279556
rect 19876 279524 19880 279556
rect 19680 279520 19880 279524
rect 17800 279400 17900 279480
rect 19680 279476 19880 279480
rect 19680 279444 19684 279476
rect 19716 279444 19844 279476
rect 19876 279444 19880 279476
rect 19680 279440 19880 279444
rect 2400 279350 17900 279400
rect 19680 279396 19880 279400
rect 19680 279364 19684 279396
rect 19716 279364 19844 279396
rect 19876 279364 19880 279396
rect 19680 279360 19880 279364
rect 2400 279250 2450 279350
rect 2550 279250 17900 279350
rect 19680 279316 19880 279320
rect 19680 279284 19684 279316
rect 19716 279284 19844 279316
rect 19876 279284 19880 279316
rect 19680 279280 19880 279284
rect 2400 279200 17900 279250
rect 19680 279236 19880 279240
rect 19680 279204 19684 279236
rect 19716 279204 19844 279236
rect 19876 279204 19880 279236
rect 19680 279200 19880 279204
rect 19680 279156 19880 279160
rect 19680 279124 19684 279156
rect 19716 279124 19844 279156
rect 19876 279124 19880 279156
rect 19680 279120 19880 279124
rect 19680 279076 19880 279080
rect 19680 279044 19684 279076
rect 19716 279044 19844 279076
rect 19876 279044 19880 279076
rect 19680 279040 19880 279044
rect 19680 278996 19880 279000
rect 19680 278964 19684 278996
rect 19716 278964 19844 278996
rect 19876 278964 19880 278996
rect 19680 278960 19880 278964
rect 19680 278916 19880 278920
rect 19680 278884 19684 278916
rect 19716 278884 19844 278916
rect 19876 278884 19880 278916
rect 19680 278880 19880 278884
rect 19680 278836 19880 278840
rect 19680 278804 19684 278836
rect 19716 278804 19844 278836
rect 19876 278804 19880 278836
rect 19680 278800 19880 278804
rect 19680 278756 19880 278760
rect 19680 278724 19684 278756
rect 19716 278724 19844 278756
rect 19876 278724 19880 278756
rect 19680 278720 19880 278724
rect 17040 278676 17240 278680
rect 17040 278644 17044 278676
rect 17076 278644 17204 278676
rect 17236 278644 17240 278676
rect 17040 278640 17240 278644
rect 17280 278676 17800 278680
rect 17280 278644 17284 278676
rect 17316 278644 17364 278676
rect 17396 278644 17444 278676
rect 17476 278644 17524 278676
rect 17556 278644 17604 278676
rect 17636 278644 17684 278676
rect 17716 278644 17764 278676
rect 17796 278644 17800 278676
rect 17280 278640 17800 278644
rect 19520 278676 19880 278680
rect 19520 278644 19524 278676
rect 19556 278644 19604 278676
rect 19636 278644 19684 278676
rect 19716 278644 19844 278676
rect 19876 278644 19880 278676
rect 19520 278640 19880 278644
rect 17040 278596 17800 278600
rect 17040 278564 17044 278596
rect 17076 278564 17204 278596
rect 17236 278564 17284 278596
rect 17316 278564 17364 278596
rect 17396 278564 17444 278596
rect 17476 278564 17524 278596
rect 17556 278564 17604 278596
rect 17636 278564 17684 278596
rect 17716 278564 17764 278596
rect 17796 278564 17800 278596
rect 17040 278560 17800 278564
rect 19520 278596 19800 278600
rect 19520 278564 19524 278596
rect 19556 278564 19604 278596
rect 19636 278564 19684 278596
rect 19716 278564 19800 278596
rect 19520 278560 19800 278564
rect 17040 278516 17240 278520
rect 17040 278484 17044 278516
rect 17076 278484 17204 278516
rect 17236 278484 17240 278516
rect 17040 278480 17240 278484
rect 17280 278516 17800 278520
rect 17280 278484 17284 278516
rect 17316 278484 17364 278516
rect 17396 278484 17444 278516
rect 17476 278484 17524 278516
rect 17556 278484 17604 278516
rect 17636 278484 17684 278516
rect 17716 278484 17764 278516
rect 17796 278484 17800 278516
rect 17280 278480 17800 278484
rect 19520 278516 19880 278520
rect 19520 278484 19524 278516
rect 19556 278484 19604 278516
rect 19636 278484 19684 278516
rect 19716 278484 19844 278516
rect 19876 278484 19880 278516
rect 19520 278480 19880 278484
rect 17040 278436 17240 278440
rect 17040 278404 17044 278436
rect 17076 278404 17204 278436
rect 17236 278404 17240 278436
rect 17040 278400 17240 278404
rect 17040 278356 17240 278360
rect 17040 278324 17044 278356
rect 17076 278324 17204 278356
rect 17236 278324 17240 278356
rect 17040 278320 17240 278324
rect 17040 278276 17240 278280
rect 17040 278244 17044 278276
rect 17076 278244 17204 278276
rect 17236 278244 17240 278276
rect 17040 278240 17240 278244
rect 17040 278196 17800 278200
rect 17040 278164 17044 278196
rect 17076 278164 17204 278196
rect 17236 278164 17800 278196
rect 17040 278116 17800 278164
rect 17040 278084 17044 278116
rect 17076 278084 17204 278116
rect 17236 278084 17800 278116
rect 17040 278036 17800 278084
rect 17040 278004 17044 278036
rect 17076 278004 17204 278036
rect 17236 278004 17800 278036
rect 17040 278000 17800 278004
rect 17040 277956 17240 277960
rect 17040 277924 17044 277956
rect 17076 277924 17204 277956
rect 17236 277924 17240 277956
rect 17040 277920 17240 277924
rect 17040 277876 17240 277880
rect 17040 277844 17044 277876
rect 17076 277844 17204 277876
rect 17236 277844 17240 277876
rect 17040 277840 17240 277844
rect 28400 275356 28760 275360
rect 28400 275324 28404 275356
rect 28436 275324 28564 275356
rect 28596 275324 28724 275356
rect 28756 275324 28760 275356
rect 28400 275320 28760 275324
rect 28400 275276 28760 275280
rect 28400 275244 28404 275276
rect 28436 275244 28564 275276
rect 28596 275244 28724 275276
rect 28756 275244 28760 275276
rect 28400 275240 28760 275244
rect 1000 275160 28760 275200
rect 1000 275040 1040 275160
rect 1160 275040 28760 275160
rect 1000 275000 28760 275040
<< metal5 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
<< comment >>
rect -50 352000 292050 352050
rect -50 0 0 352000
rect 292000 0 292050 352000
rect -50 -50 292050 0
use ESD  ESD_0 ../lib/ESD/mag
timestamp 1640909703
transform 1 0 18240 0 1 277920
box -440 80 1280 1560
use vref1v8  vref1v8_0 ../lib/vref1v8/mag
timestamp 1640958003
transform -1 0 28040 0 -1 276480
box -720 -1320 11000 1080
use sbcs1v8  sbcs1v8_1 ../lib/sbcs1v8/mag
timestamp 1640892658
transform 1 0 18720 0 1 269280
box -1520 -5880 10040 5640
use sbcs1v8  sbcs1v8_0
timestamp 1640892658
transform 1 0 4320 0 1 269280
box -1520 -5880 10040 5640
<< labels >>
flabel metal3 s 291760 134615 292400 134671 0 FreeSans 560 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -400 190932 240 190988 0 FreeSans 560 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -400 169321 240 169377 0 FreeSans 560 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -400 147710 240 147766 0 FreeSans 560 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -400 126199 240 126255 0 FreeSans 560 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -400 62388 240 62444 0 FreeSans 560 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -400 40777 240 40833 0 FreeSans 560 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -400 19166 240 19222 0 FreeSans 560 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -400 8455 240 8511 0 FreeSans 560 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 291760 156826 292400 156882 0 FreeSans 560 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 291760 179437 292400 179493 0 FreeSans 560 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 291760 202648 292400 202704 0 FreeSans 560 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 291760 224859 292400 224915 0 FreeSans 560 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 291760 247070 292400 247126 0 FreeSans 560 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 291760 291781 292400 291837 0 FreeSans 560 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -400 255765 240 255821 0 FreeSans 560 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -400 234154 240 234210 0 FreeSans 560 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -400 212543 240 212599 0 FreeSans 560 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 291760 135206 292400 135262 0 FreeSans 560 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -400 190341 240 190397 0 FreeSans 560 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -400 168730 240 168786 0 FreeSans 560 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -400 147119 240 147175 0 FreeSans 560 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -400 125608 240 125664 0 FreeSans 560 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -400 61797 240 61853 0 FreeSans 560 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -400 40186 240 40242 0 FreeSans 560 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -400 18575 240 18631 0 FreeSans 560 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -400 7864 240 7920 0 FreeSans 560 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 291760 157417 292400 157473 0 FreeSans 560 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 291760 180028 292400 180084 0 FreeSans 560 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 291760 203239 292400 203295 0 FreeSans 560 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 291760 225450 292400 225506 0 FreeSans 560 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 291760 247661 292400 247717 0 FreeSans 560 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 291760 292372 292400 292428 0 FreeSans 560 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -400 255174 240 255230 0 FreeSans 560 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -400 233563 240 233619 0 FreeSans 560 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -400 211952 240 212008 0 FreeSans 560 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 291150 338992 292400 341492 0 FreeSans 560 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 340121 850 342621 0 FreeSans 560 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 283297 351150 285797 352400 0 FreeSans 960 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 232697 351150 235197 352400 0 FreeSans 960 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 206697 351150 209197 352400 0 FreeSans 960 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 60097 351150 62597 352400 0 FreeSans 960 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 34097 351150 36597 352400 0 FreeSans 960 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 8097 351150 10597 352400 0 FreeSans 960 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 163397 351150 164497 352400 0 FreeSans 960 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 112547 351150 113647 352400 0 FreeSans 960 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 86697 351150 87797 352400 0 FreeSans 960 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 162147 351150 163247 352400 0 FreeSans 960 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 111297 351150 112397 352400 0 FreeSans 960 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 85447 351150 86547 352400 0 FreeSans 960 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 291760 1363 292400 1419 0 FreeSans 560 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 291760 204421 292400 204477 0 FreeSans 560 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 291760 226632 292400 226688 0 FreeSans 560 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 291760 248843 292400 248899 0 FreeSans 560 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 291760 293554 292400 293610 0 FreeSans 560 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -400 253992 240 254048 0 FreeSans 560 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -400 232381 240 232437 0 FreeSans 560 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -400 210770 240 210826 0 FreeSans 560 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -400 189159 240 189215 0 FreeSans 560 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -400 167548 240 167604 0 FreeSans 560 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -400 145937 240 145993 0 FreeSans 560 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 291760 3727 292400 3783 0 FreeSans 560 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -400 124426 240 124482 0 FreeSans 560 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -400 60615 240 60671 0 FreeSans 560 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -400 39004 240 39060 0 FreeSans 560 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -400 17393 240 17449 0 FreeSans 560 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -400 6682 240 6738 0 FreeSans 560 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -400 4318 240 4374 0 FreeSans 560 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -400 1954 240 2010 0 FreeSans 560 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 291760 6091 292400 6147 0 FreeSans 560 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 291760 8455 292400 8511 0 FreeSans 560 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 291760 10819 292400 10875 0 FreeSans 560 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 291760 24048 292400 24104 0 FreeSans 560 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 291760 46377 292400 46433 0 FreeSans 560 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 291760 136388 292400 136444 0 FreeSans 560 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 291760 158599 292400 158655 0 FreeSans 560 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 291760 181210 292400 181266 0 FreeSans 560 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 291760 772 292400 828 0 FreeSans 560 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 291760 203830 292400 203886 0 FreeSans 560 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 291760 226041 292400 226097 0 FreeSans 560 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 291760 248252 292400 248308 0 FreeSans 560 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 291760 292963 292400 293019 0 FreeSans 560 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -400 254583 240 254639 0 FreeSans 560 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -400 232972 240 233028 0 FreeSans 560 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -400 211361 240 211417 0 FreeSans 560 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -400 189750 240 189806 0 FreeSans 560 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -400 168139 240 168195 0 FreeSans 560 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -400 146528 240 146584 0 FreeSans 560 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 291760 3136 292400 3192 0 FreeSans 560 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -400 125017 240 125073 0 FreeSans 560 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -400 61206 240 61262 0 FreeSans 560 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -400 39595 240 39651 0 FreeSans 560 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -400 17984 240 18040 0 FreeSans 560 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -400 7273 240 7329 0 FreeSans 560 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -400 4909 240 4965 0 FreeSans 560 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -400 2545 240 2601 0 FreeSans 560 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 291760 5500 292400 5556 0 FreeSans 560 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 291760 7864 292400 7920 0 FreeSans 560 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 291760 10228 292400 10284 0 FreeSans 560 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 291760 23457 292400 23513 0 FreeSans 560 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 291760 45786 292400 45842 0 FreeSans 560 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 291760 135797 292400 135853 0 FreeSans 560 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 291760 158008 292400 158064 0 FreeSans 560 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 291760 180619 292400 180675 0 FreeSans 560 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 291760 2545 292400 2601 0 FreeSans 560 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 291760 205603 292400 205659 0 FreeSans 560 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 291760 227814 292400 227870 0 FreeSans 560 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 291760 250025 292400 250081 0 FreeSans 560 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 291760 294736 292400 294792 0 FreeSans 560 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -400 252810 240 252866 0 FreeSans 560 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -400 231199 240 231255 0 FreeSans 560 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -400 209588 240 209644 0 FreeSans 560 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -400 187977 240 188033 0 FreeSans 560 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -400 166366 240 166422 0 FreeSans 560 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -400 144755 240 144811 0 FreeSans 560 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 291760 4909 292400 4965 0 FreeSans 560 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -400 123244 240 123300 0 FreeSans 560 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -400 59433 240 59489 0 FreeSans 560 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -400 37822 240 37878 0 FreeSans 560 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -400 16211 240 16267 0 FreeSans 560 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -400 5500 240 5556 0 FreeSans 560 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -400 3136 240 3192 0 FreeSans 560 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -400 772 240 828 0 FreeSans 560 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 291760 7273 292400 7329 0 FreeSans 560 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 291760 9637 292400 9693 0 FreeSans 560 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 291760 12001 292400 12057 0 FreeSans 560 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 291760 25230 292400 25286 0 FreeSans 560 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 291760 47559 292400 47615 0 FreeSans 560 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 291760 137570 292400 137626 0 FreeSans 560 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 291760 159781 292400 159837 0 FreeSans 560 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 291760 182392 292400 182448 0 FreeSans 560 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 291760 1954 292400 2010 0 FreeSans 560 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 291760 205012 292400 205068 0 FreeSans 560 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 291760 227223 292400 227279 0 FreeSans 560 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 291760 249434 292400 249490 0 FreeSans 560 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 291760 294145 292400 294201 0 FreeSans 560 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -400 253401 240 253457 0 FreeSans 560 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -400 231790 240 231846 0 FreeSans 560 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -400 210179 240 210235 0 FreeSans 560 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -400 188568 240 188624 0 FreeSans 560 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -400 166957 240 167013 0 FreeSans 560 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -400 145346 240 145402 0 FreeSans 560 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 291760 4318 292400 4374 0 FreeSans 560 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -400 123835 240 123891 0 FreeSans 560 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -400 60024 240 60080 0 FreeSans 560 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -400 38413 240 38469 0 FreeSans 560 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -400 16802 240 16858 0 FreeSans 560 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -400 6091 240 6147 0 FreeSans 560 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -400 3727 240 3783 0 FreeSans 560 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -400 1363 240 1419 0 FreeSans 560 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 291760 6682 292400 6738 0 FreeSans 560 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 291760 9046 292400 9102 0 FreeSans 560 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 291760 11410 292400 11466 0 FreeSans 560 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 291760 24639 292400 24695 0 FreeSans 560 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 291760 46968 292400 47024 0 FreeSans 560 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 291760 136979 292400 137035 0 FreeSans 560 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 291760 159190 292400 159246 0 FreeSans 560 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 291760 181801 292400 181857 0 FreeSans 560 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 62908 -400 62964 240 0 FreeSans 560 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 240208 -400 240264 240 0 FreeSans 560 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 241981 -400 242037 240 0 FreeSans 560 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 243754 -400 243810 240 0 FreeSans 560 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 245527 -400 245583 240 0 FreeSans 560 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 247300 -400 247356 240 0 FreeSans 560 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 249073 -400 249129 240 0 FreeSans 560 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 250846 -400 250902 240 0 FreeSans 560 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 252619 -400 252675 240 0 FreeSans 560 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 254392 -400 254448 240 0 FreeSans 560 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 256165 -400 256221 240 0 FreeSans 560 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 80638 -400 80694 240 0 FreeSans 560 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 257938 -400 257994 240 0 FreeSans 560 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 259711 -400 259767 240 0 FreeSans 560 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 261484 -400 261540 240 0 FreeSans 560 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 263257 -400 263313 240 0 FreeSans 560 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 265030 -400 265086 240 0 FreeSans 560 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 266803 -400 266859 240 0 FreeSans 560 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 268576 -400 268632 240 0 FreeSans 560 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 270349 -400 270405 240 0 FreeSans 560 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 272122 -400 272178 240 0 FreeSans 560 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 273895 -400 273951 240 0 FreeSans 560 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 82411 -400 82467 240 0 FreeSans 560 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 275668 -400 275724 240 0 FreeSans 560 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 277441 -400 277497 240 0 FreeSans 560 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 279214 -400 279270 240 0 FreeSans 560 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 280987 -400 281043 240 0 FreeSans 560 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 282760 -400 282816 240 0 FreeSans 560 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 284533 -400 284589 240 0 FreeSans 560 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 286306 -400 286362 240 0 FreeSans 560 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 288079 -400 288135 240 0 FreeSans 560 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 84184 -400 84240 240 0 FreeSans 560 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 85957 -400 86013 240 0 FreeSans 560 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 87730 -400 87786 240 0 FreeSans 560 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 89503 -400 89559 240 0 FreeSans 560 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 91276 -400 91332 240 0 FreeSans 560 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 93049 -400 93105 240 0 FreeSans 560 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 94822 -400 94878 240 0 FreeSans 560 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 96595 -400 96651 240 0 FreeSans 560 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 64681 -400 64737 240 0 FreeSans 560 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 98368 -400 98424 240 0 FreeSans 560 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 100141 -400 100197 240 0 FreeSans 560 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 101914 -400 101970 240 0 FreeSans 560 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 103687 -400 103743 240 0 FreeSans 560 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 105460 -400 105516 240 0 FreeSans 560 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 107233 -400 107289 240 0 FreeSans 560 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 109006 -400 109062 240 0 FreeSans 560 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 110779 -400 110835 240 0 FreeSans 560 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 112552 -400 112608 240 0 FreeSans 560 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 114325 -400 114381 240 0 FreeSans 560 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 66454 -400 66510 240 0 FreeSans 560 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 116098 -400 116154 240 0 FreeSans 560 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 117871 -400 117927 240 0 FreeSans 560 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 119644 -400 119700 240 0 FreeSans 560 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 121417 -400 121473 240 0 FreeSans 560 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 123190 -400 123246 240 0 FreeSans 560 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 124963 -400 125019 240 0 FreeSans 560 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 126736 -400 126792 240 0 FreeSans 560 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 128509 -400 128565 240 0 FreeSans 560 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 130282 -400 130338 240 0 FreeSans 560 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 132055 -400 132111 240 0 FreeSans 560 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 68227 -400 68283 240 0 FreeSans 560 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 133828 -400 133884 240 0 FreeSans 560 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 135601 -400 135657 240 0 FreeSans 560 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 137374 -400 137430 240 0 FreeSans 560 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 139147 -400 139203 240 0 FreeSans 560 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 140920 -400 140976 240 0 FreeSans 560 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 142693 -400 142749 240 0 FreeSans 560 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 144466 -400 144522 240 0 FreeSans 560 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 146239 -400 146295 240 0 FreeSans 560 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 148012 -400 148068 240 0 FreeSans 560 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 149785 -400 149841 240 0 FreeSans 560 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 70000 -400 70056 240 0 FreeSans 560 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 151558 -400 151614 240 0 FreeSans 560 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 153331 -400 153387 240 0 FreeSans 560 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 155104 -400 155160 240 0 FreeSans 560 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 156877 -400 156933 240 0 FreeSans 560 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 158650 -400 158706 240 0 FreeSans 560 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 160423 -400 160479 240 0 FreeSans 560 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 162196 -400 162252 240 0 FreeSans 560 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 163969 -400 164025 240 0 FreeSans 560 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 165742 -400 165798 240 0 FreeSans 560 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 167515 -400 167571 240 0 FreeSans 560 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 71773 -400 71829 240 0 FreeSans 560 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 169288 -400 169344 240 0 FreeSans 560 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 171061 -400 171117 240 0 FreeSans 560 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 172834 -400 172890 240 0 FreeSans 560 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 174607 -400 174663 240 0 FreeSans 560 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 176380 -400 176436 240 0 FreeSans 560 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 178153 -400 178209 240 0 FreeSans 560 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 179926 -400 179982 240 0 FreeSans 560 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 181699 -400 181755 240 0 FreeSans 560 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 183472 -400 183528 240 0 FreeSans 560 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 185245 -400 185301 240 0 FreeSans 560 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 73546 -400 73602 240 0 FreeSans 560 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 187018 -400 187074 240 0 FreeSans 560 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 188791 -400 188847 240 0 FreeSans 560 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 190564 -400 190620 240 0 FreeSans 560 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 192337 -400 192393 240 0 FreeSans 560 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 194110 -400 194166 240 0 FreeSans 560 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 195883 -400 195939 240 0 FreeSans 560 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 197656 -400 197712 240 0 FreeSans 560 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 199429 -400 199485 240 0 FreeSans 560 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 201202 -400 201258 240 0 FreeSans 560 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 202975 -400 203031 240 0 FreeSans 560 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 75319 -400 75375 240 0 FreeSans 560 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 204748 -400 204804 240 0 FreeSans 560 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 206521 -400 206577 240 0 FreeSans 560 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 208294 -400 208350 240 0 FreeSans 560 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 210067 -400 210123 240 0 FreeSans 560 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 211840 -400 211896 240 0 FreeSans 560 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 213613 -400 213669 240 0 FreeSans 560 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 215386 -400 215442 240 0 FreeSans 560 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 217159 -400 217215 240 0 FreeSans 560 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 218932 -400 218988 240 0 FreeSans 560 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 220705 -400 220761 240 0 FreeSans 560 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 77092 -400 77148 240 0 FreeSans 560 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 222478 -400 222534 240 0 FreeSans 560 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 224251 -400 224307 240 0 FreeSans 560 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 226024 -400 226080 240 0 FreeSans 560 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 227797 -400 227853 240 0 FreeSans 560 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 229570 -400 229626 240 0 FreeSans 560 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 231343 -400 231399 240 0 FreeSans 560 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 233116 -400 233172 240 0 FreeSans 560 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 234889 -400 234945 240 0 FreeSans 560 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 236662 -400 236718 240 0 FreeSans 560 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 238435 -400 238491 240 0 FreeSans 560 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 78865 -400 78921 240 0 FreeSans 560 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 63499 -400 63555 240 0 FreeSans 560 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 240799 -400 240855 240 0 FreeSans 560 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 242572 -400 242628 240 0 FreeSans 560 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 244345 -400 244401 240 0 FreeSans 560 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 246118 -400 246174 240 0 FreeSans 560 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 247891 -400 247947 240 0 FreeSans 560 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 249664 -400 249720 240 0 FreeSans 560 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 251437 -400 251493 240 0 FreeSans 560 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 253210 -400 253266 240 0 FreeSans 560 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 254983 -400 255039 240 0 FreeSans 560 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 256756 -400 256812 240 0 FreeSans 560 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 81229 -400 81285 240 0 FreeSans 560 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 258529 -400 258585 240 0 FreeSans 560 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 260302 -400 260358 240 0 FreeSans 560 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 262075 -400 262131 240 0 FreeSans 560 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 263848 -400 263904 240 0 FreeSans 560 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 265621 -400 265677 240 0 FreeSans 560 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 267394 -400 267450 240 0 FreeSans 560 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 269167 -400 269223 240 0 FreeSans 560 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 270940 -400 270996 240 0 FreeSans 560 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 272713 -400 272769 240 0 FreeSans 560 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 274486 -400 274542 240 0 FreeSans 560 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 83002 -400 83058 240 0 FreeSans 560 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 276259 -400 276315 240 0 FreeSans 560 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 278032 -400 278088 240 0 FreeSans 560 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 279805 -400 279861 240 0 FreeSans 560 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 281578 -400 281634 240 0 FreeSans 560 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 283351 -400 283407 240 0 FreeSans 560 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 285124 -400 285180 240 0 FreeSans 560 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 286897 -400 286953 240 0 FreeSans 560 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 288670 -400 288726 240 0 FreeSans 560 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 84775 -400 84831 240 0 FreeSans 560 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 86548 -400 86604 240 0 FreeSans 560 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 88321 -400 88377 240 0 FreeSans 560 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 90094 -400 90150 240 0 FreeSans 560 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 91867 -400 91923 240 0 FreeSans 560 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 93640 -400 93696 240 0 FreeSans 560 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 95413 -400 95469 240 0 FreeSans 560 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 97186 -400 97242 240 0 FreeSans 560 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 65272 -400 65328 240 0 FreeSans 560 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 98959 -400 99015 240 0 FreeSans 560 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 100732 -400 100788 240 0 FreeSans 560 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 102505 -400 102561 240 0 FreeSans 560 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 104278 -400 104334 240 0 FreeSans 560 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 106051 -400 106107 240 0 FreeSans 560 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 107824 -400 107880 240 0 FreeSans 560 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 109597 -400 109653 240 0 FreeSans 560 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 111370 -400 111426 240 0 FreeSans 560 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 113143 -400 113199 240 0 FreeSans 560 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 114916 -400 114972 240 0 FreeSans 560 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 67045 -400 67101 240 0 FreeSans 560 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 116689 -400 116745 240 0 FreeSans 560 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 118462 -400 118518 240 0 FreeSans 560 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 120235 -400 120291 240 0 FreeSans 560 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 122008 -400 122064 240 0 FreeSans 560 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 123781 -400 123837 240 0 FreeSans 560 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 125554 -400 125610 240 0 FreeSans 560 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 127327 -400 127383 240 0 FreeSans 560 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 129100 -400 129156 240 0 FreeSans 560 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 130873 -400 130929 240 0 FreeSans 560 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 132646 -400 132702 240 0 FreeSans 560 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 68818 -400 68874 240 0 FreeSans 560 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 134419 -400 134475 240 0 FreeSans 560 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 136192 -400 136248 240 0 FreeSans 560 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 137965 -400 138021 240 0 FreeSans 560 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 139738 -400 139794 240 0 FreeSans 560 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 141511 -400 141567 240 0 FreeSans 560 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 143284 -400 143340 240 0 FreeSans 560 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 145057 -400 145113 240 0 FreeSans 560 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 146830 -400 146886 240 0 FreeSans 560 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 148603 -400 148659 240 0 FreeSans 560 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 150376 -400 150432 240 0 FreeSans 560 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 70591 -400 70647 240 0 FreeSans 560 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 152149 -400 152205 240 0 FreeSans 560 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 153922 -400 153978 240 0 FreeSans 560 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 155695 -400 155751 240 0 FreeSans 560 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 157468 -400 157524 240 0 FreeSans 560 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 159241 -400 159297 240 0 FreeSans 560 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 161014 -400 161070 240 0 FreeSans 560 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 162787 -400 162843 240 0 FreeSans 560 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 164560 -400 164616 240 0 FreeSans 560 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 166333 -400 166389 240 0 FreeSans 560 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 168106 -400 168162 240 0 FreeSans 560 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 72364 -400 72420 240 0 FreeSans 560 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 169879 -400 169935 240 0 FreeSans 560 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 171652 -400 171708 240 0 FreeSans 560 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 173425 -400 173481 240 0 FreeSans 560 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 175198 -400 175254 240 0 FreeSans 560 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 176971 -400 177027 240 0 FreeSans 560 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 178744 -400 178800 240 0 FreeSans 560 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 180517 -400 180573 240 0 FreeSans 560 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 182290 -400 182346 240 0 FreeSans 560 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 184063 -400 184119 240 0 FreeSans 560 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 185836 -400 185892 240 0 FreeSans 560 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 74137 -400 74193 240 0 FreeSans 560 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 187609 -400 187665 240 0 FreeSans 560 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 189382 -400 189438 240 0 FreeSans 560 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 191155 -400 191211 240 0 FreeSans 560 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 192928 -400 192984 240 0 FreeSans 560 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 194701 -400 194757 240 0 FreeSans 560 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 196474 -400 196530 240 0 FreeSans 560 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 198247 -400 198303 240 0 FreeSans 560 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 200020 -400 200076 240 0 FreeSans 560 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 201793 -400 201849 240 0 FreeSans 560 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 203566 -400 203622 240 0 FreeSans 560 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 75910 -400 75966 240 0 FreeSans 560 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 205339 -400 205395 240 0 FreeSans 560 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 207112 -400 207168 240 0 FreeSans 560 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 208885 -400 208941 240 0 FreeSans 560 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 210658 -400 210714 240 0 FreeSans 560 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 212431 -400 212487 240 0 FreeSans 560 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 214204 -400 214260 240 0 FreeSans 560 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 215977 -400 216033 240 0 FreeSans 560 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 217750 -400 217806 240 0 FreeSans 560 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 219523 -400 219579 240 0 FreeSans 560 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 221296 -400 221352 240 0 FreeSans 560 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 77683 -400 77739 240 0 FreeSans 560 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 223069 -400 223125 240 0 FreeSans 560 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 224842 -400 224898 240 0 FreeSans 560 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 226615 -400 226671 240 0 FreeSans 560 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 228388 -400 228444 240 0 FreeSans 560 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 230161 -400 230217 240 0 FreeSans 560 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 231934 -400 231990 240 0 FreeSans 560 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 233707 -400 233763 240 0 FreeSans 560 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 235480 -400 235536 240 0 FreeSans 560 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 237253 -400 237309 240 0 FreeSans 560 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 239026 -400 239082 240 0 FreeSans 560 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 79456 -400 79512 240 0 FreeSans 560 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 64090 -400 64146 240 0 FreeSans 560 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 241390 -400 241446 240 0 FreeSans 560 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 243163 -400 243219 240 0 FreeSans 560 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 244936 -400 244992 240 0 FreeSans 560 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 246709 -400 246765 240 0 FreeSans 560 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 248482 -400 248538 240 0 FreeSans 560 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 250255 -400 250311 240 0 FreeSans 560 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 252028 -400 252084 240 0 FreeSans 560 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 253801 -400 253857 240 0 FreeSans 560 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 255574 -400 255630 240 0 FreeSans 560 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 257347 -400 257403 240 0 FreeSans 560 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 81820 -400 81876 240 0 FreeSans 560 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 259120 -400 259176 240 0 FreeSans 560 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 260893 -400 260949 240 0 FreeSans 560 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 262666 -400 262722 240 0 FreeSans 560 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 264439 -400 264495 240 0 FreeSans 560 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 266212 -400 266268 240 0 FreeSans 560 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 267985 -400 268041 240 0 FreeSans 560 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 269758 -400 269814 240 0 FreeSans 560 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 271531 -400 271587 240 0 FreeSans 560 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 273304 -400 273360 240 0 FreeSans 560 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 275077 -400 275133 240 0 FreeSans 560 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 83593 -400 83649 240 0 FreeSans 560 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 276850 -400 276906 240 0 FreeSans 560 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 278623 -400 278679 240 0 FreeSans 560 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 280396 -400 280452 240 0 FreeSans 560 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 282169 -400 282225 240 0 FreeSans 560 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 283942 -400 283998 240 0 FreeSans 560 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 285715 -400 285771 240 0 FreeSans 560 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 287488 -400 287544 240 0 FreeSans 560 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 289261 -400 289317 240 0 FreeSans 560 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 85366 -400 85422 240 0 FreeSans 560 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 87139 -400 87195 240 0 FreeSans 560 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 88912 -400 88968 240 0 FreeSans 560 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 90685 -400 90741 240 0 FreeSans 560 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 92458 -400 92514 240 0 FreeSans 560 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 94231 -400 94287 240 0 FreeSans 560 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 96004 -400 96060 240 0 FreeSans 560 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 97777 -400 97833 240 0 FreeSans 560 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 65863 -400 65919 240 0 FreeSans 560 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 99550 -400 99606 240 0 FreeSans 560 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 101323 -400 101379 240 0 FreeSans 560 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 103096 -400 103152 240 0 FreeSans 560 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 104869 -400 104925 240 0 FreeSans 560 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 106642 -400 106698 240 0 FreeSans 560 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 108415 -400 108471 240 0 FreeSans 560 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 110188 -400 110244 240 0 FreeSans 560 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 111961 -400 112017 240 0 FreeSans 560 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 113734 -400 113790 240 0 FreeSans 560 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 115507 -400 115563 240 0 FreeSans 560 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 67636 -400 67692 240 0 FreeSans 560 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 117280 -400 117336 240 0 FreeSans 560 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 119053 -400 119109 240 0 FreeSans 560 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 120826 -400 120882 240 0 FreeSans 560 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 122599 -400 122655 240 0 FreeSans 560 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 124372 -400 124428 240 0 FreeSans 560 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 126145 -400 126201 240 0 FreeSans 560 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 127918 -400 127974 240 0 FreeSans 560 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 129691 -400 129747 240 0 FreeSans 560 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 131464 -400 131520 240 0 FreeSans 560 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 133237 -400 133293 240 0 FreeSans 560 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 69409 -400 69465 240 0 FreeSans 560 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 135010 -400 135066 240 0 FreeSans 560 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 136783 -400 136839 240 0 FreeSans 560 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 138556 -400 138612 240 0 FreeSans 560 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 140329 -400 140385 240 0 FreeSans 560 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 142102 -400 142158 240 0 FreeSans 560 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 143875 -400 143931 240 0 FreeSans 560 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 145648 -400 145704 240 0 FreeSans 560 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 147421 -400 147477 240 0 FreeSans 560 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 149194 -400 149250 240 0 FreeSans 560 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 150967 -400 151023 240 0 FreeSans 560 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 71182 -400 71238 240 0 FreeSans 560 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 152740 -400 152796 240 0 FreeSans 560 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 154513 -400 154569 240 0 FreeSans 560 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 156286 -400 156342 240 0 FreeSans 560 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 158059 -400 158115 240 0 FreeSans 560 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 159832 -400 159888 240 0 FreeSans 560 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 161605 -400 161661 240 0 FreeSans 560 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 163378 -400 163434 240 0 FreeSans 560 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 165151 -400 165207 240 0 FreeSans 560 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 166924 -400 166980 240 0 FreeSans 560 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 168697 -400 168753 240 0 FreeSans 560 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 72955 -400 73011 240 0 FreeSans 560 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 170470 -400 170526 240 0 FreeSans 560 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 172243 -400 172299 240 0 FreeSans 560 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 174016 -400 174072 240 0 FreeSans 560 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 175789 -400 175845 240 0 FreeSans 560 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 177562 -400 177618 240 0 FreeSans 560 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 179335 -400 179391 240 0 FreeSans 560 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 181108 -400 181164 240 0 FreeSans 560 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 182881 -400 182937 240 0 FreeSans 560 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 184654 -400 184710 240 0 FreeSans 560 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 186427 -400 186483 240 0 FreeSans 560 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 74728 -400 74784 240 0 FreeSans 560 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 188200 -400 188256 240 0 FreeSans 560 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 189973 -400 190029 240 0 FreeSans 560 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 191746 -400 191802 240 0 FreeSans 560 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 193519 -400 193575 240 0 FreeSans 560 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 195292 -400 195348 240 0 FreeSans 560 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 197065 -400 197121 240 0 FreeSans 560 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 198838 -400 198894 240 0 FreeSans 560 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 200611 -400 200667 240 0 FreeSans 560 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 202384 -400 202440 240 0 FreeSans 560 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 204157 -400 204213 240 0 FreeSans 560 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 76501 -400 76557 240 0 FreeSans 560 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 205930 -400 205986 240 0 FreeSans 560 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 207703 -400 207759 240 0 FreeSans 560 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 209476 -400 209532 240 0 FreeSans 560 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 211249 -400 211305 240 0 FreeSans 560 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 213022 -400 213078 240 0 FreeSans 560 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 214795 -400 214851 240 0 FreeSans 560 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 216568 -400 216624 240 0 FreeSans 560 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 218341 -400 218397 240 0 FreeSans 560 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 220114 -400 220170 240 0 FreeSans 560 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 221887 -400 221943 240 0 FreeSans 560 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 78274 -400 78330 240 0 FreeSans 560 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 223660 -400 223716 240 0 FreeSans 560 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 225433 -400 225489 240 0 FreeSans 560 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 227206 -400 227262 240 0 FreeSans 560 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 228979 -400 229035 240 0 FreeSans 560 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 230752 -400 230808 240 0 FreeSans 560 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 232525 -400 232581 240 0 FreeSans 560 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 234298 -400 234354 240 0 FreeSans 560 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 236071 -400 236127 240 0 FreeSans 560 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 237844 -400 237900 240 0 FreeSans 560 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 239617 -400 239673 240 0 FreeSans 560 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 80047 -400 80103 240 0 FreeSans 560 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 289852 -400 289908 240 0 FreeSans 560 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 290443 -400 290499 240 0 FreeSans 560 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 291034 -400 291090 240 0 FreeSans 560 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 291625 -400 291681 240 0 FreeSans 560 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 291170 319892 292400 322292 0 FreeSans 560 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 291170 314892 292400 317292 0 FreeSans 560 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 321921 830 324321 0 FreeSans 560 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 316921 830 319321 0 FreeSans 560 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 291170 270281 292400 272681 0 FreeSans 560 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 291170 275281 292400 277681 0 FreeSans 560 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 291170 117615 292400 120015 0 FreeSans 560 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 291170 112615 292400 115015 0 FreeSans 560 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 102444 830 104844 0 FreeSans 560 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 107444 830 109844 0 FreeSans 560 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 260297 351170 262697 352400 0 FreeSans 960 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 255297 351170 257697 352400 0 FreeSans 960 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 291170 73415 292400 75815 0 FreeSans 560 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 291170 68415 292400 70815 0 FreeSans 560 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 279721 830 282121 0 FreeSans 560 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 274721 830 277121 0 FreeSans 560 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 291170 95715 292400 98115 0 FreeSans 560 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 291170 90715 292400 93115 0 FreeSans 560 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 86444 830 88844 0 FreeSans 560 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 81444 830 83844 0 FreeSans 560 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 262 -400 318 240 0 FreeSans 560 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 853 -400 909 240 0 FreeSans 560 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 1444 -400 1500 240 0 FreeSans 560 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 3808 -400 3864 240 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 23902 -400 23958 240 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 25675 -400 25731 240 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 27448 -400 27504 240 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 29221 -400 29277 240 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 30994 -400 31050 240 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 32767 -400 32823 240 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 34540 -400 34596 240 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 36313 -400 36369 240 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 38086 -400 38142 240 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 39859 -400 39915 240 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 6172 -400 6228 240 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 41632 -400 41688 240 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 43405 -400 43461 240 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 45178 -400 45234 240 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 46951 -400 47007 240 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 48724 -400 48780 240 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 50497 -400 50553 240 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 52270 -400 52326 240 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 54043 -400 54099 240 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 55816 -400 55872 240 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 57589 -400 57645 240 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 8536 -400 8592 240 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 59362 -400 59418 240 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 61135 -400 61191 240 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 10900 -400 10956 240 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 13264 -400 13320 240 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 15037 -400 15093 240 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 16810 -400 16866 240 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 18583 -400 18639 240 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 20356 -400 20412 240 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 22129 -400 22185 240 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 2035 -400 2091 240 0 FreeSans 560 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 4399 -400 4455 240 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 24493 -400 24549 240 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 26266 -400 26322 240 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 28039 -400 28095 240 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 29812 -400 29868 240 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 31585 -400 31641 240 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 33358 -400 33414 240 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 35131 -400 35187 240 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 36904 -400 36960 240 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 38677 -400 38733 240 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 40450 -400 40506 240 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 6763 -400 6819 240 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 42223 -400 42279 240 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 43996 -400 44052 240 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 45769 -400 45825 240 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 47542 -400 47598 240 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 49315 -400 49371 240 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 51088 -400 51144 240 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 52861 -400 52917 240 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 54634 -400 54690 240 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 56407 -400 56463 240 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 58180 -400 58236 240 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 9127 -400 9183 240 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 59953 -400 60009 240 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 61726 -400 61782 240 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 11491 -400 11547 240 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 13855 -400 13911 240 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 15628 -400 15684 240 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 17401 -400 17457 240 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 19174 -400 19230 240 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 20947 -400 21003 240 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 22720 -400 22776 240 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 4990 -400 5046 240 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 25084 -400 25140 240 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 26857 -400 26913 240 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 28630 -400 28686 240 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 30403 -400 30459 240 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 32176 -400 32232 240 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 33949 -400 34005 240 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 35722 -400 35778 240 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 37495 -400 37551 240 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 39268 -400 39324 240 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 41041 -400 41097 240 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 7354 -400 7410 240 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 42814 -400 42870 240 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 44587 -400 44643 240 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 46360 -400 46416 240 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 48133 -400 48189 240 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 49906 -400 49962 240 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 51679 -400 51735 240 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 53452 -400 53508 240 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 55225 -400 55281 240 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 56998 -400 57054 240 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 58771 -400 58827 240 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 9718 -400 9774 240 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 60544 -400 60600 240 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 62317 -400 62373 240 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 12082 -400 12138 240 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 14446 -400 14502 240 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 16219 -400 16275 240 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 17992 -400 18048 240 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 19765 -400 19821 240 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 21538 -400 21594 240 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 23311 -400 23367 240 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 5581 -400 5637 240 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 7945 -400 8001 240 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 10309 -400 10365 240 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 12673 -400 12729 240 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 2626 -400 2682 240 0 FreeSans 560 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 3217 -400 3273 240 0 FreeSans 560 90 0 0 wbs_we_i
port 677 nsew signal input
rlabel metal3 28640 274920 28680 274960 1 ii
rlabel metal3 28560 274920 28600 274960 1 vi
rlabel metal3 17120 277800 17160 277840 1 vo
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
