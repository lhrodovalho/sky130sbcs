* Self-biased current source testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0

.include "../mag/sbcs5v0.spice"

* supply voltages
vdda	vdda 0 3.3
vssa	vssa 0 0.0

.subckt p1_2 d g s b
xd d g x b sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=1
xs x g s b sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=1
.ends

.subckt p2_2 d g s b
xl d g s b p1_2
xr d g s b p1_2
.ends

.subckt p4_2 d g s b
xl d g s b p2_2
xr d g s b p2_2
.ends

.subckt p1_4 d g s b
xd d g x b p1_2
xs x g s b p1_2
.ends

.subckt p2_4 d g s b
xl d g s b p1_4
xr d g s b p1_4
.ends

.subckt p1_8 d g s b
xd d g x b p1_4
xs x g s b p1_4
.ends

.subckt p1_12 d g s b
xd d g x b p1_4
xs x g s b p1_8
.ends

.subckt p1_16 d g s b
xd d g x b p1_8
xs x g s b p1_8
.ends


* DUT
x0 io vdda vssa x sbcs5v0
vo io y 0.0

xpa  n   x   y    y    p1_16
xpb0 ref ref y    y    sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=8
xpb1 ref ref y    y    p2_4
xna  n   n   vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=16
xnb  ref n   vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=16
.option gmin=1e-13
.control
  dc vdda 10m 5.0 10m
  plot x ref
  plot i(vo)
  
  dc temp -40 125 1
*  plot x ref
*  plot i(vo)
  meas dc r27 find ref at=27
  plot ref/r27
  
.endc

.end
