* Self-biased current source testbench - TT corner

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0

.include "../mag/sbcs5v0.spice"

* supply voltages
vdda	vdda 0 3.3 pulse(10m 3.3 0 1u 10u 10 1)
vssa	vssa 0 0.0

* DUT
x0 io vdda vssa x sbcs5v0
vo io vssa 0.0

.option method=Gear
.option gmin=1e-12
.control
  dc vdda 10m 5.0 10m
  let dc_vdd_io = i(vo)
  plot dc_vdd_io ylimit 0 300n
  wrdata ../data/tt_dc_vdd_io.txt dc_vdd_io
  let dc_vdd_psrr = abs(deriv(i(vo))/i(vo))
  plot dc_vdd_psrr ylog
  wrdata ../data/tt_dc_vdd_psrr.txt dc_vdd_psrr
  
  
  dc temp -40 125 1
  let dc_temp_io = i(vo)
  plot dc_temp_io ylimit 100n 250n
  wrdata ../data/tt_dc_temp_io.txt dc_temp_io
  
  tran 10n 20u
  let tran_io = i(vo)
  plot tran_io ylimit 0 1u
  plot vdda
  wrdata ../data/tt_tran_io.txt tran_io
  wrdata ../data/tt_tran_vdda.txt vdda
  
  reset
  op
  print i(vdda)
  print i(vo)
  
.endc

.end
