* Self-biased current source testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0

.include "../mag/sbcs5v0.spice"

* supply voltages
vdda	vdda 0 3.3
vssa	vssa 0 0.0

* DUT
x0 io vdda vssa x sbcs5v0
vo io vssa 0.0

.option gmin=1e-13
.control
  dc vdda 10m 1.8 10m
  plot i(vo)
  plot abs(deriv(i(vo))/i(vo)) ylog
  
  dc temp -40 125 1
  plot i(vo)
.endc

.end
