* NGSPICE file created from vref1v8.ext - technology: sky130A

.subckt vref1v8 ii vi vo vssa
X0 ii vo a_8080_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X1 a_4240_n2080# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X2 n n a_17360_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X3 a_12240_1320# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X4 a_400_n760# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X5 ii vo a_16080_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X6 a_400_n2080# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X7 a_16080_n760# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X8 a_10960_0# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X9 a_6160_1320# vi a_5520_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X10 a_16080_n2080# vi a_15440_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X11 vssa n a_19920_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X12 a_16720_0# n a_16080_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X13 a_19280_0# n a_18640_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X14 a_16720_n2080# vi a_16080_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X15 a_12240_n2080# vi a_11600_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X16 a_5520_0# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X17 a_8080_0# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X18 a_3600_n760# n a_2960_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X19 a_19920_n760# n a_19280_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X20 ii vo a_13520_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X21 a_1680_n760# n a_1040_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X22 a_18640_1320# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X23 ii vo a_6800_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X24 a_2960_n2080# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X25 n vi a_9360_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X26 a_9360_n760# n a_8720_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X27 ii vo a_19920_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X28 a_1040_0# n a_400_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X29 a_8080_1320# vi a_7440_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X30 ii vo a_2960_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X31 a_12240_0# n a_11600_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X32 a_11600_n760# n a_10960_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X33 vo n a_17360_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X34 ii vo a_17360_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X35 a_17360_n760# n a_16720_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X36 vo n a_12240_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X37 a_5520_n760# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X38 a_400_1320# vi ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X39 a_15440_n2080# vi a_14800_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X40 a_1040_n760# n a_400_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X41 a_6800_0# n a_6160_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X42 a_16080_1320# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X43 a_10960_n2080# vi n ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X44 a_1680_0# n a_1040_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X45 a_9360_0# n a_8720_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X46 a_400_0# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X47 a_18640_0# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X48 a_11600_n2080# vi a_10960_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X49 a_1680_n2080# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X50 n n a_6800_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X51 a_19280_n2080# vi a_18640_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X52 a_13520_n760# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X53 a_19920_n2080# vi a_19280_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X54 a_3600_1320# vi a_2960_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X55 a_2960_n760# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X56 a_19920_1320# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X57 a_19280_n760# n a_18640_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X58 n n a_1680_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X59 vo n a_6800_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X60 a_1680_1320# vi a_1040_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X61 a_11600_0# n a_10960_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X62 a_14160_0# n a_13520_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X63 a_9360_1320# vi a_8720_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X64 ii vo a_5520_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X65 a_2960_0# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X66 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X67 a_10960_n760# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X68 a_19920_0# n a_19280_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X69 a_6800_n2080# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X70 vssa n a_14800_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X71 vo n a_1680_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X72 ii vo a_1680_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X73 a_6800_n760# n a_6160_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X74 a_8720_0# n a_8080_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X75 a_17360_1320# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X76 a_5520_1320# vi a_4880_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X77 vssa n a_4240_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X78 a_1040_1320# vi a_400_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X79 a_18640_n2080# vi a_18000_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X80 a_14160_n2080# vi a_13520_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X81 a_14800_n760# n a_14160_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X82 a_13520_1320# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X83 a_14800_n2080# vi a_14160_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X84 n n a_12240_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X85 ii vo a_4240_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X86 ii vo a_400_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X87 a_4240_n760# n a_3600_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X88 a_4240_0# n a_3600_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X89 a_8720_n760# n a_8080_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X90 a_2960_1320# vi a_2320_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X91 ii vi a_19920_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X92 ii vo a_18640_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X93 a_13520_0# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X94 a_7440_1320# vi a_6800_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X95 a_5520_n2080# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X96 a_16080_0# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X97 vssa n a_9360_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X98 vssa n a_4240_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X99 a_12240_n760# n a_11600_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X100 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X101 a_16720_n760# n a_16080_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X102 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X103 a_12880_n2080# vi a_12240_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X104 a_2320_1320# vi a_1680_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X105 ii vo a_14800_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X106 a_6800_1320# vi a_6160_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X107 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X108 a_6160_n760# n a_5520_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X109 a_13520_n2080# vi a_12880_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X110 a_4880_1320# vi a_4240_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X111 a_14800_0# n a_14160_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X112 a_17360_0# n a_16720_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X113 a_14800_1320# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X114 a_17360_n2080# vi a_16720_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X115 a_14160_n760# n a_13520_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X116 a_3600_0# n a_2960_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X117 a_6160_0# n a_5520_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X118 a_18640_n760# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X119 ii vo a_12240_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X120 vssa n a_9360_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X121 vssa n a_14800_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X122 a_4240_1320# vi a_3600_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X123 a_18000_n2080# vi a_17360_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X124 vssa n a_19920_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X125 a_8720_1320# vi a_8080_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X126 a_8080_n2080# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X127 a_8080_n760# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
.ends

