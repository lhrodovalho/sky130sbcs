magic
tech sky130A
timestamp 1641013539
<< metal1 >>
rect 271860 351815 271900 351820
rect 271860 351785 271865 351815
rect 271895 351785 271900 351815
rect 271860 351780 271900 351785
rect 272020 351815 272060 351820
rect 272020 351785 272025 351815
rect 272055 351785 272060 351815
rect 272020 351780 272060 351785
rect 272100 351815 272140 351820
rect 272100 351785 272105 351815
rect 272135 351785 272140 351815
rect 272100 351780 272140 351785
rect 272180 351815 272220 351820
rect 272180 351785 272185 351815
rect 272215 351785 272220 351815
rect 272180 351780 272220 351785
rect 272260 351815 272300 351820
rect 272260 351785 272265 351815
rect 272295 351785 272300 351815
rect 272260 351780 272300 351785
rect 272340 351815 272380 351820
rect 272340 351785 272345 351815
rect 272375 351785 272380 351815
rect 272340 351780 272380 351785
rect 272420 351815 272460 351820
rect 272420 351785 272425 351815
rect 272455 351785 272460 351815
rect 272420 351780 272460 351785
rect 272500 351815 272540 351820
rect 272500 351785 272505 351815
rect 272535 351785 272540 351815
rect 272500 351780 272540 351785
rect 272580 351815 272620 351820
rect 272580 351785 272585 351815
rect 272615 351785 272620 351815
rect 272580 351780 272620 351785
rect 272660 351815 272700 351820
rect 272660 351785 272665 351815
rect 272695 351785 272700 351815
rect 272660 351780 272700 351785
rect 272740 351815 272780 351820
rect 272740 351785 272745 351815
rect 272775 351785 272780 351815
rect 272740 351780 272780 351785
rect 272820 351815 272860 351820
rect 272820 351785 272825 351815
rect 272855 351785 272860 351815
rect 272820 351780 272860 351785
rect 272900 351815 272940 351820
rect 272900 351785 272905 351815
rect 272935 351785 272940 351815
rect 272900 351780 272940 351785
rect 272980 351815 273020 351820
rect 272980 351785 272985 351815
rect 273015 351785 273020 351815
rect 272980 351780 273020 351785
rect 273060 351815 273100 351820
rect 273060 351785 273065 351815
rect 273095 351785 273100 351815
rect 273060 351780 273100 351785
rect 273140 351815 273180 351820
rect 273140 351785 273145 351815
rect 273175 351785 273180 351815
rect 273140 351780 273180 351785
rect 273220 351815 273260 351820
rect 273220 351785 273225 351815
rect 273255 351785 273260 351815
rect 273220 351780 273260 351785
rect 273300 351815 273340 351820
rect 273300 351785 273305 351815
rect 273335 351785 273340 351815
rect 273300 351780 273340 351785
rect 273380 351815 273420 351820
rect 273380 351785 273385 351815
rect 273415 351785 273420 351815
rect 273380 351780 273420 351785
rect 273460 351815 273500 351820
rect 273460 351785 273465 351815
rect 273495 351785 273500 351815
rect 273460 351780 273500 351785
rect 273540 351815 273580 351820
rect 273540 351785 273545 351815
rect 273575 351785 273580 351815
rect 273540 351780 273580 351785
rect 273620 351815 273660 351820
rect 273620 351785 273625 351815
rect 273655 351785 273660 351815
rect 273620 351780 273660 351785
rect 273700 351815 273740 351820
rect 273700 351785 273705 351815
rect 273735 351785 273740 351815
rect 273700 351780 273740 351785
rect 273780 351815 273820 351820
rect 273780 351785 273785 351815
rect 273815 351785 273820 351815
rect 273780 351780 273820 351785
rect 273860 351815 273900 351820
rect 273860 351785 273865 351815
rect 273895 351785 273900 351815
rect 273860 351780 273900 351785
rect 273940 351815 273980 351820
rect 273940 351785 273945 351815
rect 273975 351785 273980 351815
rect 273940 351780 273980 351785
rect 274020 351815 274060 351820
rect 274020 351785 274025 351815
rect 274055 351785 274060 351815
rect 274020 351780 274060 351785
rect 274100 351815 274140 351820
rect 274100 351785 274105 351815
rect 274135 351785 274140 351815
rect 274100 351780 274140 351785
rect 274180 351815 274220 351820
rect 274180 351785 274185 351815
rect 274215 351785 274220 351815
rect 274180 351780 274220 351785
rect 274260 351815 274300 351820
rect 274260 351785 274265 351815
rect 274295 351785 274300 351815
rect 274260 351780 274300 351785
rect 274340 351815 274380 351820
rect 274340 351785 274345 351815
rect 274375 351785 274380 351815
rect 274340 351780 274380 351785
rect 274420 351815 274460 351820
rect 274420 351785 274425 351815
rect 274455 351785 274460 351815
rect 274420 351780 274460 351785
rect 274500 351815 274540 351820
rect 274500 351785 274505 351815
rect 274535 351785 274540 351815
rect 274500 351780 274540 351785
rect 274580 351815 274620 351820
rect 274580 351785 274585 351815
rect 274615 351785 274620 351815
rect 274580 351780 274620 351785
rect 274660 351815 274700 351820
rect 274660 351785 274665 351815
rect 274695 351785 274700 351815
rect 274660 351780 274700 351785
rect 274740 351815 274780 351820
rect 274740 351785 274745 351815
rect 274775 351785 274780 351815
rect 274740 351780 274780 351785
rect 274820 351815 274860 351820
rect 274820 351785 274825 351815
rect 274855 351785 274860 351815
rect 274820 351780 274860 351785
rect 274900 351815 274940 351820
rect 274900 351785 274905 351815
rect 274935 351785 274940 351815
rect 274900 351780 274940 351785
rect 274980 351815 275020 351820
rect 274980 351785 274985 351815
rect 275015 351785 275020 351815
rect 274980 351780 275020 351785
rect 275060 351815 275100 351820
rect 275060 351785 275065 351815
rect 275095 351785 275100 351815
rect 275060 351780 275100 351785
rect 275140 351815 275180 351820
rect 275140 351785 275145 351815
rect 275175 351785 275180 351815
rect 275140 351780 275180 351785
rect 275220 351815 275260 351820
rect 275220 351785 275225 351815
rect 275255 351785 275260 351815
rect 275220 351780 275260 351785
rect 275300 351815 275340 351820
rect 275300 351785 275305 351815
rect 275335 351785 275340 351815
rect 275300 351780 275340 351785
rect 275380 351815 275420 351820
rect 275380 351785 275385 351815
rect 275415 351785 275420 351815
rect 275380 351780 275420 351785
rect 275460 351815 275500 351820
rect 275460 351785 275465 351815
rect 275495 351785 275500 351815
rect 275460 351780 275500 351785
rect 275540 351815 275580 351820
rect 275540 351785 275545 351815
rect 275575 351785 275580 351815
rect 275540 351780 275580 351785
rect 275620 351815 275660 351820
rect 275620 351785 275625 351815
rect 275655 351785 275660 351815
rect 275620 351780 275660 351785
rect 275700 351815 275740 351820
rect 275700 351785 275705 351815
rect 275735 351785 275740 351815
rect 275700 351780 275740 351785
rect 275780 351815 275820 351820
rect 275780 351785 275785 351815
rect 275815 351785 275820 351815
rect 275780 351780 275820 351785
rect 275860 351815 275900 351820
rect 275860 351785 275865 351815
rect 275895 351785 275900 351815
rect 275860 351780 275900 351785
rect 275940 351815 275980 351820
rect 275940 351785 275945 351815
rect 275975 351785 275980 351815
rect 275940 351780 275980 351785
rect 276020 351815 276060 351820
rect 276020 351785 276025 351815
rect 276055 351785 276060 351815
rect 276020 351780 276060 351785
rect 276100 351815 276140 351820
rect 276100 351785 276105 351815
rect 276135 351785 276140 351815
rect 276100 351780 276140 351785
rect 276180 351815 276220 351820
rect 276180 351785 276185 351815
rect 276215 351785 276220 351815
rect 276180 351780 276220 351785
rect 276260 351815 276300 351820
rect 276260 351785 276265 351815
rect 276295 351785 276300 351815
rect 276260 351780 276300 351785
rect 276340 351815 276380 351820
rect 276340 351785 276345 351815
rect 276375 351785 276380 351815
rect 276340 351780 276380 351785
rect 276420 351815 276460 351820
rect 276420 351785 276425 351815
rect 276455 351785 276460 351815
rect 276420 351780 276460 351785
rect 276500 351815 276540 351820
rect 276500 351785 276505 351815
rect 276535 351785 276540 351815
rect 276500 351780 276540 351785
rect 276580 351815 276620 351820
rect 276580 351785 276585 351815
rect 276615 351785 276620 351815
rect 276580 351780 276620 351785
rect 276660 351815 276700 351820
rect 276660 351785 276665 351815
rect 276695 351785 276700 351815
rect 276660 351780 276700 351785
rect 276740 351815 276780 351820
rect 276740 351785 276745 351815
rect 276775 351785 276780 351815
rect 276740 351780 276780 351785
rect 276820 351815 276860 351820
rect 276820 351785 276825 351815
rect 276855 351785 276860 351815
rect 276820 351780 276860 351785
rect 276900 351815 276940 351820
rect 276900 351785 276905 351815
rect 276935 351785 276940 351815
rect 276900 351780 276940 351785
rect 276980 351815 277020 351820
rect 276980 351785 276985 351815
rect 277015 351785 277020 351815
rect 276980 351780 277020 351785
rect 277060 351815 277100 351820
rect 277060 351785 277065 351815
rect 277095 351785 277100 351815
rect 277060 351780 277100 351785
rect 277140 351815 277180 351820
rect 277140 351785 277145 351815
rect 277175 351785 277180 351815
rect 277140 351780 277180 351785
rect 277220 351815 277260 351820
rect 277220 351785 277225 351815
rect 277255 351785 277260 351815
rect 277220 351780 277260 351785
rect 277300 351815 277340 351820
rect 277300 351785 277305 351815
rect 277335 351785 277340 351815
rect 277300 351780 277340 351785
rect 277380 351815 277420 351820
rect 277380 351785 277385 351815
rect 277415 351785 277420 351815
rect 277380 351780 277420 351785
rect 277460 351815 277500 351820
rect 277460 351785 277465 351815
rect 277495 351785 277500 351815
rect 277460 351780 277500 351785
rect 277540 351815 277580 351820
rect 277540 351785 277545 351815
rect 277575 351785 277580 351815
rect 277540 351780 277580 351785
rect 277620 351815 277660 351820
rect 277620 351785 277625 351815
rect 277655 351785 277660 351815
rect 277620 351780 277660 351785
rect 277700 351815 277740 351820
rect 277700 351785 277705 351815
rect 277735 351785 277740 351815
rect 277700 351780 277740 351785
rect 277780 351815 277820 351820
rect 277780 351785 277785 351815
rect 277815 351785 277820 351815
rect 277780 351780 277820 351785
rect 277860 351815 277900 351820
rect 277860 351785 277865 351815
rect 277895 351785 277900 351815
rect 277860 351780 277900 351785
rect 277940 351815 277980 351820
rect 277940 351785 277945 351815
rect 277975 351785 277980 351815
rect 277940 351780 277980 351785
rect 278020 351815 278060 351820
rect 278020 351785 278025 351815
rect 278055 351785 278060 351815
rect 278020 351780 278060 351785
rect 278100 351815 278140 351820
rect 278100 351785 278105 351815
rect 278135 351785 278140 351815
rect 278100 351780 278140 351785
rect 278180 351815 278220 351820
rect 278180 351785 278185 351815
rect 278215 351785 278220 351815
rect 278180 351780 278220 351785
rect 278260 351815 278300 351820
rect 278260 351785 278265 351815
rect 278295 351785 278300 351815
rect 278260 351780 278300 351785
rect 278340 351815 278380 351820
rect 278340 351785 278345 351815
rect 278375 351785 278380 351815
rect 278340 351780 278380 351785
rect 278420 351815 278460 351820
rect 278420 351785 278425 351815
rect 278455 351785 278460 351815
rect 278420 351780 278460 351785
rect 278500 351815 278540 351820
rect 278500 351785 278505 351815
rect 278535 351785 278540 351815
rect 278500 351780 278540 351785
rect 278580 351815 278620 351820
rect 278580 351785 278585 351815
rect 278615 351785 278620 351815
rect 278580 351780 278620 351785
rect 278660 351815 278700 351820
rect 278660 351785 278665 351815
rect 278695 351785 278700 351815
rect 278660 351780 278700 351785
rect 278740 351815 278780 351820
rect 278740 351785 278745 351815
rect 278775 351785 278780 351815
rect 278740 351780 278780 351785
rect 278820 351815 278860 351820
rect 278820 351785 278825 351815
rect 278855 351785 278860 351815
rect 278820 351780 278860 351785
rect 278900 351815 278940 351820
rect 278900 351785 278905 351815
rect 278935 351785 278940 351815
rect 278900 351780 278940 351785
rect 278980 351815 279020 351820
rect 278980 351785 278985 351815
rect 279015 351785 279020 351815
rect 278980 351780 279020 351785
rect 279060 351815 279100 351820
rect 279060 351785 279065 351815
rect 279095 351785 279100 351815
rect 279060 351780 279100 351785
rect 279140 351815 279180 351820
rect 279140 351785 279145 351815
rect 279175 351785 279180 351815
rect 279140 351780 279180 351785
rect 279220 351815 279260 351820
rect 279220 351785 279225 351815
rect 279255 351785 279260 351815
rect 279220 351780 279260 351785
rect 279300 351815 279340 351820
rect 279300 351785 279305 351815
rect 279335 351785 279340 351815
rect 279300 351780 279340 351785
rect 279380 351815 279420 351820
rect 279380 351785 279385 351815
rect 279415 351785 279420 351815
rect 279380 351780 279420 351785
rect 279460 351815 279500 351820
rect 279460 351785 279465 351815
rect 279495 351785 279500 351815
rect 279460 351780 279500 351785
rect 279540 351815 279580 351820
rect 279540 351785 279545 351815
rect 279575 351785 279580 351815
rect 279540 351780 279580 351785
rect 279620 351815 279660 351820
rect 279620 351785 279625 351815
rect 279655 351785 279660 351815
rect 279620 351780 279660 351785
rect 279700 351815 279740 351820
rect 279700 351785 279705 351815
rect 279735 351785 279740 351815
rect 279700 351780 279740 351785
rect 279780 351815 279820 351820
rect 279780 351785 279785 351815
rect 279815 351785 279820 351815
rect 279780 351780 279820 351785
rect 279860 351815 279900 351820
rect 279860 351785 279865 351815
rect 279895 351785 279900 351815
rect 279860 351780 279900 351785
rect 279940 351815 279980 351820
rect 279940 351785 279945 351815
rect 279975 351785 279980 351815
rect 279940 351780 279980 351785
rect 280020 351815 280060 351820
rect 280020 351785 280025 351815
rect 280055 351785 280060 351815
rect 280020 351780 280060 351785
rect 280100 351815 280140 351820
rect 280100 351785 280105 351815
rect 280135 351785 280140 351815
rect 280100 351780 280140 351785
rect 280180 351815 280220 351820
rect 280180 351785 280185 351815
rect 280215 351785 280220 351815
rect 280180 351780 280220 351785
rect 280260 351815 280300 351820
rect 280260 351785 280265 351815
rect 280295 351785 280300 351815
rect 280260 351780 280300 351785
rect 280340 351815 280380 351820
rect 280340 351785 280345 351815
rect 280375 351785 280380 351815
rect 280340 351780 280380 351785
rect 280420 351815 280460 351820
rect 280420 351785 280425 351815
rect 280455 351785 280460 351815
rect 280420 351780 280460 351785
rect 280500 351815 280540 351820
rect 280500 351785 280505 351815
rect 280535 351785 280540 351815
rect 280500 351780 280540 351785
rect 280580 351815 280620 351820
rect 280580 351785 280585 351815
rect 280615 351785 280620 351815
rect 280580 351780 280620 351785
rect 280660 351815 280700 351820
rect 280660 351785 280665 351815
rect 280695 351785 280700 351815
rect 280660 351780 280700 351785
rect 280740 351815 280780 351820
rect 280740 351785 280745 351815
rect 280775 351785 280780 351815
rect 280740 351780 280780 351785
rect 280820 351815 280860 351820
rect 280820 351785 280825 351815
rect 280855 351785 280860 351815
rect 280820 351780 280860 351785
rect 280900 351815 280940 351820
rect 280900 351785 280905 351815
rect 280935 351785 280940 351815
rect 280900 351780 280940 351785
rect 280980 351815 281020 351820
rect 280980 351785 280985 351815
rect 281015 351785 281020 351815
rect 280980 351780 281020 351785
rect 281060 351815 281100 351820
rect 281060 351785 281065 351815
rect 281095 351785 281100 351815
rect 281060 351780 281100 351785
rect 281140 351815 281180 351820
rect 281140 351785 281145 351815
rect 281175 351785 281180 351815
rect 281140 351780 281180 351785
rect 281220 351815 281260 351820
rect 281220 351785 281225 351815
rect 281255 351785 281260 351815
rect 281220 351780 281260 351785
rect 281300 351815 281340 351820
rect 281300 351785 281305 351815
rect 281335 351785 281340 351815
rect 281300 351780 281340 351785
rect 281380 351815 281420 351820
rect 281380 351785 281385 351815
rect 281415 351785 281420 351815
rect 281380 351780 281420 351785
rect 281460 351815 281500 351820
rect 281460 351785 281465 351815
rect 281495 351785 281500 351815
rect 281460 351780 281500 351785
rect 281540 351815 281580 351820
rect 281540 351785 281545 351815
rect 281575 351785 281580 351815
rect 281540 351780 281580 351785
rect 281620 351815 281660 351820
rect 281620 351785 281625 351815
rect 281655 351785 281660 351815
rect 281620 351780 281660 351785
rect 281700 351815 281740 351820
rect 281700 351785 281705 351815
rect 281735 351785 281740 351815
rect 281700 351780 281740 351785
rect 281780 351815 281820 351820
rect 281780 351785 281785 351815
rect 281815 351785 281820 351815
rect 281780 351780 281820 351785
rect 281860 351815 281900 351820
rect 281860 351785 281865 351815
rect 281895 351785 281900 351815
rect 281860 351780 281900 351785
rect 281940 351815 281980 351820
rect 281940 351785 281945 351815
rect 281975 351785 281980 351815
rect 281940 351780 281980 351785
rect 282020 351815 282060 351820
rect 282020 351785 282025 351815
rect 282055 351785 282060 351815
rect 282020 351780 282060 351785
rect 282100 351815 282140 351820
rect 282100 351785 282105 351815
rect 282135 351785 282140 351815
rect 282100 351780 282140 351785
rect 282180 351815 282220 351820
rect 282180 351785 282185 351815
rect 282215 351785 282220 351815
rect 282180 351780 282220 351785
rect 282260 351815 282300 351820
rect 282260 351785 282265 351815
rect 282295 351785 282300 351815
rect 282260 351780 282300 351785
rect 282340 351815 282380 351820
rect 282340 351785 282345 351815
rect 282375 351785 282380 351815
rect 282340 351780 282380 351785
rect 282420 351815 282460 351820
rect 282420 351785 282425 351815
rect 282455 351785 282460 351815
rect 282420 351780 282460 351785
rect 282500 351815 282540 351820
rect 282500 351785 282505 351815
rect 282535 351785 282540 351815
rect 282500 351780 282540 351785
rect 282580 351815 282620 351820
rect 282580 351785 282585 351815
rect 282615 351785 282620 351815
rect 282580 351780 282620 351785
rect 282660 351815 282700 351820
rect 282660 351785 282665 351815
rect 282695 351785 282700 351815
rect 282660 351780 282700 351785
rect 282740 351815 282780 351820
rect 282740 351785 282745 351815
rect 282775 351785 282780 351815
rect 282740 351780 282780 351785
rect 282820 351815 282860 351820
rect 282820 351785 282825 351815
rect 282855 351785 282860 351815
rect 282820 351780 282860 351785
rect 282900 351815 282940 351820
rect 282900 351785 282905 351815
rect 282935 351785 282940 351815
rect 282900 351780 282940 351785
rect 282980 351815 283020 351820
rect 282980 351785 282985 351815
rect 283015 351785 283020 351815
rect 282980 351780 283020 351785
rect 283060 351815 283100 351820
rect 283060 351785 283065 351815
rect 283095 351785 283100 351815
rect 283060 351780 283100 351785
rect 283140 351815 283180 351820
rect 283140 351785 283145 351815
rect 283175 351785 283180 351815
rect 283140 351780 283180 351785
rect 271860 351655 271900 351660
rect 271860 351625 271865 351655
rect 271895 351625 271900 351655
rect 271860 351620 271900 351625
rect 272020 351655 272060 351660
rect 272020 351625 272025 351655
rect 272055 351625 272060 351655
rect 272020 351620 272060 351625
rect 272100 351655 272140 351660
rect 272100 351625 272105 351655
rect 272135 351625 272140 351655
rect 272100 351620 272140 351625
rect 272180 351655 272220 351660
rect 272180 351625 272185 351655
rect 272215 351625 272220 351655
rect 272180 351620 272220 351625
rect 272260 351655 272300 351660
rect 272260 351625 272265 351655
rect 272295 351625 272300 351655
rect 272260 351620 272300 351625
rect 272340 351655 272380 351660
rect 272340 351625 272345 351655
rect 272375 351625 272380 351655
rect 272340 351620 272380 351625
rect 272420 351655 272460 351660
rect 272420 351625 272425 351655
rect 272455 351625 272460 351655
rect 272420 351620 272460 351625
rect 272500 351655 272540 351660
rect 272500 351625 272505 351655
rect 272535 351625 272540 351655
rect 272500 351620 272540 351625
rect 272580 351655 272620 351660
rect 272580 351625 272585 351655
rect 272615 351625 272620 351655
rect 272580 351620 272620 351625
rect 272660 351655 272700 351660
rect 272660 351625 272665 351655
rect 272695 351625 272700 351655
rect 272660 351620 272700 351625
rect 272740 351655 272780 351660
rect 272740 351625 272745 351655
rect 272775 351625 272780 351655
rect 272740 351620 272780 351625
rect 272820 351655 272860 351660
rect 272820 351625 272825 351655
rect 272855 351625 272860 351655
rect 272820 351620 272860 351625
rect 272900 351655 272940 351660
rect 272900 351625 272905 351655
rect 272935 351625 272940 351655
rect 272900 351620 272940 351625
rect 272980 351655 273020 351660
rect 272980 351625 272985 351655
rect 273015 351625 273020 351655
rect 272980 351620 273020 351625
rect 273060 351655 273100 351660
rect 273060 351625 273065 351655
rect 273095 351625 273100 351655
rect 273060 351620 273100 351625
rect 273140 351655 273180 351660
rect 273140 351625 273145 351655
rect 273175 351625 273180 351655
rect 273140 351620 273180 351625
rect 273220 351655 273260 351660
rect 273220 351625 273225 351655
rect 273255 351625 273260 351655
rect 273220 351620 273260 351625
rect 273300 351655 273340 351660
rect 273300 351625 273305 351655
rect 273335 351625 273340 351655
rect 273300 351620 273340 351625
rect 273380 351655 273420 351660
rect 273380 351625 273385 351655
rect 273415 351625 273420 351655
rect 273380 351620 273420 351625
rect 273460 351655 273500 351660
rect 273460 351625 273465 351655
rect 273495 351625 273500 351655
rect 273460 351620 273500 351625
rect 273540 351655 273580 351660
rect 273540 351625 273545 351655
rect 273575 351625 273580 351655
rect 273540 351620 273580 351625
rect 273620 351655 273660 351660
rect 273620 351625 273625 351655
rect 273655 351625 273660 351655
rect 273620 351620 273660 351625
rect 273700 351655 273740 351660
rect 273700 351625 273705 351655
rect 273735 351625 273740 351655
rect 273700 351620 273740 351625
rect 273780 351655 273820 351660
rect 273780 351625 273785 351655
rect 273815 351625 273820 351655
rect 273780 351620 273820 351625
rect 273860 351655 273900 351660
rect 273860 351625 273865 351655
rect 273895 351625 273900 351655
rect 273860 351620 273900 351625
rect 273940 351655 273980 351660
rect 273940 351625 273945 351655
rect 273975 351625 273980 351655
rect 273940 351620 273980 351625
rect 274020 351655 274060 351660
rect 274020 351625 274025 351655
rect 274055 351625 274060 351655
rect 274020 351620 274060 351625
rect 274100 351655 274140 351660
rect 274100 351625 274105 351655
rect 274135 351625 274140 351655
rect 274100 351620 274140 351625
rect 274180 351655 274220 351660
rect 274180 351625 274185 351655
rect 274215 351625 274220 351655
rect 274180 351620 274220 351625
rect 274260 351655 274300 351660
rect 274260 351625 274265 351655
rect 274295 351625 274300 351655
rect 274260 351620 274300 351625
rect 274340 351655 274380 351660
rect 274340 351625 274345 351655
rect 274375 351625 274380 351655
rect 274340 351620 274380 351625
rect 274420 351655 274460 351660
rect 274420 351625 274425 351655
rect 274455 351625 274460 351655
rect 274420 351620 274460 351625
rect 274500 351655 274540 351660
rect 274500 351625 274505 351655
rect 274535 351625 274540 351655
rect 274500 351620 274540 351625
rect 274580 351655 274620 351660
rect 274580 351625 274585 351655
rect 274615 351625 274620 351655
rect 274580 351620 274620 351625
rect 274660 351655 274700 351660
rect 274660 351625 274665 351655
rect 274695 351625 274700 351655
rect 274660 351620 274700 351625
rect 274740 351655 274780 351660
rect 274740 351625 274745 351655
rect 274775 351625 274780 351655
rect 274740 351620 274780 351625
rect 274820 351655 274860 351660
rect 274820 351625 274825 351655
rect 274855 351625 274860 351655
rect 274820 351620 274860 351625
rect 274900 351655 274940 351660
rect 274900 351625 274905 351655
rect 274935 351625 274940 351655
rect 274900 351620 274940 351625
rect 274980 351655 275020 351660
rect 274980 351625 274985 351655
rect 275015 351625 275020 351655
rect 274980 351620 275020 351625
rect 275060 351655 275100 351660
rect 275060 351625 275065 351655
rect 275095 351625 275100 351655
rect 275060 351620 275100 351625
rect 275140 351655 275180 351660
rect 275140 351625 275145 351655
rect 275175 351625 275180 351655
rect 275140 351620 275180 351625
rect 275220 351655 275260 351660
rect 275220 351625 275225 351655
rect 275255 351625 275260 351655
rect 275220 351620 275260 351625
rect 275300 351655 275340 351660
rect 275300 351625 275305 351655
rect 275335 351625 275340 351655
rect 275300 351620 275340 351625
rect 275380 351655 275420 351660
rect 275380 351625 275385 351655
rect 275415 351625 275420 351655
rect 275380 351620 275420 351625
rect 275460 351655 275500 351660
rect 275460 351625 275465 351655
rect 275495 351625 275500 351655
rect 275460 351620 275500 351625
rect 275540 351655 275580 351660
rect 275540 351625 275545 351655
rect 275575 351625 275580 351655
rect 275540 351620 275580 351625
rect 275620 351655 275660 351660
rect 275620 351625 275625 351655
rect 275655 351625 275660 351655
rect 275620 351620 275660 351625
rect 275700 351655 275740 351660
rect 275700 351625 275705 351655
rect 275735 351625 275740 351655
rect 275700 351620 275740 351625
rect 275780 351655 275820 351660
rect 275780 351625 275785 351655
rect 275815 351625 275820 351655
rect 275780 351620 275820 351625
rect 275860 351655 275900 351660
rect 275860 351625 275865 351655
rect 275895 351625 275900 351655
rect 275860 351620 275900 351625
rect 275940 351655 275980 351660
rect 275940 351625 275945 351655
rect 275975 351625 275980 351655
rect 275940 351620 275980 351625
rect 276020 351655 276060 351660
rect 276020 351625 276025 351655
rect 276055 351625 276060 351655
rect 276020 351620 276060 351625
rect 276100 351655 276140 351660
rect 276100 351625 276105 351655
rect 276135 351625 276140 351655
rect 276100 351620 276140 351625
rect 276180 351655 276220 351660
rect 276180 351625 276185 351655
rect 276215 351625 276220 351655
rect 276180 351620 276220 351625
rect 276260 351655 276300 351660
rect 276260 351625 276265 351655
rect 276295 351625 276300 351655
rect 276260 351620 276300 351625
rect 276340 351655 276380 351660
rect 276340 351625 276345 351655
rect 276375 351625 276380 351655
rect 276340 351620 276380 351625
rect 276420 351655 276460 351660
rect 276420 351625 276425 351655
rect 276455 351625 276460 351655
rect 276420 351620 276460 351625
rect 276500 351655 276540 351660
rect 276500 351625 276505 351655
rect 276535 351625 276540 351655
rect 276500 351620 276540 351625
rect 276580 351655 276620 351660
rect 276580 351625 276585 351655
rect 276615 351625 276620 351655
rect 276580 351620 276620 351625
rect 276660 351655 276700 351660
rect 276660 351625 276665 351655
rect 276695 351625 276700 351655
rect 276660 351620 276700 351625
rect 276740 351655 276780 351660
rect 276740 351625 276745 351655
rect 276775 351625 276780 351655
rect 276740 351620 276780 351625
rect 276820 351655 276860 351660
rect 276820 351625 276825 351655
rect 276855 351625 276860 351655
rect 276820 351620 276860 351625
rect 276900 351655 276940 351660
rect 276900 351625 276905 351655
rect 276935 351625 276940 351655
rect 276900 351620 276940 351625
rect 276980 351655 277020 351660
rect 276980 351625 276985 351655
rect 277015 351625 277020 351655
rect 276980 351620 277020 351625
rect 277060 351655 277100 351660
rect 277060 351625 277065 351655
rect 277095 351625 277100 351655
rect 277060 351620 277100 351625
rect 277140 351655 277180 351660
rect 277140 351625 277145 351655
rect 277175 351625 277180 351655
rect 277140 351620 277180 351625
rect 277220 351655 277260 351660
rect 277220 351625 277225 351655
rect 277255 351625 277260 351655
rect 277220 351620 277260 351625
rect 277300 351655 277340 351660
rect 277300 351625 277305 351655
rect 277335 351625 277340 351655
rect 277300 351620 277340 351625
rect 277380 351655 277420 351660
rect 277380 351625 277385 351655
rect 277415 351625 277420 351655
rect 277380 351620 277420 351625
rect 277460 351655 277500 351660
rect 277460 351625 277465 351655
rect 277495 351625 277500 351655
rect 277460 351620 277500 351625
rect 277540 351655 277580 351660
rect 277540 351625 277545 351655
rect 277575 351625 277580 351655
rect 277540 351620 277580 351625
rect 277620 351655 277660 351660
rect 277620 351625 277625 351655
rect 277655 351625 277660 351655
rect 277620 351620 277660 351625
rect 277700 351655 277740 351660
rect 277700 351625 277705 351655
rect 277735 351625 277740 351655
rect 277700 351620 277740 351625
rect 277780 351655 277820 351660
rect 277780 351625 277785 351655
rect 277815 351625 277820 351655
rect 277780 351620 277820 351625
rect 277860 351655 277900 351660
rect 277860 351625 277865 351655
rect 277895 351625 277900 351655
rect 277860 351620 277900 351625
rect 277940 351655 277980 351660
rect 277940 351625 277945 351655
rect 277975 351625 277980 351655
rect 277940 351620 277980 351625
rect 278020 351655 278060 351660
rect 278020 351625 278025 351655
rect 278055 351625 278060 351655
rect 278020 351620 278060 351625
rect 278100 351655 278140 351660
rect 278100 351625 278105 351655
rect 278135 351625 278140 351655
rect 278100 351620 278140 351625
rect 278180 351655 278220 351660
rect 278180 351625 278185 351655
rect 278215 351625 278220 351655
rect 278180 351620 278220 351625
rect 278260 351655 278300 351660
rect 278260 351625 278265 351655
rect 278295 351625 278300 351655
rect 278260 351620 278300 351625
rect 278340 351655 278380 351660
rect 278340 351625 278345 351655
rect 278375 351625 278380 351655
rect 278340 351620 278380 351625
rect 278420 351655 278460 351660
rect 278420 351625 278425 351655
rect 278455 351625 278460 351655
rect 278420 351620 278460 351625
rect 278500 351655 278540 351660
rect 278500 351625 278505 351655
rect 278535 351625 278540 351655
rect 278500 351620 278540 351625
rect 278580 351655 278620 351660
rect 278580 351625 278585 351655
rect 278615 351625 278620 351655
rect 278580 351620 278620 351625
rect 278660 351655 278700 351660
rect 278660 351625 278665 351655
rect 278695 351625 278700 351655
rect 278660 351620 278700 351625
rect 278740 351655 278780 351660
rect 278740 351625 278745 351655
rect 278775 351625 278780 351655
rect 278740 351620 278780 351625
rect 278820 351655 278860 351660
rect 278820 351625 278825 351655
rect 278855 351625 278860 351655
rect 278820 351620 278860 351625
rect 278900 351655 278940 351660
rect 278900 351625 278905 351655
rect 278935 351625 278940 351655
rect 278900 351620 278940 351625
rect 278980 351655 279020 351660
rect 278980 351625 278985 351655
rect 279015 351625 279020 351655
rect 278980 351620 279020 351625
rect 279060 351655 279100 351660
rect 279060 351625 279065 351655
rect 279095 351625 279100 351655
rect 279060 351620 279100 351625
rect 279140 351655 279180 351660
rect 279140 351625 279145 351655
rect 279175 351625 279180 351655
rect 279140 351620 279180 351625
rect 279220 351655 279260 351660
rect 279220 351625 279225 351655
rect 279255 351625 279260 351655
rect 279220 351620 279260 351625
rect 279300 351655 279340 351660
rect 279300 351625 279305 351655
rect 279335 351625 279340 351655
rect 279300 351620 279340 351625
rect 279380 351655 279420 351660
rect 279380 351625 279385 351655
rect 279415 351625 279420 351655
rect 279380 351620 279420 351625
rect 279460 351655 279500 351660
rect 279460 351625 279465 351655
rect 279495 351625 279500 351655
rect 279460 351620 279500 351625
rect 279540 351655 279580 351660
rect 279540 351625 279545 351655
rect 279575 351625 279580 351655
rect 279540 351620 279580 351625
rect 279620 351655 279660 351660
rect 279620 351625 279625 351655
rect 279655 351625 279660 351655
rect 279620 351620 279660 351625
rect 279700 351655 279740 351660
rect 279700 351625 279705 351655
rect 279735 351625 279740 351655
rect 279700 351620 279740 351625
rect 279780 351655 279820 351660
rect 279780 351625 279785 351655
rect 279815 351625 279820 351655
rect 279780 351620 279820 351625
rect 279860 351655 279900 351660
rect 279860 351625 279865 351655
rect 279895 351625 279900 351655
rect 279860 351620 279900 351625
rect 279940 351655 279980 351660
rect 279940 351625 279945 351655
rect 279975 351625 279980 351655
rect 279940 351620 279980 351625
rect 280020 351655 280060 351660
rect 280020 351625 280025 351655
rect 280055 351625 280060 351655
rect 280020 351620 280060 351625
rect 280100 351655 280140 351660
rect 280100 351625 280105 351655
rect 280135 351625 280140 351655
rect 280100 351620 280140 351625
rect 280180 351655 280220 351660
rect 280180 351625 280185 351655
rect 280215 351625 280220 351655
rect 280180 351620 280220 351625
rect 280260 351655 280300 351660
rect 280260 351625 280265 351655
rect 280295 351625 280300 351655
rect 280260 351620 280300 351625
rect 280340 351655 280380 351660
rect 280340 351625 280345 351655
rect 280375 351625 280380 351655
rect 280340 351620 280380 351625
rect 280420 351655 280460 351660
rect 280420 351625 280425 351655
rect 280455 351625 280460 351655
rect 280420 351620 280460 351625
rect 280500 351655 280540 351660
rect 280500 351625 280505 351655
rect 280535 351625 280540 351655
rect 280500 351620 280540 351625
rect 280580 351655 280620 351660
rect 280580 351625 280585 351655
rect 280615 351625 280620 351655
rect 280580 351620 280620 351625
rect 280660 351655 280700 351660
rect 280660 351625 280665 351655
rect 280695 351625 280700 351655
rect 280660 351620 280700 351625
rect 280740 351655 280780 351660
rect 280740 351625 280745 351655
rect 280775 351625 280780 351655
rect 280740 351620 280780 351625
rect 280820 351655 280860 351660
rect 280820 351625 280825 351655
rect 280855 351625 280860 351655
rect 280820 351620 280860 351625
rect 280900 351655 280940 351660
rect 280900 351625 280905 351655
rect 280935 351625 280940 351655
rect 280900 351620 280940 351625
rect 280980 351655 281020 351660
rect 280980 351625 280985 351655
rect 281015 351625 281020 351655
rect 280980 351620 281020 351625
rect 281060 351655 281100 351660
rect 281060 351625 281065 351655
rect 281095 351625 281100 351655
rect 281060 351620 281100 351625
rect 281140 351655 281180 351660
rect 281140 351625 281145 351655
rect 281175 351625 281180 351655
rect 281140 351620 281180 351625
rect 281220 351655 281260 351660
rect 281220 351625 281225 351655
rect 281255 351625 281260 351655
rect 281220 351620 281260 351625
rect 281300 351655 281340 351660
rect 281300 351625 281305 351655
rect 281335 351625 281340 351655
rect 281300 351620 281340 351625
rect 281380 351655 281420 351660
rect 281380 351625 281385 351655
rect 281415 351625 281420 351655
rect 281380 351620 281420 351625
rect 281460 351655 281500 351660
rect 281460 351625 281465 351655
rect 281495 351625 281500 351655
rect 281460 351620 281500 351625
rect 281540 351655 281580 351660
rect 281540 351625 281545 351655
rect 281575 351625 281580 351655
rect 281540 351620 281580 351625
rect 281620 351655 281660 351660
rect 281620 351625 281625 351655
rect 281655 351625 281660 351655
rect 281620 351620 281660 351625
rect 281700 351655 281740 351660
rect 281700 351625 281705 351655
rect 281735 351625 281740 351655
rect 281700 351620 281740 351625
rect 281780 351655 281820 351660
rect 281780 351625 281785 351655
rect 281815 351625 281820 351655
rect 281780 351620 281820 351625
rect 281860 351655 281900 351660
rect 281860 351625 281865 351655
rect 281895 351625 281900 351655
rect 281860 351620 281900 351625
rect 281940 351655 281980 351660
rect 281940 351625 281945 351655
rect 281975 351625 281980 351655
rect 281940 351620 281980 351625
rect 282020 351655 282060 351660
rect 282020 351625 282025 351655
rect 282055 351625 282060 351655
rect 282020 351620 282060 351625
rect 282100 351655 282140 351660
rect 282100 351625 282105 351655
rect 282135 351625 282140 351655
rect 282100 351620 282140 351625
rect 282180 351655 282220 351660
rect 282180 351625 282185 351655
rect 282215 351625 282220 351655
rect 282180 351620 282220 351625
rect 282260 351655 282300 351660
rect 282260 351625 282265 351655
rect 282295 351625 282300 351655
rect 282260 351620 282300 351625
rect 282340 351655 282380 351660
rect 282340 351625 282345 351655
rect 282375 351625 282380 351655
rect 282340 351620 282380 351625
rect 282420 351655 282460 351660
rect 282420 351625 282425 351655
rect 282455 351625 282460 351655
rect 282420 351620 282460 351625
rect 282500 351655 282540 351660
rect 282500 351625 282505 351655
rect 282535 351625 282540 351655
rect 282500 351620 282540 351625
rect 282580 351655 282620 351660
rect 282580 351625 282585 351655
rect 282615 351625 282620 351655
rect 282580 351620 282620 351625
rect 282660 351655 282700 351660
rect 282660 351625 282665 351655
rect 282695 351625 282700 351655
rect 282660 351620 282700 351625
rect 282740 351655 282780 351660
rect 282740 351625 282745 351655
rect 282775 351625 282780 351655
rect 282740 351620 282780 351625
rect 282820 351655 282860 351660
rect 282820 351625 282825 351655
rect 282855 351625 282860 351655
rect 282820 351620 282860 351625
rect 282900 351655 282940 351660
rect 282900 351625 282905 351655
rect 282935 351625 282940 351655
rect 282900 351620 282940 351625
rect 282980 351655 283020 351660
rect 282980 351625 282985 351655
rect 283015 351625 283020 351655
rect 282980 351620 283020 351625
rect 283060 351655 283100 351660
rect 283060 351625 283065 351655
rect 283095 351625 283100 351655
rect 283060 351620 283100 351625
rect 283140 351655 283180 351660
rect 283140 351625 283145 351655
rect 283175 351625 283180 351655
rect 283140 351620 283180 351625
rect 16720 275475 16760 275480
rect 16720 275445 16725 275475
rect 16755 275445 16760 275475
rect 16720 275440 16760 275445
rect 16880 275475 16920 275480
rect 16880 275445 16885 275475
rect 16915 275445 16920 275475
rect 16880 275440 16920 275445
rect 16960 275475 17000 275480
rect 16960 275445 16965 275475
rect 16995 275445 17000 275475
rect 16960 275440 17000 275445
rect 17040 275475 17080 275480
rect 17040 275445 17045 275475
rect 17075 275445 17080 275475
rect 17040 275440 17080 275445
rect 17120 275475 17160 275480
rect 17120 275445 17125 275475
rect 17155 275445 17160 275475
rect 17120 275440 17160 275445
rect 17200 275475 17240 275480
rect 17200 275445 17205 275475
rect 17235 275445 17240 275475
rect 17200 275440 17240 275445
rect 16720 275315 16760 275320
rect 16720 275285 16725 275315
rect 16755 275285 16760 275315
rect 16720 275280 16760 275285
rect 16880 275315 16920 275320
rect 16880 275285 16885 275315
rect 16915 275285 16920 275315
rect 16880 275280 16920 275285
rect 16960 275315 17000 275320
rect 16960 275285 16965 275315
rect 16995 275285 17000 275315
rect 16960 275280 17000 275285
rect 17040 275315 17080 275320
rect 17040 275285 17045 275315
rect 17075 275285 17080 275315
rect 17040 275280 17080 275285
rect 17200 275315 17240 275320
rect 17200 275285 17205 275315
rect 17235 275285 17240 275315
rect 17200 275280 17240 275285
rect 16720 274955 16760 274960
rect 16720 274925 16725 274955
rect 16755 274925 16760 274955
rect 16720 274920 16760 274925
rect 16880 274955 16920 274960
rect 16880 274925 16885 274955
rect 16915 274925 16920 274955
rect 16880 274920 16920 274925
rect 16720 274875 16760 274880
rect 16720 274845 16725 274875
rect 16755 274845 16760 274875
rect 16720 274840 16760 274845
rect 16880 274875 16920 274880
rect 16880 274845 16885 274875
rect 16915 274845 16920 274875
rect 16880 274840 16920 274845
rect 16720 274795 16760 274800
rect 16720 274765 16725 274795
rect 16755 274765 16760 274795
rect 16720 274760 16760 274765
rect 16880 274795 16920 274800
rect 16880 274765 16885 274795
rect 16915 274765 16920 274795
rect 16880 274760 16920 274765
rect 16720 274715 16760 274720
rect 16720 274685 16725 274715
rect 16755 274685 16760 274715
rect 16720 274680 16760 274685
rect 16880 274715 16920 274720
rect 16880 274685 16885 274715
rect 16915 274685 16920 274715
rect 16880 274680 16920 274685
rect 16720 274635 16760 274640
rect 16720 274605 16725 274635
rect 16755 274605 16760 274635
rect 16720 274600 16760 274605
rect 16880 274635 16920 274640
rect 16880 274605 16885 274635
rect 16915 274605 16920 274635
rect 16880 274600 16920 274605
rect 16720 274555 16760 274560
rect 16720 274525 16725 274555
rect 16755 274525 16760 274555
rect 16720 274520 16760 274525
rect 16880 274555 16920 274560
rect 16880 274525 16885 274555
rect 16915 274525 16920 274555
rect 16880 274520 16920 274525
rect 16720 274475 16760 274480
rect 16720 274445 16725 274475
rect 16755 274445 16760 274475
rect 16720 274440 16760 274445
rect 16880 274475 16920 274480
rect 16880 274445 16885 274475
rect 16915 274445 16920 274475
rect 16880 274440 16920 274445
rect 16720 274395 16760 274400
rect 16720 274365 16725 274395
rect 16755 274365 16760 274395
rect 16720 274360 16760 274365
rect 16880 274395 16920 274400
rect 16880 274365 16885 274395
rect 16915 274365 16920 274395
rect 16880 274360 16920 274365
rect 16720 274315 16760 274320
rect 16720 274285 16725 274315
rect 16755 274285 16760 274315
rect 16720 274280 16760 274285
rect 16880 274315 16920 274320
rect 16880 274285 16885 274315
rect 16915 274285 16920 274315
rect 16880 274280 16920 274285
rect 16720 274235 16760 274240
rect 16720 274205 16725 274235
rect 16755 274205 16760 274235
rect 16720 274200 16760 274205
rect 16880 274235 16920 274240
rect 16880 274205 16885 274235
rect 16915 274205 16920 274235
rect 16880 274200 16920 274205
rect 16720 274155 16760 274160
rect 16720 274125 16725 274155
rect 16755 274125 16760 274155
rect 16720 274120 16760 274125
rect 16880 274155 16920 274160
rect 16880 274125 16885 274155
rect 16915 274125 16920 274155
rect 16880 274120 16920 274125
rect 16720 274075 16760 274080
rect 16720 274045 16725 274075
rect 16755 274045 16760 274075
rect 16720 274040 16760 274045
rect 16880 274075 16920 274080
rect 16880 274045 16885 274075
rect 16915 274045 16920 274075
rect 16880 274040 16920 274045
rect 16720 273995 16760 274000
rect 16720 273965 16725 273995
rect 16755 273965 16760 273995
rect 16720 273960 16760 273965
rect 16880 273995 16920 274000
rect 16880 273965 16885 273995
rect 16915 273965 16920 273995
rect 16880 273960 16920 273965
rect 16720 273915 16760 273920
rect 16720 273885 16725 273915
rect 16755 273885 16760 273915
rect 16720 273880 16760 273885
rect 16880 273915 16920 273920
rect 16880 273885 16885 273915
rect 16915 273885 16920 273915
rect 16880 273880 16920 273885
rect 16720 273835 16760 273840
rect 16720 273805 16725 273835
rect 16755 273805 16760 273835
rect 16720 273800 16760 273805
rect 16880 273835 16920 273840
rect 16880 273805 16885 273835
rect 16915 273805 16920 273835
rect 16880 273800 16920 273805
rect 16720 273755 16760 273760
rect 16720 273725 16725 273755
rect 16755 273725 16760 273755
rect 16720 273720 16760 273725
rect 16880 273755 16920 273760
rect 16880 273725 16885 273755
rect 16915 273725 16920 273755
rect 16880 273720 16920 273725
rect 16720 273675 16760 273680
rect 16720 273645 16725 273675
rect 16755 273645 16760 273675
rect 16720 273640 16760 273645
rect 16880 273675 16920 273680
rect 16880 273645 16885 273675
rect 16915 273645 16920 273675
rect 16880 273640 16920 273645
rect 16720 273595 16760 273600
rect 16720 273565 16725 273595
rect 16755 273565 16760 273595
rect 16720 273560 16760 273565
rect 16880 273595 16920 273600
rect 16880 273565 16885 273595
rect 16915 273565 16920 273595
rect 16880 273560 16920 273565
rect 16720 273515 16760 273520
rect 16720 273485 16725 273515
rect 16755 273485 16760 273515
rect 16720 273480 16760 273485
rect 16880 273515 16920 273520
rect 16880 273485 16885 273515
rect 16915 273485 16920 273515
rect 16880 273480 16920 273485
rect 16720 273435 16760 273440
rect 16720 273405 16725 273435
rect 16755 273405 16760 273435
rect 16720 273400 16760 273405
rect 16880 273435 16920 273440
rect 16880 273405 16885 273435
rect 16915 273405 16920 273435
rect 16880 273400 16920 273405
rect 16720 273355 16760 273360
rect 16720 273325 16725 273355
rect 16755 273325 16760 273355
rect 16720 273320 16760 273325
rect 16880 273355 16920 273360
rect 16880 273325 16885 273355
rect 16915 273325 16920 273355
rect 16880 273320 16920 273325
rect 16720 273275 16760 273280
rect 16720 273245 16725 273275
rect 16755 273245 16760 273275
rect 16720 273240 16760 273245
rect 16880 273275 16920 273280
rect 16880 273245 16885 273275
rect 16915 273245 16920 273275
rect 16880 273240 16920 273245
rect 16720 273195 16760 273200
rect 16720 273165 16725 273195
rect 16755 273165 16760 273195
rect 16720 273160 16760 273165
rect 16880 273195 16920 273200
rect 16880 273165 16885 273195
rect 16915 273165 16920 273195
rect 16880 273160 16920 273165
rect 16720 273115 16760 273120
rect 16720 273085 16725 273115
rect 16755 273085 16760 273115
rect 16720 273080 16760 273085
rect 16880 273115 16920 273120
rect 16880 273085 16885 273115
rect 16915 273085 16920 273115
rect 16880 273080 16920 273085
rect 16720 273035 16760 273040
rect 16720 273005 16725 273035
rect 16755 273005 16760 273035
rect 16720 273000 16760 273005
rect 16880 273035 16920 273040
rect 16880 273005 16885 273035
rect 16915 273005 16920 273035
rect 16880 273000 16920 273005
rect 16720 272955 16760 272960
rect 16720 272925 16725 272955
rect 16755 272925 16760 272955
rect 16720 272920 16760 272925
rect 16880 272955 16920 272960
rect 16880 272925 16885 272955
rect 16915 272925 16920 272955
rect 16880 272920 16920 272925
rect 16720 272875 16760 272880
rect 16720 272845 16725 272875
rect 16755 272845 16760 272875
rect 16720 272840 16760 272845
rect 16880 272875 16920 272880
rect 16880 272845 16885 272875
rect 16915 272845 16920 272875
rect 16880 272840 16920 272845
rect 16720 272795 16760 272800
rect 16720 272765 16725 272795
rect 16755 272765 16760 272795
rect 16720 272760 16760 272765
rect 16880 272795 16920 272800
rect 16880 272765 16885 272795
rect 16915 272765 16920 272795
rect 16880 272760 16920 272765
rect 16720 272715 16760 272720
rect 16720 272685 16725 272715
rect 16755 272685 16760 272715
rect 16720 272680 16760 272685
rect 16880 272715 16920 272720
rect 16880 272685 16885 272715
rect 16915 272685 16920 272715
rect 16880 272680 16920 272685
rect 16720 272635 16760 272640
rect 16720 272605 16725 272635
rect 16755 272605 16760 272635
rect 16720 272600 16760 272605
rect 16880 272635 16920 272640
rect 16880 272605 16885 272635
rect 16915 272605 16920 272635
rect 16880 272600 16920 272605
rect 16720 272555 16760 272560
rect 16720 272525 16725 272555
rect 16755 272525 16760 272555
rect 16720 272520 16760 272525
rect 16880 272555 16920 272560
rect 16880 272525 16885 272555
rect 16915 272525 16920 272555
rect 16880 272520 16920 272525
rect 16720 272475 16760 272480
rect 16720 272445 16725 272475
rect 16755 272445 16760 272475
rect 16720 272440 16760 272445
rect 16880 272475 16920 272480
rect 16880 272445 16885 272475
rect 16915 272445 16920 272475
rect 16880 272440 16920 272445
rect 16720 272395 16760 272400
rect 16720 272365 16725 272395
rect 16755 272365 16760 272395
rect 16720 272360 16760 272365
rect 16880 272395 16920 272400
rect 16880 272365 16885 272395
rect 16915 272365 16920 272395
rect 16880 272360 16920 272365
rect 16720 272315 16760 272320
rect 16720 272285 16725 272315
rect 16755 272285 16760 272315
rect 16720 272280 16760 272285
rect 16880 272315 16920 272320
rect 16880 272285 16885 272315
rect 16915 272285 16920 272315
rect 16880 272280 16920 272285
rect 16720 272235 16760 272240
rect 16720 272205 16725 272235
rect 16755 272205 16760 272235
rect 16720 272200 16760 272205
rect 16880 272235 16920 272240
rect 16880 272205 16885 272235
rect 16915 272205 16920 272235
rect 16880 272200 16920 272205
rect 16720 272155 16760 272160
rect 16720 272125 16725 272155
rect 16755 272125 16760 272155
rect 16720 272120 16760 272125
rect 16880 272155 16920 272160
rect 16880 272125 16885 272155
rect 16915 272125 16920 272155
rect 16880 272120 16920 272125
rect 16720 272075 16760 272080
rect 16720 272045 16725 272075
rect 16755 272045 16760 272075
rect 16720 272040 16760 272045
rect 16880 272075 16920 272080
rect 16880 272045 16885 272075
rect 16915 272045 16920 272075
rect 16880 272040 16920 272045
rect 16720 271995 16760 272000
rect 16720 271965 16725 271995
rect 16755 271965 16760 271995
rect 16720 271960 16760 271965
rect 16880 271995 16920 272000
rect 16880 271965 16885 271995
rect 16915 271965 16920 271995
rect 16880 271960 16920 271965
rect 16720 271915 16760 271920
rect 16720 271885 16725 271915
rect 16755 271885 16760 271915
rect 16720 271880 16760 271885
rect 16880 271915 16920 271920
rect 16880 271885 16885 271915
rect 16915 271885 16920 271915
rect 16880 271880 16920 271885
rect 16720 271835 16760 271840
rect 16720 271805 16725 271835
rect 16755 271805 16760 271835
rect 16720 271800 16760 271805
rect 16880 271835 16920 271840
rect 16880 271805 16885 271835
rect 16915 271805 16920 271835
rect 16880 271800 16920 271805
rect 16720 271755 16760 271760
rect 16720 271725 16725 271755
rect 16755 271725 16760 271755
rect 16720 271720 16760 271725
rect 16880 271755 16920 271760
rect 16880 271725 16885 271755
rect 16915 271725 16920 271755
rect 16880 271720 16920 271725
rect 16720 271675 16760 271680
rect 16720 271645 16725 271675
rect 16755 271645 16760 271675
rect 16720 271640 16760 271645
rect 16880 271675 16920 271680
rect 16880 271645 16885 271675
rect 16915 271645 16920 271675
rect 16880 271640 16920 271645
rect 16720 271595 16760 271600
rect 16720 271565 16725 271595
rect 16755 271565 16760 271595
rect 16720 271560 16760 271565
rect 16880 271595 16920 271600
rect 16880 271565 16885 271595
rect 16915 271565 16920 271595
rect 16880 271560 16920 271565
rect 16720 271515 16760 271520
rect 16720 271485 16725 271515
rect 16755 271485 16760 271515
rect 16720 271480 16760 271485
rect 16880 271515 16920 271520
rect 16880 271485 16885 271515
rect 16915 271485 16920 271515
rect 16880 271480 16920 271485
rect 16720 271435 16760 271440
rect 16720 271405 16725 271435
rect 16755 271405 16760 271435
rect 16720 271400 16760 271405
rect 16880 271435 16920 271440
rect 16880 271405 16885 271435
rect 16915 271405 16920 271435
rect 16880 271400 16920 271405
rect 16720 271355 16760 271360
rect 16720 271325 16725 271355
rect 16755 271325 16760 271355
rect 16720 271320 16760 271325
rect 16880 271355 16920 271360
rect 16880 271325 16885 271355
rect 16915 271325 16920 271355
rect 16880 271320 16920 271325
rect 16720 271275 16760 271280
rect 16720 271245 16725 271275
rect 16755 271245 16760 271275
rect 16720 271240 16760 271245
rect 16880 271275 16920 271280
rect 16880 271245 16885 271275
rect 16915 271245 16920 271275
rect 16880 271240 16920 271245
rect 16720 271195 16760 271200
rect 16720 271165 16725 271195
rect 16755 271165 16760 271195
rect 16720 271160 16760 271165
rect 16880 271195 16920 271200
rect 16880 271165 16885 271195
rect 16915 271165 16920 271195
rect 16880 271160 16920 271165
rect 16720 271115 16760 271120
rect 16720 271085 16725 271115
rect 16755 271085 16760 271115
rect 16720 271080 16760 271085
rect 16880 271115 16920 271120
rect 16880 271085 16885 271115
rect 16915 271085 16920 271115
rect 16880 271080 16920 271085
rect 16720 271035 16760 271040
rect 16720 271005 16725 271035
rect 16755 271005 16760 271035
rect 16720 271000 16760 271005
rect 16880 271035 16920 271040
rect 16880 271005 16885 271035
rect 16915 271005 16920 271035
rect 16880 271000 16920 271005
rect 16720 270955 16760 270960
rect 16720 270925 16725 270955
rect 16755 270925 16760 270955
rect 16720 270920 16760 270925
rect 16880 270955 16920 270960
rect 16880 270925 16885 270955
rect 16915 270925 16920 270955
rect 16880 270920 16920 270925
rect 16720 270875 16760 270880
rect 16720 270845 16725 270875
rect 16755 270845 16760 270875
rect 16720 270840 16760 270845
rect 16880 270875 16920 270880
rect 16880 270845 16885 270875
rect 16915 270845 16920 270875
rect 16880 270840 16920 270845
rect 16720 270795 16760 270800
rect 16720 270765 16725 270795
rect 16755 270765 16760 270795
rect 16720 270760 16760 270765
rect 16880 270795 16920 270800
rect 16880 270765 16885 270795
rect 16915 270765 16920 270795
rect 16880 270760 16920 270765
rect 16720 270715 16760 270720
rect 16720 270685 16725 270715
rect 16755 270685 16760 270715
rect 16720 270680 16760 270685
rect 16880 270715 16920 270720
rect 16880 270685 16885 270715
rect 16915 270685 16920 270715
rect 16880 270680 16920 270685
rect 16720 270635 16760 270640
rect 16720 270605 16725 270635
rect 16755 270605 16760 270635
rect 16720 270600 16760 270605
rect 16880 270635 16920 270640
rect 16880 270605 16885 270635
rect 16915 270605 16920 270635
rect 16880 270600 16920 270605
rect 16720 270555 16760 270560
rect 16720 270525 16725 270555
rect 16755 270525 16760 270555
rect 16720 270520 16760 270525
rect 16880 270555 16920 270560
rect 16880 270525 16885 270555
rect 16915 270525 16920 270555
rect 16880 270520 16920 270525
rect 16720 270475 16760 270480
rect 16720 270445 16725 270475
rect 16755 270445 16760 270475
rect 16720 270440 16760 270445
rect 16880 270475 16920 270480
rect 16880 270445 16885 270475
rect 16915 270445 16920 270475
rect 16880 270440 16920 270445
rect 16720 270395 16760 270400
rect 16720 270365 16725 270395
rect 16755 270365 16760 270395
rect 16720 270360 16760 270365
rect 16880 270395 16920 270400
rect 16880 270365 16885 270395
rect 16915 270365 16920 270395
rect 16880 270360 16920 270365
rect 16720 270315 16760 270320
rect 16720 270285 16725 270315
rect 16755 270285 16760 270315
rect 16720 270280 16760 270285
rect 16880 270315 16920 270320
rect 16880 270285 16885 270315
rect 16915 270285 16920 270315
rect 16880 270280 16920 270285
rect 16720 270235 16760 270240
rect 16720 270205 16725 270235
rect 16755 270205 16760 270235
rect 16720 270200 16760 270205
rect 16880 270235 16920 270240
rect 16880 270205 16885 270235
rect 16915 270205 16920 270235
rect 16880 270200 16920 270205
rect 16720 270155 16760 270160
rect 16720 270125 16725 270155
rect 16755 270125 16760 270155
rect 16720 270120 16760 270125
rect 16880 270155 16920 270160
rect 16880 270125 16885 270155
rect 16915 270125 16920 270155
rect 16880 270120 16920 270125
rect 16720 270075 16760 270080
rect 16720 270045 16725 270075
rect 16755 270045 16760 270075
rect 16720 270040 16760 270045
rect 16880 270075 16920 270080
rect 16880 270045 16885 270075
rect 16915 270045 16920 270075
rect 16880 270040 16920 270045
rect 16720 269995 16760 270000
rect 16720 269965 16725 269995
rect 16755 269965 16760 269995
rect 16720 269960 16760 269965
rect 16880 269995 16920 270000
rect 16880 269965 16885 269995
rect 16915 269965 16920 269995
rect 16880 269960 16920 269965
rect 16720 269915 16760 269920
rect 16720 269885 16725 269915
rect 16755 269885 16760 269915
rect 16720 269880 16760 269885
rect 16880 269915 16920 269920
rect 16880 269885 16885 269915
rect 16915 269885 16920 269915
rect 16880 269880 16920 269885
rect 16720 269835 16760 269840
rect 16720 269805 16725 269835
rect 16755 269805 16760 269835
rect 16720 269800 16760 269805
rect 16880 269835 16920 269840
rect 16880 269805 16885 269835
rect 16915 269805 16920 269835
rect 16880 269800 16920 269805
rect 16720 269755 16760 269760
rect 16720 269725 16725 269755
rect 16755 269725 16760 269755
rect 16720 269720 16760 269725
rect 16880 269755 16920 269760
rect 16880 269725 16885 269755
rect 16915 269725 16920 269755
rect 16880 269720 16920 269725
rect 16720 269675 16760 269680
rect 16720 269645 16725 269675
rect 16755 269645 16760 269675
rect 16720 269640 16760 269645
rect 16880 269675 16920 269680
rect 16880 269645 16885 269675
rect 16915 269645 16920 269675
rect 16880 269640 16920 269645
rect 16720 269595 16760 269600
rect 16720 269565 16725 269595
rect 16755 269565 16760 269595
rect 16720 269560 16760 269565
rect 16880 269595 16920 269600
rect 16880 269565 16885 269595
rect 16915 269565 16920 269595
rect 16880 269560 16920 269565
rect 16720 269515 16760 269520
rect 16720 269485 16725 269515
rect 16755 269485 16760 269515
rect 16720 269480 16760 269485
rect 16880 269515 16920 269520
rect 16880 269485 16885 269515
rect 16915 269485 16920 269515
rect 16880 269480 16920 269485
rect 16720 269435 16760 269440
rect 16720 269405 16725 269435
rect 16755 269405 16760 269435
rect 16720 269400 16760 269405
rect 16880 269435 16920 269440
rect 16880 269405 16885 269435
rect 16915 269405 16920 269435
rect 16880 269400 16920 269405
rect 16720 269355 16760 269360
rect 16720 269325 16725 269355
rect 16755 269325 16760 269355
rect 16720 269320 16760 269325
rect 16880 269355 16920 269360
rect 16880 269325 16885 269355
rect 16915 269325 16920 269355
rect 16880 269320 16920 269325
rect 16720 269275 16760 269280
rect 16720 269245 16725 269275
rect 16755 269245 16760 269275
rect 16720 269240 16760 269245
rect 16880 269275 16920 269280
rect 16880 269245 16885 269275
rect 16915 269245 16920 269275
rect 16880 269240 16920 269245
rect 16720 269195 16760 269200
rect 16720 269165 16725 269195
rect 16755 269165 16760 269195
rect 16720 269160 16760 269165
rect 16880 269195 16920 269200
rect 16880 269165 16885 269195
rect 16915 269165 16920 269195
rect 16880 269160 16920 269165
rect 16720 269115 16760 269120
rect 16720 269085 16725 269115
rect 16755 269085 16760 269115
rect 16720 269080 16760 269085
rect 16880 269115 16920 269120
rect 16880 269085 16885 269115
rect 16915 269085 16920 269115
rect 16880 269080 16920 269085
rect 16720 269035 16760 269040
rect 16720 269005 16725 269035
rect 16755 269005 16760 269035
rect 16720 269000 16760 269005
rect 16880 269035 16920 269040
rect 16880 269005 16885 269035
rect 16915 269005 16920 269035
rect 16880 269000 16920 269005
rect 16720 268955 16760 268960
rect 16720 268925 16725 268955
rect 16755 268925 16760 268955
rect 16720 268920 16760 268925
rect 16880 268955 16920 268960
rect 16880 268925 16885 268955
rect 16915 268925 16920 268955
rect 16880 268920 16920 268925
rect 16720 268875 16760 268880
rect 16720 268845 16725 268875
rect 16755 268845 16760 268875
rect 16720 268840 16760 268845
rect 16880 268875 16920 268880
rect 16880 268845 16885 268875
rect 16915 268845 16920 268875
rect 16880 268840 16920 268845
rect 16720 268795 16760 268800
rect 16720 268765 16725 268795
rect 16755 268765 16760 268795
rect 16720 268760 16760 268765
rect 16880 268795 16920 268800
rect 16880 268765 16885 268795
rect 16915 268765 16920 268795
rect 16880 268760 16920 268765
rect 16720 268715 16760 268720
rect 16720 268685 16725 268715
rect 16755 268685 16760 268715
rect 16720 268680 16760 268685
rect 16880 268715 16920 268720
rect 16880 268685 16885 268715
rect 16915 268685 16920 268715
rect 16880 268680 16920 268685
rect 16720 268635 16760 268640
rect 16720 268605 16725 268635
rect 16755 268605 16760 268635
rect 16720 268600 16760 268605
rect 16880 268635 16920 268640
rect 16880 268605 16885 268635
rect 16915 268605 16920 268635
rect 16880 268600 16920 268605
rect 16720 268555 16760 268560
rect 16720 268525 16725 268555
rect 16755 268525 16760 268555
rect 16720 268520 16760 268525
rect 16880 268555 16920 268560
rect 16880 268525 16885 268555
rect 16915 268525 16920 268555
rect 16880 268520 16920 268525
rect 16720 268475 16760 268480
rect 16720 268445 16725 268475
rect 16755 268445 16760 268475
rect 16720 268440 16760 268445
rect 16880 268475 16920 268480
rect 16880 268445 16885 268475
rect 16915 268445 16920 268475
rect 16880 268440 16920 268445
rect 16720 268395 16760 268400
rect 16720 268365 16725 268395
rect 16755 268365 16760 268395
rect 16720 268360 16760 268365
rect 16880 268395 16920 268400
rect 16880 268365 16885 268395
rect 16915 268365 16920 268395
rect 16880 268360 16920 268365
rect 16720 268315 16760 268320
rect 16720 268285 16725 268315
rect 16755 268285 16760 268315
rect 16720 268280 16760 268285
rect 16880 268315 16920 268320
rect 16880 268285 16885 268315
rect 16915 268285 16920 268315
rect 16880 268280 16920 268285
rect 16720 268235 16760 268240
rect 16720 268205 16725 268235
rect 16755 268205 16760 268235
rect 16720 268200 16760 268205
rect 16880 268235 16920 268240
rect 16880 268205 16885 268235
rect 16915 268205 16920 268235
rect 16880 268200 16920 268205
rect 16720 268155 16760 268160
rect 16720 268125 16725 268155
rect 16755 268125 16760 268155
rect 16720 268120 16760 268125
rect 16880 268155 16920 268160
rect 16880 268125 16885 268155
rect 16915 268125 16920 268155
rect 16880 268120 16920 268125
rect 16720 268075 16760 268080
rect 16720 268045 16725 268075
rect 16755 268045 16760 268075
rect 16720 268040 16760 268045
rect 16880 268075 16920 268080
rect 16880 268045 16885 268075
rect 16915 268045 16920 268075
rect 16880 268040 16920 268045
rect 16720 267995 16760 268000
rect 16720 267965 16725 267995
rect 16755 267965 16760 267995
rect 16720 267960 16760 267965
rect 16880 267995 16920 268000
rect 16880 267965 16885 267995
rect 16915 267965 16920 267995
rect 16880 267960 16920 267965
rect 16720 267915 16760 267920
rect 16720 267885 16725 267915
rect 16755 267885 16760 267915
rect 16720 267880 16760 267885
rect 16880 267915 16920 267920
rect 16880 267885 16885 267915
rect 16915 267885 16920 267915
rect 16880 267880 16920 267885
rect 16720 267835 16760 267840
rect 16720 267805 16725 267835
rect 16755 267805 16760 267835
rect 16720 267800 16760 267805
rect 16880 267835 16920 267840
rect 16880 267805 16885 267835
rect 16915 267805 16920 267835
rect 16880 267800 16920 267805
rect 16720 267755 16760 267760
rect 16720 267725 16725 267755
rect 16755 267725 16760 267755
rect 16720 267720 16760 267725
rect 16880 267755 16920 267760
rect 16880 267725 16885 267755
rect 16915 267725 16920 267755
rect 16880 267720 16920 267725
rect 16720 267675 16760 267680
rect 16720 267645 16725 267675
rect 16755 267645 16760 267675
rect 16720 267640 16760 267645
rect 16880 267675 16920 267680
rect 16880 267645 16885 267675
rect 16915 267645 16920 267675
rect 16880 267640 16920 267645
rect 16720 267595 16760 267600
rect 16720 267565 16725 267595
rect 16755 267565 16760 267595
rect 16720 267560 16760 267565
rect 16880 267595 16920 267600
rect 16880 267565 16885 267595
rect 16915 267565 16920 267595
rect 16880 267560 16920 267565
rect 16720 267515 16760 267520
rect 16720 267485 16725 267515
rect 16755 267485 16760 267515
rect 16720 267480 16760 267485
rect 16880 267515 16920 267520
rect 16880 267485 16885 267515
rect 16915 267485 16920 267515
rect 16880 267480 16920 267485
rect 16720 267435 16760 267440
rect 16720 267405 16725 267435
rect 16755 267405 16760 267435
rect 16720 267400 16760 267405
rect 16880 267435 16920 267440
rect 16880 267405 16885 267435
rect 16915 267405 16920 267435
rect 16880 267400 16920 267405
rect 16720 267355 16760 267360
rect 16720 267325 16725 267355
rect 16755 267325 16760 267355
rect 16720 267320 16760 267325
rect 16880 267355 16920 267360
rect 16880 267325 16885 267355
rect 16915 267325 16920 267355
rect 16880 267320 16920 267325
rect 16720 267275 16760 267280
rect 16720 267245 16725 267275
rect 16755 267245 16760 267275
rect 16720 267240 16760 267245
rect 16880 267275 16920 267280
rect 16880 267245 16885 267275
rect 16915 267245 16920 267275
rect 16880 267240 16920 267245
rect 16720 267195 16760 267200
rect 16720 267165 16725 267195
rect 16755 267165 16760 267195
rect 16720 267160 16760 267165
rect 16880 267195 16920 267200
rect 16880 267165 16885 267195
rect 16915 267165 16920 267195
rect 16880 267160 16920 267165
rect 16720 267115 16760 267120
rect 16720 267085 16725 267115
rect 16755 267085 16760 267115
rect 16720 267080 16760 267085
rect 16880 267115 16920 267120
rect 16880 267085 16885 267115
rect 16915 267085 16920 267115
rect 16880 267080 16920 267085
rect 16720 267035 16760 267040
rect 16720 267005 16725 267035
rect 16755 267005 16760 267035
rect 16720 267000 16760 267005
rect 16880 267035 16920 267040
rect 16880 267005 16885 267035
rect 16915 267005 16920 267035
rect 16880 267000 16920 267005
rect 16720 266955 16760 266960
rect 16720 266925 16725 266955
rect 16755 266925 16760 266955
rect 16720 266920 16760 266925
rect 16880 266955 16920 266960
rect 16880 266925 16885 266955
rect 16915 266925 16920 266955
rect 16880 266920 16920 266925
rect 16720 266875 16760 266880
rect 16720 266845 16725 266875
rect 16755 266845 16760 266875
rect 16720 266840 16760 266845
rect 16880 266875 16920 266880
rect 16880 266845 16885 266875
rect 16915 266845 16920 266875
rect 16880 266840 16920 266845
rect 16720 266795 16760 266800
rect 16720 266765 16725 266795
rect 16755 266765 16760 266795
rect 16720 266760 16760 266765
rect 16880 266795 16920 266800
rect 16880 266765 16885 266795
rect 16915 266765 16920 266795
rect 16880 266760 16920 266765
rect 16720 266715 16760 266720
rect 16720 266685 16725 266715
rect 16755 266685 16760 266715
rect 16720 266680 16760 266685
rect 16880 266715 16920 266720
rect 16880 266685 16885 266715
rect 16915 266685 16920 266715
rect 16880 266680 16920 266685
rect 16720 266635 16760 266640
rect 16720 266605 16725 266635
rect 16755 266605 16760 266635
rect 16720 266600 16760 266605
rect 16880 266635 16920 266640
rect 16880 266605 16885 266635
rect 16915 266605 16920 266635
rect 16880 266600 16920 266605
rect 16720 266555 16760 266560
rect 16720 266525 16725 266555
rect 16755 266525 16760 266555
rect 16720 266520 16760 266525
rect 16880 266555 16920 266560
rect 16880 266525 16885 266555
rect 16915 266525 16920 266555
rect 16880 266520 16920 266525
rect 16720 266475 16760 266480
rect 16720 266445 16725 266475
rect 16755 266445 16760 266475
rect 16720 266440 16760 266445
rect 16880 266475 16920 266480
rect 16880 266445 16885 266475
rect 16915 266445 16920 266475
rect 16880 266440 16920 266445
rect 16720 266395 16760 266400
rect 16720 266365 16725 266395
rect 16755 266365 16760 266395
rect 16720 266360 16760 266365
rect 16880 266395 16920 266400
rect 16880 266365 16885 266395
rect 16915 266365 16920 266395
rect 16880 266360 16920 266365
rect 16720 266315 16760 266320
rect 16720 266285 16725 266315
rect 16755 266285 16760 266315
rect 16720 266280 16760 266285
rect 16880 266315 16920 266320
rect 16880 266285 16885 266315
rect 16915 266285 16920 266315
rect 16880 266280 16920 266285
rect 16720 266235 16760 266240
rect 16720 266205 16725 266235
rect 16755 266205 16760 266235
rect 16720 266200 16760 266205
rect 16880 266235 16920 266240
rect 16880 266205 16885 266235
rect 16915 266205 16920 266235
rect 16880 266200 16920 266205
rect 16720 266155 16760 266160
rect 16720 266125 16725 266155
rect 16755 266125 16760 266155
rect 16720 266120 16760 266125
rect 16880 266155 16920 266160
rect 16880 266125 16885 266155
rect 16915 266125 16920 266155
rect 16880 266120 16920 266125
rect 16720 266075 16760 266080
rect 16720 266045 16725 266075
rect 16755 266045 16760 266075
rect 16720 266040 16760 266045
rect 16880 266075 16920 266080
rect 16880 266045 16885 266075
rect 16915 266045 16920 266075
rect 16880 266040 16920 266045
rect 16720 265995 16760 266000
rect 16720 265965 16725 265995
rect 16755 265965 16760 265995
rect 16720 265960 16760 265965
rect 16880 265995 16920 266000
rect 16880 265965 16885 265995
rect 16915 265965 16920 265995
rect 16880 265960 16920 265965
rect 16720 265915 16760 265920
rect 16720 265885 16725 265915
rect 16755 265885 16760 265915
rect 16720 265880 16760 265885
rect 16880 265915 16920 265920
rect 16880 265885 16885 265915
rect 16915 265885 16920 265915
rect 16880 265880 16920 265885
rect 16720 265835 16760 265840
rect 16720 265805 16725 265835
rect 16755 265805 16760 265835
rect 16720 265800 16760 265805
rect 16880 265835 16920 265840
rect 16880 265805 16885 265835
rect 16915 265805 16920 265835
rect 16880 265800 16920 265805
rect 16720 265755 16760 265760
rect 16720 265725 16725 265755
rect 16755 265725 16760 265755
rect 16720 265720 16760 265725
rect 16880 265755 16920 265760
rect 16880 265725 16885 265755
rect 16915 265725 16920 265755
rect 16880 265720 16920 265725
rect 16720 265675 16760 265680
rect 16720 265645 16725 265675
rect 16755 265645 16760 265675
rect 16720 265640 16760 265645
rect 16880 265675 16920 265680
rect 16880 265645 16885 265675
rect 16915 265645 16920 265675
rect 16880 265640 16920 265645
rect 16720 265595 16760 265600
rect 16720 265565 16725 265595
rect 16755 265565 16760 265595
rect 16720 265560 16760 265565
rect 16880 265595 16920 265600
rect 16880 265565 16885 265595
rect 16915 265565 16920 265595
rect 16880 265560 16920 265565
rect 16720 265515 16760 265520
rect 16720 265485 16725 265515
rect 16755 265485 16760 265515
rect 16720 265480 16760 265485
rect 16880 265515 16920 265520
rect 16880 265485 16885 265515
rect 16915 265485 16920 265515
rect 16880 265480 16920 265485
rect 16720 265435 16760 265440
rect 16720 265405 16725 265435
rect 16755 265405 16760 265435
rect 16720 265400 16760 265405
rect 16880 265435 16920 265440
rect 16880 265405 16885 265435
rect 16915 265405 16920 265435
rect 16880 265400 16920 265405
rect 16720 265355 16760 265360
rect 16720 265325 16725 265355
rect 16755 265325 16760 265355
rect 16720 265320 16760 265325
rect 16880 265355 16920 265360
rect 16880 265325 16885 265355
rect 16915 265325 16920 265355
rect 16880 265320 16920 265325
rect 16720 265275 16760 265280
rect 16720 265245 16725 265275
rect 16755 265245 16760 265275
rect 16720 265240 16760 265245
rect 16880 265275 16920 265280
rect 16880 265245 16885 265275
rect 16915 265245 16920 265275
rect 16880 265240 16920 265245
rect 16720 265195 16760 265200
rect 16720 265165 16725 265195
rect 16755 265165 16760 265195
rect 16720 265160 16760 265165
rect 16880 265195 16920 265200
rect 16880 265165 16885 265195
rect 16915 265165 16920 265195
rect 16880 265160 16920 265165
rect 16720 265115 16760 265120
rect 16720 265085 16725 265115
rect 16755 265085 16760 265115
rect 16720 265080 16760 265085
rect 16880 265115 16920 265120
rect 16880 265085 16885 265115
rect 16915 265085 16920 265115
rect 16880 265080 16920 265085
rect 16720 265035 16760 265040
rect 16720 265005 16725 265035
rect 16755 265005 16760 265035
rect 16720 265000 16760 265005
rect 16880 265035 16920 265040
rect 16880 265005 16885 265035
rect 16915 265005 16920 265035
rect 16880 265000 16920 265005
rect 16720 264955 16760 264960
rect 16720 264925 16725 264955
rect 16755 264925 16760 264955
rect 16720 264920 16760 264925
rect 16880 264955 16920 264960
rect 16880 264925 16885 264955
rect 16915 264925 16920 264955
rect 16880 264920 16920 264925
rect 16720 264875 16760 264880
rect 16720 264845 16725 264875
rect 16755 264845 16760 264875
rect 16720 264840 16760 264845
rect 16880 264875 16920 264880
rect 16880 264845 16885 264875
rect 16915 264845 16920 264875
rect 16880 264840 16920 264845
rect 16720 264795 16760 264800
rect 16720 264765 16725 264795
rect 16755 264765 16760 264795
rect 16720 264760 16760 264765
rect 16880 264795 16920 264800
rect 16880 264765 16885 264795
rect 16915 264765 16920 264795
rect 16880 264760 16920 264765
rect 16720 264715 16760 264720
rect 16720 264685 16725 264715
rect 16755 264685 16760 264715
rect 16720 264680 16760 264685
rect 16880 264715 16920 264720
rect 16880 264685 16885 264715
rect 16915 264685 16920 264715
rect 16880 264680 16920 264685
rect 16720 264635 16760 264640
rect 16720 264605 16725 264635
rect 16755 264605 16760 264635
rect 16720 264600 16760 264605
rect 16880 264635 16920 264640
rect 16880 264605 16885 264635
rect 16915 264605 16920 264635
rect 16880 264600 16920 264605
rect 16720 264555 16760 264560
rect 16720 264525 16725 264555
rect 16755 264525 16760 264555
rect 16720 264520 16760 264525
rect 16880 264555 16920 264560
rect 16880 264525 16885 264555
rect 16915 264525 16920 264555
rect 16880 264520 16920 264525
rect 16720 264475 16760 264480
rect 16720 264445 16725 264475
rect 16755 264445 16760 264475
rect 16720 264440 16760 264445
rect 16880 264475 16920 264480
rect 16880 264445 16885 264475
rect 16915 264445 16920 264475
rect 16880 264440 16920 264445
rect 16720 264395 16760 264400
rect 16720 264365 16725 264395
rect 16755 264365 16760 264395
rect 16720 264360 16760 264365
rect 16880 264395 16920 264400
rect 16880 264365 16885 264395
rect 16915 264365 16920 264395
rect 16880 264360 16920 264365
rect 16720 264315 16760 264320
rect 16720 264285 16725 264315
rect 16755 264285 16760 264315
rect 16720 264280 16760 264285
rect 16880 264315 16920 264320
rect 16880 264285 16885 264315
rect 16915 264285 16920 264315
rect 16880 264280 16920 264285
rect 16720 264235 16760 264240
rect 16720 264205 16725 264235
rect 16755 264205 16760 264235
rect 16720 264200 16760 264205
rect 16880 264235 16920 264240
rect 16880 264205 16885 264235
rect 16915 264205 16920 264235
rect 16880 264200 16920 264205
rect 16720 264155 16760 264160
rect 16720 264125 16725 264155
rect 16755 264125 16760 264155
rect 16720 264120 16760 264125
rect 16880 264155 16920 264160
rect 16880 264125 16885 264155
rect 16915 264125 16920 264155
rect 16880 264120 16920 264125
rect 16720 264075 16760 264080
rect 16720 264045 16725 264075
rect 16755 264045 16760 264075
rect 16720 264040 16760 264045
rect 16880 264075 16920 264080
rect 16880 264045 16885 264075
rect 16915 264045 16920 264075
rect 16880 264040 16920 264045
rect 16720 263995 16760 264000
rect 16720 263965 16725 263995
rect 16755 263965 16760 263995
rect 16720 263960 16760 263965
rect 16880 263995 16920 264000
rect 16880 263965 16885 263995
rect 16915 263965 16920 263995
rect 16880 263960 16920 263965
rect 16720 263915 16760 263920
rect 16720 263885 16725 263915
rect 16755 263885 16760 263915
rect 16720 263880 16760 263885
rect 16880 263915 16920 263920
rect 16880 263885 16885 263915
rect 16915 263885 16920 263915
rect 16880 263880 16920 263885
rect 16720 263835 16760 263840
rect 16720 263805 16725 263835
rect 16755 263805 16760 263835
rect 16720 263800 16760 263805
rect 16880 263835 16920 263840
rect 16880 263805 16885 263835
rect 16915 263805 16920 263835
rect 16880 263800 16920 263805
rect 16720 263755 16760 263760
rect 16720 263725 16725 263755
rect 16755 263725 16760 263755
rect 16720 263720 16760 263725
rect 16880 263755 16920 263760
rect 16880 263725 16885 263755
rect 16915 263725 16920 263755
rect 16880 263720 16920 263725
rect 16720 263675 16760 263680
rect 16720 263645 16725 263675
rect 16755 263645 16760 263675
rect 16720 263640 16760 263645
rect 16880 263675 16920 263680
rect 16880 263645 16885 263675
rect 16915 263645 16920 263675
rect 16880 263640 16920 263645
rect 16720 263595 16760 263600
rect 16720 263565 16725 263595
rect 16755 263565 16760 263595
rect 16720 263560 16760 263565
rect 16880 263595 16920 263600
rect 16880 263565 16885 263595
rect 16915 263565 16920 263595
rect 16880 263560 16920 263565
rect 16720 263515 16760 263520
rect 16720 263485 16725 263515
rect 16755 263485 16760 263515
rect 16720 263480 16760 263485
rect 16880 263515 16920 263520
rect 16880 263485 16885 263515
rect 16915 263485 16920 263515
rect 16880 263480 16920 263485
rect 16720 263435 16760 263440
rect 16720 263405 16725 263435
rect 16755 263405 16760 263435
rect 16720 263400 16760 263405
rect 16880 263435 16920 263440
rect 16880 263405 16885 263435
rect 16915 263405 16920 263435
rect 16880 263400 16920 263405
rect 16720 263355 16760 263360
rect 16720 263325 16725 263355
rect 16755 263325 16760 263355
rect 16720 263320 16760 263325
rect 16880 263355 16920 263360
rect 16880 263325 16885 263355
rect 16915 263325 16920 263355
rect 16880 263320 16920 263325
rect 16720 263275 16760 263280
rect 16720 263245 16725 263275
rect 16755 263245 16760 263275
rect 16720 263240 16760 263245
rect 16880 263275 16920 263280
rect 16880 263245 16885 263275
rect 16915 263245 16920 263275
rect 16880 263240 16920 263245
rect 16720 263195 16760 263200
rect 16720 263165 16725 263195
rect 16755 263165 16760 263195
rect 16720 263160 16760 263165
rect 16880 263195 16920 263200
rect 16880 263165 16885 263195
rect 16915 263165 16920 263195
rect 16880 263160 16920 263165
rect 16720 263115 16760 263120
rect 16720 263085 16725 263115
rect 16755 263085 16760 263115
rect 16720 263080 16760 263085
rect 16880 263115 16920 263120
rect 16880 263085 16885 263115
rect 16915 263085 16920 263115
rect 16880 263080 16920 263085
rect 16720 263035 16760 263040
rect 16720 263005 16725 263035
rect 16755 263005 16760 263035
rect 16720 263000 16760 263005
rect 16880 263035 16920 263040
rect 16880 263005 16885 263035
rect 16915 263005 16920 263035
rect 16880 263000 16920 263005
rect 16720 262955 16760 262960
rect 16720 262925 16725 262955
rect 16755 262925 16760 262955
rect 16720 262920 16760 262925
rect 16880 262955 16920 262960
rect 16880 262925 16885 262955
rect 16915 262925 16920 262955
rect 16880 262920 16920 262925
rect 16720 262875 16760 262880
rect 16720 262845 16725 262875
rect 16755 262845 16760 262875
rect 16720 262840 16760 262845
rect 16880 262875 16920 262880
rect 16880 262845 16885 262875
rect 16915 262845 16920 262875
rect 16880 262840 16920 262845
rect 16720 262795 16760 262800
rect 16720 262765 16725 262795
rect 16755 262765 16760 262795
rect 16720 262760 16760 262765
rect 16880 262795 16920 262800
rect 16880 262765 16885 262795
rect 16915 262765 16920 262795
rect 16880 262760 16920 262765
rect 16720 262715 16760 262720
rect 16720 262685 16725 262715
rect 16755 262685 16760 262715
rect 16720 262680 16760 262685
rect 16880 262715 16920 262720
rect 16880 262685 16885 262715
rect 16915 262685 16920 262715
rect 16880 262680 16920 262685
rect 16720 262635 16760 262640
rect 16720 262605 16725 262635
rect 16755 262605 16760 262635
rect 16720 262600 16760 262605
rect 16880 262635 16920 262640
rect 16880 262605 16885 262635
rect 16915 262605 16920 262635
rect 16880 262600 16920 262605
rect 16720 262555 16760 262560
rect 16720 262525 16725 262555
rect 16755 262525 16760 262555
rect 16720 262520 16760 262525
rect 16880 262555 16920 262560
rect 16880 262525 16885 262555
rect 16915 262525 16920 262555
rect 16880 262520 16920 262525
rect 16720 262475 16760 262480
rect 16720 262445 16725 262475
rect 16755 262445 16760 262475
rect 16720 262440 16760 262445
rect 16880 262475 16920 262480
rect 16880 262445 16885 262475
rect 16915 262445 16920 262475
rect 16880 262440 16920 262445
rect 16720 262395 16760 262400
rect 16720 262365 16725 262395
rect 16755 262365 16760 262395
rect 16720 262360 16760 262365
rect 16880 262395 16920 262400
rect 16880 262365 16885 262395
rect 16915 262365 16920 262395
rect 16880 262360 16920 262365
rect 16720 262315 16760 262320
rect 16720 262285 16725 262315
rect 16755 262285 16760 262315
rect 16720 262280 16760 262285
rect 16880 262315 16920 262320
rect 16880 262285 16885 262315
rect 16915 262285 16920 262315
rect 16880 262280 16920 262285
rect 16720 262235 16760 262240
rect 16720 262205 16725 262235
rect 16755 262205 16760 262235
rect 16720 262200 16760 262205
rect 16880 262235 16920 262240
rect 16880 262205 16885 262235
rect 16915 262205 16920 262235
rect 16880 262200 16920 262205
rect 16720 262155 16760 262160
rect 16720 262125 16725 262155
rect 16755 262125 16760 262155
rect 16720 262120 16760 262125
rect 16880 262155 16920 262160
rect 16880 262125 16885 262155
rect 16915 262125 16920 262155
rect 16880 262120 16920 262125
rect 16720 262075 16760 262080
rect 16720 262045 16725 262075
rect 16755 262045 16760 262075
rect 16720 262040 16760 262045
rect 16880 262075 16920 262080
rect 16880 262045 16885 262075
rect 16915 262045 16920 262075
rect 16880 262040 16920 262045
rect 16720 261995 16760 262000
rect 16720 261965 16725 261995
rect 16755 261965 16760 261995
rect 16720 261960 16760 261965
rect 16880 261995 16920 262000
rect 16880 261965 16885 261995
rect 16915 261965 16920 261995
rect 16880 261960 16920 261965
rect 16720 261915 16760 261920
rect 16720 261885 16725 261915
rect 16755 261885 16760 261915
rect 16720 261880 16760 261885
rect 16880 261915 16920 261920
rect 16880 261885 16885 261915
rect 16915 261885 16920 261915
rect 16880 261880 16920 261885
rect 16720 261835 16760 261840
rect 16720 261805 16725 261835
rect 16755 261805 16760 261835
rect 16720 261800 16760 261805
rect 16880 261835 16920 261840
rect 16880 261805 16885 261835
rect 16915 261805 16920 261835
rect 16880 261800 16920 261805
rect 16720 261755 16760 261760
rect 16720 261725 16725 261755
rect 16755 261725 16760 261755
rect 16720 261720 16760 261725
rect 16880 261755 16920 261760
rect 16880 261725 16885 261755
rect 16915 261725 16920 261755
rect 16880 261720 16920 261725
rect 16720 261675 16760 261680
rect 16720 261645 16725 261675
rect 16755 261645 16760 261675
rect 16720 261640 16760 261645
rect 16880 261675 16920 261680
rect 16880 261645 16885 261675
rect 16915 261645 16920 261675
rect 16880 261640 16920 261645
rect 16720 261595 16760 261600
rect 16720 261565 16725 261595
rect 16755 261565 16760 261595
rect 16720 261560 16760 261565
rect 16880 261595 16920 261600
rect 16880 261565 16885 261595
rect 16915 261565 16920 261595
rect 16880 261560 16920 261565
rect 16720 261515 16760 261520
rect 16720 261485 16725 261515
rect 16755 261485 16760 261515
rect 16720 261480 16760 261485
rect 16880 261515 16920 261520
rect 16880 261485 16885 261515
rect 16915 261485 16920 261515
rect 16880 261480 16920 261485
rect 16720 261435 16760 261440
rect 16720 261405 16725 261435
rect 16755 261405 16760 261435
rect 16720 261400 16760 261405
rect 16880 261435 16920 261440
rect 16880 261405 16885 261435
rect 16915 261405 16920 261435
rect 16880 261400 16920 261405
rect 16720 261355 16760 261360
rect 16720 261325 16725 261355
rect 16755 261325 16760 261355
rect 16720 261320 16760 261325
rect 16880 261355 16920 261360
rect 16880 261325 16885 261355
rect 16915 261325 16920 261355
rect 16880 261320 16920 261325
rect 16720 261275 16760 261280
rect 16720 261245 16725 261275
rect 16755 261245 16760 261275
rect 16720 261240 16760 261245
rect 16880 261275 16920 261280
rect 16880 261245 16885 261275
rect 16915 261245 16920 261275
rect 16880 261240 16920 261245
rect 16720 261195 16760 261200
rect 16720 261165 16725 261195
rect 16755 261165 16760 261195
rect 16720 261160 16760 261165
rect 16880 261195 16920 261200
rect 16880 261165 16885 261195
rect 16915 261165 16920 261195
rect 16880 261160 16920 261165
rect 16720 261115 16760 261120
rect 16720 261085 16725 261115
rect 16755 261085 16760 261115
rect 16720 261080 16760 261085
rect 16880 261115 16920 261120
rect 16880 261085 16885 261115
rect 16915 261085 16920 261115
rect 16880 261080 16920 261085
rect 16720 261035 16760 261040
rect 16720 261005 16725 261035
rect 16755 261005 16760 261035
rect 16720 261000 16760 261005
rect 16880 261035 16920 261040
rect 16880 261005 16885 261035
rect 16915 261005 16920 261035
rect 16880 261000 16920 261005
rect 16720 260955 16760 260960
rect 16720 260925 16725 260955
rect 16755 260925 16760 260955
rect 16720 260920 16760 260925
rect 16880 260955 16920 260960
rect 16880 260925 16885 260955
rect 16915 260925 16920 260955
rect 16880 260920 16920 260925
rect 16720 260875 16760 260880
rect 16720 260845 16725 260875
rect 16755 260845 16760 260875
rect 16720 260840 16760 260845
rect 16880 260875 16920 260880
rect 16880 260845 16885 260875
rect 16915 260845 16920 260875
rect 16880 260840 16920 260845
rect 16720 260795 16760 260800
rect 16720 260765 16725 260795
rect 16755 260765 16760 260795
rect 16720 260760 16760 260765
rect 16880 260795 16920 260800
rect 16880 260765 16885 260795
rect 16915 260765 16920 260795
rect 16880 260760 16920 260765
rect 16720 260715 16760 260720
rect 16720 260685 16725 260715
rect 16755 260685 16760 260715
rect 16720 260680 16760 260685
rect 16880 260715 16920 260720
rect 16880 260685 16885 260715
rect 16915 260685 16920 260715
rect 16880 260680 16920 260685
rect 16720 260635 16760 260640
rect 16720 260605 16725 260635
rect 16755 260605 16760 260635
rect 16720 260600 16760 260605
rect 16880 260635 16920 260640
rect 16880 260605 16885 260635
rect 16915 260605 16920 260635
rect 16880 260600 16920 260605
rect 16720 260555 16760 260560
rect 16720 260525 16725 260555
rect 16755 260525 16760 260555
rect 16720 260520 16760 260525
rect 16880 260555 16920 260560
rect 16880 260525 16885 260555
rect 16915 260525 16920 260555
rect 16880 260520 16920 260525
rect 16720 260475 16760 260480
rect 16720 260445 16725 260475
rect 16755 260445 16760 260475
rect 16720 260440 16760 260445
rect 16880 260475 16920 260480
rect 16880 260445 16885 260475
rect 16915 260445 16920 260475
rect 16880 260440 16920 260445
rect 16720 260395 16760 260400
rect 16720 260365 16725 260395
rect 16755 260365 16760 260395
rect 16720 260360 16760 260365
rect 16880 260395 16920 260400
rect 16880 260365 16885 260395
rect 16915 260365 16920 260395
rect 16880 260360 16920 260365
rect 16720 260315 16760 260320
rect 16720 260285 16725 260315
rect 16755 260285 16760 260315
rect 16720 260280 16760 260285
rect 16880 260315 16920 260320
rect 16880 260285 16885 260315
rect 16915 260285 16920 260315
rect 16880 260280 16920 260285
rect 16720 260235 16760 260240
rect 16720 260205 16725 260235
rect 16755 260205 16760 260235
rect 16720 260200 16760 260205
rect 16880 260235 16920 260240
rect 16880 260205 16885 260235
rect 16915 260205 16920 260235
rect 16880 260200 16920 260205
rect 16720 260155 16760 260160
rect 16720 260125 16725 260155
rect 16755 260125 16760 260155
rect 16720 260120 16760 260125
rect 16880 260155 16920 260160
rect 16880 260125 16885 260155
rect 16915 260125 16920 260155
rect 16880 260120 16920 260125
rect 16720 260075 16760 260080
rect 16720 260045 16725 260075
rect 16755 260045 16760 260075
rect 16720 260040 16760 260045
rect 16880 260075 16920 260080
rect 16880 260045 16885 260075
rect 16915 260045 16920 260075
rect 16880 260040 16920 260045
rect 16720 259995 16760 260000
rect 16720 259965 16725 259995
rect 16755 259965 16760 259995
rect 16720 259960 16760 259965
rect 16880 259995 16920 260000
rect 16880 259965 16885 259995
rect 16915 259965 16920 259995
rect 16880 259960 16920 259965
rect 16720 259915 16760 259920
rect 16720 259885 16725 259915
rect 16755 259885 16760 259915
rect 16720 259880 16760 259885
rect 16880 259915 16920 259920
rect 16880 259885 16885 259915
rect 16915 259885 16920 259915
rect 16880 259880 16920 259885
rect 16720 259835 16760 259840
rect 16720 259805 16725 259835
rect 16755 259805 16760 259835
rect 16720 259800 16760 259805
rect 16880 259835 16920 259840
rect 16880 259805 16885 259835
rect 16915 259805 16920 259835
rect 16880 259800 16920 259805
rect 16720 259755 16760 259760
rect 16720 259725 16725 259755
rect 16755 259725 16760 259755
rect 16720 259720 16760 259725
rect 16880 259755 16920 259760
rect 16880 259725 16885 259755
rect 16915 259725 16920 259755
rect 16880 259720 16920 259725
rect 16720 259675 16760 259680
rect 16720 259645 16725 259675
rect 16755 259645 16760 259675
rect 16720 259640 16760 259645
rect 16880 259675 16920 259680
rect 16880 259645 16885 259675
rect 16915 259645 16920 259675
rect 16880 259640 16920 259645
rect 16720 259595 16760 259600
rect 16720 259565 16725 259595
rect 16755 259565 16760 259595
rect 16720 259560 16760 259565
rect 16880 259595 16920 259600
rect 16880 259565 16885 259595
rect 16915 259565 16920 259595
rect 16880 259560 16920 259565
rect 16720 259515 16760 259520
rect 16720 259485 16725 259515
rect 16755 259485 16760 259515
rect 16720 259480 16760 259485
rect 16880 259515 16920 259520
rect 16880 259485 16885 259515
rect 16915 259485 16920 259515
rect 16880 259480 16920 259485
rect 16720 259435 16760 259440
rect 16720 259405 16725 259435
rect 16755 259405 16760 259435
rect 16720 259400 16760 259405
rect 16880 259435 16920 259440
rect 16880 259405 16885 259435
rect 16915 259405 16920 259435
rect 16880 259400 16920 259405
rect 16720 259355 16760 259360
rect 16720 259325 16725 259355
rect 16755 259325 16760 259355
rect 16720 259320 16760 259325
rect 16880 259355 16920 259360
rect 16880 259325 16885 259355
rect 16915 259325 16920 259355
rect 16880 259320 16920 259325
rect 16720 259275 16760 259280
rect 16720 259245 16725 259275
rect 16755 259245 16760 259275
rect 16720 259240 16760 259245
rect 16880 259275 16920 259280
rect 16880 259245 16885 259275
rect 16915 259245 16920 259275
rect 16880 259240 16920 259245
rect 16720 259195 16760 259200
rect 16720 259165 16725 259195
rect 16755 259165 16760 259195
rect 16720 259160 16760 259165
rect 16880 259195 16920 259200
rect 16880 259165 16885 259195
rect 16915 259165 16920 259195
rect 16880 259160 16920 259165
rect 16720 259115 16760 259120
rect 16720 259085 16725 259115
rect 16755 259085 16760 259115
rect 16720 259080 16760 259085
rect 16880 259115 16920 259120
rect 16880 259085 16885 259115
rect 16915 259085 16920 259115
rect 16880 259080 16920 259085
rect 16720 259035 16760 259040
rect 16720 259005 16725 259035
rect 16755 259005 16760 259035
rect 16720 259000 16760 259005
rect 16880 259035 16920 259040
rect 16880 259005 16885 259035
rect 16915 259005 16920 259035
rect 16880 259000 16920 259005
rect 16720 258955 16760 258960
rect 16720 258925 16725 258955
rect 16755 258925 16760 258955
rect 16720 258920 16760 258925
rect 16880 258955 16920 258960
rect 16880 258925 16885 258955
rect 16915 258925 16920 258955
rect 16880 258920 16920 258925
rect 16720 258875 16760 258880
rect 16720 258845 16725 258875
rect 16755 258845 16760 258875
rect 16720 258840 16760 258845
rect 16880 258875 16920 258880
rect 16880 258845 16885 258875
rect 16915 258845 16920 258875
rect 16880 258840 16920 258845
rect 16720 258795 16760 258800
rect 16720 258765 16725 258795
rect 16755 258765 16760 258795
rect 16720 258760 16760 258765
rect 16880 258795 16920 258800
rect 16880 258765 16885 258795
rect 16915 258765 16920 258795
rect 16880 258760 16920 258765
rect 16720 258715 16760 258720
rect 16720 258685 16725 258715
rect 16755 258685 16760 258715
rect 16720 258680 16760 258685
rect 16880 258715 16920 258720
rect 16880 258685 16885 258715
rect 16915 258685 16920 258715
rect 16880 258680 16920 258685
rect 16720 258635 16760 258640
rect 16720 258605 16725 258635
rect 16755 258605 16760 258635
rect 16720 258600 16760 258605
rect 16880 258635 16920 258640
rect 16880 258605 16885 258635
rect 16915 258605 16920 258635
rect 16880 258600 16920 258605
rect 16720 258555 16760 258560
rect 16720 258525 16725 258555
rect 16755 258525 16760 258555
rect 16720 258520 16760 258525
rect 16880 258555 16920 258560
rect 16880 258525 16885 258555
rect 16915 258525 16920 258555
rect 16880 258520 16920 258525
rect 16720 258475 16760 258480
rect 16720 258445 16725 258475
rect 16755 258445 16760 258475
rect 16720 258440 16760 258445
rect 16880 258475 16920 258480
rect 16880 258445 16885 258475
rect 16915 258445 16920 258475
rect 16880 258440 16920 258445
rect 16720 258395 16760 258400
rect 16720 258365 16725 258395
rect 16755 258365 16760 258395
rect 16720 258360 16760 258365
rect 16880 258395 16920 258400
rect 16880 258365 16885 258395
rect 16915 258365 16920 258395
rect 16880 258360 16920 258365
rect 16720 258315 16760 258320
rect 16720 258285 16725 258315
rect 16755 258285 16760 258315
rect 16720 258280 16760 258285
rect 16880 258315 16920 258320
rect 16880 258285 16885 258315
rect 16915 258285 16920 258315
rect 16880 258280 16920 258285
rect 16720 258235 16760 258240
rect 16720 258205 16725 258235
rect 16755 258205 16760 258235
rect 16720 258200 16760 258205
rect 16880 258235 16920 258240
rect 16880 258205 16885 258235
rect 16915 258205 16920 258235
rect 16880 258200 16920 258205
rect 16720 258155 16760 258160
rect 16720 258125 16725 258155
rect 16755 258125 16760 258155
rect 16720 258120 16760 258125
rect 16880 258155 16920 258160
rect 16880 258125 16885 258155
rect 16915 258125 16920 258155
rect 16880 258120 16920 258125
rect 16720 258075 16760 258080
rect 16720 258045 16725 258075
rect 16755 258045 16760 258075
rect 16720 258040 16760 258045
rect 16880 258075 16920 258080
rect 16880 258045 16885 258075
rect 16915 258045 16920 258075
rect 16880 258040 16920 258045
rect 16720 257995 16760 258000
rect 16720 257965 16725 257995
rect 16755 257965 16760 257995
rect 16720 257960 16760 257965
rect 16880 257995 16920 258000
rect 16880 257965 16885 257995
rect 16915 257965 16920 257995
rect 16880 257960 16920 257965
rect 16720 257915 16760 257920
rect 16720 257885 16725 257915
rect 16755 257885 16760 257915
rect 16720 257880 16760 257885
rect 16880 257915 16920 257920
rect 16880 257885 16885 257915
rect 16915 257885 16920 257915
rect 16880 257880 16920 257885
rect 16720 257835 16760 257840
rect 16720 257805 16725 257835
rect 16755 257805 16760 257835
rect 16720 257800 16760 257805
rect 16880 257835 16920 257840
rect 16880 257805 16885 257835
rect 16915 257805 16920 257835
rect 16880 257800 16920 257805
rect 16720 257755 16760 257760
rect 16720 257725 16725 257755
rect 16755 257725 16760 257755
rect 16720 257720 16760 257725
rect 16880 257755 16920 257760
rect 16880 257725 16885 257755
rect 16915 257725 16920 257755
rect 16880 257720 16920 257725
rect 16720 257675 16760 257680
rect 16720 257645 16725 257675
rect 16755 257645 16760 257675
rect 16720 257640 16760 257645
rect 16880 257675 16920 257680
rect 16880 257645 16885 257675
rect 16915 257645 16920 257675
rect 16880 257640 16920 257645
rect 16720 257595 16760 257600
rect 16720 257565 16725 257595
rect 16755 257565 16760 257595
rect 16720 257560 16760 257565
rect 16880 257595 16920 257600
rect 16880 257565 16885 257595
rect 16915 257565 16920 257595
rect 16880 257560 16920 257565
rect 16720 257515 16760 257520
rect 16720 257485 16725 257515
rect 16755 257485 16760 257515
rect 16720 257480 16760 257485
rect 16880 257515 16920 257520
rect 16880 257485 16885 257515
rect 16915 257485 16920 257515
rect 16880 257480 16920 257485
rect 16720 257435 16760 257440
rect 16720 257405 16725 257435
rect 16755 257405 16760 257435
rect 16720 257400 16760 257405
rect 16880 257435 16920 257440
rect 16880 257405 16885 257435
rect 16915 257405 16920 257435
rect 16880 257400 16920 257405
rect 16720 257355 16760 257360
rect 16720 257325 16725 257355
rect 16755 257325 16760 257355
rect 16720 257320 16760 257325
rect 16880 257355 16920 257360
rect 16880 257325 16885 257355
rect 16915 257325 16920 257355
rect 16880 257320 16920 257325
rect 16720 257275 16760 257280
rect 16720 257245 16725 257275
rect 16755 257245 16760 257275
rect 16720 257240 16760 257245
rect 16880 257275 16920 257280
rect 16880 257245 16885 257275
rect 16915 257245 16920 257275
rect 16880 257240 16920 257245
rect 16720 257195 16760 257200
rect 16720 257165 16725 257195
rect 16755 257165 16760 257195
rect 16720 257160 16760 257165
rect 16880 257195 16920 257200
rect 16880 257165 16885 257195
rect 16915 257165 16920 257195
rect 16880 257160 16920 257165
rect 16720 257115 16760 257120
rect 16720 257085 16725 257115
rect 16755 257085 16760 257115
rect 16720 257080 16760 257085
rect 16880 257115 16920 257120
rect 16880 257085 16885 257115
rect 16915 257085 16920 257115
rect 16880 257080 16920 257085
rect 16720 257035 16760 257040
rect 16720 257005 16725 257035
rect 16755 257005 16760 257035
rect 16720 257000 16760 257005
rect 16880 257035 16920 257040
rect 16880 257005 16885 257035
rect 16915 257005 16920 257035
rect 16880 257000 16920 257005
rect 16720 256955 16760 256960
rect 16720 256925 16725 256955
rect 16755 256925 16760 256955
rect 16720 256920 16760 256925
rect 16880 256955 16920 256960
rect 16880 256925 16885 256955
rect 16915 256925 16920 256955
rect 16880 256920 16920 256925
rect 16720 256875 16760 256880
rect 16720 256845 16725 256875
rect 16755 256845 16760 256875
rect 16720 256840 16760 256845
rect 16880 256875 16920 256880
rect 16880 256845 16885 256875
rect 16915 256845 16920 256875
rect 16880 256840 16920 256845
rect 16720 256795 16760 256800
rect 16720 256765 16725 256795
rect 16755 256765 16760 256795
rect 16720 256760 16760 256765
rect 16880 256795 16920 256800
rect 16880 256765 16885 256795
rect 16915 256765 16920 256795
rect 16880 256760 16920 256765
rect 16720 256715 16760 256720
rect 16720 256685 16725 256715
rect 16755 256685 16760 256715
rect 16720 256680 16760 256685
rect 16880 256715 16920 256720
rect 16880 256685 16885 256715
rect 16915 256685 16920 256715
rect 16880 256680 16920 256685
rect 16720 256635 16760 256640
rect 16720 256605 16725 256635
rect 16755 256605 16760 256635
rect 16720 256600 16760 256605
rect 16880 256635 16920 256640
rect 16880 256605 16885 256635
rect 16915 256605 16920 256635
rect 16880 256600 16920 256605
rect 16720 256555 16760 256560
rect 16720 256525 16725 256555
rect 16755 256525 16760 256555
rect 16720 256520 16760 256525
rect 16880 256555 16920 256560
rect 16880 256525 16885 256555
rect 16915 256525 16920 256555
rect 16880 256520 16920 256525
rect 16720 256475 16760 256480
rect 16720 256445 16725 256475
rect 16755 256445 16760 256475
rect 16720 256440 16760 256445
rect 16880 256475 16920 256480
rect 16880 256445 16885 256475
rect 16915 256445 16920 256475
rect 16880 256440 16920 256445
rect 16720 256395 16760 256400
rect 16720 256365 16725 256395
rect 16755 256365 16760 256395
rect 16720 256360 16760 256365
rect 16880 256395 16920 256400
rect 16880 256365 16885 256395
rect 16915 256365 16920 256395
rect 16880 256360 16920 256365
rect 16720 256315 16760 256320
rect 16720 256285 16725 256315
rect 16755 256285 16760 256315
rect 16720 256280 16760 256285
rect 16880 256315 16920 256320
rect 16880 256285 16885 256315
rect 16915 256285 16920 256315
rect 16880 256280 16920 256285
rect 16720 256235 16760 256240
rect 16720 256205 16725 256235
rect 16755 256205 16760 256235
rect 16720 256200 16760 256205
rect 16880 256235 16920 256240
rect 16880 256205 16885 256235
rect 16915 256205 16920 256235
rect 16880 256200 16920 256205
rect 16720 256155 16760 256160
rect 16720 256125 16725 256155
rect 16755 256125 16760 256155
rect 16720 256120 16760 256125
rect 16880 256155 16920 256160
rect 16880 256125 16885 256155
rect 16915 256125 16920 256155
rect 16880 256120 16920 256125
rect 16720 256075 16760 256080
rect 16720 256045 16725 256075
rect 16755 256045 16760 256075
rect 16720 256040 16760 256045
rect 16880 256075 16920 256080
rect 16880 256045 16885 256075
rect 16915 256045 16920 256075
rect 16880 256040 16920 256045
rect 16720 255995 16760 256000
rect 16720 255965 16725 255995
rect 16755 255965 16760 255995
rect 16720 255960 16760 255965
rect 16880 255995 16920 256000
rect 16880 255965 16885 255995
rect 16915 255965 16920 255995
rect 16880 255960 16920 255965
rect 400 255875 440 255880
rect 400 255845 405 255875
rect 435 255845 440 255875
rect 400 255840 440 255845
rect 480 255875 520 255880
rect 480 255845 485 255875
rect 515 255845 520 255875
rect 480 255840 520 255845
rect 560 255875 600 255880
rect 560 255845 565 255875
rect 595 255845 600 255875
rect 560 255840 600 255845
rect 640 255875 680 255880
rect 640 255845 645 255875
rect 675 255845 680 255875
rect 640 255840 680 255845
rect 720 255875 760 255880
rect 720 255845 725 255875
rect 755 255845 760 255875
rect 720 255840 760 255845
rect 800 255875 840 255880
rect 800 255845 805 255875
rect 835 255845 840 255875
rect 800 255840 840 255845
rect 880 255875 920 255880
rect 880 255845 885 255875
rect 915 255845 920 255875
rect 880 255840 920 255845
rect 960 255875 1000 255880
rect 960 255845 965 255875
rect 995 255845 1000 255875
rect 960 255840 1000 255845
rect 1040 255875 1080 255880
rect 1040 255845 1045 255875
rect 1075 255845 1080 255875
rect 1040 255840 1080 255845
rect 1120 255875 1160 255880
rect 1120 255845 1125 255875
rect 1155 255845 1160 255875
rect 1120 255840 1160 255845
rect 1200 255875 1240 255880
rect 1200 255845 1205 255875
rect 1235 255845 1240 255875
rect 1200 255840 1240 255845
rect 1280 255875 1320 255880
rect 1280 255845 1285 255875
rect 1315 255845 1320 255875
rect 1280 255840 1320 255845
rect 1360 255875 1400 255880
rect 1360 255845 1365 255875
rect 1395 255845 1400 255875
rect 1360 255840 1400 255845
rect 1440 255875 1480 255880
rect 1440 255845 1445 255875
rect 1475 255845 1480 255875
rect 1440 255840 1480 255845
rect 1520 255875 1560 255880
rect 1520 255845 1525 255875
rect 1555 255845 1560 255875
rect 1520 255840 1560 255845
rect 1600 255875 1640 255880
rect 1600 255845 1605 255875
rect 1635 255845 1640 255875
rect 1600 255840 1640 255845
rect 1680 255875 1720 255880
rect 1680 255845 1685 255875
rect 1715 255845 1720 255875
rect 1680 255840 1720 255845
rect 1760 255875 1800 255880
rect 1760 255845 1765 255875
rect 1795 255845 1800 255875
rect 1760 255840 1800 255845
rect 1840 255875 1880 255880
rect 1840 255845 1845 255875
rect 1875 255845 1880 255875
rect 1840 255840 1880 255845
rect 1920 255875 1960 255880
rect 1920 255845 1925 255875
rect 1955 255845 1960 255875
rect 1920 255840 1960 255845
rect 2000 255875 2040 255880
rect 2000 255845 2005 255875
rect 2035 255845 2040 255875
rect 2000 255840 2040 255845
rect 2080 255875 2120 255880
rect 2080 255845 2085 255875
rect 2115 255845 2120 255875
rect 2080 255840 2120 255845
rect 2160 255875 2200 255880
rect 2160 255845 2165 255875
rect 2195 255845 2200 255875
rect 2160 255840 2200 255845
rect 2240 255875 2280 255880
rect 2240 255845 2245 255875
rect 2275 255845 2280 255875
rect 2240 255840 2280 255845
rect 2320 255875 2360 255880
rect 2320 255845 2325 255875
rect 2355 255845 2360 255875
rect 2320 255840 2360 255845
rect 2400 255875 2440 255880
rect 2400 255845 2405 255875
rect 2435 255845 2440 255875
rect 2400 255840 2440 255845
rect 2480 255875 2520 255880
rect 2480 255845 2485 255875
rect 2515 255845 2520 255875
rect 2480 255840 2520 255845
rect 2560 255875 2600 255880
rect 2560 255845 2565 255875
rect 2595 255845 2600 255875
rect 2560 255840 2600 255845
rect 2640 255875 2680 255880
rect 2640 255845 2645 255875
rect 2675 255845 2680 255875
rect 2640 255840 2680 255845
rect 2720 255875 2760 255880
rect 2720 255845 2725 255875
rect 2755 255845 2760 255875
rect 2720 255840 2760 255845
rect 3040 255875 3080 255880
rect 3040 255845 3045 255875
rect 3075 255845 3080 255875
rect 3040 255840 3080 255845
rect 3120 255875 3160 255880
rect 3120 255845 3125 255875
rect 3155 255845 3160 255875
rect 3120 255840 3160 255845
rect 3200 255875 3240 255880
rect 3200 255845 3205 255875
rect 3235 255845 3240 255875
rect 3200 255840 3240 255845
rect 3280 255875 3320 255880
rect 3280 255845 3285 255875
rect 3315 255845 3320 255875
rect 3280 255840 3320 255845
rect 3360 255875 3400 255880
rect 3360 255845 3365 255875
rect 3395 255845 3400 255875
rect 3360 255840 3400 255845
rect 3440 255875 3480 255880
rect 3440 255845 3445 255875
rect 3475 255845 3480 255875
rect 3440 255840 3480 255845
rect 3520 255875 3560 255880
rect 3520 255845 3525 255875
rect 3555 255845 3560 255875
rect 3520 255840 3560 255845
rect 3600 255875 3640 255880
rect 3600 255845 3605 255875
rect 3635 255845 3640 255875
rect 3600 255840 3640 255845
rect 3680 255875 3720 255880
rect 3680 255845 3685 255875
rect 3715 255845 3720 255875
rect 3680 255840 3720 255845
rect 3760 255875 3800 255880
rect 3760 255845 3765 255875
rect 3795 255845 3800 255875
rect 3760 255840 3800 255845
rect 3840 255875 3880 255880
rect 3840 255845 3845 255875
rect 3875 255845 3880 255875
rect 3840 255840 3880 255845
rect 3920 255875 3960 255880
rect 3920 255845 3925 255875
rect 3955 255845 3960 255875
rect 3920 255840 3960 255845
rect 4000 255875 4040 255880
rect 4000 255845 4005 255875
rect 4035 255845 4040 255875
rect 4000 255840 4040 255845
rect 4080 255875 4120 255880
rect 4080 255845 4085 255875
rect 4115 255845 4120 255875
rect 4080 255840 4120 255845
rect 4160 255875 4200 255880
rect 4160 255845 4165 255875
rect 4195 255845 4200 255875
rect 4160 255840 4200 255845
rect 4240 255875 4280 255880
rect 4240 255845 4245 255875
rect 4275 255845 4280 255875
rect 4240 255840 4280 255845
rect 4320 255875 4360 255880
rect 4320 255845 4325 255875
rect 4355 255845 4360 255875
rect 4320 255840 4360 255845
rect 4400 255875 4440 255880
rect 4400 255845 4405 255875
rect 4435 255845 4440 255875
rect 4400 255840 4440 255845
rect 4480 255875 4520 255880
rect 4480 255845 4485 255875
rect 4515 255845 4520 255875
rect 4480 255840 4520 255845
rect 4560 255875 4600 255880
rect 4560 255845 4565 255875
rect 4595 255845 4600 255875
rect 4560 255840 4600 255845
rect 4640 255875 4680 255880
rect 4640 255845 4645 255875
rect 4675 255845 4680 255875
rect 4640 255840 4680 255845
rect 4720 255875 4760 255880
rect 4720 255845 4725 255875
rect 4755 255845 4760 255875
rect 4720 255840 4760 255845
rect 4800 255875 4840 255880
rect 4800 255845 4805 255875
rect 4835 255845 4840 255875
rect 4800 255840 4840 255845
rect 4880 255875 4920 255880
rect 4880 255845 4885 255875
rect 4915 255845 4920 255875
rect 4880 255840 4920 255845
rect 4960 255875 5000 255880
rect 4960 255845 4965 255875
rect 4995 255845 5000 255875
rect 4960 255840 5000 255845
rect 5040 255875 5080 255880
rect 5040 255845 5045 255875
rect 5075 255845 5080 255875
rect 5040 255840 5080 255845
rect 5120 255875 5160 255880
rect 5120 255845 5125 255875
rect 5155 255845 5160 255875
rect 5120 255840 5160 255845
rect 5200 255875 5240 255880
rect 5200 255845 5205 255875
rect 5235 255845 5240 255875
rect 5200 255840 5240 255845
rect 5280 255875 5320 255880
rect 5280 255845 5285 255875
rect 5315 255845 5320 255875
rect 5280 255840 5320 255845
rect 5360 255875 5400 255880
rect 5360 255845 5365 255875
rect 5395 255845 5400 255875
rect 5360 255840 5400 255845
rect 5440 255875 5480 255880
rect 5440 255845 5445 255875
rect 5475 255845 5480 255875
rect 5440 255840 5480 255845
rect 5520 255875 5560 255880
rect 5520 255845 5525 255875
rect 5555 255845 5560 255875
rect 5520 255840 5560 255845
rect 5600 255875 5640 255880
rect 5600 255845 5605 255875
rect 5635 255845 5640 255875
rect 5600 255840 5640 255845
rect 5680 255875 5720 255880
rect 5680 255845 5685 255875
rect 5715 255845 5720 255875
rect 5680 255840 5720 255845
rect 5760 255875 5800 255880
rect 5760 255845 5765 255875
rect 5795 255845 5800 255875
rect 5760 255840 5800 255845
rect 5840 255875 5880 255880
rect 5840 255845 5845 255875
rect 5875 255845 5880 255875
rect 5840 255840 5880 255845
rect 5920 255875 5960 255880
rect 5920 255845 5925 255875
rect 5955 255845 5960 255875
rect 5920 255840 5960 255845
rect 6000 255875 6040 255880
rect 6000 255845 6005 255875
rect 6035 255845 6040 255875
rect 6000 255840 6040 255845
rect 6080 255875 6120 255880
rect 6080 255845 6085 255875
rect 6115 255845 6120 255875
rect 6080 255840 6120 255845
rect 6160 255875 6200 255880
rect 6160 255845 6165 255875
rect 6195 255845 6200 255875
rect 6160 255840 6200 255845
rect 6240 255875 6280 255880
rect 6240 255845 6245 255875
rect 6275 255845 6280 255875
rect 6240 255840 6280 255845
rect 6320 255875 6360 255880
rect 6320 255845 6325 255875
rect 6355 255845 6360 255875
rect 6320 255840 6360 255845
rect 6400 255875 6440 255880
rect 6400 255845 6405 255875
rect 6435 255845 6440 255875
rect 6400 255840 6440 255845
rect 6480 255875 6520 255880
rect 6480 255845 6485 255875
rect 6515 255845 6520 255875
rect 6480 255840 6520 255845
rect 6560 255875 6600 255880
rect 6560 255845 6565 255875
rect 6595 255845 6600 255875
rect 6560 255840 6600 255845
rect 6640 255875 6680 255880
rect 6640 255845 6645 255875
rect 6675 255845 6680 255875
rect 6640 255840 6680 255845
rect 6720 255875 6760 255880
rect 6720 255845 6725 255875
rect 6755 255845 6760 255875
rect 6720 255840 6760 255845
rect 6800 255875 6840 255880
rect 6800 255845 6805 255875
rect 6835 255845 6840 255875
rect 6800 255840 6840 255845
rect 6880 255875 6920 255880
rect 6880 255845 6885 255875
rect 6915 255845 6920 255875
rect 6880 255840 6920 255845
rect 6960 255875 7000 255880
rect 6960 255845 6965 255875
rect 6995 255845 7000 255875
rect 6960 255840 7000 255845
rect 7040 255875 7080 255880
rect 7040 255845 7045 255875
rect 7075 255845 7080 255875
rect 7040 255840 7080 255845
rect 7120 255875 7160 255880
rect 7120 255845 7125 255875
rect 7155 255845 7160 255875
rect 7120 255840 7160 255845
rect 7200 255875 7240 255880
rect 7200 255845 7205 255875
rect 7235 255845 7240 255875
rect 7200 255840 7240 255845
rect 7280 255875 7320 255880
rect 7280 255845 7285 255875
rect 7315 255845 7320 255875
rect 7280 255840 7320 255845
rect 7360 255875 7400 255880
rect 7360 255845 7365 255875
rect 7395 255845 7400 255875
rect 7360 255840 7400 255845
rect 7440 255875 7480 255880
rect 7440 255845 7445 255875
rect 7475 255845 7480 255875
rect 7440 255840 7480 255845
rect 7520 255875 7560 255880
rect 7520 255845 7525 255875
rect 7555 255845 7560 255875
rect 7520 255840 7560 255845
rect 7600 255875 7640 255880
rect 7600 255845 7605 255875
rect 7635 255845 7640 255875
rect 7600 255840 7640 255845
rect 7680 255875 7720 255880
rect 7680 255845 7685 255875
rect 7715 255845 7720 255875
rect 7680 255840 7720 255845
rect 7760 255875 7800 255880
rect 7760 255845 7765 255875
rect 7795 255845 7800 255875
rect 7760 255840 7800 255845
rect 7840 255875 7880 255880
rect 7840 255845 7845 255875
rect 7875 255845 7880 255875
rect 7840 255840 7880 255845
rect 7920 255875 7960 255880
rect 7920 255845 7925 255875
rect 7955 255845 7960 255875
rect 7920 255840 7960 255845
rect 8000 255875 8040 255880
rect 8000 255845 8005 255875
rect 8035 255845 8040 255875
rect 8000 255840 8040 255845
rect 8080 255875 8120 255880
rect 8080 255845 8085 255875
rect 8115 255845 8120 255875
rect 8080 255840 8120 255845
rect 8160 255875 8200 255880
rect 8160 255845 8165 255875
rect 8195 255845 8200 255875
rect 8160 255840 8200 255845
rect 8240 255875 8280 255880
rect 8240 255845 8245 255875
rect 8275 255845 8280 255875
rect 8240 255840 8280 255845
rect 8320 255875 8360 255880
rect 8320 255845 8325 255875
rect 8355 255845 8360 255875
rect 8320 255840 8360 255845
rect 8400 255875 8440 255880
rect 8400 255845 8405 255875
rect 8435 255845 8440 255875
rect 8400 255840 8440 255845
rect 8480 255875 8520 255880
rect 8480 255845 8485 255875
rect 8515 255845 8520 255875
rect 8480 255840 8520 255845
rect 8560 255875 8600 255880
rect 8560 255845 8565 255875
rect 8595 255845 8600 255875
rect 8560 255840 8600 255845
rect 8640 255875 8680 255880
rect 8640 255845 8645 255875
rect 8675 255845 8680 255875
rect 8640 255840 8680 255845
rect 8720 255875 8760 255880
rect 8720 255845 8725 255875
rect 8755 255845 8760 255875
rect 8720 255840 8760 255845
rect 8800 255875 8840 255880
rect 8800 255845 8805 255875
rect 8835 255845 8840 255875
rect 8800 255840 8840 255845
rect 8880 255875 8920 255880
rect 8880 255845 8885 255875
rect 8915 255845 8920 255875
rect 8880 255840 8920 255845
rect 8960 255875 9000 255880
rect 8960 255845 8965 255875
rect 8995 255845 9000 255875
rect 8960 255840 9000 255845
rect 9040 255875 9080 255880
rect 9040 255845 9045 255875
rect 9075 255845 9080 255875
rect 9040 255840 9080 255845
rect 9120 255875 9160 255880
rect 9120 255845 9125 255875
rect 9155 255845 9160 255875
rect 9120 255840 9160 255845
rect 9200 255875 9240 255880
rect 9200 255845 9205 255875
rect 9235 255845 9240 255875
rect 9200 255840 9240 255845
rect 9280 255875 9320 255880
rect 9280 255845 9285 255875
rect 9315 255845 9320 255875
rect 9280 255840 9320 255845
rect 9360 255875 9400 255880
rect 9360 255845 9365 255875
rect 9395 255845 9400 255875
rect 9360 255840 9400 255845
rect 9440 255875 9480 255880
rect 9440 255845 9445 255875
rect 9475 255845 9480 255875
rect 9440 255840 9480 255845
rect 9520 255875 9560 255880
rect 9520 255845 9525 255875
rect 9555 255845 9560 255875
rect 9520 255840 9560 255845
rect 9600 255875 9640 255880
rect 9600 255845 9605 255875
rect 9635 255845 9640 255875
rect 9600 255840 9640 255845
rect 9680 255875 9720 255880
rect 9680 255845 9685 255875
rect 9715 255845 9720 255875
rect 9680 255840 9720 255845
rect 9760 255875 9800 255880
rect 9760 255845 9765 255875
rect 9795 255845 9800 255875
rect 9760 255840 9800 255845
rect 9840 255875 9880 255880
rect 9840 255845 9845 255875
rect 9875 255845 9880 255875
rect 9840 255840 9880 255845
rect 9920 255875 9960 255880
rect 9920 255845 9925 255875
rect 9955 255845 9960 255875
rect 9920 255840 9960 255845
rect 10000 255875 10040 255880
rect 10000 255845 10005 255875
rect 10035 255845 10040 255875
rect 10000 255840 10040 255845
rect 10080 255875 10120 255880
rect 10080 255845 10085 255875
rect 10115 255845 10120 255875
rect 10080 255840 10120 255845
rect 10160 255875 10200 255880
rect 10160 255845 10165 255875
rect 10195 255845 10200 255875
rect 10160 255840 10200 255845
rect 10240 255875 10280 255880
rect 10240 255845 10245 255875
rect 10275 255845 10280 255875
rect 10240 255840 10280 255845
rect 10320 255875 10360 255880
rect 10320 255845 10325 255875
rect 10355 255845 10360 255875
rect 10320 255840 10360 255845
rect 10400 255875 10440 255880
rect 10400 255845 10405 255875
rect 10435 255845 10440 255875
rect 10400 255840 10440 255845
rect 10480 255875 10520 255880
rect 10480 255845 10485 255875
rect 10515 255845 10520 255875
rect 10480 255840 10520 255845
rect 10560 255875 10600 255880
rect 10560 255845 10565 255875
rect 10595 255845 10600 255875
rect 10560 255840 10600 255845
rect 10640 255875 10680 255880
rect 10640 255845 10645 255875
rect 10675 255845 10680 255875
rect 10640 255840 10680 255845
rect 10720 255875 10760 255880
rect 10720 255845 10725 255875
rect 10755 255845 10760 255875
rect 10720 255840 10760 255845
rect 10800 255875 10840 255880
rect 10800 255845 10805 255875
rect 10835 255845 10840 255875
rect 10800 255840 10840 255845
rect 10880 255875 10920 255880
rect 10880 255845 10885 255875
rect 10915 255845 10920 255875
rect 10880 255840 10920 255845
rect 10960 255875 11000 255880
rect 10960 255845 10965 255875
rect 10995 255845 11000 255875
rect 10960 255840 11000 255845
rect 11040 255875 11080 255880
rect 11040 255845 11045 255875
rect 11075 255845 11080 255875
rect 11040 255840 11080 255845
rect 11120 255875 11160 255880
rect 11120 255845 11125 255875
rect 11155 255845 11160 255875
rect 11120 255840 11160 255845
rect 11200 255875 11240 255880
rect 11200 255845 11205 255875
rect 11235 255845 11240 255875
rect 11200 255840 11240 255845
rect 11280 255875 11320 255880
rect 11280 255845 11285 255875
rect 11315 255845 11320 255875
rect 11280 255840 11320 255845
rect 11360 255875 11400 255880
rect 11360 255845 11365 255875
rect 11395 255845 11400 255875
rect 11360 255840 11400 255845
rect 11440 255875 11480 255880
rect 11440 255845 11445 255875
rect 11475 255845 11480 255875
rect 11440 255840 11480 255845
rect 11520 255875 11560 255880
rect 11520 255845 11525 255875
rect 11555 255845 11560 255875
rect 11520 255840 11560 255845
rect 11600 255875 11640 255880
rect 11600 255845 11605 255875
rect 11635 255845 11640 255875
rect 11600 255840 11640 255845
rect 11680 255875 11720 255880
rect 11680 255845 11685 255875
rect 11715 255845 11720 255875
rect 11680 255840 11720 255845
rect 11760 255875 11800 255880
rect 11760 255845 11765 255875
rect 11795 255845 11800 255875
rect 11760 255840 11800 255845
rect 11840 255875 11880 255880
rect 11840 255845 11845 255875
rect 11875 255845 11880 255875
rect 11840 255840 11880 255845
rect 11920 255875 11960 255880
rect 11920 255845 11925 255875
rect 11955 255845 11960 255875
rect 11920 255840 11960 255845
rect 12000 255875 12040 255880
rect 12000 255845 12005 255875
rect 12035 255845 12040 255875
rect 12000 255840 12040 255845
rect 12080 255875 12120 255880
rect 12080 255845 12085 255875
rect 12115 255845 12120 255875
rect 12080 255840 12120 255845
rect 12160 255875 12200 255880
rect 12160 255845 12165 255875
rect 12195 255845 12200 255875
rect 12160 255840 12200 255845
rect 12240 255875 12280 255880
rect 12240 255845 12245 255875
rect 12275 255845 12280 255875
rect 12240 255840 12280 255845
rect 12320 255875 12360 255880
rect 12320 255845 12325 255875
rect 12355 255845 12360 255875
rect 12320 255840 12360 255845
rect 12400 255875 12440 255880
rect 12400 255845 12405 255875
rect 12435 255845 12440 255875
rect 12400 255840 12440 255845
rect 12480 255875 12520 255880
rect 12480 255845 12485 255875
rect 12515 255845 12520 255875
rect 12480 255840 12520 255845
rect 12560 255875 12600 255880
rect 12560 255845 12565 255875
rect 12595 255845 12600 255875
rect 12560 255840 12600 255845
rect 12640 255875 12680 255880
rect 12640 255845 12645 255875
rect 12675 255845 12680 255875
rect 12640 255840 12680 255845
rect 12720 255875 12760 255880
rect 12720 255845 12725 255875
rect 12755 255845 12760 255875
rect 12720 255840 12760 255845
rect 12800 255875 12840 255880
rect 12800 255845 12805 255875
rect 12835 255845 12840 255875
rect 12800 255840 12840 255845
rect 12880 255875 12920 255880
rect 12880 255845 12885 255875
rect 12915 255845 12920 255875
rect 12880 255840 12920 255845
rect 12960 255875 13000 255880
rect 12960 255845 12965 255875
rect 12995 255845 13000 255875
rect 12960 255840 13000 255845
rect 13040 255875 13080 255880
rect 13040 255845 13045 255875
rect 13075 255845 13080 255875
rect 13040 255840 13080 255845
rect 13120 255875 13160 255880
rect 13120 255845 13125 255875
rect 13155 255845 13160 255875
rect 13120 255840 13160 255845
rect 13200 255875 13240 255880
rect 13200 255845 13205 255875
rect 13235 255845 13240 255875
rect 13200 255840 13240 255845
rect 13280 255875 13320 255880
rect 13280 255845 13285 255875
rect 13315 255845 13320 255875
rect 13280 255840 13320 255845
rect 13360 255875 13400 255880
rect 13360 255845 13365 255875
rect 13395 255845 13400 255875
rect 13360 255840 13400 255845
rect 13440 255875 13480 255880
rect 13440 255845 13445 255875
rect 13475 255845 13480 255875
rect 13440 255840 13480 255845
rect 13520 255875 13560 255880
rect 13520 255845 13525 255875
rect 13555 255845 13560 255875
rect 13520 255840 13560 255845
rect 13600 255875 13640 255880
rect 13600 255845 13605 255875
rect 13635 255845 13640 255875
rect 13600 255840 13640 255845
rect 13680 255875 13720 255880
rect 13680 255845 13685 255875
rect 13715 255845 13720 255875
rect 13680 255840 13720 255845
rect 13760 255875 13800 255880
rect 13760 255845 13765 255875
rect 13795 255845 13800 255875
rect 13760 255840 13800 255845
rect 13840 255875 13880 255880
rect 13840 255845 13845 255875
rect 13875 255845 13880 255875
rect 13840 255840 13880 255845
rect 13920 255875 13960 255880
rect 13920 255845 13925 255875
rect 13955 255845 13960 255875
rect 13920 255840 13960 255845
rect 14000 255875 14040 255880
rect 14000 255845 14005 255875
rect 14035 255845 14040 255875
rect 14000 255840 14040 255845
rect 14080 255875 14120 255880
rect 14080 255845 14085 255875
rect 14115 255845 14120 255875
rect 14080 255840 14120 255845
rect 14160 255875 14200 255880
rect 14160 255845 14165 255875
rect 14195 255845 14200 255875
rect 14160 255840 14200 255845
rect 14240 255875 14280 255880
rect 14240 255845 14245 255875
rect 14275 255845 14280 255875
rect 14240 255840 14280 255845
rect 14320 255875 14360 255880
rect 14320 255845 14325 255875
rect 14355 255845 14360 255875
rect 14320 255840 14360 255845
rect 14400 255875 14440 255880
rect 14400 255845 14405 255875
rect 14435 255845 14440 255875
rect 14400 255840 14440 255845
rect 14480 255875 14520 255880
rect 14480 255845 14485 255875
rect 14515 255845 14520 255875
rect 14480 255840 14520 255845
rect 14560 255875 14600 255880
rect 14560 255845 14565 255875
rect 14595 255845 14600 255875
rect 14560 255840 14600 255845
rect 14640 255875 14680 255880
rect 14640 255845 14645 255875
rect 14675 255845 14680 255875
rect 14640 255840 14680 255845
rect 14720 255875 14760 255880
rect 14720 255845 14725 255875
rect 14755 255845 14760 255875
rect 14720 255840 14760 255845
rect 14800 255875 14840 255880
rect 14800 255845 14805 255875
rect 14835 255845 14840 255875
rect 14800 255840 14840 255845
rect 14880 255875 14920 255880
rect 14880 255845 14885 255875
rect 14915 255845 14920 255875
rect 14880 255840 14920 255845
rect 14960 255875 15000 255880
rect 14960 255845 14965 255875
rect 14995 255845 15000 255875
rect 14960 255840 15000 255845
rect 15040 255875 15080 255880
rect 15040 255845 15045 255875
rect 15075 255845 15080 255875
rect 15040 255840 15080 255845
rect 15120 255875 15160 255880
rect 15120 255845 15125 255875
rect 15155 255845 15160 255875
rect 15120 255840 15160 255845
rect 15200 255875 15240 255880
rect 15200 255845 15205 255875
rect 15235 255845 15240 255875
rect 15200 255840 15240 255845
rect 15280 255875 15320 255880
rect 15280 255845 15285 255875
rect 15315 255845 15320 255875
rect 15280 255840 15320 255845
rect 15360 255875 15400 255880
rect 15360 255845 15365 255875
rect 15395 255845 15400 255875
rect 15360 255840 15400 255845
rect 15440 255875 15480 255880
rect 15440 255845 15445 255875
rect 15475 255845 15480 255875
rect 15440 255840 15480 255845
rect 15520 255875 15560 255880
rect 15520 255845 15525 255875
rect 15555 255845 15560 255875
rect 15520 255840 15560 255845
rect 15600 255875 15640 255880
rect 15600 255845 15605 255875
rect 15635 255845 15640 255875
rect 15600 255840 15640 255845
rect 15680 255875 15720 255880
rect 15680 255845 15685 255875
rect 15715 255845 15720 255875
rect 15680 255840 15720 255845
rect 15760 255875 15800 255880
rect 15760 255845 15765 255875
rect 15795 255845 15800 255875
rect 15760 255840 15800 255845
rect 15840 255875 15880 255880
rect 15840 255845 15845 255875
rect 15875 255845 15880 255875
rect 15840 255840 15880 255845
rect 15920 255875 15960 255880
rect 15920 255845 15925 255875
rect 15955 255845 15960 255875
rect 15920 255840 15960 255845
rect 16000 255875 16040 255880
rect 16000 255845 16005 255875
rect 16035 255845 16040 255875
rect 16000 255840 16040 255845
rect 16080 255875 16120 255880
rect 16080 255845 16085 255875
rect 16115 255845 16120 255875
rect 16080 255840 16120 255845
rect 16160 255875 16200 255880
rect 16160 255845 16165 255875
rect 16195 255845 16200 255875
rect 16160 255840 16200 255845
rect 16240 255875 16280 255880
rect 16240 255845 16245 255875
rect 16275 255845 16280 255875
rect 16240 255840 16280 255845
rect 16320 255875 16360 255880
rect 16320 255845 16325 255875
rect 16355 255845 16360 255875
rect 16320 255840 16360 255845
rect 16400 255875 16440 255880
rect 16400 255845 16405 255875
rect 16435 255845 16440 255875
rect 16400 255840 16440 255845
rect 16480 255875 16520 255880
rect 16480 255845 16485 255875
rect 16515 255845 16520 255875
rect 16480 255840 16520 255845
rect 16560 255875 16600 255880
rect 16560 255845 16565 255875
rect 16595 255845 16600 255875
rect 16560 255840 16600 255845
rect 16640 255875 16680 255880
rect 16640 255845 16645 255875
rect 16675 255845 16680 255875
rect 16640 255840 16680 255845
rect 16720 255875 16760 255880
rect 16720 255845 16725 255875
rect 16755 255845 16760 255875
rect 16720 255840 16760 255845
rect 16880 255875 16920 255880
rect 16880 255845 16885 255875
rect 16915 255845 16920 255875
rect 16880 255840 16920 255845
rect 400 255715 440 255720
rect 400 255685 405 255715
rect 435 255685 440 255715
rect 400 255680 440 255685
rect 480 255715 520 255720
rect 480 255685 485 255715
rect 515 255685 520 255715
rect 480 255680 520 255685
rect 560 255715 600 255720
rect 560 255685 565 255715
rect 595 255685 600 255715
rect 560 255680 600 255685
rect 640 255715 680 255720
rect 640 255685 645 255715
rect 675 255685 680 255715
rect 640 255680 680 255685
rect 720 255715 760 255720
rect 720 255685 725 255715
rect 755 255685 760 255715
rect 720 255680 760 255685
rect 800 255715 840 255720
rect 800 255685 805 255715
rect 835 255685 840 255715
rect 800 255680 840 255685
rect 880 255715 920 255720
rect 880 255685 885 255715
rect 915 255685 920 255715
rect 880 255680 920 255685
rect 960 255715 1000 255720
rect 960 255685 965 255715
rect 995 255685 1000 255715
rect 960 255680 1000 255685
rect 1040 255715 1080 255720
rect 1040 255685 1045 255715
rect 1075 255685 1080 255715
rect 1040 255680 1080 255685
rect 1120 255715 1160 255720
rect 1120 255685 1125 255715
rect 1155 255685 1160 255715
rect 1120 255680 1160 255685
rect 1200 255715 1240 255720
rect 1200 255685 1205 255715
rect 1235 255685 1240 255715
rect 1200 255680 1240 255685
rect 1280 255715 1320 255720
rect 1280 255685 1285 255715
rect 1315 255685 1320 255715
rect 1280 255680 1320 255685
rect 1360 255715 1400 255720
rect 1360 255685 1365 255715
rect 1395 255685 1400 255715
rect 1360 255680 1400 255685
rect 1440 255715 1480 255720
rect 1440 255685 1445 255715
rect 1475 255685 1480 255715
rect 1440 255680 1480 255685
rect 1520 255715 1560 255720
rect 1520 255685 1525 255715
rect 1555 255685 1560 255715
rect 1520 255680 1560 255685
rect 1600 255715 1640 255720
rect 1600 255685 1605 255715
rect 1635 255685 1640 255715
rect 1600 255680 1640 255685
rect 1680 255715 1720 255720
rect 1680 255685 1685 255715
rect 1715 255685 1720 255715
rect 1680 255680 1720 255685
rect 1760 255715 1800 255720
rect 1760 255685 1765 255715
rect 1795 255685 1800 255715
rect 1760 255680 1800 255685
rect 1840 255715 1880 255720
rect 1840 255685 1845 255715
rect 1875 255685 1880 255715
rect 1840 255680 1880 255685
rect 1920 255715 1960 255720
rect 1920 255685 1925 255715
rect 1955 255685 1960 255715
rect 1920 255680 1960 255685
rect 2000 255715 2040 255720
rect 2000 255685 2005 255715
rect 2035 255685 2040 255715
rect 2000 255680 2040 255685
rect 2080 255715 2120 255720
rect 2080 255685 2085 255715
rect 2115 255685 2120 255715
rect 2080 255680 2120 255685
rect 2160 255715 2200 255720
rect 2160 255685 2165 255715
rect 2195 255685 2200 255715
rect 2160 255680 2200 255685
rect 2240 255715 2280 255720
rect 2240 255685 2245 255715
rect 2275 255685 2280 255715
rect 2240 255680 2280 255685
rect 2320 255715 2360 255720
rect 2320 255685 2325 255715
rect 2355 255685 2360 255715
rect 2320 255680 2360 255685
rect 2400 255715 2440 255720
rect 2400 255685 2405 255715
rect 2435 255685 2440 255715
rect 2400 255680 2440 255685
rect 2480 255715 2520 255720
rect 2480 255685 2485 255715
rect 2515 255685 2520 255715
rect 2480 255680 2520 255685
rect 2560 255715 2600 255720
rect 2560 255685 2565 255715
rect 2595 255685 2600 255715
rect 2560 255680 2600 255685
rect 2640 255715 2680 255720
rect 2640 255685 2645 255715
rect 2675 255685 2680 255715
rect 2640 255680 2680 255685
rect 2720 255715 2760 255720
rect 2720 255685 2725 255715
rect 2755 255685 2760 255715
rect 2720 255680 2760 255685
rect 3040 255715 3080 255720
rect 3040 255685 3045 255715
rect 3075 255685 3080 255715
rect 3040 255680 3080 255685
rect 3120 255715 3160 255720
rect 3120 255685 3125 255715
rect 3155 255685 3160 255715
rect 3120 255680 3160 255685
rect 3200 255715 3240 255720
rect 3200 255685 3205 255715
rect 3235 255685 3240 255715
rect 3200 255680 3240 255685
rect 3280 255715 3320 255720
rect 3280 255685 3285 255715
rect 3315 255685 3320 255715
rect 3280 255680 3320 255685
rect 3360 255715 3400 255720
rect 3360 255685 3365 255715
rect 3395 255685 3400 255715
rect 3360 255680 3400 255685
rect 3440 255715 3480 255720
rect 3440 255685 3445 255715
rect 3475 255685 3480 255715
rect 3440 255680 3480 255685
rect 3520 255715 3560 255720
rect 3520 255685 3525 255715
rect 3555 255685 3560 255715
rect 3520 255680 3560 255685
rect 3600 255715 3640 255720
rect 3600 255685 3605 255715
rect 3635 255685 3640 255715
rect 3600 255680 3640 255685
rect 3680 255715 3720 255720
rect 3680 255685 3685 255715
rect 3715 255685 3720 255715
rect 3680 255680 3720 255685
rect 3760 255715 3800 255720
rect 3760 255685 3765 255715
rect 3795 255685 3800 255715
rect 3760 255680 3800 255685
rect 3840 255715 3880 255720
rect 3840 255685 3845 255715
rect 3875 255685 3880 255715
rect 3840 255680 3880 255685
rect 3920 255715 3960 255720
rect 3920 255685 3925 255715
rect 3955 255685 3960 255715
rect 3920 255680 3960 255685
rect 4000 255715 4040 255720
rect 4000 255685 4005 255715
rect 4035 255685 4040 255715
rect 4000 255680 4040 255685
rect 4080 255715 4120 255720
rect 4080 255685 4085 255715
rect 4115 255685 4120 255715
rect 4080 255680 4120 255685
rect 4160 255715 4200 255720
rect 4160 255685 4165 255715
rect 4195 255685 4200 255715
rect 4160 255680 4200 255685
rect 4240 255715 4280 255720
rect 4240 255685 4245 255715
rect 4275 255685 4280 255715
rect 4240 255680 4280 255685
rect 4320 255715 4360 255720
rect 4320 255685 4325 255715
rect 4355 255685 4360 255715
rect 4320 255680 4360 255685
rect 4400 255715 4440 255720
rect 4400 255685 4405 255715
rect 4435 255685 4440 255715
rect 4400 255680 4440 255685
rect 4480 255715 4520 255720
rect 4480 255685 4485 255715
rect 4515 255685 4520 255715
rect 4480 255680 4520 255685
rect 4560 255715 4600 255720
rect 4560 255685 4565 255715
rect 4595 255685 4600 255715
rect 4560 255680 4600 255685
rect 4640 255715 4680 255720
rect 4640 255685 4645 255715
rect 4675 255685 4680 255715
rect 4640 255680 4680 255685
rect 4720 255715 4760 255720
rect 4720 255685 4725 255715
rect 4755 255685 4760 255715
rect 4720 255680 4760 255685
rect 4800 255715 4840 255720
rect 4800 255685 4805 255715
rect 4835 255685 4840 255715
rect 4800 255680 4840 255685
rect 4880 255715 4920 255720
rect 4880 255685 4885 255715
rect 4915 255685 4920 255715
rect 4880 255680 4920 255685
rect 4960 255715 5000 255720
rect 4960 255685 4965 255715
rect 4995 255685 5000 255715
rect 4960 255680 5000 255685
rect 5040 255715 5080 255720
rect 5040 255685 5045 255715
rect 5075 255685 5080 255715
rect 5040 255680 5080 255685
rect 5120 255715 5160 255720
rect 5120 255685 5125 255715
rect 5155 255685 5160 255715
rect 5120 255680 5160 255685
rect 5200 255715 5240 255720
rect 5200 255685 5205 255715
rect 5235 255685 5240 255715
rect 5200 255680 5240 255685
rect 5280 255715 5320 255720
rect 5280 255685 5285 255715
rect 5315 255685 5320 255715
rect 5280 255680 5320 255685
rect 5360 255715 5400 255720
rect 5360 255685 5365 255715
rect 5395 255685 5400 255715
rect 5360 255680 5400 255685
rect 5440 255715 5480 255720
rect 5440 255685 5445 255715
rect 5475 255685 5480 255715
rect 5440 255680 5480 255685
rect 5520 255715 5560 255720
rect 5520 255685 5525 255715
rect 5555 255685 5560 255715
rect 5520 255680 5560 255685
rect 5600 255715 5640 255720
rect 5600 255685 5605 255715
rect 5635 255685 5640 255715
rect 5600 255680 5640 255685
rect 5680 255715 5720 255720
rect 5680 255685 5685 255715
rect 5715 255685 5720 255715
rect 5680 255680 5720 255685
rect 5760 255715 5800 255720
rect 5760 255685 5765 255715
rect 5795 255685 5800 255715
rect 5760 255680 5800 255685
rect 5840 255715 5880 255720
rect 5840 255685 5845 255715
rect 5875 255685 5880 255715
rect 5840 255680 5880 255685
rect 5920 255715 5960 255720
rect 5920 255685 5925 255715
rect 5955 255685 5960 255715
rect 5920 255680 5960 255685
rect 6000 255715 6040 255720
rect 6000 255685 6005 255715
rect 6035 255685 6040 255715
rect 6000 255680 6040 255685
rect 6080 255715 6120 255720
rect 6080 255685 6085 255715
rect 6115 255685 6120 255715
rect 6080 255680 6120 255685
rect 6160 255715 6200 255720
rect 6160 255685 6165 255715
rect 6195 255685 6200 255715
rect 6160 255680 6200 255685
rect 6240 255715 6280 255720
rect 6240 255685 6245 255715
rect 6275 255685 6280 255715
rect 6240 255680 6280 255685
rect 6320 255715 6360 255720
rect 6320 255685 6325 255715
rect 6355 255685 6360 255715
rect 6320 255680 6360 255685
rect 6400 255715 6440 255720
rect 6400 255685 6405 255715
rect 6435 255685 6440 255715
rect 6400 255680 6440 255685
rect 6480 255715 6520 255720
rect 6480 255685 6485 255715
rect 6515 255685 6520 255715
rect 6480 255680 6520 255685
rect 6560 255715 6600 255720
rect 6560 255685 6565 255715
rect 6595 255685 6600 255715
rect 6560 255680 6600 255685
rect 6640 255715 6680 255720
rect 6640 255685 6645 255715
rect 6675 255685 6680 255715
rect 6640 255680 6680 255685
rect 6720 255715 6760 255720
rect 6720 255685 6725 255715
rect 6755 255685 6760 255715
rect 6720 255680 6760 255685
rect 6800 255715 6840 255720
rect 6800 255685 6805 255715
rect 6835 255685 6840 255715
rect 6800 255680 6840 255685
rect 6880 255715 6920 255720
rect 6880 255685 6885 255715
rect 6915 255685 6920 255715
rect 6880 255680 6920 255685
rect 6960 255715 7000 255720
rect 6960 255685 6965 255715
rect 6995 255685 7000 255715
rect 6960 255680 7000 255685
rect 7040 255715 7080 255720
rect 7040 255685 7045 255715
rect 7075 255685 7080 255715
rect 7040 255680 7080 255685
rect 7120 255715 7160 255720
rect 7120 255685 7125 255715
rect 7155 255685 7160 255715
rect 7120 255680 7160 255685
rect 7200 255715 7240 255720
rect 7200 255685 7205 255715
rect 7235 255685 7240 255715
rect 7200 255680 7240 255685
rect 7280 255715 7320 255720
rect 7280 255685 7285 255715
rect 7315 255685 7320 255715
rect 7280 255680 7320 255685
rect 7360 255715 7400 255720
rect 7360 255685 7365 255715
rect 7395 255685 7400 255715
rect 7360 255680 7400 255685
rect 7440 255715 7480 255720
rect 7440 255685 7445 255715
rect 7475 255685 7480 255715
rect 7440 255680 7480 255685
rect 7520 255715 7560 255720
rect 7520 255685 7525 255715
rect 7555 255685 7560 255715
rect 7520 255680 7560 255685
rect 7600 255715 7640 255720
rect 7600 255685 7605 255715
rect 7635 255685 7640 255715
rect 7600 255680 7640 255685
rect 7680 255715 7720 255720
rect 7680 255685 7685 255715
rect 7715 255685 7720 255715
rect 7680 255680 7720 255685
rect 7760 255715 7800 255720
rect 7760 255685 7765 255715
rect 7795 255685 7800 255715
rect 7760 255680 7800 255685
rect 7840 255715 7880 255720
rect 7840 255685 7845 255715
rect 7875 255685 7880 255715
rect 7840 255680 7880 255685
rect 7920 255715 7960 255720
rect 7920 255685 7925 255715
rect 7955 255685 7960 255715
rect 7920 255680 7960 255685
rect 8000 255715 8040 255720
rect 8000 255685 8005 255715
rect 8035 255685 8040 255715
rect 8000 255680 8040 255685
rect 8080 255715 8120 255720
rect 8080 255685 8085 255715
rect 8115 255685 8120 255715
rect 8080 255680 8120 255685
rect 8160 255715 8200 255720
rect 8160 255685 8165 255715
rect 8195 255685 8200 255715
rect 8160 255680 8200 255685
rect 8240 255715 8280 255720
rect 8240 255685 8245 255715
rect 8275 255685 8280 255715
rect 8240 255680 8280 255685
rect 8320 255715 8360 255720
rect 8320 255685 8325 255715
rect 8355 255685 8360 255715
rect 8320 255680 8360 255685
rect 8400 255715 8440 255720
rect 8400 255685 8405 255715
rect 8435 255685 8440 255715
rect 8400 255680 8440 255685
rect 8480 255715 8520 255720
rect 8480 255685 8485 255715
rect 8515 255685 8520 255715
rect 8480 255680 8520 255685
rect 8560 255715 8600 255720
rect 8560 255685 8565 255715
rect 8595 255685 8600 255715
rect 8560 255680 8600 255685
rect 8640 255715 8680 255720
rect 8640 255685 8645 255715
rect 8675 255685 8680 255715
rect 8640 255680 8680 255685
rect 8720 255715 8760 255720
rect 8720 255685 8725 255715
rect 8755 255685 8760 255715
rect 8720 255680 8760 255685
rect 8800 255715 8840 255720
rect 8800 255685 8805 255715
rect 8835 255685 8840 255715
rect 8800 255680 8840 255685
rect 8880 255715 8920 255720
rect 8880 255685 8885 255715
rect 8915 255685 8920 255715
rect 8880 255680 8920 255685
rect 8960 255715 9000 255720
rect 8960 255685 8965 255715
rect 8995 255685 9000 255715
rect 8960 255680 9000 255685
rect 9040 255715 9080 255720
rect 9040 255685 9045 255715
rect 9075 255685 9080 255715
rect 9040 255680 9080 255685
rect 9120 255715 9160 255720
rect 9120 255685 9125 255715
rect 9155 255685 9160 255715
rect 9120 255680 9160 255685
rect 9200 255715 9240 255720
rect 9200 255685 9205 255715
rect 9235 255685 9240 255715
rect 9200 255680 9240 255685
rect 9280 255715 9320 255720
rect 9280 255685 9285 255715
rect 9315 255685 9320 255715
rect 9280 255680 9320 255685
rect 9360 255715 9400 255720
rect 9360 255685 9365 255715
rect 9395 255685 9400 255715
rect 9360 255680 9400 255685
rect 9440 255715 9480 255720
rect 9440 255685 9445 255715
rect 9475 255685 9480 255715
rect 9440 255680 9480 255685
rect 9520 255715 9560 255720
rect 9520 255685 9525 255715
rect 9555 255685 9560 255715
rect 9520 255680 9560 255685
rect 9600 255715 9640 255720
rect 9600 255685 9605 255715
rect 9635 255685 9640 255715
rect 9600 255680 9640 255685
rect 9680 255715 9720 255720
rect 9680 255685 9685 255715
rect 9715 255685 9720 255715
rect 9680 255680 9720 255685
rect 9760 255715 9800 255720
rect 9760 255685 9765 255715
rect 9795 255685 9800 255715
rect 9760 255680 9800 255685
rect 9840 255715 9880 255720
rect 9840 255685 9845 255715
rect 9875 255685 9880 255715
rect 9840 255680 9880 255685
rect 9920 255715 9960 255720
rect 9920 255685 9925 255715
rect 9955 255685 9960 255715
rect 9920 255680 9960 255685
rect 10000 255715 10040 255720
rect 10000 255685 10005 255715
rect 10035 255685 10040 255715
rect 10000 255680 10040 255685
rect 10080 255715 10120 255720
rect 10080 255685 10085 255715
rect 10115 255685 10120 255715
rect 10080 255680 10120 255685
rect 10160 255715 10200 255720
rect 10160 255685 10165 255715
rect 10195 255685 10200 255715
rect 10160 255680 10200 255685
rect 10240 255715 10280 255720
rect 10240 255685 10245 255715
rect 10275 255685 10280 255715
rect 10240 255680 10280 255685
rect 10320 255715 10360 255720
rect 10320 255685 10325 255715
rect 10355 255685 10360 255715
rect 10320 255680 10360 255685
rect 10400 255715 10440 255720
rect 10400 255685 10405 255715
rect 10435 255685 10440 255715
rect 10400 255680 10440 255685
rect 10480 255715 10520 255720
rect 10480 255685 10485 255715
rect 10515 255685 10520 255715
rect 10480 255680 10520 255685
rect 10560 255715 10600 255720
rect 10560 255685 10565 255715
rect 10595 255685 10600 255715
rect 10560 255680 10600 255685
rect 10640 255715 10680 255720
rect 10640 255685 10645 255715
rect 10675 255685 10680 255715
rect 10640 255680 10680 255685
rect 10720 255715 10760 255720
rect 10720 255685 10725 255715
rect 10755 255685 10760 255715
rect 10720 255680 10760 255685
rect 10800 255715 10840 255720
rect 10800 255685 10805 255715
rect 10835 255685 10840 255715
rect 10800 255680 10840 255685
rect 10880 255715 10920 255720
rect 10880 255685 10885 255715
rect 10915 255685 10920 255715
rect 10880 255680 10920 255685
rect 10960 255715 11000 255720
rect 10960 255685 10965 255715
rect 10995 255685 11000 255715
rect 10960 255680 11000 255685
rect 11040 255715 11080 255720
rect 11040 255685 11045 255715
rect 11075 255685 11080 255715
rect 11040 255680 11080 255685
rect 11120 255715 11160 255720
rect 11120 255685 11125 255715
rect 11155 255685 11160 255715
rect 11120 255680 11160 255685
rect 11200 255715 11240 255720
rect 11200 255685 11205 255715
rect 11235 255685 11240 255715
rect 11200 255680 11240 255685
rect 11280 255715 11320 255720
rect 11280 255685 11285 255715
rect 11315 255685 11320 255715
rect 11280 255680 11320 255685
rect 11360 255715 11400 255720
rect 11360 255685 11365 255715
rect 11395 255685 11400 255715
rect 11360 255680 11400 255685
rect 11440 255715 11480 255720
rect 11440 255685 11445 255715
rect 11475 255685 11480 255715
rect 11440 255680 11480 255685
rect 11520 255715 11560 255720
rect 11520 255685 11525 255715
rect 11555 255685 11560 255715
rect 11520 255680 11560 255685
rect 11600 255715 11640 255720
rect 11600 255685 11605 255715
rect 11635 255685 11640 255715
rect 11600 255680 11640 255685
rect 11680 255715 11720 255720
rect 11680 255685 11685 255715
rect 11715 255685 11720 255715
rect 11680 255680 11720 255685
rect 11760 255715 11800 255720
rect 11760 255685 11765 255715
rect 11795 255685 11800 255715
rect 11760 255680 11800 255685
rect 11840 255715 11880 255720
rect 11840 255685 11845 255715
rect 11875 255685 11880 255715
rect 11840 255680 11880 255685
rect 11920 255715 11960 255720
rect 11920 255685 11925 255715
rect 11955 255685 11960 255715
rect 11920 255680 11960 255685
rect 12000 255715 12040 255720
rect 12000 255685 12005 255715
rect 12035 255685 12040 255715
rect 12000 255680 12040 255685
rect 12080 255715 12120 255720
rect 12080 255685 12085 255715
rect 12115 255685 12120 255715
rect 12080 255680 12120 255685
rect 12160 255715 12200 255720
rect 12160 255685 12165 255715
rect 12195 255685 12200 255715
rect 12160 255680 12200 255685
rect 12240 255715 12280 255720
rect 12240 255685 12245 255715
rect 12275 255685 12280 255715
rect 12240 255680 12280 255685
rect 12320 255715 12360 255720
rect 12320 255685 12325 255715
rect 12355 255685 12360 255715
rect 12320 255680 12360 255685
rect 12400 255715 12440 255720
rect 12400 255685 12405 255715
rect 12435 255685 12440 255715
rect 12400 255680 12440 255685
rect 12480 255715 12520 255720
rect 12480 255685 12485 255715
rect 12515 255685 12520 255715
rect 12480 255680 12520 255685
rect 12560 255715 12600 255720
rect 12560 255685 12565 255715
rect 12595 255685 12600 255715
rect 12560 255680 12600 255685
rect 12640 255715 12680 255720
rect 12640 255685 12645 255715
rect 12675 255685 12680 255715
rect 12640 255680 12680 255685
rect 12720 255715 12760 255720
rect 12720 255685 12725 255715
rect 12755 255685 12760 255715
rect 12720 255680 12760 255685
rect 12800 255715 12840 255720
rect 12800 255685 12805 255715
rect 12835 255685 12840 255715
rect 12800 255680 12840 255685
rect 12880 255715 12920 255720
rect 12880 255685 12885 255715
rect 12915 255685 12920 255715
rect 12880 255680 12920 255685
rect 12960 255715 13000 255720
rect 12960 255685 12965 255715
rect 12995 255685 13000 255715
rect 12960 255680 13000 255685
rect 13040 255715 13080 255720
rect 13040 255685 13045 255715
rect 13075 255685 13080 255715
rect 13040 255680 13080 255685
rect 13120 255715 13160 255720
rect 13120 255685 13125 255715
rect 13155 255685 13160 255715
rect 13120 255680 13160 255685
rect 13200 255715 13240 255720
rect 13200 255685 13205 255715
rect 13235 255685 13240 255715
rect 13200 255680 13240 255685
rect 13280 255715 13320 255720
rect 13280 255685 13285 255715
rect 13315 255685 13320 255715
rect 13280 255680 13320 255685
rect 13360 255715 13400 255720
rect 13360 255685 13365 255715
rect 13395 255685 13400 255715
rect 13360 255680 13400 255685
rect 13440 255715 13480 255720
rect 13440 255685 13445 255715
rect 13475 255685 13480 255715
rect 13440 255680 13480 255685
rect 13520 255715 13560 255720
rect 13520 255685 13525 255715
rect 13555 255685 13560 255715
rect 13520 255680 13560 255685
rect 13600 255715 13640 255720
rect 13600 255685 13605 255715
rect 13635 255685 13640 255715
rect 13600 255680 13640 255685
rect 13680 255715 13720 255720
rect 13680 255685 13685 255715
rect 13715 255685 13720 255715
rect 13680 255680 13720 255685
rect 13760 255715 13800 255720
rect 13760 255685 13765 255715
rect 13795 255685 13800 255715
rect 13760 255680 13800 255685
rect 13840 255715 13880 255720
rect 13840 255685 13845 255715
rect 13875 255685 13880 255715
rect 13840 255680 13880 255685
rect 13920 255715 13960 255720
rect 13920 255685 13925 255715
rect 13955 255685 13960 255715
rect 13920 255680 13960 255685
rect 14000 255715 14040 255720
rect 14000 255685 14005 255715
rect 14035 255685 14040 255715
rect 14000 255680 14040 255685
rect 14080 255715 14120 255720
rect 14080 255685 14085 255715
rect 14115 255685 14120 255715
rect 14080 255680 14120 255685
rect 14160 255715 14200 255720
rect 14160 255685 14165 255715
rect 14195 255685 14200 255715
rect 14160 255680 14200 255685
rect 14240 255715 14280 255720
rect 14240 255685 14245 255715
rect 14275 255685 14280 255715
rect 14240 255680 14280 255685
rect 14320 255715 14360 255720
rect 14320 255685 14325 255715
rect 14355 255685 14360 255715
rect 14320 255680 14360 255685
rect 14400 255715 14440 255720
rect 14400 255685 14405 255715
rect 14435 255685 14440 255715
rect 14400 255680 14440 255685
rect 14480 255715 14520 255720
rect 14480 255685 14485 255715
rect 14515 255685 14520 255715
rect 14480 255680 14520 255685
rect 14560 255715 14600 255720
rect 14560 255685 14565 255715
rect 14595 255685 14600 255715
rect 14560 255680 14600 255685
rect 14640 255715 14680 255720
rect 14640 255685 14645 255715
rect 14675 255685 14680 255715
rect 14640 255680 14680 255685
rect 14720 255715 14760 255720
rect 14720 255685 14725 255715
rect 14755 255685 14760 255715
rect 14720 255680 14760 255685
rect 14800 255715 14840 255720
rect 14800 255685 14805 255715
rect 14835 255685 14840 255715
rect 14800 255680 14840 255685
rect 14880 255715 14920 255720
rect 14880 255685 14885 255715
rect 14915 255685 14920 255715
rect 14880 255680 14920 255685
rect 14960 255715 15000 255720
rect 14960 255685 14965 255715
rect 14995 255685 15000 255715
rect 14960 255680 15000 255685
rect 15040 255715 15080 255720
rect 15040 255685 15045 255715
rect 15075 255685 15080 255715
rect 15040 255680 15080 255685
rect 15120 255715 15160 255720
rect 15120 255685 15125 255715
rect 15155 255685 15160 255715
rect 15120 255680 15160 255685
rect 15200 255715 15240 255720
rect 15200 255685 15205 255715
rect 15235 255685 15240 255715
rect 15200 255680 15240 255685
rect 15280 255715 15320 255720
rect 15280 255685 15285 255715
rect 15315 255685 15320 255715
rect 15280 255680 15320 255685
rect 15360 255715 15400 255720
rect 15360 255685 15365 255715
rect 15395 255685 15400 255715
rect 15360 255680 15400 255685
rect 15440 255715 15480 255720
rect 15440 255685 15445 255715
rect 15475 255685 15480 255715
rect 15440 255680 15480 255685
rect 15520 255715 15560 255720
rect 15520 255685 15525 255715
rect 15555 255685 15560 255715
rect 15520 255680 15560 255685
rect 15600 255715 15640 255720
rect 15600 255685 15605 255715
rect 15635 255685 15640 255715
rect 15600 255680 15640 255685
rect 15680 255715 15720 255720
rect 15680 255685 15685 255715
rect 15715 255685 15720 255715
rect 15680 255680 15720 255685
rect 15760 255715 15800 255720
rect 15760 255685 15765 255715
rect 15795 255685 15800 255715
rect 15760 255680 15800 255685
rect 15840 255715 15880 255720
rect 15840 255685 15845 255715
rect 15875 255685 15880 255715
rect 15840 255680 15880 255685
rect 15920 255715 15960 255720
rect 15920 255685 15925 255715
rect 15955 255685 15960 255715
rect 15920 255680 15960 255685
rect 16000 255715 16040 255720
rect 16000 255685 16005 255715
rect 16035 255685 16040 255715
rect 16000 255680 16040 255685
rect 16080 255715 16120 255720
rect 16080 255685 16085 255715
rect 16115 255685 16120 255715
rect 16080 255680 16120 255685
rect 16160 255715 16200 255720
rect 16160 255685 16165 255715
rect 16195 255685 16200 255715
rect 16160 255680 16200 255685
rect 16240 255715 16280 255720
rect 16240 255685 16245 255715
rect 16275 255685 16280 255715
rect 16240 255680 16280 255685
rect 16320 255715 16360 255720
rect 16320 255685 16325 255715
rect 16355 255685 16360 255715
rect 16320 255680 16360 255685
rect 16400 255715 16440 255720
rect 16400 255685 16405 255715
rect 16435 255685 16440 255715
rect 16400 255680 16440 255685
rect 16480 255715 16520 255720
rect 16480 255685 16485 255715
rect 16515 255685 16520 255715
rect 16480 255680 16520 255685
rect 16560 255715 16600 255720
rect 16560 255685 16565 255715
rect 16595 255685 16600 255715
rect 16560 255680 16600 255685
rect 16640 255715 16680 255720
rect 16640 255685 16645 255715
rect 16675 255685 16680 255715
rect 16640 255680 16680 255685
rect 16720 255715 16760 255720
rect 16720 255685 16725 255715
rect 16755 255685 16760 255715
rect 16720 255680 16760 255685
rect 16880 255715 16920 255720
rect 16880 255685 16885 255715
rect 16915 255685 16920 255715
rect 16880 255680 16920 255685
<< via1 >>
rect 271865 351785 271895 351815
rect 272025 351785 272055 351815
rect 272105 351785 272135 351815
rect 272185 351785 272215 351815
rect 272265 351785 272295 351815
rect 272345 351785 272375 351815
rect 272425 351785 272455 351815
rect 272505 351785 272535 351815
rect 272585 351785 272615 351815
rect 272665 351785 272695 351815
rect 272745 351785 272775 351815
rect 272825 351785 272855 351815
rect 272905 351785 272935 351815
rect 272985 351785 273015 351815
rect 273065 351785 273095 351815
rect 273145 351785 273175 351815
rect 273225 351785 273255 351815
rect 273305 351785 273335 351815
rect 273385 351785 273415 351815
rect 273465 351785 273495 351815
rect 273545 351785 273575 351815
rect 273625 351785 273655 351815
rect 273705 351785 273735 351815
rect 273785 351785 273815 351815
rect 273865 351785 273895 351815
rect 273945 351785 273975 351815
rect 274025 351785 274055 351815
rect 274105 351785 274135 351815
rect 274185 351785 274215 351815
rect 274265 351785 274295 351815
rect 274345 351785 274375 351815
rect 274425 351785 274455 351815
rect 274505 351785 274535 351815
rect 274585 351785 274615 351815
rect 274665 351785 274695 351815
rect 274745 351785 274775 351815
rect 274825 351785 274855 351815
rect 274905 351785 274935 351815
rect 274985 351785 275015 351815
rect 275065 351785 275095 351815
rect 275145 351785 275175 351815
rect 275225 351785 275255 351815
rect 275305 351785 275335 351815
rect 275385 351785 275415 351815
rect 275465 351785 275495 351815
rect 275545 351785 275575 351815
rect 275625 351785 275655 351815
rect 275705 351785 275735 351815
rect 275785 351785 275815 351815
rect 275865 351785 275895 351815
rect 275945 351785 275975 351815
rect 276025 351785 276055 351815
rect 276105 351785 276135 351815
rect 276185 351785 276215 351815
rect 276265 351785 276295 351815
rect 276345 351785 276375 351815
rect 276425 351785 276455 351815
rect 276505 351785 276535 351815
rect 276585 351785 276615 351815
rect 276665 351785 276695 351815
rect 276745 351785 276775 351815
rect 276825 351785 276855 351815
rect 276905 351785 276935 351815
rect 276985 351785 277015 351815
rect 277065 351785 277095 351815
rect 277145 351785 277175 351815
rect 277225 351785 277255 351815
rect 277305 351785 277335 351815
rect 277385 351785 277415 351815
rect 277465 351785 277495 351815
rect 277545 351785 277575 351815
rect 277625 351785 277655 351815
rect 277705 351785 277735 351815
rect 277785 351785 277815 351815
rect 277865 351785 277895 351815
rect 277945 351785 277975 351815
rect 278025 351785 278055 351815
rect 278105 351785 278135 351815
rect 278185 351785 278215 351815
rect 278265 351785 278295 351815
rect 278345 351785 278375 351815
rect 278425 351785 278455 351815
rect 278505 351785 278535 351815
rect 278585 351785 278615 351815
rect 278665 351785 278695 351815
rect 278745 351785 278775 351815
rect 278825 351785 278855 351815
rect 278905 351785 278935 351815
rect 278985 351785 279015 351815
rect 279065 351785 279095 351815
rect 279145 351785 279175 351815
rect 279225 351785 279255 351815
rect 279305 351785 279335 351815
rect 279385 351785 279415 351815
rect 279465 351785 279495 351815
rect 279545 351785 279575 351815
rect 279625 351785 279655 351815
rect 279705 351785 279735 351815
rect 279785 351785 279815 351815
rect 279865 351785 279895 351815
rect 279945 351785 279975 351815
rect 280025 351785 280055 351815
rect 280105 351785 280135 351815
rect 280185 351785 280215 351815
rect 280265 351785 280295 351815
rect 280345 351785 280375 351815
rect 280425 351785 280455 351815
rect 280505 351785 280535 351815
rect 280585 351785 280615 351815
rect 280665 351785 280695 351815
rect 280745 351785 280775 351815
rect 280825 351785 280855 351815
rect 280905 351785 280935 351815
rect 280985 351785 281015 351815
rect 281065 351785 281095 351815
rect 281145 351785 281175 351815
rect 281225 351785 281255 351815
rect 281305 351785 281335 351815
rect 281385 351785 281415 351815
rect 281465 351785 281495 351815
rect 281545 351785 281575 351815
rect 281625 351785 281655 351815
rect 281705 351785 281735 351815
rect 281785 351785 281815 351815
rect 281865 351785 281895 351815
rect 281945 351785 281975 351815
rect 282025 351785 282055 351815
rect 282105 351785 282135 351815
rect 282185 351785 282215 351815
rect 282265 351785 282295 351815
rect 282345 351785 282375 351815
rect 282425 351785 282455 351815
rect 282505 351785 282535 351815
rect 282585 351785 282615 351815
rect 282665 351785 282695 351815
rect 282745 351785 282775 351815
rect 282825 351785 282855 351815
rect 282905 351785 282935 351815
rect 282985 351785 283015 351815
rect 283065 351785 283095 351815
rect 283145 351785 283175 351815
rect 271865 351625 271895 351655
rect 272025 351625 272055 351655
rect 272105 351625 272135 351655
rect 272185 351625 272215 351655
rect 272265 351625 272295 351655
rect 272345 351625 272375 351655
rect 272425 351625 272455 351655
rect 272505 351625 272535 351655
rect 272585 351625 272615 351655
rect 272665 351625 272695 351655
rect 272745 351625 272775 351655
rect 272825 351625 272855 351655
rect 272905 351625 272935 351655
rect 272985 351625 273015 351655
rect 273065 351625 273095 351655
rect 273145 351625 273175 351655
rect 273225 351625 273255 351655
rect 273305 351625 273335 351655
rect 273385 351625 273415 351655
rect 273465 351625 273495 351655
rect 273545 351625 273575 351655
rect 273625 351625 273655 351655
rect 273705 351625 273735 351655
rect 273785 351625 273815 351655
rect 273865 351625 273895 351655
rect 273945 351625 273975 351655
rect 274025 351625 274055 351655
rect 274105 351625 274135 351655
rect 274185 351625 274215 351655
rect 274265 351625 274295 351655
rect 274345 351625 274375 351655
rect 274425 351625 274455 351655
rect 274505 351625 274535 351655
rect 274585 351625 274615 351655
rect 274665 351625 274695 351655
rect 274745 351625 274775 351655
rect 274825 351625 274855 351655
rect 274905 351625 274935 351655
rect 274985 351625 275015 351655
rect 275065 351625 275095 351655
rect 275145 351625 275175 351655
rect 275225 351625 275255 351655
rect 275305 351625 275335 351655
rect 275385 351625 275415 351655
rect 275465 351625 275495 351655
rect 275545 351625 275575 351655
rect 275625 351625 275655 351655
rect 275705 351625 275735 351655
rect 275785 351625 275815 351655
rect 275865 351625 275895 351655
rect 275945 351625 275975 351655
rect 276025 351625 276055 351655
rect 276105 351625 276135 351655
rect 276185 351625 276215 351655
rect 276265 351625 276295 351655
rect 276345 351625 276375 351655
rect 276425 351625 276455 351655
rect 276505 351625 276535 351655
rect 276585 351625 276615 351655
rect 276665 351625 276695 351655
rect 276745 351625 276775 351655
rect 276825 351625 276855 351655
rect 276905 351625 276935 351655
rect 276985 351625 277015 351655
rect 277065 351625 277095 351655
rect 277145 351625 277175 351655
rect 277225 351625 277255 351655
rect 277305 351625 277335 351655
rect 277385 351625 277415 351655
rect 277465 351625 277495 351655
rect 277545 351625 277575 351655
rect 277625 351625 277655 351655
rect 277705 351625 277735 351655
rect 277785 351625 277815 351655
rect 277865 351625 277895 351655
rect 277945 351625 277975 351655
rect 278025 351625 278055 351655
rect 278105 351625 278135 351655
rect 278185 351625 278215 351655
rect 278265 351625 278295 351655
rect 278345 351625 278375 351655
rect 278425 351625 278455 351655
rect 278505 351625 278535 351655
rect 278585 351625 278615 351655
rect 278665 351625 278695 351655
rect 278745 351625 278775 351655
rect 278825 351625 278855 351655
rect 278905 351625 278935 351655
rect 278985 351625 279015 351655
rect 279065 351625 279095 351655
rect 279145 351625 279175 351655
rect 279225 351625 279255 351655
rect 279305 351625 279335 351655
rect 279385 351625 279415 351655
rect 279465 351625 279495 351655
rect 279545 351625 279575 351655
rect 279625 351625 279655 351655
rect 279705 351625 279735 351655
rect 279785 351625 279815 351655
rect 279865 351625 279895 351655
rect 279945 351625 279975 351655
rect 280025 351625 280055 351655
rect 280105 351625 280135 351655
rect 280185 351625 280215 351655
rect 280265 351625 280295 351655
rect 280345 351625 280375 351655
rect 280425 351625 280455 351655
rect 280505 351625 280535 351655
rect 280585 351625 280615 351655
rect 280665 351625 280695 351655
rect 280745 351625 280775 351655
rect 280825 351625 280855 351655
rect 280905 351625 280935 351655
rect 280985 351625 281015 351655
rect 281065 351625 281095 351655
rect 281145 351625 281175 351655
rect 281225 351625 281255 351655
rect 281305 351625 281335 351655
rect 281385 351625 281415 351655
rect 281465 351625 281495 351655
rect 281545 351625 281575 351655
rect 281625 351625 281655 351655
rect 281705 351625 281735 351655
rect 281785 351625 281815 351655
rect 281865 351625 281895 351655
rect 281945 351625 281975 351655
rect 282025 351625 282055 351655
rect 282105 351625 282135 351655
rect 282185 351625 282215 351655
rect 282265 351625 282295 351655
rect 282345 351625 282375 351655
rect 282425 351625 282455 351655
rect 282505 351625 282535 351655
rect 282585 351625 282615 351655
rect 282665 351625 282695 351655
rect 282745 351625 282775 351655
rect 282825 351625 282855 351655
rect 282905 351625 282935 351655
rect 282985 351625 283015 351655
rect 283065 351625 283095 351655
rect 283145 351625 283175 351655
rect 16725 275445 16755 275475
rect 16885 275445 16915 275475
rect 16965 275445 16995 275475
rect 17045 275445 17075 275475
rect 17125 275445 17155 275475
rect 17205 275445 17235 275475
rect 16725 275285 16755 275315
rect 16885 275285 16915 275315
rect 16965 275285 16995 275315
rect 17045 275285 17075 275315
rect 17205 275285 17235 275315
rect 16725 274925 16755 274955
rect 16885 274925 16915 274955
rect 16725 274845 16755 274875
rect 16885 274845 16915 274875
rect 16725 274765 16755 274795
rect 16885 274765 16915 274795
rect 16725 274685 16755 274715
rect 16885 274685 16915 274715
rect 16725 274605 16755 274635
rect 16885 274605 16915 274635
rect 16725 274525 16755 274555
rect 16885 274525 16915 274555
rect 16725 274445 16755 274475
rect 16885 274445 16915 274475
rect 16725 274365 16755 274395
rect 16885 274365 16915 274395
rect 16725 274285 16755 274315
rect 16885 274285 16915 274315
rect 16725 274205 16755 274235
rect 16885 274205 16915 274235
rect 16725 274125 16755 274155
rect 16885 274125 16915 274155
rect 16725 274045 16755 274075
rect 16885 274045 16915 274075
rect 16725 273965 16755 273995
rect 16885 273965 16915 273995
rect 16725 273885 16755 273915
rect 16885 273885 16915 273915
rect 16725 273805 16755 273835
rect 16885 273805 16915 273835
rect 16725 273725 16755 273755
rect 16885 273725 16915 273755
rect 16725 273645 16755 273675
rect 16885 273645 16915 273675
rect 16725 273565 16755 273595
rect 16885 273565 16915 273595
rect 16725 273485 16755 273515
rect 16885 273485 16915 273515
rect 16725 273405 16755 273435
rect 16885 273405 16915 273435
rect 16725 273325 16755 273355
rect 16885 273325 16915 273355
rect 16725 273245 16755 273275
rect 16885 273245 16915 273275
rect 16725 273165 16755 273195
rect 16885 273165 16915 273195
rect 16725 273085 16755 273115
rect 16885 273085 16915 273115
rect 16725 273005 16755 273035
rect 16885 273005 16915 273035
rect 16725 272925 16755 272955
rect 16885 272925 16915 272955
rect 16725 272845 16755 272875
rect 16885 272845 16915 272875
rect 16725 272765 16755 272795
rect 16885 272765 16915 272795
rect 16725 272685 16755 272715
rect 16885 272685 16915 272715
rect 16725 272605 16755 272635
rect 16885 272605 16915 272635
rect 16725 272525 16755 272555
rect 16885 272525 16915 272555
rect 16725 272445 16755 272475
rect 16885 272445 16915 272475
rect 16725 272365 16755 272395
rect 16885 272365 16915 272395
rect 16725 272285 16755 272315
rect 16885 272285 16915 272315
rect 16725 272205 16755 272235
rect 16885 272205 16915 272235
rect 16725 272125 16755 272155
rect 16885 272125 16915 272155
rect 16725 272045 16755 272075
rect 16885 272045 16915 272075
rect 16725 271965 16755 271995
rect 16885 271965 16915 271995
rect 16725 271885 16755 271915
rect 16885 271885 16915 271915
rect 16725 271805 16755 271835
rect 16885 271805 16915 271835
rect 16725 271725 16755 271755
rect 16885 271725 16915 271755
rect 16725 271645 16755 271675
rect 16885 271645 16915 271675
rect 16725 271565 16755 271595
rect 16885 271565 16915 271595
rect 16725 271485 16755 271515
rect 16885 271485 16915 271515
rect 16725 271405 16755 271435
rect 16885 271405 16915 271435
rect 16725 271325 16755 271355
rect 16885 271325 16915 271355
rect 16725 271245 16755 271275
rect 16885 271245 16915 271275
rect 16725 271165 16755 271195
rect 16885 271165 16915 271195
rect 16725 271085 16755 271115
rect 16885 271085 16915 271115
rect 16725 271005 16755 271035
rect 16885 271005 16915 271035
rect 16725 270925 16755 270955
rect 16885 270925 16915 270955
rect 16725 270845 16755 270875
rect 16885 270845 16915 270875
rect 16725 270765 16755 270795
rect 16885 270765 16915 270795
rect 16725 270685 16755 270715
rect 16885 270685 16915 270715
rect 16725 270605 16755 270635
rect 16885 270605 16915 270635
rect 16725 270525 16755 270555
rect 16885 270525 16915 270555
rect 16725 270445 16755 270475
rect 16885 270445 16915 270475
rect 16725 270365 16755 270395
rect 16885 270365 16915 270395
rect 16725 270285 16755 270315
rect 16885 270285 16915 270315
rect 16725 270205 16755 270235
rect 16885 270205 16915 270235
rect 16725 270125 16755 270155
rect 16885 270125 16915 270155
rect 16725 270045 16755 270075
rect 16885 270045 16915 270075
rect 16725 269965 16755 269995
rect 16885 269965 16915 269995
rect 16725 269885 16755 269915
rect 16885 269885 16915 269915
rect 16725 269805 16755 269835
rect 16885 269805 16915 269835
rect 16725 269725 16755 269755
rect 16885 269725 16915 269755
rect 16725 269645 16755 269675
rect 16885 269645 16915 269675
rect 16725 269565 16755 269595
rect 16885 269565 16915 269595
rect 16725 269485 16755 269515
rect 16885 269485 16915 269515
rect 16725 269405 16755 269435
rect 16885 269405 16915 269435
rect 16725 269325 16755 269355
rect 16885 269325 16915 269355
rect 16725 269245 16755 269275
rect 16885 269245 16915 269275
rect 16725 269165 16755 269195
rect 16885 269165 16915 269195
rect 16725 269085 16755 269115
rect 16885 269085 16915 269115
rect 16725 269005 16755 269035
rect 16885 269005 16915 269035
rect 16725 268925 16755 268955
rect 16885 268925 16915 268955
rect 16725 268845 16755 268875
rect 16885 268845 16915 268875
rect 16725 268765 16755 268795
rect 16885 268765 16915 268795
rect 16725 268685 16755 268715
rect 16885 268685 16915 268715
rect 16725 268605 16755 268635
rect 16885 268605 16915 268635
rect 16725 268525 16755 268555
rect 16885 268525 16915 268555
rect 16725 268445 16755 268475
rect 16885 268445 16915 268475
rect 16725 268365 16755 268395
rect 16885 268365 16915 268395
rect 16725 268285 16755 268315
rect 16885 268285 16915 268315
rect 16725 268205 16755 268235
rect 16885 268205 16915 268235
rect 16725 268125 16755 268155
rect 16885 268125 16915 268155
rect 16725 268045 16755 268075
rect 16885 268045 16915 268075
rect 16725 267965 16755 267995
rect 16885 267965 16915 267995
rect 16725 267885 16755 267915
rect 16885 267885 16915 267915
rect 16725 267805 16755 267835
rect 16885 267805 16915 267835
rect 16725 267725 16755 267755
rect 16885 267725 16915 267755
rect 16725 267645 16755 267675
rect 16885 267645 16915 267675
rect 16725 267565 16755 267595
rect 16885 267565 16915 267595
rect 16725 267485 16755 267515
rect 16885 267485 16915 267515
rect 16725 267405 16755 267435
rect 16885 267405 16915 267435
rect 16725 267325 16755 267355
rect 16885 267325 16915 267355
rect 16725 267245 16755 267275
rect 16885 267245 16915 267275
rect 16725 267165 16755 267195
rect 16885 267165 16915 267195
rect 16725 267085 16755 267115
rect 16885 267085 16915 267115
rect 16725 267005 16755 267035
rect 16885 267005 16915 267035
rect 16725 266925 16755 266955
rect 16885 266925 16915 266955
rect 16725 266845 16755 266875
rect 16885 266845 16915 266875
rect 16725 266765 16755 266795
rect 16885 266765 16915 266795
rect 16725 266685 16755 266715
rect 16885 266685 16915 266715
rect 16725 266605 16755 266635
rect 16885 266605 16915 266635
rect 16725 266525 16755 266555
rect 16885 266525 16915 266555
rect 16725 266445 16755 266475
rect 16885 266445 16915 266475
rect 16725 266365 16755 266395
rect 16885 266365 16915 266395
rect 16725 266285 16755 266315
rect 16885 266285 16915 266315
rect 16725 266205 16755 266235
rect 16885 266205 16915 266235
rect 16725 266125 16755 266155
rect 16885 266125 16915 266155
rect 16725 266045 16755 266075
rect 16885 266045 16915 266075
rect 16725 265965 16755 265995
rect 16885 265965 16915 265995
rect 16725 265885 16755 265915
rect 16885 265885 16915 265915
rect 16725 265805 16755 265835
rect 16885 265805 16915 265835
rect 16725 265725 16755 265755
rect 16885 265725 16915 265755
rect 16725 265645 16755 265675
rect 16885 265645 16915 265675
rect 16725 265565 16755 265595
rect 16885 265565 16915 265595
rect 16725 265485 16755 265515
rect 16885 265485 16915 265515
rect 16725 265405 16755 265435
rect 16885 265405 16915 265435
rect 16725 265325 16755 265355
rect 16885 265325 16915 265355
rect 16725 265245 16755 265275
rect 16885 265245 16915 265275
rect 16725 265165 16755 265195
rect 16885 265165 16915 265195
rect 16725 265085 16755 265115
rect 16885 265085 16915 265115
rect 16725 265005 16755 265035
rect 16885 265005 16915 265035
rect 16725 264925 16755 264955
rect 16885 264925 16915 264955
rect 16725 264845 16755 264875
rect 16885 264845 16915 264875
rect 16725 264765 16755 264795
rect 16885 264765 16915 264795
rect 16725 264685 16755 264715
rect 16885 264685 16915 264715
rect 16725 264605 16755 264635
rect 16885 264605 16915 264635
rect 16725 264525 16755 264555
rect 16885 264525 16915 264555
rect 16725 264445 16755 264475
rect 16885 264445 16915 264475
rect 16725 264365 16755 264395
rect 16885 264365 16915 264395
rect 16725 264285 16755 264315
rect 16885 264285 16915 264315
rect 16725 264205 16755 264235
rect 16885 264205 16915 264235
rect 16725 264125 16755 264155
rect 16885 264125 16915 264155
rect 16725 264045 16755 264075
rect 16885 264045 16915 264075
rect 16725 263965 16755 263995
rect 16885 263965 16915 263995
rect 16725 263885 16755 263915
rect 16885 263885 16915 263915
rect 16725 263805 16755 263835
rect 16885 263805 16915 263835
rect 16725 263725 16755 263755
rect 16885 263725 16915 263755
rect 16725 263645 16755 263675
rect 16885 263645 16915 263675
rect 16725 263565 16755 263595
rect 16885 263565 16915 263595
rect 16725 263485 16755 263515
rect 16885 263485 16915 263515
rect 16725 263405 16755 263435
rect 16885 263405 16915 263435
rect 16725 263325 16755 263355
rect 16885 263325 16915 263355
rect 16725 263245 16755 263275
rect 16885 263245 16915 263275
rect 16725 263165 16755 263195
rect 16885 263165 16915 263195
rect 16725 263085 16755 263115
rect 16885 263085 16915 263115
rect 16725 263005 16755 263035
rect 16885 263005 16915 263035
rect 16725 262925 16755 262955
rect 16885 262925 16915 262955
rect 16725 262845 16755 262875
rect 16885 262845 16915 262875
rect 16725 262765 16755 262795
rect 16885 262765 16915 262795
rect 16725 262685 16755 262715
rect 16885 262685 16915 262715
rect 16725 262605 16755 262635
rect 16885 262605 16915 262635
rect 16725 262525 16755 262555
rect 16885 262525 16915 262555
rect 16725 262445 16755 262475
rect 16885 262445 16915 262475
rect 16725 262365 16755 262395
rect 16885 262365 16915 262395
rect 16725 262285 16755 262315
rect 16885 262285 16915 262315
rect 16725 262205 16755 262235
rect 16885 262205 16915 262235
rect 16725 262125 16755 262155
rect 16885 262125 16915 262155
rect 16725 262045 16755 262075
rect 16885 262045 16915 262075
rect 16725 261965 16755 261995
rect 16885 261965 16915 261995
rect 16725 261885 16755 261915
rect 16885 261885 16915 261915
rect 16725 261805 16755 261835
rect 16885 261805 16915 261835
rect 16725 261725 16755 261755
rect 16885 261725 16915 261755
rect 16725 261645 16755 261675
rect 16885 261645 16915 261675
rect 16725 261565 16755 261595
rect 16885 261565 16915 261595
rect 16725 261485 16755 261515
rect 16885 261485 16915 261515
rect 16725 261405 16755 261435
rect 16885 261405 16915 261435
rect 16725 261325 16755 261355
rect 16885 261325 16915 261355
rect 16725 261245 16755 261275
rect 16885 261245 16915 261275
rect 16725 261165 16755 261195
rect 16885 261165 16915 261195
rect 16725 261085 16755 261115
rect 16885 261085 16915 261115
rect 16725 261005 16755 261035
rect 16885 261005 16915 261035
rect 16725 260925 16755 260955
rect 16885 260925 16915 260955
rect 16725 260845 16755 260875
rect 16885 260845 16915 260875
rect 16725 260765 16755 260795
rect 16885 260765 16915 260795
rect 16725 260685 16755 260715
rect 16885 260685 16915 260715
rect 16725 260605 16755 260635
rect 16885 260605 16915 260635
rect 16725 260525 16755 260555
rect 16885 260525 16915 260555
rect 16725 260445 16755 260475
rect 16885 260445 16915 260475
rect 16725 260365 16755 260395
rect 16885 260365 16915 260395
rect 16725 260285 16755 260315
rect 16885 260285 16915 260315
rect 16725 260205 16755 260235
rect 16885 260205 16915 260235
rect 16725 260125 16755 260155
rect 16885 260125 16915 260155
rect 16725 260045 16755 260075
rect 16885 260045 16915 260075
rect 16725 259965 16755 259995
rect 16885 259965 16915 259995
rect 16725 259885 16755 259915
rect 16885 259885 16915 259915
rect 16725 259805 16755 259835
rect 16885 259805 16915 259835
rect 16725 259725 16755 259755
rect 16885 259725 16915 259755
rect 16725 259645 16755 259675
rect 16885 259645 16915 259675
rect 16725 259565 16755 259595
rect 16885 259565 16915 259595
rect 16725 259485 16755 259515
rect 16885 259485 16915 259515
rect 16725 259405 16755 259435
rect 16885 259405 16915 259435
rect 16725 259325 16755 259355
rect 16885 259325 16915 259355
rect 16725 259245 16755 259275
rect 16885 259245 16915 259275
rect 16725 259165 16755 259195
rect 16885 259165 16915 259195
rect 16725 259085 16755 259115
rect 16885 259085 16915 259115
rect 16725 259005 16755 259035
rect 16885 259005 16915 259035
rect 16725 258925 16755 258955
rect 16885 258925 16915 258955
rect 16725 258845 16755 258875
rect 16885 258845 16915 258875
rect 16725 258765 16755 258795
rect 16885 258765 16915 258795
rect 16725 258685 16755 258715
rect 16885 258685 16915 258715
rect 16725 258605 16755 258635
rect 16885 258605 16915 258635
rect 16725 258525 16755 258555
rect 16885 258525 16915 258555
rect 16725 258445 16755 258475
rect 16885 258445 16915 258475
rect 16725 258365 16755 258395
rect 16885 258365 16915 258395
rect 16725 258285 16755 258315
rect 16885 258285 16915 258315
rect 16725 258205 16755 258235
rect 16885 258205 16915 258235
rect 16725 258125 16755 258155
rect 16885 258125 16915 258155
rect 16725 258045 16755 258075
rect 16885 258045 16915 258075
rect 16725 257965 16755 257995
rect 16885 257965 16915 257995
rect 16725 257885 16755 257915
rect 16885 257885 16915 257915
rect 16725 257805 16755 257835
rect 16885 257805 16915 257835
rect 16725 257725 16755 257755
rect 16885 257725 16915 257755
rect 16725 257645 16755 257675
rect 16885 257645 16915 257675
rect 16725 257565 16755 257595
rect 16885 257565 16915 257595
rect 16725 257485 16755 257515
rect 16885 257485 16915 257515
rect 16725 257405 16755 257435
rect 16885 257405 16915 257435
rect 16725 257325 16755 257355
rect 16885 257325 16915 257355
rect 16725 257245 16755 257275
rect 16885 257245 16915 257275
rect 16725 257165 16755 257195
rect 16885 257165 16915 257195
rect 16725 257085 16755 257115
rect 16885 257085 16915 257115
rect 16725 257005 16755 257035
rect 16885 257005 16915 257035
rect 16725 256925 16755 256955
rect 16885 256925 16915 256955
rect 16725 256845 16755 256875
rect 16885 256845 16915 256875
rect 16725 256765 16755 256795
rect 16885 256765 16915 256795
rect 16725 256685 16755 256715
rect 16885 256685 16915 256715
rect 16725 256605 16755 256635
rect 16885 256605 16915 256635
rect 16725 256525 16755 256555
rect 16885 256525 16915 256555
rect 16725 256445 16755 256475
rect 16885 256445 16915 256475
rect 16725 256365 16755 256395
rect 16885 256365 16915 256395
rect 16725 256285 16755 256315
rect 16885 256285 16915 256315
rect 16725 256205 16755 256235
rect 16885 256205 16915 256235
rect 16725 256125 16755 256155
rect 16885 256125 16915 256155
rect 16725 256045 16755 256075
rect 16885 256045 16915 256075
rect 16725 255965 16755 255995
rect 16885 255965 16915 255995
rect 405 255845 435 255875
rect 485 255845 515 255875
rect 565 255845 595 255875
rect 645 255845 675 255875
rect 725 255845 755 255875
rect 805 255845 835 255875
rect 885 255845 915 255875
rect 965 255845 995 255875
rect 1045 255845 1075 255875
rect 1125 255845 1155 255875
rect 1205 255845 1235 255875
rect 1285 255845 1315 255875
rect 1365 255845 1395 255875
rect 1445 255845 1475 255875
rect 1525 255845 1555 255875
rect 1605 255845 1635 255875
rect 1685 255845 1715 255875
rect 1765 255845 1795 255875
rect 1845 255845 1875 255875
rect 1925 255845 1955 255875
rect 2005 255845 2035 255875
rect 2085 255845 2115 255875
rect 2165 255845 2195 255875
rect 2245 255845 2275 255875
rect 2325 255845 2355 255875
rect 2405 255845 2435 255875
rect 2485 255845 2515 255875
rect 2565 255845 2595 255875
rect 2645 255845 2675 255875
rect 2725 255845 2755 255875
rect 3045 255845 3075 255875
rect 3125 255845 3155 255875
rect 3205 255845 3235 255875
rect 3285 255845 3315 255875
rect 3365 255845 3395 255875
rect 3445 255845 3475 255875
rect 3525 255845 3555 255875
rect 3605 255845 3635 255875
rect 3685 255845 3715 255875
rect 3765 255845 3795 255875
rect 3845 255845 3875 255875
rect 3925 255845 3955 255875
rect 4005 255845 4035 255875
rect 4085 255845 4115 255875
rect 4165 255845 4195 255875
rect 4245 255845 4275 255875
rect 4325 255845 4355 255875
rect 4405 255845 4435 255875
rect 4485 255845 4515 255875
rect 4565 255845 4595 255875
rect 4645 255845 4675 255875
rect 4725 255845 4755 255875
rect 4805 255845 4835 255875
rect 4885 255845 4915 255875
rect 4965 255845 4995 255875
rect 5045 255845 5075 255875
rect 5125 255845 5155 255875
rect 5205 255845 5235 255875
rect 5285 255845 5315 255875
rect 5365 255845 5395 255875
rect 5445 255845 5475 255875
rect 5525 255845 5555 255875
rect 5605 255845 5635 255875
rect 5685 255845 5715 255875
rect 5765 255845 5795 255875
rect 5845 255845 5875 255875
rect 5925 255845 5955 255875
rect 6005 255845 6035 255875
rect 6085 255845 6115 255875
rect 6165 255845 6195 255875
rect 6245 255845 6275 255875
rect 6325 255845 6355 255875
rect 6405 255845 6435 255875
rect 6485 255845 6515 255875
rect 6565 255845 6595 255875
rect 6645 255845 6675 255875
rect 6725 255845 6755 255875
rect 6805 255845 6835 255875
rect 6885 255845 6915 255875
rect 6965 255845 6995 255875
rect 7045 255845 7075 255875
rect 7125 255845 7155 255875
rect 7205 255845 7235 255875
rect 7285 255845 7315 255875
rect 7365 255845 7395 255875
rect 7445 255845 7475 255875
rect 7525 255845 7555 255875
rect 7605 255845 7635 255875
rect 7685 255845 7715 255875
rect 7765 255845 7795 255875
rect 7845 255845 7875 255875
rect 7925 255845 7955 255875
rect 8005 255845 8035 255875
rect 8085 255845 8115 255875
rect 8165 255845 8195 255875
rect 8245 255845 8275 255875
rect 8325 255845 8355 255875
rect 8405 255845 8435 255875
rect 8485 255845 8515 255875
rect 8565 255845 8595 255875
rect 8645 255845 8675 255875
rect 8725 255845 8755 255875
rect 8805 255845 8835 255875
rect 8885 255845 8915 255875
rect 8965 255845 8995 255875
rect 9045 255845 9075 255875
rect 9125 255845 9155 255875
rect 9205 255845 9235 255875
rect 9285 255845 9315 255875
rect 9365 255845 9395 255875
rect 9445 255845 9475 255875
rect 9525 255845 9555 255875
rect 9605 255845 9635 255875
rect 9685 255845 9715 255875
rect 9765 255845 9795 255875
rect 9845 255845 9875 255875
rect 9925 255845 9955 255875
rect 10005 255845 10035 255875
rect 10085 255845 10115 255875
rect 10165 255845 10195 255875
rect 10245 255845 10275 255875
rect 10325 255845 10355 255875
rect 10405 255845 10435 255875
rect 10485 255845 10515 255875
rect 10565 255845 10595 255875
rect 10645 255845 10675 255875
rect 10725 255845 10755 255875
rect 10805 255845 10835 255875
rect 10885 255845 10915 255875
rect 10965 255845 10995 255875
rect 11045 255845 11075 255875
rect 11125 255845 11155 255875
rect 11205 255845 11235 255875
rect 11285 255845 11315 255875
rect 11365 255845 11395 255875
rect 11445 255845 11475 255875
rect 11525 255845 11555 255875
rect 11605 255845 11635 255875
rect 11685 255845 11715 255875
rect 11765 255845 11795 255875
rect 11845 255845 11875 255875
rect 11925 255845 11955 255875
rect 12005 255845 12035 255875
rect 12085 255845 12115 255875
rect 12165 255845 12195 255875
rect 12245 255845 12275 255875
rect 12325 255845 12355 255875
rect 12405 255845 12435 255875
rect 12485 255845 12515 255875
rect 12565 255845 12595 255875
rect 12645 255845 12675 255875
rect 12725 255845 12755 255875
rect 12805 255845 12835 255875
rect 12885 255845 12915 255875
rect 12965 255845 12995 255875
rect 13045 255845 13075 255875
rect 13125 255845 13155 255875
rect 13205 255845 13235 255875
rect 13285 255845 13315 255875
rect 13365 255845 13395 255875
rect 13445 255845 13475 255875
rect 13525 255845 13555 255875
rect 13605 255845 13635 255875
rect 13685 255845 13715 255875
rect 13765 255845 13795 255875
rect 13845 255845 13875 255875
rect 13925 255845 13955 255875
rect 14005 255845 14035 255875
rect 14085 255845 14115 255875
rect 14165 255845 14195 255875
rect 14245 255845 14275 255875
rect 14325 255845 14355 255875
rect 14405 255845 14435 255875
rect 14485 255845 14515 255875
rect 14565 255845 14595 255875
rect 14645 255845 14675 255875
rect 14725 255845 14755 255875
rect 14805 255845 14835 255875
rect 14885 255845 14915 255875
rect 14965 255845 14995 255875
rect 15045 255845 15075 255875
rect 15125 255845 15155 255875
rect 15205 255845 15235 255875
rect 15285 255845 15315 255875
rect 15365 255845 15395 255875
rect 15445 255845 15475 255875
rect 15525 255845 15555 255875
rect 15605 255845 15635 255875
rect 15685 255845 15715 255875
rect 15765 255845 15795 255875
rect 15845 255845 15875 255875
rect 15925 255845 15955 255875
rect 16005 255845 16035 255875
rect 16085 255845 16115 255875
rect 16165 255845 16195 255875
rect 16245 255845 16275 255875
rect 16325 255845 16355 255875
rect 16405 255845 16435 255875
rect 16485 255845 16515 255875
rect 16565 255845 16595 255875
rect 16645 255845 16675 255875
rect 16725 255845 16755 255875
rect 16885 255845 16915 255875
rect 405 255685 435 255715
rect 485 255685 515 255715
rect 565 255685 595 255715
rect 645 255685 675 255715
rect 725 255685 755 255715
rect 805 255685 835 255715
rect 885 255685 915 255715
rect 965 255685 995 255715
rect 1045 255685 1075 255715
rect 1125 255685 1155 255715
rect 1205 255685 1235 255715
rect 1285 255685 1315 255715
rect 1365 255685 1395 255715
rect 1445 255685 1475 255715
rect 1525 255685 1555 255715
rect 1605 255685 1635 255715
rect 1685 255685 1715 255715
rect 1765 255685 1795 255715
rect 1845 255685 1875 255715
rect 1925 255685 1955 255715
rect 2005 255685 2035 255715
rect 2085 255685 2115 255715
rect 2165 255685 2195 255715
rect 2245 255685 2275 255715
rect 2325 255685 2355 255715
rect 2405 255685 2435 255715
rect 2485 255685 2515 255715
rect 2565 255685 2595 255715
rect 2645 255685 2675 255715
rect 2725 255685 2755 255715
rect 3045 255685 3075 255715
rect 3125 255685 3155 255715
rect 3205 255685 3235 255715
rect 3285 255685 3315 255715
rect 3365 255685 3395 255715
rect 3445 255685 3475 255715
rect 3525 255685 3555 255715
rect 3605 255685 3635 255715
rect 3685 255685 3715 255715
rect 3765 255685 3795 255715
rect 3845 255685 3875 255715
rect 3925 255685 3955 255715
rect 4005 255685 4035 255715
rect 4085 255685 4115 255715
rect 4165 255685 4195 255715
rect 4245 255685 4275 255715
rect 4325 255685 4355 255715
rect 4405 255685 4435 255715
rect 4485 255685 4515 255715
rect 4565 255685 4595 255715
rect 4645 255685 4675 255715
rect 4725 255685 4755 255715
rect 4805 255685 4835 255715
rect 4885 255685 4915 255715
rect 4965 255685 4995 255715
rect 5045 255685 5075 255715
rect 5125 255685 5155 255715
rect 5205 255685 5235 255715
rect 5285 255685 5315 255715
rect 5365 255685 5395 255715
rect 5445 255685 5475 255715
rect 5525 255685 5555 255715
rect 5605 255685 5635 255715
rect 5685 255685 5715 255715
rect 5765 255685 5795 255715
rect 5845 255685 5875 255715
rect 5925 255685 5955 255715
rect 6005 255685 6035 255715
rect 6085 255685 6115 255715
rect 6165 255685 6195 255715
rect 6245 255685 6275 255715
rect 6325 255685 6355 255715
rect 6405 255685 6435 255715
rect 6485 255685 6515 255715
rect 6565 255685 6595 255715
rect 6645 255685 6675 255715
rect 6725 255685 6755 255715
rect 6805 255685 6835 255715
rect 6885 255685 6915 255715
rect 6965 255685 6995 255715
rect 7045 255685 7075 255715
rect 7125 255685 7155 255715
rect 7205 255685 7235 255715
rect 7285 255685 7315 255715
rect 7365 255685 7395 255715
rect 7445 255685 7475 255715
rect 7525 255685 7555 255715
rect 7605 255685 7635 255715
rect 7685 255685 7715 255715
rect 7765 255685 7795 255715
rect 7845 255685 7875 255715
rect 7925 255685 7955 255715
rect 8005 255685 8035 255715
rect 8085 255685 8115 255715
rect 8165 255685 8195 255715
rect 8245 255685 8275 255715
rect 8325 255685 8355 255715
rect 8405 255685 8435 255715
rect 8485 255685 8515 255715
rect 8565 255685 8595 255715
rect 8645 255685 8675 255715
rect 8725 255685 8755 255715
rect 8805 255685 8835 255715
rect 8885 255685 8915 255715
rect 8965 255685 8995 255715
rect 9045 255685 9075 255715
rect 9125 255685 9155 255715
rect 9205 255685 9235 255715
rect 9285 255685 9315 255715
rect 9365 255685 9395 255715
rect 9445 255685 9475 255715
rect 9525 255685 9555 255715
rect 9605 255685 9635 255715
rect 9685 255685 9715 255715
rect 9765 255685 9795 255715
rect 9845 255685 9875 255715
rect 9925 255685 9955 255715
rect 10005 255685 10035 255715
rect 10085 255685 10115 255715
rect 10165 255685 10195 255715
rect 10245 255685 10275 255715
rect 10325 255685 10355 255715
rect 10405 255685 10435 255715
rect 10485 255685 10515 255715
rect 10565 255685 10595 255715
rect 10645 255685 10675 255715
rect 10725 255685 10755 255715
rect 10805 255685 10835 255715
rect 10885 255685 10915 255715
rect 10965 255685 10995 255715
rect 11045 255685 11075 255715
rect 11125 255685 11155 255715
rect 11205 255685 11235 255715
rect 11285 255685 11315 255715
rect 11365 255685 11395 255715
rect 11445 255685 11475 255715
rect 11525 255685 11555 255715
rect 11605 255685 11635 255715
rect 11685 255685 11715 255715
rect 11765 255685 11795 255715
rect 11845 255685 11875 255715
rect 11925 255685 11955 255715
rect 12005 255685 12035 255715
rect 12085 255685 12115 255715
rect 12165 255685 12195 255715
rect 12245 255685 12275 255715
rect 12325 255685 12355 255715
rect 12405 255685 12435 255715
rect 12485 255685 12515 255715
rect 12565 255685 12595 255715
rect 12645 255685 12675 255715
rect 12725 255685 12755 255715
rect 12805 255685 12835 255715
rect 12885 255685 12915 255715
rect 12965 255685 12995 255715
rect 13045 255685 13075 255715
rect 13125 255685 13155 255715
rect 13205 255685 13235 255715
rect 13285 255685 13315 255715
rect 13365 255685 13395 255715
rect 13445 255685 13475 255715
rect 13525 255685 13555 255715
rect 13605 255685 13635 255715
rect 13685 255685 13715 255715
rect 13765 255685 13795 255715
rect 13845 255685 13875 255715
rect 13925 255685 13955 255715
rect 14005 255685 14035 255715
rect 14085 255685 14115 255715
rect 14165 255685 14195 255715
rect 14245 255685 14275 255715
rect 14325 255685 14355 255715
rect 14405 255685 14435 255715
rect 14485 255685 14515 255715
rect 14565 255685 14595 255715
rect 14645 255685 14675 255715
rect 14725 255685 14755 255715
rect 14805 255685 14835 255715
rect 14885 255685 14915 255715
rect 14965 255685 14995 255715
rect 15045 255685 15075 255715
rect 15125 255685 15155 255715
rect 15205 255685 15235 255715
rect 15285 255685 15315 255715
rect 15365 255685 15395 255715
rect 15445 255685 15475 255715
rect 15525 255685 15555 255715
rect 15605 255685 15635 255715
rect 15685 255685 15715 255715
rect 15765 255685 15795 255715
rect 15845 255685 15875 255715
rect 15925 255685 15955 255715
rect 16005 255685 16035 255715
rect 16085 255685 16115 255715
rect 16165 255685 16195 255715
rect 16245 255685 16275 255715
rect 16325 255685 16355 255715
rect 16405 255685 16435 255715
rect 16485 255685 16515 255715
rect 16565 255685 16595 255715
rect 16645 255685 16675 255715
rect 16725 255685 16755 255715
rect 16885 255685 16915 255715
<< metal2 >>
rect 271860 351815 283220 351820
rect 271860 351785 271865 351815
rect 271895 351785 272025 351815
rect 272055 351785 272105 351815
rect 272135 351785 272185 351815
rect 272215 351785 272265 351815
rect 272295 351785 272345 351815
rect 272375 351785 272425 351815
rect 272455 351785 272505 351815
rect 272535 351785 272585 351815
rect 272615 351785 272665 351815
rect 272695 351785 272745 351815
rect 272775 351785 272825 351815
rect 272855 351785 272905 351815
rect 272935 351785 272985 351815
rect 273015 351785 273065 351815
rect 273095 351785 273145 351815
rect 273175 351785 273225 351815
rect 273255 351785 273305 351815
rect 273335 351785 273385 351815
rect 273415 351785 273465 351815
rect 273495 351785 273545 351815
rect 273575 351785 273625 351815
rect 273655 351785 273705 351815
rect 273735 351785 273785 351815
rect 273815 351785 273865 351815
rect 273895 351785 273945 351815
rect 273975 351785 274025 351815
rect 274055 351785 274105 351815
rect 274135 351785 274185 351815
rect 274215 351785 274265 351815
rect 274295 351785 274345 351815
rect 274375 351785 274425 351815
rect 274455 351785 274505 351815
rect 274535 351785 274585 351815
rect 274615 351785 274665 351815
rect 274695 351785 274745 351815
rect 274775 351785 274825 351815
rect 274855 351785 274905 351815
rect 274935 351785 274985 351815
rect 275015 351785 275065 351815
rect 275095 351785 275145 351815
rect 275175 351785 275225 351815
rect 275255 351785 275305 351815
rect 275335 351785 275385 351815
rect 275415 351785 275465 351815
rect 275495 351785 275545 351815
rect 275575 351785 275625 351815
rect 275655 351785 275705 351815
rect 275735 351785 275785 351815
rect 275815 351785 275865 351815
rect 275895 351785 275945 351815
rect 275975 351785 276025 351815
rect 276055 351785 276105 351815
rect 276135 351785 276185 351815
rect 276215 351785 276265 351815
rect 276295 351785 276345 351815
rect 276375 351785 276425 351815
rect 276455 351785 276505 351815
rect 276535 351785 276585 351815
rect 276615 351785 276665 351815
rect 276695 351785 276745 351815
rect 276775 351785 276825 351815
rect 276855 351785 276905 351815
rect 276935 351785 276985 351815
rect 277015 351785 277065 351815
rect 277095 351785 277145 351815
rect 277175 351785 277225 351815
rect 277255 351785 277305 351815
rect 277335 351785 277385 351815
rect 277415 351785 277465 351815
rect 277495 351785 277545 351815
rect 277575 351785 277625 351815
rect 277655 351785 277705 351815
rect 277735 351785 277785 351815
rect 277815 351785 277865 351815
rect 277895 351785 277945 351815
rect 277975 351785 278025 351815
rect 278055 351785 278105 351815
rect 278135 351785 278185 351815
rect 278215 351785 278265 351815
rect 278295 351785 278345 351815
rect 278375 351785 278425 351815
rect 278455 351785 278505 351815
rect 278535 351785 278585 351815
rect 278615 351785 278665 351815
rect 278695 351785 278745 351815
rect 278775 351785 278825 351815
rect 278855 351785 278905 351815
rect 278935 351785 278985 351815
rect 279015 351785 279065 351815
rect 279095 351785 279145 351815
rect 279175 351785 279225 351815
rect 279255 351785 279305 351815
rect 279335 351785 279385 351815
rect 279415 351785 279465 351815
rect 279495 351785 279545 351815
rect 279575 351785 279625 351815
rect 279655 351785 279705 351815
rect 279735 351785 279785 351815
rect 279815 351785 279865 351815
rect 279895 351785 279945 351815
rect 279975 351785 280025 351815
rect 280055 351785 280105 351815
rect 280135 351785 280185 351815
rect 280215 351785 280265 351815
rect 280295 351785 280345 351815
rect 280375 351785 280425 351815
rect 280455 351785 280505 351815
rect 280535 351785 280585 351815
rect 280615 351785 280665 351815
rect 280695 351785 280745 351815
rect 280775 351785 280825 351815
rect 280855 351785 280905 351815
rect 280935 351785 280985 351815
rect 281015 351785 281065 351815
rect 281095 351785 281145 351815
rect 281175 351785 281225 351815
rect 281255 351785 281305 351815
rect 281335 351785 281385 351815
rect 281415 351785 281465 351815
rect 281495 351785 281545 351815
rect 281575 351785 281625 351815
rect 281655 351785 281705 351815
rect 281735 351785 281785 351815
rect 281815 351785 281865 351815
rect 281895 351785 281945 351815
rect 281975 351785 282025 351815
rect 282055 351785 282105 351815
rect 282135 351785 282185 351815
rect 282215 351785 282265 351815
rect 282295 351785 282345 351815
rect 282375 351785 282425 351815
rect 282455 351785 282505 351815
rect 282535 351785 282585 351815
rect 282615 351785 282665 351815
rect 282695 351785 282745 351815
rect 282775 351785 282825 351815
rect 282855 351785 282905 351815
rect 282935 351785 282985 351815
rect 283015 351785 283065 351815
rect 283095 351785 283145 351815
rect 283175 351785 283220 351815
rect 271860 351780 283220 351785
rect 271940 351735 283260 351740
rect 271940 351705 271945 351735
rect 271975 351705 283225 351735
rect 283255 351705 283260 351735
rect 271940 351700 283260 351705
rect 271860 351655 283220 351660
rect 271860 351625 271865 351655
rect 271895 351625 272025 351655
rect 272055 351625 272105 351655
rect 272135 351625 272185 351655
rect 272215 351625 272265 351655
rect 272295 351625 272345 351655
rect 272375 351625 272425 351655
rect 272455 351625 272505 351655
rect 272535 351625 272585 351655
rect 272615 351625 272665 351655
rect 272695 351625 272745 351655
rect 272775 351625 272825 351655
rect 272855 351625 272905 351655
rect 272935 351625 272985 351655
rect 273015 351625 273065 351655
rect 273095 351625 273145 351655
rect 273175 351625 273225 351655
rect 273255 351625 273305 351655
rect 273335 351625 273385 351655
rect 273415 351625 273465 351655
rect 273495 351625 273545 351655
rect 273575 351625 273625 351655
rect 273655 351625 273705 351655
rect 273735 351625 273785 351655
rect 273815 351625 273865 351655
rect 273895 351625 273945 351655
rect 273975 351625 274025 351655
rect 274055 351625 274105 351655
rect 274135 351625 274185 351655
rect 274215 351625 274265 351655
rect 274295 351625 274345 351655
rect 274375 351625 274425 351655
rect 274455 351625 274505 351655
rect 274535 351625 274585 351655
rect 274615 351625 274665 351655
rect 274695 351625 274745 351655
rect 274775 351625 274825 351655
rect 274855 351625 274905 351655
rect 274935 351625 274985 351655
rect 275015 351625 275065 351655
rect 275095 351625 275145 351655
rect 275175 351625 275225 351655
rect 275255 351625 275305 351655
rect 275335 351625 275385 351655
rect 275415 351625 275465 351655
rect 275495 351625 275545 351655
rect 275575 351625 275625 351655
rect 275655 351625 275705 351655
rect 275735 351625 275785 351655
rect 275815 351625 275865 351655
rect 275895 351625 275945 351655
rect 275975 351625 276025 351655
rect 276055 351625 276105 351655
rect 276135 351625 276185 351655
rect 276215 351625 276265 351655
rect 276295 351625 276345 351655
rect 276375 351625 276425 351655
rect 276455 351625 276505 351655
rect 276535 351625 276585 351655
rect 276615 351625 276665 351655
rect 276695 351625 276745 351655
rect 276775 351625 276825 351655
rect 276855 351625 276905 351655
rect 276935 351625 276985 351655
rect 277015 351625 277065 351655
rect 277095 351625 277145 351655
rect 277175 351625 277225 351655
rect 277255 351625 277305 351655
rect 277335 351625 277385 351655
rect 277415 351625 277465 351655
rect 277495 351625 277545 351655
rect 277575 351625 277625 351655
rect 277655 351625 277705 351655
rect 277735 351625 277785 351655
rect 277815 351625 277865 351655
rect 277895 351625 277945 351655
rect 277975 351625 278025 351655
rect 278055 351625 278105 351655
rect 278135 351625 278185 351655
rect 278215 351625 278265 351655
rect 278295 351625 278345 351655
rect 278375 351625 278425 351655
rect 278455 351625 278505 351655
rect 278535 351625 278585 351655
rect 278615 351625 278665 351655
rect 278695 351625 278745 351655
rect 278775 351625 278825 351655
rect 278855 351625 278905 351655
rect 278935 351625 278985 351655
rect 279015 351625 279065 351655
rect 279095 351625 279145 351655
rect 279175 351625 279225 351655
rect 279255 351625 279305 351655
rect 279335 351625 279385 351655
rect 279415 351625 279465 351655
rect 279495 351625 279545 351655
rect 279575 351625 279625 351655
rect 279655 351625 279705 351655
rect 279735 351625 279785 351655
rect 279815 351625 279865 351655
rect 279895 351625 279945 351655
rect 279975 351625 280025 351655
rect 280055 351625 280105 351655
rect 280135 351625 280185 351655
rect 280215 351625 280265 351655
rect 280295 351625 280345 351655
rect 280375 351625 280425 351655
rect 280455 351625 280505 351655
rect 280535 351625 280585 351655
rect 280615 351625 280665 351655
rect 280695 351625 280745 351655
rect 280775 351625 280825 351655
rect 280855 351625 280905 351655
rect 280935 351625 280985 351655
rect 281015 351625 281065 351655
rect 281095 351625 281145 351655
rect 281175 351625 281225 351655
rect 281255 351625 281305 351655
rect 281335 351625 281385 351655
rect 281415 351625 281465 351655
rect 281495 351625 281545 351655
rect 281575 351625 281625 351655
rect 281655 351625 281705 351655
rect 281735 351625 281785 351655
rect 281815 351625 281865 351655
rect 281895 351625 281945 351655
rect 281975 351625 282025 351655
rect 282055 351625 282105 351655
rect 282135 351625 282185 351655
rect 282215 351625 282265 351655
rect 282295 351625 282345 351655
rect 282375 351625 282425 351655
rect 282455 351625 282505 351655
rect 282535 351625 282585 351655
rect 282615 351625 282665 351655
rect 282695 351625 282745 351655
rect 282775 351625 282825 351655
rect 282855 351625 282905 351655
rect 282935 351625 282985 351655
rect 283015 351625 283065 351655
rect 283095 351625 283145 351655
rect 283175 351625 283220 351655
rect 271860 351620 283220 351625
rect 271860 351575 272060 351580
rect 271860 351545 271865 351575
rect 271895 351545 272025 351575
rect 272055 351545 272060 351575
rect 271860 351540 272060 351545
rect 271860 351495 272060 351500
rect 271860 351465 271865 351495
rect 271895 351465 272025 351495
rect 272055 351465 272060 351495
rect 271860 351460 272060 351465
rect 271860 351415 272060 351420
rect 271860 351385 271865 351415
rect 271895 351385 272025 351415
rect 272055 351385 272060 351415
rect 271860 351380 272060 351385
rect 271860 351335 272060 351340
rect 271860 351305 271865 351335
rect 271895 351305 272025 351335
rect 272055 351305 272060 351335
rect 271860 351300 272060 351305
rect 271860 351255 272060 351260
rect 271860 351225 271865 351255
rect 271895 351225 272025 351255
rect 272055 351225 272060 351255
rect 271860 351220 272060 351225
rect 271860 351175 272060 351180
rect 271860 351145 271865 351175
rect 271895 351145 272025 351175
rect 272055 351145 272060 351175
rect 271860 351140 272060 351145
rect 271860 351095 272060 351100
rect 271860 351065 271865 351095
rect 271895 351065 272025 351095
rect 272055 351065 272060 351095
rect 271860 351060 272060 351065
rect 271860 351015 272060 351020
rect 271860 350985 271865 351015
rect 271895 350985 272025 351015
rect 272055 350985 272060 351015
rect 271860 350980 272060 350985
rect 271860 350935 272060 350940
rect 271860 350905 271865 350935
rect 271895 350905 272025 350935
rect 272055 350905 272060 350935
rect 271860 350900 272060 350905
rect 271860 350855 272060 350860
rect 271860 350825 271865 350855
rect 271895 350825 272025 350855
rect 272055 350825 272060 350855
rect 271860 350820 272060 350825
rect 271860 350775 272060 350780
rect 271860 350745 271865 350775
rect 271895 350745 272025 350775
rect 272055 350745 272060 350775
rect 271860 350740 272060 350745
rect 271860 350695 272060 350700
rect 271860 350665 271865 350695
rect 271895 350665 272025 350695
rect 272055 350665 272060 350695
rect 271860 350660 272060 350665
rect 271860 350615 272060 350620
rect 271860 350585 271865 350615
rect 271895 350585 272025 350615
rect 272055 350585 272060 350615
rect 271860 350580 272060 350585
rect 271860 350535 272060 350540
rect 271860 350505 271865 350535
rect 271895 350505 272025 350535
rect 272055 350505 272060 350535
rect 271860 350500 272060 350505
rect 271860 350455 272060 350460
rect 271860 350425 271865 350455
rect 271895 350425 272025 350455
rect 272055 350425 272060 350455
rect 271860 350420 272060 350425
rect 271860 350375 272060 350380
rect 271860 350345 271865 350375
rect 271895 350345 272025 350375
rect 272055 350345 272060 350375
rect 271860 350340 272060 350345
rect 271860 350295 272060 350300
rect 271860 350265 271865 350295
rect 271895 350265 272025 350295
rect 272055 350265 272060 350295
rect 271860 350260 272060 350265
rect 271860 350215 272060 350220
rect 271860 350185 271865 350215
rect 271895 350185 272025 350215
rect 272055 350185 272060 350215
rect 271860 350180 272060 350185
rect 271860 350135 272060 350140
rect 271860 350105 271865 350135
rect 271895 350105 272025 350135
rect 272055 350105 272060 350135
rect 271860 350100 272060 350105
rect 271860 350055 272060 350060
rect 271860 350025 271865 350055
rect 271895 350025 272025 350055
rect 272055 350025 272060 350055
rect 271860 350020 272060 350025
rect 16720 275475 17240 275480
rect 16720 275445 16725 275475
rect 16755 275445 16885 275475
rect 16915 275445 16965 275475
rect 16995 275445 17045 275475
rect 17075 275445 17125 275475
rect 17155 275445 17205 275475
rect 17235 275445 17240 275475
rect 16720 275440 17240 275445
rect 16720 275395 17240 275400
rect 16720 275365 16805 275395
rect 16835 275365 17125 275395
rect 17155 275365 17240 275395
rect 16720 275360 17240 275365
rect 28400 275355 28760 275360
rect 28400 275325 28405 275355
rect 28435 275325 28565 275355
rect 28595 275325 28725 275355
rect 28755 275325 28760 275355
rect 28400 275320 28760 275325
rect 16720 275315 17240 275320
rect 16720 275285 16725 275315
rect 16755 275285 16885 275315
rect 16915 275285 16965 275315
rect 16995 275285 17045 275315
rect 17075 275285 17205 275315
rect 17235 275285 17240 275315
rect 16720 275280 17240 275285
rect 28400 275275 28760 275280
rect 28400 275245 28405 275275
rect 28435 275245 28565 275275
rect 28595 275245 28725 275275
rect 28755 275245 28760 275275
rect 28400 275240 28760 275245
rect 1000 275195 259100 275200
rect 1000 275160 13525 275195
rect 1000 275040 1040 275160
rect 1160 275040 13525 275160
rect 1000 275005 13525 275040
rect 13555 275005 13685 275195
rect 13715 275005 13845 275195
rect 13875 275005 14005 275195
rect 14035 275005 14165 275195
rect 14195 275005 14325 275195
rect 14355 275005 27925 275195
rect 27955 275005 28085 275195
rect 28115 275005 28245 275195
rect 28275 275005 28405 275195
rect 28435 275005 28565 275195
rect 28595 275005 28725 275195
rect 28755 275190 259100 275195
rect 28755 275010 258910 275190
rect 259090 275010 259100 275190
rect 28755 275005 259100 275010
rect 1000 275000 259100 275005
rect 16720 274955 16920 274960
rect 16720 274925 16725 274955
rect 16755 274925 16885 274955
rect 16915 274925 16920 274955
rect 16720 274920 16920 274925
rect 16720 274875 16920 274880
rect 16720 274845 16725 274875
rect 16755 274845 16885 274875
rect 16915 274845 16920 274875
rect 16720 274840 16920 274845
rect 16720 274795 16920 274800
rect 16720 274765 16725 274795
rect 16755 274765 16885 274795
rect 16915 274765 16920 274795
rect 16720 274760 16920 274765
rect 16720 274715 16920 274720
rect 16720 274685 16725 274715
rect 16755 274685 16885 274715
rect 16915 274685 16920 274715
rect 16720 274680 16920 274685
rect 16720 274635 16920 274640
rect 16720 274605 16725 274635
rect 16755 274605 16885 274635
rect 16915 274605 16920 274635
rect 16720 274600 16920 274605
rect 16720 274555 16920 274560
rect 16720 274525 16725 274555
rect 16755 274525 16885 274555
rect 16915 274525 16920 274555
rect 16720 274520 16920 274525
rect 16720 274475 16920 274480
rect 16720 274445 16725 274475
rect 16755 274445 16885 274475
rect 16915 274445 16920 274475
rect 16720 274440 16920 274445
rect 16720 274395 16920 274400
rect 16720 274365 16725 274395
rect 16755 274365 16885 274395
rect 16915 274365 16920 274395
rect 16720 274360 16920 274365
rect 16720 274315 16920 274320
rect 16720 274285 16725 274315
rect 16755 274285 16885 274315
rect 16915 274285 16920 274315
rect 16720 274280 16920 274285
rect 16720 274235 16920 274240
rect 16720 274205 16725 274235
rect 16755 274205 16885 274235
rect 16915 274205 16920 274235
rect 16720 274200 16920 274205
rect 16720 274155 16920 274160
rect 16720 274125 16725 274155
rect 16755 274125 16885 274155
rect 16915 274125 16920 274155
rect 16720 274120 16920 274125
rect 16720 274075 16920 274080
rect 16720 274045 16725 274075
rect 16755 274045 16885 274075
rect 16915 274045 16920 274075
rect 16720 274040 16920 274045
rect 16720 273995 16920 274000
rect 16720 273965 16725 273995
rect 16755 273965 16885 273995
rect 16915 273965 16920 273995
rect 16720 273960 16920 273965
rect 16720 273915 16920 273920
rect 16720 273885 16725 273915
rect 16755 273885 16885 273915
rect 16915 273885 16920 273915
rect 16720 273880 16920 273885
rect 16720 273835 16920 273840
rect 16720 273805 16725 273835
rect 16755 273805 16885 273835
rect 16915 273805 16920 273835
rect 16720 273800 16920 273805
rect 16720 273755 16920 273760
rect 16720 273725 16725 273755
rect 16755 273725 16885 273755
rect 16915 273725 16920 273755
rect 16720 273720 16920 273725
rect 16720 273675 16920 273680
rect 16720 273645 16725 273675
rect 16755 273645 16885 273675
rect 16915 273645 16920 273675
rect 16720 273640 16920 273645
rect 16720 273595 16920 273600
rect 16720 273565 16725 273595
rect 16755 273565 16885 273595
rect 16915 273565 16920 273595
rect 16720 273560 16920 273565
rect 16720 273515 16920 273520
rect 16720 273485 16725 273515
rect 16755 273485 16885 273515
rect 16915 273485 16920 273515
rect 16720 273480 16920 273485
rect 16720 273435 16920 273440
rect 16720 273405 16725 273435
rect 16755 273405 16885 273435
rect 16915 273405 16920 273435
rect 16720 273400 16920 273405
rect 16720 273355 16920 273360
rect 16720 273325 16725 273355
rect 16755 273325 16885 273355
rect 16915 273325 16920 273355
rect 16720 273320 16920 273325
rect 16720 273275 16920 273280
rect 16720 273245 16725 273275
rect 16755 273245 16885 273275
rect 16915 273245 16920 273275
rect 16720 273240 16920 273245
rect 16720 273195 16920 273200
rect 16720 273165 16725 273195
rect 16755 273165 16885 273195
rect 16915 273165 16920 273195
rect 16720 273160 16920 273165
rect 16720 273115 16920 273120
rect 16720 273085 16725 273115
rect 16755 273085 16885 273115
rect 16915 273085 16920 273115
rect 16720 273080 16920 273085
rect 16720 273035 16920 273040
rect 16720 273005 16725 273035
rect 16755 273005 16885 273035
rect 16915 273005 16920 273035
rect 16720 273000 16920 273005
rect 16720 272955 16920 272960
rect 16720 272925 16725 272955
rect 16755 272925 16885 272955
rect 16915 272925 16920 272955
rect 16720 272920 16920 272925
rect 16720 272875 16920 272880
rect 16720 272845 16725 272875
rect 16755 272845 16885 272875
rect 16915 272845 16920 272875
rect 16720 272840 16920 272845
rect 16720 272795 16920 272800
rect 16720 272765 16725 272795
rect 16755 272765 16885 272795
rect 16915 272765 16920 272795
rect 16720 272760 16920 272765
rect 16720 272715 16920 272720
rect 16720 272685 16725 272715
rect 16755 272685 16885 272715
rect 16915 272685 16920 272715
rect 16720 272680 16920 272685
rect 16720 272635 16920 272640
rect 16720 272605 16725 272635
rect 16755 272605 16885 272635
rect 16915 272605 16920 272635
rect 16720 272600 16920 272605
rect 16720 272555 16920 272560
rect 16720 272525 16725 272555
rect 16755 272525 16885 272555
rect 16915 272525 16920 272555
rect 16720 272520 16920 272525
rect 16720 272475 16920 272480
rect 16720 272445 16725 272475
rect 16755 272445 16885 272475
rect 16915 272445 16920 272475
rect 16720 272440 16920 272445
rect 16720 272395 16920 272400
rect 16720 272365 16725 272395
rect 16755 272365 16885 272395
rect 16915 272365 16920 272395
rect 16720 272360 16920 272365
rect 16720 272315 16920 272320
rect 16720 272285 16725 272315
rect 16755 272285 16885 272315
rect 16915 272285 16920 272315
rect 16720 272280 16920 272285
rect 16720 272235 16920 272240
rect 16720 272205 16725 272235
rect 16755 272205 16885 272235
rect 16915 272205 16920 272235
rect 16720 272200 16920 272205
rect 16720 272155 16920 272160
rect 16720 272125 16725 272155
rect 16755 272125 16885 272155
rect 16915 272125 16920 272155
rect 16720 272120 16920 272125
rect 16720 272075 16920 272080
rect 16720 272045 16725 272075
rect 16755 272045 16885 272075
rect 16915 272045 16920 272075
rect 16720 272040 16920 272045
rect 16720 271995 16920 272000
rect 16720 271965 16725 271995
rect 16755 271965 16885 271995
rect 16915 271965 16920 271995
rect 16720 271960 16920 271965
rect 16720 271915 16920 271920
rect 16720 271885 16725 271915
rect 16755 271885 16885 271915
rect 16915 271885 16920 271915
rect 16720 271880 16920 271885
rect 16720 271835 16920 271840
rect 16720 271805 16725 271835
rect 16755 271805 16885 271835
rect 16915 271805 16920 271835
rect 16720 271800 16920 271805
rect 16720 271755 16920 271760
rect 16720 271725 16725 271755
rect 16755 271725 16885 271755
rect 16915 271725 16920 271755
rect 16720 271720 16920 271725
rect 16720 271675 16920 271680
rect 16720 271645 16725 271675
rect 16755 271645 16885 271675
rect 16915 271645 16920 271675
rect 16720 271640 16920 271645
rect 16720 271595 16920 271600
rect 16720 271565 16725 271595
rect 16755 271565 16885 271595
rect 16915 271565 16920 271595
rect 16720 271560 16920 271565
rect 16720 271515 16920 271520
rect 16720 271485 16725 271515
rect 16755 271485 16885 271515
rect 16915 271485 16920 271515
rect 16720 271480 16920 271485
rect 16720 271435 16920 271440
rect 16720 271405 16725 271435
rect 16755 271405 16885 271435
rect 16915 271405 16920 271435
rect 16720 271400 16920 271405
rect 16720 271355 16920 271360
rect 16720 271325 16725 271355
rect 16755 271325 16885 271355
rect 16915 271325 16920 271355
rect 16720 271320 16920 271325
rect 16720 271275 16920 271280
rect 16720 271245 16725 271275
rect 16755 271245 16885 271275
rect 16915 271245 16920 271275
rect 16720 271240 16920 271245
rect 16720 271195 16920 271200
rect 16720 271165 16725 271195
rect 16755 271165 16885 271195
rect 16915 271165 16920 271195
rect 16720 271160 16920 271165
rect 16720 271115 16920 271120
rect 16720 271085 16725 271115
rect 16755 271085 16885 271115
rect 16915 271085 16920 271115
rect 16720 271080 16920 271085
rect 16720 271035 16920 271040
rect 16720 271005 16725 271035
rect 16755 271005 16885 271035
rect 16915 271005 16920 271035
rect 16720 271000 16920 271005
rect 16720 270955 16920 270960
rect 16720 270925 16725 270955
rect 16755 270925 16885 270955
rect 16915 270925 16920 270955
rect 16720 270920 16920 270925
rect 16720 270875 16920 270880
rect 16720 270845 16725 270875
rect 16755 270845 16885 270875
rect 16915 270845 16920 270875
rect 16720 270840 16920 270845
rect 16720 270795 16920 270800
rect 16720 270765 16725 270795
rect 16755 270765 16885 270795
rect 16915 270765 16920 270795
rect 16720 270760 16920 270765
rect 16720 270715 16920 270720
rect 16720 270685 16725 270715
rect 16755 270685 16885 270715
rect 16915 270685 16920 270715
rect 16720 270680 16920 270685
rect 16720 270635 16920 270640
rect 16720 270605 16725 270635
rect 16755 270605 16885 270635
rect 16915 270605 16920 270635
rect 16720 270600 16920 270605
rect 16720 270555 16920 270560
rect 16720 270525 16725 270555
rect 16755 270525 16885 270555
rect 16915 270525 16920 270555
rect 16720 270520 16920 270525
rect 16720 270475 16920 270480
rect 16720 270445 16725 270475
rect 16755 270445 16885 270475
rect 16915 270445 16920 270475
rect 16720 270440 16920 270445
rect 16720 270395 16920 270400
rect 16720 270365 16725 270395
rect 16755 270365 16885 270395
rect 16915 270365 16920 270395
rect 16720 270360 16920 270365
rect 16720 270315 16920 270320
rect 16720 270285 16725 270315
rect 16755 270285 16885 270315
rect 16915 270285 16920 270315
rect 16720 270280 16920 270285
rect 16720 270235 16920 270240
rect 16720 270205 16725 270235
rect 16755 270205 16885 270235
rect 16915 270205 16920 270235
rect 16720 270200 16920 270205
rect 16720 270155 16920 270160
rect 16720 270125 16725 270155
rect 16755 270125 16885 270155
rect 16915 270125 16920 270155
rect 16720 270120 16920 270125
rect 16720 270075 16920 270080
rect 16720 270045 16725 270075
rect 16755 270045 16885 270075
rect 16915 270045 16920 270075
rect 16720 270040 16920 270045
rect 16720 269995 16920 270000
rect 16720 269965 16725 269995
rect 16755 269965 16885 269995
rect 16915 269965 16920 269995
rect 16720 269960 16920 269965
rect 16720 269915 16920 269920
rect 16720 269885 16725 269915
rect 16755 269885 16885 269915
rect 16915 269885 16920 269915
rect 16720 269880 16920 269885
rect 16720 269835 16920 269840
rect 16720 269805 16725 269835
rect 16755 269805 16885 269835
rect 16915 269805 16920 269835
rect 16720 269800 16920 269805
rect 16720 269755 16920 269760
rect 16720 269725 16725 269755
rect 16755 269725 16885 269755
rect 16915 269725 16920 269755
rect 16720 269720 16920 269725
rect 16720 269675 16920 269680
rect 16720 269645 16725 269675
rect 16755 269645 16885 269675
rect 16915 269645 16920 269675
rect 16720 269640 16920 269645
rect 16720 269595 16920 269600
rect 16720 269565 16725 269595
rect 16755 269565 16885 269595
rect 16915 269565 16920 269595
rect 16720 269560 16920 269565
rect 16720 269515 16920 269520
rect 16720 269485 16725 269515
rect 16755 269485 16885 269515
rect 16915 269485 16920 269515
rect 16720 269480 16920 269485
rect 16720 269435 16920 269440
rect 16720 269405 16725 269435
rect 16755 269405 16885 269435
rect 16915 269405 16920 269435
rect 16720 269400 16920 269405
rect 16720 269355 16920 269360
rect 16720 269325 16725 269355
rect 16755 269325 16885 269355
rect 16915 269325 16920 269355
rect 16720 269320 16920 269325
rect 16720 269275 16920 269280
rect 16720 269245 16725 269275
rect 16755 269245 16885 269275
rect 16915 269245 16920 269275
rect 16720 269240 16920 269245
rect 16720 269195 16920 269200
rect 16720 269165 16725 269195
rect 16755 269165 16885 269195
rect 16915 269165 16920 269195
rect 16720 269160 16920 269165
rect 16720 269115 16920 269120
rect 16720 269085 16725 269115
rect 16755 269085 16885 269115
rect 16915 269085 16920 269115
rect 16720 269080 16920 269085
rect 16720 269035 16920 269040
rect 16720 269005 16725 269035
rect 16755 269005 16885 269035
rect 16915 269005 16920 269035
rect 16720 269000 16920 269005
rect 16720 268955 16920 268960
rect 16720 268925 16725 268955
rect 16755 268925 16885 268955
rect 16915 268925 16920 268955
rect 16720 268920 16920 268925
rect 16720 268875 16920 268880
rect 16720 268845 16725 268875
rect 16755 268845 16885 268875
rect 16915 268845 16920 268875
rect 16720 268840 16920 268845
rect 16720 268795 16920 268800
rect 16720 268765 16725 268795
rect 16755 268765 16885 268795
rect 16915 268765 16920 268795
rect 16720 268760 16920 268765
rect 16720 268715 16920 268720
rect 16720 268685 16725 268715
rect 16755 268685 16885 268715
rect 16915 268685 16920 268715
rect 16720 268680 16920 268685
rect 16720 268635 16920 268640
rect 16720 268605 16725 268635
rect 16755 268605 16885 268635
rect 16915 268605 16920 268635
rect 16720 268600 16920 268605
rect 16720 268555 16920 268560
rect 16720 268525 16725 268555
rect 16755 268525 16885 268555
rect 16915 268525 16920 268555
rect 16720 268520 16920 268525
rect 16720 268475 16920 268480
rect 16720 268445 16725 268475
rect 16755 268445 16885 268475
rect 16915 268445 16920 268475
rect 16720 268440 16920 268445
rect 16720 268395 16920 268400
rect 16720 268365 16725 268395
rect 16755 268365 16885 268395
rect 16915 268365 16920 268395
rect 16720 268360 16920 268365
rect 16720 268315 16920 268320
rect 16720 268285 16725 268315
rect 16755 268285 16885 268315
rect 16915 268285 16920 268315
rect 16720 268280 16920 268285
rect 16720 268235 16920 268240
rect 16720 268205 16725 268235
rect 16755 268205 16885 268235
rect 16915 268205 16920 268235
rect 16720 268200 16920 268205
rect 16720 268155 16920 268160
rect 16720 268125 16725 268155
rect 16755 268125 16885 268155
rect 16915 268125 16920 268155
rect 16720 268120 16920 268125
rect 16720 268075 16920 268080
rect 16720 268045 16725 268075
rect 16755 268045 16885 268075
rect 16915 268045 16920 268075
rect 16720 268040 16920 268045
rect 16720 267995 16920 268000
rect 16720 267965 16725 267995
rect 16755 267965 16885 267995
rect 16915 267965 16920 267995
rect 16720 267960 16920 267965
rect 16720 267915 16920 267920
rect 16720 267885 16725 267915
rect 16755 267885 16885 267915
rect 16915 267885 16920 267915
rect 16720 267880 16920 267885
rect 16720 267835 16920 267840
rect 16720 267805 16725 267835
rect 16755 267805 16885 267835
rect 16915 267805 16920 267835
rect 16720 267800 16920 267805
rect 16720 267755 16920 267760
rect 16720 267725 16725 267755
rect 16755 267725 16885 267755
rect 16915 267725 16920 267755
rect 16720 267720 16920 267725
rect 16720 267675 16920 267680
rect 16720 267645 16725 267675
rect 16755 267645 16885 267675
rect 16915 267645 16920 267675
rect 16720 267640 16920 267645
rect 16720 267595 16920 267600
rect 16720 267565 16725 267595
rect 16755 267565 16885 267595
rect 16915 267565 16920 267595
rect 16720 267560 16920 267565
rect 16720 267515 16920 267520
rect 16720 267485 16725 267515
rect 16755 267485 16885 267515
rect 16915 267485 16920 267515
rect 16720 267480 16920 267485
rect 16720 267435 16920 267440
rect 16720 267405 16725 267435
rect 16755 267405 16885 267435
rect 16915 267405 16920 267435
rect 16720 267400 16920 267405
rect 16720 267355 16920 267360
rect 16720 267325 16725 267355
rect 16755 267325 16885 267355
rect 16915 267325 16920 267355
rect 16720 267320 16920 267325
rect 16720 267275 16920 267280
rect 16720 267245 16725 267275
rect 16755 267245 16885 267275
rect 16915 267245 16920 267275
rect 16720 267240 16920 267245
rect 16720 267195 16920 267200
rect 16720 267165 16725 267195
rect 16755 267165 16885 267195
rect 16915 267165 16920 267195
rect 16720 267160 16920 267165
rect 16720 267115 16920 267120
rect 16720 267085 16725 267115
rect 16755 267085 16885 267115
rect 16915 267085 16920 267115
rect 16720 267080 16920 267085
rect 16720 267035 16920 267040
rect 16720 267005 16725 267035
rect 16755 267005 16885 267035
rect 16915 267005 16920 267035
rect 16720 267000 16920 267005
rect 16720 266955 16920 266960
rect 16720 266925 16725 266955
rect 16755 266925 16885 266955
rect 16915 266925 16920 266955
rect 16720 266920 16920 266925
rect 16720 266875 16920 266880
rect 16720 266845 16725 266875
rect 16755 266845 16885 266875
rect 16915 266845 16920 266875
rect 16720 266840 16920 266845
rect 16720 266795 16920 266800
rect 16720 266765 16725 266795
rect 16755 266765 16885 266795
rect 16915 266765 16920 266795
rect 16720 266760 16920 266765
rect 16720 266715 16920 266720
rect 16720 266685 16725 266715
rect 16755 266685 16885 266715
rect 16915 266685 16920 266715
rect 16720 266680 16920 266685
rect 16720 266635 16920 266640
rect 16720 266605 16725 266635
rect 16755 266605 16885 266635
rect 16915 266605 16920 266635
rect 16720 266600 16920 266605
rect 16720 266555 16920 266560
rect 16720 266525 16725 266555
rect 16755 266525 16885 266555
rect 16915 266525 16920 266555
rect 16720 266520 16920 266525
rect 16720 266475 16920 266480
rect 16720 266445 16725 266475
rect 16755 266445 16885 266475
rect 16915 266445 16920 266475
rect 16720 266440 16920 266445
rect 16720 266395 16920 266400
rect 16720 266365 16725 266395
rect 16755 266365 16885 266395
rect 16915 266365 16920 266395
rect 16720 266360 16920 266365
rect 16720 266315 16920 266320
rect 16720 266285 16725 266315
rect 16755 266285 16885 266315
rect 16915 266285 16920 266315
rect 16720 266280 16920 266285
rect 16720 266235 16920 266240
rect 16720 266205 16725 266235
rect 16755 266205 16885 266235
rect 16915 266205 16920 266235
rect 16720 266200 16920 266205
rect 16720 266155 16920 266160
rect 16720 266125 16725 266155
rect 16755 266125 16885 266155
rect 16915 266125 16920 266155
rect 16720 266120 16920 266125
rect 16720 266075 16920 266080
rect 16720 266045 16725 266075
rect 16755 266045 16885 266075
rect 16915 266045 16920 266075
rect 16720 266040 16920 266045
rect 16720 265995 16920 266000
rect 16720 265965 16725 265995
rect 16755 265965 16885 265995
rect 16915 265965 16920 265995
rect 16720 265960 16920 265965
rect 16720 265915 16920 265920
rect 16720 265885 16725 265915
rect 16755 265885 16885 265915
rect 16915 265885 16920 265915
rect 16720 265880 16920 265885
rect 16720 265835 16920 265840
rect 16720 265805 16725 265835
rect 16755 265805 16885 265835
rect 16915 265805 16920 265835
rect 16720 265800 16920 265805
rect 16720 265755 16920 265760
rect 16720 265725 16725 265755
rect 16755 265725 16885 265755
rect 16915 265725 16920 265755
rect 16720 265720 16920 265725
rect 16720 265675 16920 265680
rect 16720 265645 16725 265675
rect 16755 265645 16885 265675
rect 16915 265645 16920 265675
rect 16720 265640 16920 265645
rect 16720 265595 16920 265600
rect 16720 265565 16725 265595
rect 16755 265565 16885 265595
rect 16915 265565 16920 265595
rect 16720 265560 16920 265565
rect 16720 265515 16920 265520
rect 16720 265485 16725 265515
rect 16755 265485 16885 265515
rect 16915 265485 16920 265515
rect 16720 265480 16920 265485
rect 16720 265435 16920 265440
rect 16720 265405 16725 265435
rect 16755 265405 16885 265435
rect 16915 265405 16920 265435
rect 16720 265400 16920 265405
rect 16720 265355 16920 265360
rect 16720 265325 16725 265355
rect 16755 265325 16885 265355
rect 16915 265325 16920 265355
rect 16720 265320 16920 265325
rect 16720 265275 16920 265280
rect 16720 265245 16725 265275
rect 16755 265245 16885 265275
rect 16915 265245 16920 265275
rect 16720 265240 16920 265245
rect 16720 265195 16920 265200
rect 16720 265165 16725 265195
rect 16755 265165 16885 265195
rect 16915 265165 16920 265195
rect 16720 265160 16920 265165
rect 16720 265115 16920 265120
rect 16720 265085 16725 265115
rect 16755 265085 16885 265115
rect 16915 265085 16920 265115
rect 16720 265080 16920 265085
rect 16720 265035 16920 265040
rect 16720 265005 16725 265035
rect 16755 265005 16885 265035
rect 16915 265005 16920 265035
rect 16720 265000 16920 265005
rect 16720 264955 16920 264960
rect 16720 264925 16725 264955
rect 16755 264925 16885 264955
rect 16915 264925 16920 264955
rect 16720 264920 16920 264925
rect 16720 264875 16920 264880
rect 16720 264845 16725 264875
rect 16755 264845 16885 264875
rect 16915 264845 16920 264875
rect 16720 264840 16920 264845
rect 16720 264795 16920 264800
rect 16720 264765 16725 264795
rect 16755 264765 16885 264795
rect 16915 264765 16920 264795
rect 16720 264760 16920 264765
rect 16720 264715 16920 264720
rect 16720 264685 16725 264715
rect 16755 264685 16885 264715
rect 16915 264685 16920 264715
rect 16720 264680 16920 264685
rect 16720 264635 16920 264640
rect 16720 264605 16725 264635
rect 16755 264605 16885 264635
rect 16915 264605 16920 264635
rect 16720 264600 16920 264605
rect 16720 264555 16920 264560
rect 16720 264525 16725 264555
rect 16755 264525 16885 264555
rect 16915 264525 16920 264555
rect 16720 264520 16920 264525
rect 16720 264475 16920 264480
rect 16720 264445 16725 264475
rect 16755 264445 16885 264475
rect 16915 264445 16920 264475
rect 16720 264440 16920 264445
rect 16720 264395 16920 264400
rect 16720 264365 16725 264395
rect 16755 264365 16885 264395
rect 16915 264365 16920 264395
rect 16720 264360 16920 264365
rect 16720 264315 16920 264320
rect 16720 264285 16725 264315
rect 16755 264285 16885 264315
rect 16915 264285 16920 264315
rect 16720 264280 16920 264285
rect 16720 264235 16920 264240
rect 16720 264205 16725 264235
rect 16755 264205 16885 264235
rect 16915 264205 16920 264235
rect 16720 264200 16920 264205
rect 16720 264155 16920 264160
rect 16720 264125 16725 264155
rect 16755 264125 16885 264155
rect 16915 264125 16920 264155
rect 16720 264120 16920 264125
rect 16720 264075 16920 264080
rect 16720 264045 16725 264075
rect 16755 264045 16885 264075
rect 16915 264045 16920 264075
rect 16720 264040 16920 264045
rect 16720 263995 16920 264000
rect 16720 263965 16725 263995
rect 16755 263965 16885 263995
rect 16915 263965 16920 263995
rect 16720 263960 16920 263965
rect 16720 263915 16920 263920
rect 16720 263885 16725 263915
rect 16755 263885 16885 263915
rect 16915 263885 16920 263915
rect 16720 263880 16920 263885
rect 16720 263835 16920 263840
rect 16720 263805 16725 263835
rect 16755 263805 16885 263835
rect 16915 263805 16920 263835
rect 16720 263800 16920 263805
rect 16720 263755 16920 263760
rect 16720 263725 16725 263755
rect 16755 263725 16885 263755
rect 16915 263725 16920 263755
rect 16720 263720 16920 263725
rect 16720 263675 16920 263680
rect 16720 263645 16725 263675
rect 16755 263645 16885 263675
rect 16915 263645 16920 263675
rect 16720 263640 16920 263645
rect 16720 263595 16920 263600
rect 16720 263565 16725 263595
rect 16755 263565 16885 263595
rect 16915 263565 16920 263595
rect 16720 263560 16920 263565
rect 16720 263515 16920 263520
rect 16720 263485 16725 263515
rect 16755 263485 16885 263515
rect 16915 263485 16920 263515
rect 16720 263480 16920 263485
rect 16720 263435 16920 263440
rect 16720 263405 16725 263435
rect 16755 263405 16885 263435
rect 16915 263405 16920 263435
rect 16720 263400 16920 263405
rect 16720 263355 16920 263360
rect 16720 263325 16725 263355
rect 16755 263325 16885 263355
rect 16915 263325 16920 263355
rect 16720 263320 16920 263325
rect 16720 263275 16920 263280
rect 16720 263245 16725 263275
rect 16755 263245 16885 263275
rect 16915 263245 16920 263275
rect 16720 263240 16920 263245
rect 16720 263195 16920 263200
rect 16720 263165 16725 263195
rect 16755 263165 16885 263195
rect 16915 263165 16920 263195
rect 16720 263160 16920 263165
rect 16720 263115 16920 263120
rect 16720 263085 16725 263115
rect 16755 263085 16885 263115
rect 16915 263085 16920 263115
rect 16720 263080 16920 263085
rect 16720 263035 16920 263040
rect 16720 263005 16725 263035
rect 16755 263005 16885 263035
rect 16915 263005 16920 263035
rect 16720 263000 16920 263005
rect 16720 262955 16920 262960
rect 16720 262925 16725 262955
rect 16755 262925 16885 262955
rect 16915 262925 16920 262955
rect 16720 262920 16920 262925
rect 16720 262875 16920 262880
rect 16720 262845 16725 262875
rect 16755 262845 16885 262875
rect 16915 262845 16920 262875
rect 16720 262840 16920 262845
rect 16720 262795 16920 262800
rect 16720 262765 16725 262795
rect 16755 262765 16885 262795
rect 16915 262765 16920 262795
rect 16720 262760 16920 262765
rect 16720 262715 16920 262720
rect 16720 262685 16725 262715
rect 16755 262685 16885 262715
rect 16915 262685 16920 262715
rect 16720 262680 16920 262685
rect 16720 262635 16920 262640
rect 16720 262605 16725 262635
rect 16755 262605 16885 262635
rect 16915 262605 16920 262635
rect 16720 262600 16920 262605
rect 16720 262555 16920 262560
rect 16720 262525 16725 262555
rect 16755 262525 16885 262555
rect 16915 262525 16920 262555
rect 16720 262520 16920 262525
rect 16720 262475 16920 262480
rect 16720 262445 16725 262475
rect 16755 262445 16885 262475
rect 16915 262445 16920 262475
rect 16720 262440 16920 262445
rect 16720 262395 16920 262400
rect 16720 262365 16725 262395
rect 16755 262365 16885 262395
rect 16915 262365 16920 262395
rect 16720 262360 16920 262365
rect 16720 262315 16920 262320
rect 16720 262285 16725 262315
rect 16755 262285 16885 262315
rect 16915 262285 16920 262315
rect 16720 262280 16920 262285
rect 16720 262235 16920 262240
rect 16720 262205 16725 262235
rect 16755 262205 16885 262235
rect 16915 262205 16920 262235
rect 16720 262200 16920 262205
rect 16720 262155 16920 262160
rect 16720 262125 16725 262155
rect 16755 262125 16885 262155
rect 16915 262125 16920 262155
rect 16720 262120 16920 262125
rect 16720 262075 16920 262080
rect 16720 262045 16725 262075
rect 16755 262045 16885 262075
rect 16915 262045 16920 262075
rect 16720 262040 16920 262045
rect 16720 261995 16920 262000
rect 16720 261965 16725 261995
rect 16755 261965 16885 261995
rect 16915 261965 16920 261995
rect 16720 261960 16920 261965
rect 16720 261915 16920 261920
rect 16720 261885 16725 261915
rect 16755 261885 16885 261915
rect 16915 261885 16920 261915
rect 16720 261880 16920 261885
rect 16720 261835 16920 261840
rect 16720 261805 16725 261835
rect 16755 261805 16885 261835
rect 16915 261805 16920 261835
rect 16720 261800 16920 261805
rect 16720 261755 16920 261760
rect 16720 261725 16725 261755
rect 16755 261725 16885 261755
rect 16915 261725 16920 261755
rect 16720 261720 16920 261725
rect 16720 261675 16920 261680
rect 16720 261645 16725 261675
rect 16755 261645 16885 261675
rect 16915 261645 16920 261675
rect 16720 261640 16920 261645
rect 16720 261595 16920 261600
rect 16720 261565 16725 261595
rect 16755 261565 16885 261595
rect 16915 261565 16920 261595
rect 16720 261560 16920 261565
rect 16720 261515 16920 261520
rect 16720 261485 16725 261515
rect 16755 261485 16885 261515
rect 16915 261485 16920 261515
rect 16720 261480 16920 261485
rect 16720 261435 16920 261440
rect 16720 261405 16725 261435
rect 16755 261405 16885 261435
rect 16915 261405 16920 261435
rect 16720 261400 16920 261405
rect 16720 261355 16920 261360
rect 16720 261325 16725 261355
rect 16755 261325 16885 261355
rect 16915 261325 16920 261355
rect 16720 261320 16920 261325
rect 16720 261275 16920 261280
rect 16720 261245 16725 261275
rect 16755 261245 16885 261275
rect 16915 261245 16920 261275
rect 16720 261240 16920 261245
rect 16720 261195 16920 261200
rect 16720 261165 16725 261195
rect 16755 261165 16885 261195
rect 16915 261165 16920 261195
rect 16720 261160 16920 261165
rect 16720 261115 16920 261120
rect 16720 261085 16725 261115
rect 16755 261085 16885 261115
rect 16915 261085 16920 261115
rect 16720 261080 16920 261085
rect 16720 261035 16920 261040
rect 16720 261005 16725 261035
rect 16755 261005 16885 261035
rect 16915 261005 16920 261035
rect 16720 261000 16920 261005
rect 16720 260955 16920 260960
rect 16720 260925 16725 260955
rect 16755 260925 16885 260955
rect 16915 260925 16920 260955
rect 16720 260920 16920 260925
rect 16720 260875 16920 260880
rect 16720 260845 16725 260875
rect 16755 260845 16885 260875
rect 16915 260845 16920 260875
rect 16720 260840 16920 260845
rect 16720 260795 16920 260800
rect 16720 260765 16725 260795
rect 16755 260765 16885 260795
rect 16915 260765 16920 260795
rect 16720 260760 16920 260765
rect 16720 260715 16920 260720
rect 16720 260685 16725 260715
rect 16755 260685 16885 260715
rect 16915 260685 16920 260715
rect 16720 260680 16920 260685
rect 16720 260635 16920 260640
rect 16720 260605 16725 260635
rect 16755 260605 16885 260635
rect 16915 260605 16920 260635
rect 16720 260600 16920 260605
rect 16720 260555 16920 260560
rect 16720 260525 16725 260555
rect 16755 260525 16885 260555
rect 16915 260525 16920 260555
rect 16720 260520 16920 260525
rect 16720 260475 16920 260480
rect 16720 260445 16725 260475
rect 16755 260445 16885 260475
rect 16915 260445 16920 260475
rect 16720 260440 16920 260445
rect 16720 260395 16920 260400
rect 16720 260365 16725 260395
rect 16755 260365 16885 260395
rect 16915 260365 16920 260395
rect 16720 260360 16920 260365
rect 16720 260315 16920 260320
rect 16720 260285 16725 260315
rect 16755 260285 16885 260315
rect 16915 260285 16920 260315
rect 16720 260280 16920 260285
rect 16720 260235 16920 260240
rect 16720 260205 16725 260235
rect 16755 260205 16885 260235
rect 16915 260205 16920 260235
rect 16720 260200 16920 260205
rect 16720 260155 16920 260160
rect 16720 260125 16725 260155
rect 16755 260125 16885 260155
rect 16915 260125 16920 260155
rect 16720 260120 16920 260125
rect 16720 260075 16920 260080
rect 16720 260045 16725 260075
rect 16755 260045 16885 260075
rect 16915 260045 16920 260075
rect 16720 260040 16920 260045
rect 16720 259995 16920 260000
rect 16720 259965 16725 259995
rect 16755 259965 16885 259995
rect 16915 259965 16920 259995
rect 16720 259960 16920 259965
rect 16720 259915 16920 259920
rect 16720 259885 16725 259915
rect 16755 259885 16885 259915
rect 16915 259885 16920 259915
rect 16720 259880 16920 259885
rect 16720 259835 16920 259840
rect 16720 259805 16725 259835
rect 16755 259805 16885 259835
rect 16915 259805 16920 259835
rect 16720 259800 16920 259805
rect 16720 259755 16920 259760
rect 16720 259725 16725 259755
rect 16755 259725 16885 259755
rect 16915 259725 16920 259755
rect 16720 259720 16920 259725
rect 16720 259675 16920 259680
rect 16720 259645 16725 259675
rect 16755 259645 16885 259675
rect 16915 259645 16920 259675
rect 16720 259640 16920 259645
rect 16720 259595 16920 259600
rect 16720 259565 16725 259595
rect 16755 259565 16885 259595
rect 16915 259565 16920 259595
rect 16720 259560 16920 259565
rect 16720 259515 16920 259520
rect 16720 259485 16725 259515
rect 16755 259485 16885 259515
rect 16915 259485 16920 259515
rect 16720 259480 16920 259485
rect 16720 259435 16920 259440
rect 16720 259405 16725 259435
rect 16755 259405 16885 259435
rect 16915 259405 16920 259435
rect 16720 259400 16920 259405
rect 16720 259355 16920 259360
rect 16720 259325 16725 259355
rect 16755 259325 16885 259355
rect 16915 259325 16920 259355
rect 16720 259320 16920 259325
rect 16720 259275 16920 259280
rect 16720 259245 16725 259275
rect 16755 259245 16885 259275
rect 16915 259245 16920 259275
rect 16720 259240 16920 259245
rect 16720 259195 16920 259200
rect 16720 259165 16725 259195
rect 16755 259165 16885 259195
rect 16915 259165 16920 259195
rect 16720 259160 16920 259165
rect 16720 259115 16920 259120
rect 16720 259085 16725 259115
rect 16755 259085 16885 259115
rect 16915 259085 16920 259115
rect 16720 259080 16920 259085
rect 16720 259035 16920 259040
rect 16720 259005 16725 259035
rect 16755 259005 16885 259035
rect 16915 259005 16920 259035
rect 16720 259000 16920 259005
rect 16720 258955 16920 258960
rect 16720 258925 16725 258955
rect 16755 258925 16885 258955
rect 16915 258925 16920 258955
rect 16720 258920 16920 258925
rect 16720 258875 16920 258880
rect 16720 258845 16725 258875
rect 16755 258845 16885 258875
rect 16915 258845 16920 258875
rect 16720 258840 16920 258845
rect 16720 258795 16920 258800
rect 16720 258765 16725 258795
rect 16755 258765 16885 258795
rect 16915 258765 16920 258795
rect 16720 258760 16920 258765
rect 16720 258715 16920 258720
rect 16720 258685 16725 258715
rect 16755 258685 16885 258715
rect 16915 258685 16920 258715
rect 16720 258680 16920 258685
rect 16720 258635 16920 258640
rect 16720 258605 16725 258635
rect 16755 258605 16885 258635
rect 16915 258605 16920 258635
rect 16720 258600 16920 258605
rect 16720 258555 16920 258560
rect 16720 258525 16725 258555
rect 16755 258525 16885 258555
rect 16915 258525 16920 258555
rect 16720 258520 16920 258525
rect 16720 258475 16920 258480
rect 16720 258445 16725 258475
rect 16755 258445 16885 258475
rect 16915 258445 16920 258475
rect 16720 258440 16920 258445
rect 16720 258395 16920 258400
rect 16720 258365 16725 258395
rect 16755 258365 16885 258395
rect 16915 258365 16920 258395
rect 16720 258360 16920 258365
rect 16720 258315 16920 258320
rect 16720 258285 16725 258315
rect 16755 258285 16885 258315
rect 16915 258285 16920 258315
rect 16720 258280 16920 258285
rect 16720 258235 16920 258240
rect 16720 258205 16725 258235
rect 16755 258205 16885 258235
rect 16915 258205 16920 258235
rect 16720 258200 16920 258205
rect 16720 258155 16920 258160
rect 16720 258125 16725 258155
rect 16755 258125 16885 258155
rect 16915 258125 16920 258155
rect 16720 258120 16920 258125
rect 16720 258075 16920 258080
rect 16720 258045 16725 258075
rect 16755 258045 16885 258075
rect 16915 258045 16920 258075
rect 16720 258040 16920 258045
rect 16720 257995 16920 258000
rect 16720 257965 16725 257995
rect 16755 257965 16885 257995
rect 16915 257965 16920 257995
rect 16720 257960 16920 257965
rect 16720 257915 16920 257920
rect 16720 257885 16725 257915
rect 16755 257885 16885 257915
rect 16915 257885 16920 257915
rect 16720 257880 16920 257885
rect 16720 257835 16920 257840
rect 16720 257805 16725 257835
rect 16755 257805 16885 257835
rect 16915 257805 16920 257835
rect 16720 257800 16920 257805
rect 16720 257755 16920 257760
rect 16720 257725 16725 257755
rect 16755 257725 16885 257755
rect 16915 257725 16920 257755
rect 16720 257720 16920 257725
rect 16720 257675 16920 257680
rect 16720 257645 16725 257675
rect 16755 257645 16885 257675
rect 16915 257645 16920 257675
rect 16720 257640 16920 257645
rect 16720 257595 16920 257600
rect 16720 257565 16725 257595
rect 16755 257565 16885 257595
rect 16915 257565 16920 257595
rect 16720 257560 16920 257565
rect 16720 257515 16920 257520
rect 16720 257485 16725 257515
rect 16755 257485 16885 257515
rect 16915 257485 16920 257515
rect 16720 257480 16920 257485
rect 16720 257435 16920 257440
rect 16720 257405 16725 257435
rect 16755 257405 16885 257435
rect 16915 257405 16920 257435
rect 16720 257400 16920 257405
rect 16720 257355 16920 257360
rect 16720 257325 16725 257355
rect 16755 257325 16885 257355
rect 16915 257325 16920 257355
rect 16720 257320 16920 257325
rect 16720 257275 16920 257280
rect 16720 257245 16725 257275
rect 16755 257245 16885 257275
rect 16915 257245 16920 257275
rect 16720 257240 16920 257245
rect 16720 257195 16920 257200
rect 16720 257165 16725 257195
rect 16755 257165 16885 257195
rect 16915 257165 16920 257195
rect 16720 257160 16920 257165
rect 16720 257115 16920 257120
rect 16720 257085 16725 257115
rect 16755 257085 16885 257115
rect 16915 257085 16920 257115
rect 16720 257080 16920 257085
rect 16720 257035 16920 257040
rect 16720 257005 16725 257035
rect 16755 257005 16885 257035
rect 16915 257005 16920 257035
rect 16720 257000 16920 257005
rect 16720 256955 16920 256960
rect 16720 256925 16725 256955
rect 16755 256925 16885 256955
rect 16915 256925 16920 256955
rect 16720 256920 16920 256925
rect 16720 256875 16920 256880
rect 16720 256845 16725 256875
rect 16755 256845 16885 256875
rect 16915 256845 16920 256875
rect 16720 256840 16920 256845
rect 16720 256795 16920 256800
rect 16720 256765 16725 256795
rect 16755 256765 16885 256795
rect 16915 256765 16920 256795
rect 16720 256760 16920 256765
rect 16720 256715 16920 256720
rect 16720 256685 16725 256715
rect 16755 256685 16885 256715
rect 16915 256685 16920 256715
rect 16720 256680 16920 256685
rect 16720 256635 16920 256640
rect 16720 256605 16725 256635
rect 16755 256605 16885 256635
rect 16915 256605 16920 256635
rect 16720 256600 16920 256605
rect 16720 256555 16920 256560
rect 16720 256525 16725 256555
rect 16755 256525 16885 256555
rect 16915 256525 16920 256555
rect 16720 256520 16920 256525
rect 16720 256475 16920 256480
rect 16720 256445 16725 256475
rect 16755 256445 16885 256475
rect 16915 256445 16920 256475
rect 16720 256440 16920 256445
rect 16720 256395 16920 256400
rect 16720 256365 16725 256395
rect 16755 256365 16885 256395
rect 16915 256365 16920 256395
rect 16720 256360 16920 256365
rect 16720 256315 16920 256320
rect 16720 256285 16725 256315
rect 16755 256285 16885 256315
rect 16915 256285 16920 256315
rect 16720 256280 16920 256285
rect 16720 256235 16920 256240
rect 16720 256205 16725 256235
rect 16755 256205 16885 256235
rect 16915 256205 16920 256235
rect 16720 256200 16920 256205
rect 16720 256155 16920 256160
rect 16720 256125 16725 256155
rect 16755 256125 16885 256155
rect 16915 256125 16920 256155
rect 16720 256120 16920 256125
rect 16720 256075 16920 256080
rect 16720 256045 16725 256075
rect 16755 256045 16885 256075
rect 16915 256045 16920 256075
rect 16720 256040 16920 256045
rect 16720 255995 16920 256000
rect 16720 255965 16725 255995
rect 16755 255965 16885 255995
rect 16915 255965 16920 255995
rect 16720 255960 16920 255965
rect 400 255875 16920 255880
rect 400 255845 405 255875
rect 435 255845 485 255875
rect 515 255845 565 255875
rect 595 255845 645 255875
rect 675 255845 725 255875
rect 755 255845 805 255875
rect 835 255845 885 255875
rect 915 255845 965 255875
rect 995 255845 1045 255875
rect 1075 255845 1125 255875
rect 1155 255845 1205 255875
rect 1235 255845 1285 255875
rect 1315 255845 1365 255875
rect 1395 255845 1445 255875
rect 1475 255845 1525 255875
rect 1555 255845 1605 255875
rect 1635 255845 1685 255875
rect 1715 255845 1765 255875
rect 1795 255845 1845 255875
rect 1875 255845 1925 255875
rect 1955 255845 2005 255875
rect 2035 255845 2085 255875
rect 2115 255845 2165 255875
rect 2195 255845 2245 255875
rect 2275 255845 2325 255875
rect 2355 255845 2405 255875
rect 2435 255845 2485 255875
rect 2515 255845 2565 255875
rect 2595 255845 2645 255875
rect 2675 255845 2725 255875
rect 2755 255845 3045 255875
rect 3075 255845 3125 255875
rect 3155 255845 3205 255875
rect 3235 255845 3285 255875
rect 3315 255845 3365 255875
rect 3395 255845 3445 255875
rect 3475 255845 3525 255875
rect 3555 255845 3605 255875
rect 3635 255845 3685 255875
rect 3715 255845 3765 255875
rect 3795 255845 3845 255875
rect 3875 255845 3925 255875
rect 3955 255845 4005 255875
rect 4035 255845 4085 255875
rect 4115 255845 4165 255875
rect 4195 255845 4245 255875
rect 4275 255845 4325 255875
rect 4355 255845 4405 255875
rect 4435 255845 4485 255875
rect 4515 255845 4565 255875
rect 4595 255845 4645 255875
rect 4675 255845 4725 255875
rect 4755 255845 4805 255875
rect 4835 255845 4885 255875
rect 4915 255845 4965 255875
rect 4995 255845 5045 255875
rect 5075 255845 5125 255875
rect 5155 255845 5205 255875
rect 5235 255845 5285 255875
rect 5315 255845 5365 255875
rect 5395 255845 5445 255875
rect 5475 255845 5525 255875
rect 5555 255845 5605 255875
rect 5635 255845 5685 255875
rect 5715 255845 5765 255875
rect 5795 255845 5845 255875
rect 5875 255845 5925 255875
rect 5955 255845 6005 255875
rect 6035 255845 6085 255875
rect 6115 255845 6165 255875
rect 6195 255845 6245 255875
rect 6275 255845 6325 255875
rect 6355 255845 6405 255875
rect 6435 255845 6485 255875
rect 6515 255845 6565 255875
rect 6595 255845 6645 255875
rect 6675 255845 6725 255875
rect 6755 255845 6805 255875
rect 6835 255845 6885 255875
rect 6915 255845 6965 255875
rect 6995 255845 7045 255875
rect 7075 255845 7125 255875
rect 7155 255845 7205 255875
rect 7235 255845 7285 255875
rect 7315 255845 7365 255875
rect 7395 255845 7445 255875
rect 7475 255845 7525 255875
rect 7555 255845 7605 255875
rect 7635 255845 7685 255875
rect 7715 255845 7765 255875
rect 7795 255845 7845 255875
rect 7875 255845 7925 255875
rect 7955 255845 8005 255875
rect 8035 255845 8085 255875
rect 8115 255845 8165 255875
rect 8195 255845 8245 255875
rect 8275 255845 8325 255875
rect 8355 255845 8405 255875
rect 8435 255845 8485 255875
rect 8515 255845 8565 255875
rect 8595 255845 8645 255875
rect 8675 255845 8725 255875
rect 8755 255845 8805 255875
rect 8835 255845 8885 255875
rect 8915 255845 8965 255875
rect 8995 255845 9045 255875
rect 9075 255845 9125 255875
rect 9155 255845 9205 255875
rect 9235 255845 9285 255875
rect 9315 255845 9365 255875
rect 9395 255845 9445 255875
rect 9475 255845 9525 255875
rect 9555 255845 9605 255875
rect 9635 255845 9685 255875
rect 9715 255845 9765 255875
rect 9795 255845 9845 255875
rect 9875 255845 9925 255875
rect 9955 255845 10005 255875
rect 10035 255845 10085 255875
rect 10115 255845 10165 255875
rect 10195 255845 10245 255875
rect 10275 255845 10325 255875
rect 10355 255845 10405 255875
rect 10435 255845 10485 255875
rect 10515 255845 10565 255875
rect 10595 255845 10645 255875
rect 10675 255845 10725 255875
rect 10755 255845 10805 255875
rect 10835 255845 10885 255875
rect 10915 255845 10965 255875
rect 10995 255845 11045 255875
rect 11075 255845 11125 255875
rect 11155 255845 11205 255875
rect 11235 255845 11285 255875
rect 11315 255845 11365 255875
rect 11395 255845 11445 255875
rect 11475 255845 11525 255875
rect 11555 255845 11605 255875
rect 11635 255845 11685 255875
rect 11715 255845 11765 255875
rect 11795 255845 11845 255875
rect 11875 255845 11925 255875
rect 11955 255845 12005 255875
rect 12035 255845 12085 255875
rect 12115 255845 12165 255875
rect 12195 255845 12245 255875
rect 12275 255845 12325 255875
rect 12355 255845 12405 255875
rect 12435 255845 12485 255875
rect 12515 255845 12565 255875
rect 12595 255845 12645 255875
rect 12675 255845 12725 255875
rect 12755 255845 12805 255875
rect 12835 255845 12885 255875
rect 12915 255845 12965 255875
rect 12995 255845 13045 255875
rect 13075 255845 13125 255875
rect 13155 255845 13205 255875
rect 13235 255845 13285 255875
rect 13315 255845 13365 255875
rect 13395 255845 13445 255875
rect 13475 255845 13525 255875
rect 13555 255845 13605 255875
rect 13635 255845 13685 255875
rect 13715 255845 13765 255875
rect 13795 255845 13845 255875
rect 13875 255845 13925 255875
rect 13955 255845 14005 255875
rect 14035 255845 14085 255875
rect 14115 255845 14165 255875
rect 14195 255845 14245 255875
rect 14275 255845 14325 255875
rect 14355 255845 14405 255875
rect 14435 255845 14485 255875
rect 14515 255845 14565 255875
rect 14595 255845 14645 255875
rect 14675 255845 14725 255875
rect 14755 255845 14805 255875
rect 14835 255845 14885 255875
rect 14915 255845 14965 255875
rect 14995 255845 15045 255875
rect 15075 255845 15125 255875
rect 15155 255845 15205 255875
rect 15235 255845 15285 255875
rect 15315 255845 15365 255875
rect 15395 255845 15445 255875
rect 15475 255845 15525 255875
rect 15555 255845 15605 255875
rect 15635 255845 15685 255875
rect 15715 255845 15765 255875
rect 15795 255845 15845 255875
rect 15875 255845 15925 255875
rect 15955 255845 16005 255875
rect 16035 255845 16085 255875
rect 16115 255845 16165 255875
rect 16195 255845 16245 255875
rect 16275 255845 16325 255875
rect 16355 255845 16405 255875
rect 16435 255845 16485 255875
rect 16515 255845 16565 255875
rect 16595 255845 16645 255875
rect 16675 255845 16725 255875
rect 16755 255845 16885 255875
rect 16915 255845 16920 255875
rect 400 255840 16920 255845
rect 320 255795 16840 255800
rect 320 255765 325 255795
rect 355 255765 16805 255795
rect 16835 255765 16840 255795
rect 320 255760 16840 255765
rect 400 255715 16920 255720
rect 400 255685 405 255715
rect 435 255685 485 255715
rect 515 255685 565 255715
rect 595 255685 645 255715
rect 675 255685 725 255715
rect 755 255685 805 255715
rect 835 255685 885 255715
rect 915 255685 965 255715
rect 995 255685 1045 255715
rect 1075 255685 1125 255715
rect 1155 255685 1205 255715
rect 1235 255685 1285 255715
rect 1315 255685 1365 255715
rect 1395 255685 1445 255715
rect 1475 255685 1525 255715
rect 1555 255685 1605 255715
rect 1635 255685 1685 255715
rect 1715 255685 1765 255715
rect 1795 255685 1845 255715
rect 1875 255685 1925 255715
rect 1955 255685 2005 255715
rect 2035 255685 2085 255715
rect 2115 255685 2165 255715
rect 2195 255685 2245 255715
rect 2275 255685 2325 255715
rect 2355 255685 2405 255715
rect 2435 255685 2485 255715
rect 2515 255685 2565 255715
rect 2595 255685 2645 255715
rect 2675 255685 2725 255715
rect 2755 255685 3045 255715
rect 3075 255685 3125 255715
rect 3155 255685 3205 255715
rect 3235 255685 3285 255715
rect 3315 255685 3365 255715
rect 3395 255685 3445 255715
rect 3475 255685 3525 255715
rect 3555 255685 3605 255715
rect 3635 255685 3685 255715
rect 3715 255685 3765 255715
rect 3795 255685 3845 255715
rect 3875 255685 3925 255715
rect 3955 255685 4005 255715
rect 4035 255685 4085 255715
rect 4115 255685 4165 255715
rect 4195 255685 4245 255715
rect 4275 255685 4325 255715
rect 4355 255685 4405 255715
rect 4435 255685 4485 255715
rect 4515 255685 4565 255715
rect 4595 255685 4645 255715
rect 4675 255685 4725 255715
rect 4755 255685 4805 255715
rect 4835 255685 4885 255715
rect 4915 255685 4965 255715
rect 4995 255685 5045 255715
rect 5075 255685 5125 255715
rect 5155 255685 5205 255715
rect 5235 255685 5285 255715
rect 5315 255685 5365 255715
rect 5395 255685 5445 255715
rect 5475 255685 5525 255715
rect 5555 255685 5605 255715
rect 5635 255685 5685 255715
rect 5715 255685 5765 255715
rect 5795 255685 5845 255715
rect 5875 255685 5925 255715
rect 5955 255685 6005 255715
rect 6035 255685 6085 255715
rect 6115 255685 6165 255715
rect 6195 255685 6245 255715
rect 6275 255685 6325 255715
rect 6355 255685 6405 255715
rect 6435 255685 6485 255715
rect 6515 255685 6565 255715
rect 6595 255685 6645 255715
rect 6675 255685 6725 255715
rect 6755 255685 6805 255715
rect 6835 255685 6885 255715
rect 6915 255685 6965 255715
rect 6995 255685 7045 255715
rect 7075 255685 7125 255715
rect 7155 255685 7205 255715
rect 7235 255685 7285 255715
rect 7315 255685 7365 255715
rect 7395 255685 7445 255715
rect 7475 255685 7525 255715
rect 7555 255685 7605 255715
rect 7635 255685 7685 255715
rect 7715 255685 7765 255715
rect 7795 255685 7845 255715
rect 7875 255685 7925 255715
rect 7955 255685 8005 255715
rect 8035 255685 8085 255715
rect 8115 255685 8165 255715
rect 8195 255685 8245 255715
rect 8275 255685 8325 255715
rect 8355 255685 8405 255715
rect 8435 255685 8485 255715
rect 8515 255685 8565 255715
rect 8595 255685 8645 255715
rect 8675 255685 8725 255715
rect 8755 255685 8805 255715
rect 8835 255685 8885 255715
rect 8915 255685 8965 255715
rect 8995 255685 9045 255715
rect 9075 255685 9125 255715
rect 9155 255685 9205 255715
rect 9235 255685 9285 255715
rect 9315 255685 9365 255715
rect 9395 255685 9445 255715
rect 9475 255685 9525 255715
rect 9555 255685 9605 255715
rect 9635 255685 9685 255715
rect 9715 255685 9765 255715
rect 9795 255685 9845 255715
rect 9875 255685 9925 255715
rect 9955 255685 10005 255715
rect 10035 255685 10085 255715
rect 10115 255685 10165 255715
rect 10195 255685 10245 255715
rect 10275 255685 10325 255715
rect 10355 255685 10405 255715
rect 10435 255685 10485 255715
rect 10515 255685 10565 255715
rect 10595 255685 10645 255715
rect 10675 255685 10725 255715
rect 10755 255685 10805 255715
rect 10835 255685 10885 255715
rect 10915 255685 10965 255715
rect 10995 255685 11045 255715
rect 11075 255685 11125 255715
rect 11155 255685 11205 255715
rect 11235 255685 11285 255715
rect 11315 255685 11365 255715
rect 11395 255685 11445 255715
rect 11475 255685 11525 255715
rect 11555 255685 11605 255715
rect 11635 255685 11685 255715
rect 11715 255685 11765 255715
rect 11795 255685 11845 255715
rect 11875 255685 11925 255715
rect 11955 255685 12005 255715
rect 12035 255685 12085 255715
rect 12115 255685 12165 255715
rect 12195 255685 12245 255715
rect 12275 255685 12325 255715
rect 12355 255685 12405 255715
rect 12435 255685 12485 255715
rect 12515 255685 12565 255715
rect 12595 255685 12645 255715
rect 12675 255685 12725 255715
rect 12755 255685 12805 255715
rect 12835 255685 12885 255715
rect 12915 255685 12965 255715
rect 12995 255685 13045 255715
rect 13075 255685 13125 255715
rect 13155 255685 13205 255715
rect 13235 255685 13285 255715
rect 13315 255685 13365 255715
rect 13395 255685 13445 255715
rect 13475 255685 13525 255715
rect 13555 255685 13605 255715
rect 13635 255685 13685 255715
rect 13715 255685 13765 255715
rect 13795 255685 13845 255715
rect 13875 255685 13925 255715
rect 13955 255685 14005 255715
rect 14035 255685 14085 255715
rect 14115 255685 14165 255715
rect 14195 255685 14245 255715
rect 14275 255685 14325 255715
rect 14355 255685 14405 255715
rect 14435 255685 14485 255715
rect 14515 255685 14565 255715
rect 14595 255685 14645 255715
rect 14675 255685 14725 255715
rect 14755 255685 14805 255715
rect 14835 255685 14885 255715
rect 14915 255685 14965 255715
rect 14995 255685 15045 255715
rect 15075 255685 15125 255715
rect 15155 255685 15205 255715
rect 15235 255685 15285 255715
rect 15315 255685 15365 255715
rect 15395 255685 15445 255715
rect 15475 255685 15525 255715
rect 15555 255685 15605 255715
rect 15635 255685 15685 255715
rect 15715 255685 15765 255715
rect 15795 255685 15845 255715
rect 15875 255685 15925 255715
rect 15955 255685 16005 255715
rect 16035 255685 16085 255715
rect 16115 255685 16165 255715
rect 16195 255685 16245 255715
rect 16275 255685 16325 255715
rect 16355 255685 16405 255715
rect 16435 255685 16485 255715
rect 16515 255685 16565 255715
rect 16595 255685 16645 255715
rect 16675 255685 16725 255715
rect 16755 255685 16885 255715
rect 16915 255685 16920 255715
rect 400 255680 16920 255685
rect 262 -400 318 240
rect 853 -400 909 240
rect 1444 -400 1500 240
rect 2035 -400 2091 240
rect 2626 -400 2682 240
rect 3217 -400 3273 240
rect 3808 -400 3864 240
rect 4399 -400 4455 240
rect 4990 -400 5046 240
rect 5581 -400 5637 240
rect 6172 -400 6228 240
rect 6763 -400 6819 240
rect 7354 -400 7410 240
rect 7945 -400 8001 240
rect 8536 -400 8592 240
rect 9127 -400 9183 240
rect 9718 -400 9774 240
rect 10309 -400 10365 240
rect 10900 -400 10956 240
rect 11491 -400 11547 240
rect 12082 -400 12138 240
rect 12673 -400 12729 240
rect 13264 -400 13320 240
rect 13855 -400 13911 240
rect 14446 -400 14502 240
rect 15037 -400 15093 240
rect 15628 -400 15684 240
rect 16219 -400 16275 240
rect 16810 -400 16866 240
rect 17401 -400 17457 240
rect 17992 -400 18048 240
rect 18583 -400 18639 240
rect 19174 -400 19230 240
rect 19765 -400 19821 240
rect 20356 -400 20412 240
rect 20947 -400 21003 240
rect 21538 -400 21594 240
rect 22129 -400 22185 240
rect 22720 -400 22776 240
rect 23311 -400 23367 240
rect 23902 -400 23958 240
rect 24493 -400 24549 240
rect 25084 -400 25140 240
rect 25675 -400 25731 240
rect 26266 -400 26322 240
rect 26857 -400 26913 240
rect 27448 -400 27504 240
rect 28039 -400 28095 240
rect 28630 -400 28686 240
rect 29221 -400 29277 240
rect 29812 -400 29868 240
rect 30403 -400 30459 240
rect 30994 -400 31050 240
rect 31585 -400 31641 240
rect 32176 -400 32232 240
rect 32767 -400 32823 240
rect 33358 -400 33414 240
rect 33949 -400 34005 240
rect 34540 -400 34596 240
rect 35131 -400 35187 240
rect 35722 -400 35778 240
rect 36313 -400 36369 240
rect 36904 -400 36960 240
rect 37495 -400 37551 240
rect 38086 -400 38142 240
rect 38677 -400 38733 240
rect 39268 -400 39324 240
rect 39859 -400 39915 240
rect 40450 -400 40506 240
rect 41041 -400 41097 240
rect 41632 -400 41688 240
rect 42223 -400 42279 240
rect 42814 -400 42870 240
rect 43405 -400 43461 240
rect 43996 -400 44052 240
rect 44587 -400 44643 240
rect 45178 -400 45234 240
rect 45769 -400 45825 240
rect 46360 -400 46416 240
rect 46951 -400 47007 240
rect 47542 -400 47598 240
rect 48133 -400 48189 240
rect 48724 -400 48780 240
rect 49315 -400 49371 240
rect 49906 -400 49962 240
rect 50497 -400 50553 240
rect 51088 -400 51144 240
rect 51679 -400 51735 240
rect 52270 -400 52326 240
rect 52861 -400 52917 240
rect 53452 -400 53508 240
rect 54043 -400 54099 240
rect 54634 -400 54690 240
rect 55225 -400 55281 240
rect 55816 -400 55872 240
rect 56407 -400 56463 240
rect 56998 -400 57054 240
rect 57589 -400 57645 240
rect 58180 -400 58236 240
rect 58771 -400 58827 240
rect 59362 -400 59418 240
rect 59953 -400 60009 240
rect 60544 -400 60600 240
rect 61135 -400 61191 240
rect 61726 -400 61782 240
rect 62317 -400 62373 240
rect 62908 -400 62964 240
rect 63499 -400 63555 240
rect 64090 -400 64146 240
rect 64681 -400 64737 240
rect 65272 -400 65328 240
rect 65863 -400 65919 240
rect 66454 -400 66510 240
rect 67045 -400 67101 240
rect 67636 -400 67692 240
rect 68227 -400 68283 240
rect 68818 -400 68874 240
rect 69409 -400 69465 240
rect 70000 -400 70056 240
rect 70591 -400 70647 240
rect 71182 -400 71238 240
rect 71773 -400 71829 240
rect 72364 -400 72420 240
rect 72955 -400 73011 240
rect 73546 -400 73602 240
rect 74137 -400 74193 240
rect 74728 -400 74784 240
rect 75319 -400 75375 240
rect 75910 -400 75966 240
rect 76501 -400 76557 240
rect 77092 -400 77148 240
rect 77683 -400 77739 240
rect 78274 -400 78330 240
rect 78865 -400 78921 240
rect 79456 -400 79512 240
rect 80047 -400 80103 240
rect 80638 -400 80694 240
rect 81229 -400 81285 240
rect 81820 -400 81876 240
rect 82411 -400 82467 240
rect 83002 -400 83058 240
rect 83593 -400 83649 240
rect 84184 -400 84240 240
rect 84775 -400 84831 240
rect 85366 -400 85422 240
rect 85957 -400 86013 240
rect 86548 -400 86604 240
rect 87139 -400 87195 240
rect 87730 -400 87786 240
rect 88321 -400 88377 240
rect 88912 -400 88968 240
rect 89503 -400 89559 240
rect 90094 -400 90150 240
rect 90685 -400 90741 240
rect 91276 -400 91332 240
rect 91867 -400 91923 240
rect 92458 -400 92514 240
rect 93049 -400 93105 240
rect 93640 -400 93696 240
rect 94231 -400 94287 240
rect 94822 -400 94878 240
rect 95413 -400 95469 240
rect 96004 -400 96060 240
rect 96595 -400 96651 240
rect 97186 -400 97242 240
rect 97777 -400 97833 240
rect 98368 -400 98424 240
rect 98959 -400 99015 240
rect 99550 -400 99606 240
rect 100141 -400 100197 240
rect 100732 -400 100788 240
rect 101323 -400 101379 240
rect 101914 -400 101970 240
rect 102505 -400 102561 240
rect 103096 -400 103152 240
rect 103687 -400 103743 240
rect 104278 -400 104334 240
rect 104869 -400 104925 240
rect 105460 -400 105516 240
rect 106051 -400 106107 240
rect 106642 -400 106698 240
rect 107233 -400 107289 240
rect 107824 -400 107880 240
rect 108415 -400 108471 240
rect 109006 -400 109062 240
rect 109597 -400 109653 240
rect 110188 -400 110244 240
rect 110779 -400 110835 240
rect 111370 -400 111426 240
rect 111961 -400 112017 240
rect 112552 -400 112608 240
rect 113143 -400 113199 240
rect 113734 -400 113790 240
rect 114325 -400 114381 240
rect 114916 -400 114972 240
rect 115507 -400 115563 240
rect 116098 -400 116154 240
rect 116689 -400 116745 240
rect 117280 -400 117336 240
rect 117871 -400 117927 240
rect 118462 -400 118518 240
rect 119053 -400 119109 240
rect 119644 -400 119700 240
rect 120235 -400 120291 240
rect 120826 -400 120882 240
rect 121417 -400 121473 240
rect 122008 -400 122064 240
rect 122599 -400 122655 240
rect 123190 -400 123246 240
rect 123781 -400 123837 240
rect 124372 -400 124428 240
rect 124963 -400 125019 240
rect 125554 -400 125610 240
rect 126145 -400 126201 240
rect 126736 -400 126792 240
rect 127327 -400 127383 240
rect 127918 -400 127974 240
rect 128509 -400 128565 240
rect 129100 -400 129156 240
rect 129691 -400 129747 240
rect 130282 -400 130338 240
rect 130873 -400 130929 240
rect 131464 -400 131520 240
rect 132055 -400 132111 240
rect 132646 -400 132702 240
rect 133237 -400 133293 240
rect 133828 -400 133884 240
rect 134419 -400 134475 240
rect 135010 -400 135066 240
rect 135601 -400 135657 240
rect 136192 -400 136248 240
rect 136783 -400 136839 240
rect 137374 -400 137430 240
rect 137965 -400 138021 240
rect 138556 -400 138612 240
rect 139147 -400 139203 240
rect 139738 -400 139794 240
rect 140329 -400 140385 240
rect 140920 -400 140976 240
rect 141511 -400 141567 240
rect 142102 -400 142158 240
rect 142693 -400 142749 240
rect 143284 -400 143340 240
rect 143875 -400 143931 240
rect 144466 -400 144522 240
rect 145057 -400 145113 240
rect 145648 -400 145704 240
rect 146239 -400 146295 240
rect 146830 -400 146886 240
rect 147421 -400 147477 240
rect 148012 -400 148068 240
rect 148603 -400 148659 240
rect 149194 -400 149250 240
rect 149785 -400 149841 240
rect 150376 -400 150432 240
rect 150967 -400 151023 240
rect 151558 -400 151614 240
rect 152149 -400 152205 240
rect 152740 -400 152796 240
rect 153331 -400 153387 240
rect 153922 -400 153978 240
rect 154513 -400 154569 240
rect 155104 -400 155160 240
rect 155695 -400 155751 240
rect 156286 -400 156342 240
rect 156877 -400 156933 240
rect 157468 -400 157524 240
rect 158059 -400 158115 240
rect 158650 -400 158706 240
rect 159241 -400 159297 240
rect 159832 -400 159888 240
rect 160423 -400 160479 240
rect 161014 -400 161070 240
rect 161605 -400 161661 240
rect 162196 -400 162252 240
rect 162787 -400 162843 240
rect 163378 -400 163434 240
rect 163969 -400 164025 240
rect 164560 -400 164616 240
rect 165151 -400 165207 240
rect 165742 -400 165798 240
rect 166333 -400 166389 240
rect 166924 -400 166980 240
rect 167515 -400 167571 240
rect 168106 -400 168162 240
rect 168697 -400 168753 240
rect 169288 -400 169344 240
rect 169879 -400 169935 240
rect 170470 -400 170526 240
rect 171061 -400 171117 240
rect 171652 -400 171708 240
rect 172243 -400 172299 240
rect 172834 -400 172890 240
rect 173425 -400 173481 240
rect 174016 -400 174072 240
rect 174607 -400 174663 240
rect 175198 -400 175254 240
rect 175789 -400 175845 240
rect 176380 -400 176436 240
rect 176971 -400 177027 240
rect 177562 -400 177618 240
rect 178153 -400 178209 240
rect 178744 -400 178800 240
rect 179335 -400 179391 240
rect 179926 -400 179982 240
rect 180517 -400 180573 240
rect 181108 -400 181164 240
rect 181699 -400 181755 240
rect 182290 -400 182346 240
rect 182881 -400 182937 240
rect 183472 -400 183528 240
rect 184063 -400 184119 240
rect 184654 -400 184710 240
rect 185245 -400 185301 240
rect 185836 -400 185892 240
rect 186427 -400 186483 240
rect 187018 -400 187074 240
rect 187609 -400 187665 240
rect 188200 -400 188256 240
rect 188791 -400 188847 240
rect 189382 -400 189438 240
rect 189973 -400 190029 240
rect 190564 -400 190620 240
rect 191155 -400 191211 240
rect 191746 -400 191802 240
rect 192337 -400 192393 240
rect 192928 -400 192984 240
rect 193519 -400 193575 240
rect 194110 -400 194166 240
rect 194701 -400 194757 240
rect 195292 -400 195348 240
rect 195883 -400 195939 240
rect 196474 -400 196530 240
rect 197065 -400 197121 240
rect 197656 -400 197712 240
rect 198247 -400 198303 240
rect 198838 -400 198894 240
rect 199429 -400 199485 240
rect 200020 -400 200076 240
rect 200611 -400 200667 240
rect 201202 -400 201258 240
rect 201793 -400 201849 240
rect 202384 -400 202440 240
rect 202975 -400 203031 240
rect 203566 -400 203622 240
rect 204157 -400 204213 240
rect 204748 -400 204804 240
rect 205339 -400 205395 240
rect 205930 -400 205986 240
rect 206521 -400 206577 240
rect 207112 -400 207168 240
rect 207703 -400 207759 240
rect 208294 -400 208350 240
rect 208885 -400 208941 240
rect 209476 -400 209532 240
rect 210067 -400 210123 240
rect 210658 -400 210714 240
rect 211249 -400 211305 240
rect 211840 -400 211896 240
rect 212431 -400 212487 240
rect 213022 -400 213078 240
rect 213613 -400 213669 240
rect 214204 -400 214260 240
rect 214795 -400 214851 240
rect 215386 -400 215442 240
rect 215977 -400 216033 240
rect 216568 -400 216624 240
rect 217159 -400 217215 240
rect 217750 -400 217806 240
rect 218341 -400 218397 240
rect 218932 -400 218988 240
rect 219523 -400 219579 240
rect 220114 -400 220170 240
rect 220705 -400 220761 240
rect 221296 -400 221352 240
rect 221887 -400 221943 240
rect 222478 -400 222534 240
rect 223069 -400 223125 240
rect 223660 -400 223716 240
rect 224251 -400 224307 240
rect 224842 -400 224898 240
rect 225433 -400 225489 240
rect 226024 -400 226080 240
rect 226615 -400 226671 240
rect 227206 -400 227262 240
rect 227797 -400 227853 240
rect 228388 -400 228444 240
rect 228979 -400 229035 240
rect 229570 -400 229626 240
rect 230161 -400 230217 240
rect 230752 -400 230808 240
rect 231343 -400 231399 240
rect 231934 -400 231990 240
rect 232525 -400 232581 240
rect 233116 -400 233172 240
rect 233707 -400 233763 240
rect 234298 -400 234354 240
rect 234889 -400 234945 240
rect 235480 -400 235536 240
rect 236071 -400 236127 240
rect 236662 -400 236718 240
rect 237253 -400 237309 240
rect 237844 -400 237900 240
rect 238435 -400 238491 240
rect 239026 -400 239082 240
rect 239617 -400 239673 240
rect 240208 -400 240264 240
rect 240799 -400 240855 240
rect 241390 -400 241446 240
rect 241981 -400 242037 240
rect 242572 -400 242628 240
rect 243163 -400 243219 240
rect 243754 -400 243810 240
rect 244345 -400 244401 240
rect 244936 -400 244992 240
rect 245527 -400 245583 240
rect 246118 -400 246174 240
rect 246709 -400 246765 240
rect 247300 -400 247356 240
rect 247891 -400 247947 240
rect 248482 -400 248538 240
rect 249073 -400 249129 240
rect 249664 -400 249720 240
rect 250255 -400 250311 240
rect 250846 -400 250902 240
rect 251437 -400 251493 240
rect 252028 -400 252084 240
rect 252619 -400 252675 240
rect 253210 -400 253266 240
rect 253801 -400 253857 240
rect 254392 -400 254448 240
rect 254983 -400 255039 240
rect 255574 -400 255630 240
rect 256165 -400 256221 240
rect 256756 -400 256812 240
rect 257347 -400 257403 240
rect 257938 -400 257994 240
rect 258529 -400 258585 240
rect 259120 -400 259176 240
rect 259711 -400 259767 240
rect 260302 -400 260358 240
rect 260893 -400 260949 240
rect 261484 -400 261540 240
rect 262075 -400 262131 240
rect 262666 -400 262722 240
rect 263257 -400 263313 240
rect 263848 -400 263904 240
rect 264439 -400 264495 240
rect 265030 -400 265086 240
rect 265621 -400 265677 240
rect 266212 -400 266268 240
rect 266803 -400 266859 240
rect 267394 -400 267450 240
rect 267985 -400 268041 240
rect 268576 -400 268632 240
rect 269167 -400 269223 240
rect 269758 -400 269814 240
rect 270349 -400 270405 240
rect 270940 -400 270996 240
rect 271531 -400 271587 240
rect 272122 -400 272178 240
rect 272713 -400 272769 240
rect 273304 -400 273360 240
rect 273895 -400 273951 240
rect 274486 -400 274542 240
rect 275077 -400 275133 240
rect 275668 -400 275724 240
rect 276259 -400 276315 240
rect 276850 -400 276906 240
rect 277441 -400 277497 240
rect 278032 -400 278088 240
rect 278623 -400 278679 240
rect 279214 -400 279270 240
rect 279805 -400 279861 240
rect 280396 -400 280452 240
rect 280987 -400 281043 240
rect 281578 -400 281634 240
rect 282169 -400 282225 240
rect 282760 -400 282816 240
rect 283351 -400 283407 240
rect 283942 -400 283998 240
rect 284533 -400 284589 240
rect 285124 -400 285180 240
rect 285715 -400 285771 240
rect 286306 -400 286362 240
rect 286897 -400 286953 240
rect 287488 -400 287544 240
rect 288079 -400 288135 240
rect 288670 -400 288726 240
rect 289261 -400 289317 240
rect 289852 -400 289908 240
rect 290443 -400 290499 240
rect 291034 -400 291090 240
rect 291625 -400 291681 240
<< via2 >>
rect 271865 351785 271895 351815
rect 272025 351785 272055 351815
rect 272105 351785 272135 351815
rect 272185 351785 272215 351815
rect 272265 351785 272295 351815
rect 272345 351785 272375 351815
rect 272425 351785 272455 351815
rect 272505 351785 272535 351815
rect 272585 351785 272615 351815
rect 272665 351785 272695 351815
rect 272745 351785 272775 351815
rect 272825 351785 272855 351815
rect 272905 351785 272935 351815
rect 272985 351785 273015 351815
rect 273065 351785 273095 351815
rect 273145 351785 273175 351815
rect 273225 351785 273255 351815
rect 273305 351785 273335 351815
rect 273385 351785 273415 351815
rect 273465 351785 273495 351815
rect 273545 351785 273575 351815
rect 273625 351785 273655 351815
rect 273705 351785 273735 351815
rect 273785 351785 273815 351815
rect 273865 351785 273895 351815
rect 273945 351785 273975 351815
rect 274025 351785 274055 351815
rect 274105 351785 274135 351815
rect 274185 351785 274215 351815
rect 274265 351785 274295 351815
rect 274345 351785 274375 351815
rect 274425 351785 274455 351815
rect 274505 351785 274535 351815
rect 274585 351785 274615 351815
rect 274665 351785 274695 351815
rect 274745 351785 274775 351815
rect 274825 351785 274855 351815
rect 274905 351785 274935 351815
rect 274985 351785 275015 351815
rect 275065 351785 275095 351815
rect 275145 351785 275175 351815
rect 275225 351785 275255 351815
rect 275305 351785 275335 351815
rect 275385 351785 275415 351815
rect 275465 351785 275495 351815
rect 275545 351785 275575 351815
rect 275625 351785 275655 351815
rect 275705 351785 275735 351815
rect 275785 351785 275815 351815
rect 275865 351785 275895 351815
rect 275945 351785 275975 351815
rect 276025 351785 276055 351815
rect 276105 351785 276135 351815
rect 276185 351785 276215 351815
rect 276265 351785 276295 351815
rect 276345 351785 276375 351815
rect 276425 351785 276455 351815
rect 276505 351785 276535 351815
rect 276585 351785 276615 351815
rect 276665 351785 276695 351815
rect 276745 351785 276775 351815
rect 276825 351785 276855 351815
rect 276905 351785 276935 351815
rect 276985 351785 277015 351815
rect 277065 351785 277095 351815
rect 277145 351785 277175 351815
rect 277225 351785 277255 351815
rect 277305 351785 277335 351815
rect 277385 351785 277415 351815
rect 277465 351785 277495 351815
rect 277545 351785 277575 351815
rect 277625 351785 277655 351815
rect 277705 351785 277735 351815
rect 277785 351785 277815 351815
rect 277865 351785 277895 351815
rect 277945 351785 277975 351815
rect 278025 351785 278055 351815
rect 278105 351785 278135 351815
rect 278185 351785 278215 351815
rect 278265 351785 278295 351815
rect 278345 351785 278375 351815
rect 278425 351785 278455 351815
rect 278505 351785 278535 351815
rect 278585 351785 278615 351815
rect 278665 351785 278695 351815
rect 278745 351785 278775 351815
rect 278825 351785 278855 351815
rect 278905 351785 278935 351815
rect 278985 351785 279015 351815
rect 279065 351785 279095 351815
rect 279145 351785 279175 351815
rect 279225 351785 279255 351815
rect 279305 351785 279335 351815
rect 279385 351785 279415 351815
rect 279465 351785 279495 351815
rect 279545 351785 279575 351815
rect 279625 351785 279655 351815
rect 279705 351785 279735 351815
rect 279785 351785 279815 351815
rect 279865 351785 279895 351815
rect 279945 351785 279975 351815
rect 280025 351785 280055 351815
rect 280105 351785 280135 351815
rect 280185 351785 280215 351815
rect 280265 351785 280295 351815
rect 280345 351785 280375 351815
rect 280425 351785 280455 351815
rect 280505 351785 280535 351815
rect 280585 351785 280615 351815
rect 280665 351785 280695 351815
rect 280745 351785 280775 351815
rect 280825 351785 280855 351815
rect 280905 351785 280935 351815
rect 280985 351785 281015 351815
rect 281065 351785 281095 351815
rect 281145 351785 281175 351815
rect 281225 351785 281255 351815
rect 281305 351785 281335 351815
rect 281385 351785 281415 351815
rect 281465 351785 281495 351815
rect 281545 351785 281575 351815
rect 281625 351785 281655 351815
rect 281705 351785 281735 351815
rect 281785 351785 281815 351815
rect 281865 351785 281895 351815
rect 281945 351785 281975 351815
rect 282025 351785 282055 351815
rect 282105 351785 282135 351815
rect 282185 351785 282215 351815
rect 282265 351785 282295 351815
rect 282345 351785 282375 351815
rect 282425 351785 282455 351815
rect 282505 351785 282535 351815
rect 282585 351785 282615 351815
rect 282665 351785 282695 351815
rect 282745 351785 282775 351815
rect 282825 351785 282855 351815
rect 282905 351785 282935 351815
rect 282985 351785 283015 351815
rect 283065 351785 283095 351815
rect 283145 351785 283175 351815
rect 271945 351705 271975 351735
rect 283225 351705 283255 351735
rect 271865 351625 271895 351655
rect 272025 351625 272055 351655
rect 272105 351625 272135 351655
rect 272185 351625 272215 351655
rect 272265 351625 272295 351655
rect 272345 351625 272375 351655
rect 272425 351625 272455 351655
rect 272505 351625 272535 351655
rect 272585 351625 272615 351655
rect 272665 351625 272695 351655
rect 272745 351625 272775 351655
rect 272825 351625 272855 351655
rect 272905 351625 272935 351655
rect 272985 351625 273015 351655
rect 273065 351625 273095 351655
rect 273145 351625 273175 351655
rect 273225 351625 273255 351655
rect 273305 351625 273335 351655
rect 273385 351625 273415 351655
rect 273465 351625 273495 351655
rect 273545 351625 273575 351655
rect 273625 351625 273655 351655
rect 273705 351625 273735 351655
rect 273785 351625 273815 351655
rect 273865 351625 273895 351655
rect 273945 351625 273975 351655
rect 274025 351625 274055 351655
rect 274105 351625 274135 351655
rect 274185 351625 274215 351655
rect 274265 351625 274295 351655
rect 274345 351625 274375 351655
rect 274425 351625 274455 351655
rect 274505 351625 274535 351655
rect 274585 351625 274615 351655
rect 274665 351625 274695 351655
rect 274745 351625 274775 351655
rect 274825 351625 274855 351655
rect 274905 351625 274935 351655
rect 274985 351625 275015 351655
rect 275065 351625 275095 351655
rect 275145 351625 275175 351655
rect 275225 351625 275255 351655
rect 275305 351625 275335 351655
rect 275385 351625 275415 351655
rect 275465 351625 275495 351655
rect 275545 351625 275575 351655
rect 275625 351625 275655 351655
rect 275705 351625 275735 351655
rect 275785 351625 275815 351655
rect 275865 351625 275895 351655
rect 275945 351625 275975 351655
rect 276025 351625 276055 351655
rect 276105 351625 276135 351655
rect 276185 351625 276215 351655
rect 276265 351625 276295 351655
rect 276345 351625 276375 351655
rect 276425 351625 276455 351655
rect 276505 351625 276535 351655
rect 276585 351625 276615 351655
rect 276665 351625 276695 351655
rect 276745 351625 276775 351655
rect 276825 351625 276855 351655
rect 276905 351625 276935 351655
rect 276985 351625 277015 351655
rect 277065 351625 277095 351655
rect 277145 351625 277175 351655
rect 277225 351625 277255 351655
rect 277305 351625 277335 351655
rect 277385 351625 277415 351655
rect 277465 351625 277495 351655
rect 277545 351625 277575 351655
rect 277625 351625 277655 351655
rect 277705 351625 277735 351655
rect 277785 351625 277815 351655
rect 277865 351625 277895 351655
rect 277945 351625 277975 351655
rect 278025 351625 278055 351655
rect 278105 351625 278135 351655
rect 278185 351625 278215 351655
rect 278265 351625 278295 351655
rect 278345 351625 278375 351655
rect 278425 351625 278455 351655
rect 278505 351625 278535 351655
rect 278585 351625 278615 351655
rect 278665 351625 278695 351655
rect 278745 351625 278775 351655
rect 278825 351625 278855 351655
rect 278905 351625 278935 351655
rect 278985 351625 279015 351655
rect 279065 351625 279095 351655
rect 279145 351625 279175 351655
rect 279225 351625 279255 351655
rect 279305 351625 279335 351655
rect 279385 351625 279415 351655
rect 279465 351625 279495 351655
rect 279545 351625 279575 351655
rect 279625 351625 279655 351655
rect 279705 351625 279735 351655
rect 279785 351625 279815 351655
rect 279865 351625 279895 351655
rect 279945 351625 279975 351655
rect 280025 351625 280055 351655
rect 280105 351625 280135 351655
rect 280185 351625 280215 351655
rect 280265 351625 280295 351655
rect 280345 351625 280375 351655
rect 280425 351625 280455 351655
rect 280505 351625 280535 351655
rect 280585 351625 280615 351655
rect 280665 351625 280695 351655
rect 280745 351625 280775 351655
rect 280825 351625 280855 351655
rect 280905 351625 280935 351655
rect 280985 351625 281015 351655
rect 281065 351625 281095 351655
rect 281145 351625 281175 351655
rect 281225 351625 281255 351655
rect 281305 351625 281335 351655
rect 281385 351625 281415 351655
rect 281465 351625 281495 351655
rect 281545 351625 281575 351655
rect 281625 351625 281655 351655
rect 281705 351625 281735 351655
rect 281785 351625 281815 351655
rect 281865 351625 281895 351655
rect 281945 351625 281975 351655
rect 282025 351625 282055 351655
rect 282105 351625 282135 351655
rect 282185 351625 282215 351655
rect 282265 351625 282295 351655
rect 282345 351625 282375 351655
rect 282425 351625 282455 351655
rect 282505 351625 282535 351655
rect 282585 351625 282615 351655
rect 282665 351625 282695 351655
rect 282745 351625 282775 351655
rect 282825 351625 282855 351655
rect 282905 351625 282935 351655
rect 282985 351625 283015 351655
rect 283065 351625 283095 351655
rect 283145 351625 283175 351655
rect 271865 351545 271895 351575
rect 272025 351545 272055 351575
rect 271865 351465 271895 351495
rect 272025 351465 272055 351495
rect 271865 351385 271895 351415
rect 272025 351385 272055 351415
rect 271865 351305 271895 351335
rect 272025 351305 272055 351335
rect 271865 351225 271895 351255
rect 272025 351225 272055 351255
rect 271865 351145 271895 351175
rect 272025 351145 272055 351175
rect 271865 351065 271895 351095
rect 272025 351065 272055 351095
rect 271865 350985 271895 351015
rect 272025 350985 272055 351015
rect 271865 350905 271895 350935
rect 272025 350905 272055 350935
rect 271865 350825 271895 350855
rect 272025 350825 272055 350855
rect 271865 350745 271895 350775
rect 272025 350745 272055 350775
rect 271865 350665 271895 350695
rect 272025 350665 272055 350695
rect 271865 350585 271895 350615
rect 272025 350585 272055 350615
rect 271865 350505 271895 350535
rect 272025 350505 272055 350535
rect 271865 350425 271895 350455
rect 272025 350425 272055 350455
rect 271865 350345 271895 350375
rect 272025 350345 272055 350375
rect 271865 350265 271895 350295
rect 272025 350265 272055 350295
rect 271865 350185 271895 350215
rect 272025 350185 272055 350215
rect 271865 350105 271895 350135
rect 272025 350105 272055 350135
rect 271865 350025 271895 350055
rect 272025 350025 272055 350055
rect 16725 275445 16755 275475
rect 16885 275445 16915 275475
rect 16965 275445 16995 275475
rect 17045 275445 17075 275475
rect 17125 275445 17155 275475
rect 17205 275445 17235 275475
rect 16805 275365 16835 275395
rect 17125 275365 17155 275395
rect 28405 275325 28435 275355
rect 28565 275325 28595 275355
rect 28725 275325 28755 275355
rect 16725 275285 16755 275315
rect 16885 275285 16915 275315
rect 16965 275285 16995 275315
rect 17045 275285 17075 275315
rect 17205 275285 17235 275315
rect 28405 275245 28435 275275
rect 28565 275245 28595 275275
rect 28725 275245 28755 275275
rect 1040 275040 1160 275160
rect 13525 275005 13555 275195
rect 13685 275005 13715 275195
rect 13845 275005 13875 275195
rect 14005 275005 14035 275195
rect 14165 275005 14195 275195
rect 14325 275005 14355 275195
rect 27925 275005 27955 275195
rect 28085 275005 28115 275195
rect 28245 275005 28275 275195
rect 28405 275005 28435 275195
rect 28565 275005 28595 275195
rect 28725 275005 28755 275195
rect 258910 275010 259090 275190
rect 16725 274925 16755 274955
rect 16885 274925 16915 274955
rect 16725 274845 16755 274875
rect 16885 274845 16915 274875
rect 16725 274765 16755 274795
rect 16885 274765 16915 274795
rect 16725 274685 16755 274715
rect 16885 274685 16915 274715
rect 16725 274605 16755 274635
rect 16885 274605 16915 274635
rect 16725 274525 16755 274555
rect 16885 274525 16915 274555
rect 16725 274445 16755 274475
rect 16885 274445 16915 274475
rect 16725 274365 16755 274395
rect 16885 274365 16915 274395
rect 16725 274285 16755 274315
rect 16885 274285 16915 274315
rect 16725 274205 16755 274235
rect 16885 274205 16915 274235
rect 16725 274125 16755 274155
rect 16885 274125 16915 274155
rect 16725 274045 16755 274075
rect 16885 274045 16915 274075
rect 16725 273965 16755 273995
rect 16885 273965 16915 273995
rect 16725 273885 16755 273915
rect 16885 273885 16915 273915
rect 16725 273805 16755 273835
rect 16885 273805 16915 273835
rect 16725 273725 16755 273755
rect 16885 273725 16915 273755
rect 16725 273645 16755 273675
rect 16885 273645 16915 273675
rect 16725 273565 16755 273595
rect 16885 273565 16915 273595
rect 16725 273485 16755 273515
rect 16885 273485 16915 273515
rect 16725 273405 16755 273435
rect 16885 273405 16915 273435
rect 16725 273325 16755 273355
rect 16885 273325 16915 273355
rect 16725 273245 16755 273275
rect 16885 273245 16915 273275
rect 16725 273165 16755 273195
rect 16885 273165 16915 273195
rect 16725 273085 16755 273115
rect 16885 273085 16915 273115
rect 16725 273005 16755 273035
rect 16885 273005 16915 273035
rect 16725 272925 16755 272955
rect 16885 272925 16915 272955
rect 16725 272845 16755 272875
rect 16885 272845 16915 272875
rect 16725 272765 16755 272795
rect 16885 272765 16915 272795
rect 16725 272685 16755 272715
rect 16885 272685 16915 272715
rect 16725 272605 16755 272635
rect 16885 272605 16915 272635
rect 16725 272525 16755 272555
rect 16885 272525 16915 272555
rect 16725 272445 16755 272475
rect 16885 272445 16915 272475
rect 16725 272365 16755 272395
rect 16885 272365 16915 272395
rect 16725 272285 16755 272315
rect 16885 272285 16915 272315
rect 16725 272205 16755 272235
rect 16885 272205 16915 272235
rect 16725 272125 16755 272155
rect 16885 272125 16915 272155
rect 16725 272045 16755 272075
rect 16885 272045 16915 272075
rect 16725 271965 16755 271995
rect 16885 271965 16915 271995
rect 16725 271885 16755 271915
rect 16885 271885 16915 271915
rect 16725 271805 16755 271835
rect 16885 271805 16915 271835
rect 16725 271725 16755 271755
rect 16885 271725 16915 271755
rect 16725 271645 16755 271675
rect 16885 271645 16915 271675
rect 16725 271565 16755 271595
rect 16885 271565 16915 271595
rect 16725 271485 16755 271515
rect 16885 271485 16915 271515
rect 16725 271405 16755 271435
rect 16885 271405 16915 271435
rect 16725 271325 16755 271355
rect 16885 271325 16915 271355
rect 16725 271245 16755 271275
rect 16885 271245 16915 271275
rect 16725 271165 16755 271195
rect 16885 271165 16915 271195
rect 16725 271085 16755 271115
rect 16885 271085 16915 271115
rect 16725 271005 16755 271035
rect 16885 271005 16915 271035
rect 16725 270925 16755 270955
rect 16885 270925 16915 270955
rect 16725 270845 16755 270875
rect 16885 270845 16915 270875
rect 16725 270765 16755 270795
rect 16885 270765 16915 270795
rect 16725 270685 16755 270715
rect 16885 270685 16915 270715
rect 16725 270605 16755 270635
rect 16885 270605 16915 270635
rect 16725 270525 16755 270555
rect 16885 270525 16915 270555
rect 16725 270445 16755 270475
rect 16885 270445 16915 270475
rect 16725 270365 16755 270395
rect 16885 270365 16915 270395
rect 16725 270285 16755 270315
rect 16885 270285 16915 270315
rect 16725 270205 16755 270235
rect 16885 270205 16915 270235
rect 16725 270125 16755 270155
rect 16885 270125 16915 270155
rect 16725 270045 16755 270075
rect 16885 270045 16915 270075
rect 16725 269965 16755 269995
rect 16885 269965 16915 269995
rect 16725 269885 16755 269915
rect 16885 269885 16915 269915
rect 16725 269805 16755 269835
rect 16885 269805 16915 269835
rect 16725 269725 16755 269755
rect 16885 269725 16915 269755
rect 16725 269645 16755 269675
rect 16885 269645 16915 269675
rect 16725 269565 16755 269595
rect 16885 269565 16915 269595
rect 16725 269485 16755 269515
rect 16885 269485 16915 269515
rect 16725 269405 16755 269435
rect 16885 269405 16915 269435
rect 16725 269325 16755 269355
rect 16885 269325 16915 269355
rect 16725 269245 16755 269275
rect 16885 269245 16915 269275
rect 16725 269165 16755 269195
rect 16885 269165 16915 269195
rect 16725 269085 16755 269115
rect 16885 269085 16915 269115
rect 16725 269005 16755 269035
rect 16885 269005 16915 269035
rect 16725 268925 16755 268955
rect 16885 268925 16915 268955
rect 16725 268845 16755 268875
rect 16885 268845 16915 268875
rect 16725 268765 16755 268795
rect 16885 268765 16915 268795
rect 16725 268685 16755 268715
rect 16885 268685 16915 268715
rect 16725 268605 16755 268635
rect 16885 268605 16915 268635
rect 16725 268525 16755 268555
rect 16885 268525 16915 268555
rect 16725 268445 16755 268475
rect 16885 268445 16915 268475
rect 16725 268365 16755 268395
rect 16885 268365 16915 268395
rect 16725 268285 16755 268315
rect 16885 268285 16915 268315
rect 16725 268205 16755 268235
rect 16885 268205 16915 268235
rect 16725 268125 16755 268155
rect 16885 268125 16915 268155
rect 16725 268045 16755 268075
rect 16885 268045 16915 268075
rect 16725 267965 16755 267995
rect 16885 267965 16915 267995
rect 16725 267885 16755 267915
rect 16885 267885 16915 267915
rect 16725 267805 16755 267835
rect 16885 267805 16915 267835
rect 16725 267725 16755 267755
rect 16885 267725 16915 267755
rect 16725 267645 16755 267675
rect 16885 267645 16915 267675
rect 16725 267565 16755 267595
rect 16885 267565 16915 267595
rect 16725 267485 16755 267515
rect 16885 267485 16915 267515
rect 16725 267405 16755 267435
rect 16885 267405 16915 267435
rect 16725 267325 16755 267355
rect 16885 267325 16915 267355
rect 16725 267245 16755 267275
rect 16885 267245 16915 267275
rect 16725 267165 16755 267195
rect 16885 267165 16915 267195
rect 16725 267085 16755 267115
rect 16885 267085 16915 267115
rect 16725 267005 16755 267035
rect 16885 267005 16915 267035
rect 16725 266925 16755 266955
rect 16885 266925 16915 266955
rect 16725 266845 16755 266875
rect 16885 266845 16915 266875
rect 16725 266765 16755 266795
rect 16885 266765 16915 266795
rect 16725 266685 16755 266715
rect 16885 266685 16915 266715
rect 16725 266605 16755 266635
rect 16885 266605 16915 266635
rect 16725 266525 16755 266555
rect 16885 266525 16915 266555
rect 16725 266445 16755 266475
rect 16885 266445 16915 266475
rect 16725 266365 16755 266395
rect 16885 266365 16915 266395
rect 16725 266285 16755 266315
rect 16885 266285 16915 266315
rect 16725 266205 16755 266235
rect 16885 266205 16915 266235
rect 16725 266125 16755 266155
rect 16885 266125 16915 266155
rect 16725 266045 16755 266075
rect 16885 266045 16915 266075
rect 16725 265965 16755 265995
rect 16885 265965 16915 265995
rect 16725 265885 16755 265915
rect 16885 265885 16915 265915
rect 16725 265805 16755 265835
rect 16885 265805 16915 265835
rect 16725 265725 16755 265755
rect 16885 265725 16915 265755
rect 16725 265645 16755 265675
rect 16885 265645 16915 265675
rect 16725 265565 16755 265595
rect 16885 265565 16915 265595
rect 16725 265485 16755 265515
rect 16885 265485 16915 265515
rect 16725 265405 16755 265435
rect 16885 265405 16915 265435
rect 16725 265325 16755 265355
rect 16885 265325 16915 265355
rect 16725 265245 16755 265275
rect 16885 265245 16915 265275
rect 16725 265165 16755 265195
rect 16885 265165 16915 265195
rect 16725 265085 16755 265115
rect 16885 265085 16915 265115
rect 16725 265005 16755 265035
rect 16885 265005 16915 265035
rect 16725 264925 16755 264955
rect 16885 264925 16915 264955
rect 16725 264845 16755 264875
rect 16885 264845 16915 264875
rect 16725 264765 16755 264795
rect 16885 264765 16915 264795
rect 16725 264685 16755 264715
rect 16885 264685 16915 264715
rect 16725 264605 16755 264635
rect 16885 264605 16915 264635
rect 16725 264525 16755 264555
rect 16885 264525 16915 264555
rect 16725 264445 16755 264475
rect 16885 264445 16915 264475
rect 16725 264365 16755 264395
rect 16885 264365 16915 264395
rect 16725 264285 16755 264315
rect 16885 264285 16915 264315
rect 16725 264205 16755 264235
rect 16885 264205 16915 264235
rect 16725 264125 16755 264155
rect 16885 264125 16915 264155
rect 16725 264045 16755 264075
rect 16885 264045 16915 264075
rect 16725 263965 16755 263995
rect 16885 263965 16915 263995
rect 16725 263885 16755 263915
rect 16885 263885 16915 263915
rect 16725 263805 16755 263835
rect 16885 263805 16915 263835
rect 16725 263725 16755 263755
rect 16885 263725 16915 263755
rect 16725 263645 16755 263675
rect 16885 263645 16915 263675
rect 16725 263565 16755 263595
rect 16885 263565 16915 263595
rect 16725 263485 16755 263515
rect 16885 263485 16915 263515
rect 16725 263405 16755 263435
rect 16885 263405 16915 263435
rect 16725 263325 16755 263355
rect 16885 263325 16915 263355
rect 16725 263245 16755 263275
rect 16885 263245 16915 263275
rect 16725 263165 16755 263195
rect 16885 263165 16915 263195
rect 16725 263085 16755 263115
rect 16885 263085 16915 263115
rect 16725 263005 16755 263035
rect 16885 263005 16915 263035
rect 16725 262925 16755 262955
rect 16885 262925 16915 262955
rect 16725 262845 16755 262875
rect 16885 262845 16915 262875
rect 16725 262765 16755 262795
rect 16885 262765 16915 262795
rect 16725 262685 16755 262715
rect 16885 262685 16915 262715
rect 16725 262605 16755 262635
rect 16885 262605 16915 262635
rect 16725 262525 16755 262555
rect 16885 262525 16915 262555
rect 16725 262445 16755 262475
rect 16885 262445 16915 262475
rect 16725 262365 16755 262395
rect 16885 262365 16915 262395
rect 16725 262285 16755 262315
rect 16885 262285 16915 262315
rect 16725 262205 16755 262235
rect 16885 262205 16915 262235
rect 16725 262125 16755 262155
rect 16885 262125 16915 262155
rect 16725 262045 16755 262075
rect 16885 262045 16915 262075
rect 16725 261965 16755 261995
rect 16885 261965 16915 261995
rect 16725 261885 16755 261915
rect 16885 261885 16915 261915
rect 16725 261805 16755 261835
rect 16885 261805 16915 261835
rect 16725 261725 16755 261755
rect 16885 261725 16915 261755
rect 16725 261645 16755 261675
rect 16885 261645 16915 261675
rect 16725 261565 16755 261595
rect 16885 261565 16915 261595
rect 16725 261485 16755 261515
rect 16885 261485 16915 261515
rect 16725 261405 16755 261435
rect 16885 261405 16915 261435
rect 16725 261325 16755 261355
rect 16885 261325 16915 261355
rect 16725 261245 16755 261275
rect 16885 261245 16915 261275
rect 16725 261165 16755 261195
rect 16885 261165 16915 261195
rect 16725 261085 16755 261115
rect 16885 261085 16915 261115
rect 16725 261005 16755 261035
rect 16885 261005 16915 261035
rect 16725 260925 16755 260955
rect 16885 260925 16915 260955
rect 16725 260845 16755 260875
rect 16885 260845 16915 260875
rect 16725 260765 16755 260795
rect 16885 260765 16915 260795
rect 16725 260685 16755 260715
rect 16885 260685 16915 260715
rect 16725 260605 16755 260635
rect 16885 260605 16915 260635
rect 16725 260525 16755 260555
rect 16885 260525 16915 260555
rect 16725 260445 16755 260475
rect 16885 260445 16915 260475
rect 16725 260365 16755 260395
rect 16885 260365 16915 260395
rect 16725 260285 16755 260315
rect 16885 260285 16915 260315
rect 16725 260205 16755 260235
rect 16885 260205 16915 260235
rect 16725 260125 16755 260155
rect 16885 260125 16915 260155
rect 16725 260045 16755 260075
rect 16885 260045 16915 260075
rect 16725 259965 16755 259995
rect 16885 259965 16915 259995
rect 16725 259885 16755 259915
rect 16885 259885 16915 259915
rect 16725 259805 16755 259835
rect 16885 259805 16915 259835
rect 16725 259725 16755 259755
rect 16885 259725 16915 259755
rect 16725 259645 16755 259675
rect 16885 259645 16915 259675
rect 16725 259565 16755 259595
rect 16885 259565 16915 259595
rect 16725 259485 16755 259515
rect 16885 259485 16915 259515
rect 16725 259405 16755 259435
rect 16885 259405 16915 259435
rect 16725 259325 16755 259355
rect 16885 259325 16915 259355
rect 16725 259245 16755 259275
rect 16885 259245 16915 259275
rect 16725 259165 16755 259195
rect 16885 259165 16915 259195
rect 16725 259085 16755 259115
rect 16885 259085 16915 259115
rect 16725 259005 16755 259035
rect 16885 259005 16915 259035
rect 16725 258925 16755 258955
rect 16885 258925 16915 258955
rect 16725 258845 16755 258875
rect 16885 258845 16915 258875
rect 16725 258765 16755 258795
rect 16885 258765 16915 258795
rect 16725 258685 16755 258715
rect 16885 258685 16915 258715
rect 16725 258605 16755 258635
rect 16885 258605 16915 258635
rect 16725 258525 16755 258555
rect 16885 258525 16915 258555
rect 16725 258445 16755 258475
rect 16885 258445 16915 258475
rect 16725 258365 16755 258395
rect 16885 258365 16915 258395
rect 16725 258285 16755 258315
rect 16885 258285 16915 258315
rect 16725 258205 16755 258235
rect 16885 258205 16915 258235
rect 16725 258125 16755 258155
rect 16885 258125 16915 258155
rect 16725 258045 16755 258075
rect 16885 258045 16915 258075
rect 16725 257965 16755 257995
rect 16885 257965 16915 257995
rect 16725 257885 16755 257915
rect 16885 257885 16915 257915
rect 16725 257805 16755 257835
rect 16885 257805 16915 257835
rect 16725 257725 16755 257755
rect 16885 257725 16915 257755
rect 16725 257645 16755 257675
rect 16885 257645 16915 257675
rect 16725 257565 16755 257595
rect 16885 257565 16915 257595
rect 16725 257485 16755 257515
rect 16885 257485 16915 257515
rect 16725 257405 16755 257435
rect 16885 257405 16915 257435
rect 16725 257325 16755 257355
rect 16885 257325 16915 257355
rect 16725 257245 16755 257275
rect 16885 257245 16915 257275
rect 16725 257165 16755 257195
rect 16885 257165 16915 257195
rect 16725 257085 16755 257115
rect 16885 257085 16915 257115
rect 16725 257005 16755 257035
rect 16885 257005 16915 257035
rect 16725 256925 16755 256955
rect 16885 256925 16915 256955
rect 16725 256845 16755 256875
rect 16885 256845 16915 256875
rect 16725 256765 16755 256795
rect 16885 256765 16915 256795
rect 16725 256685 16755 256715
rect 16885 256685 16915 256715
rect 16725 256605 16755 256635
rect 16885 256605 16915 256635
rect 16725 256525 16755 256555
rect 16885 256525 16915 256555
rect 16725 256445 16755 256475
rect 16885 256445 16915 256475
rect 16725 256365 16755 256395
rect 16885 256365 16915 256395
rect 16725 256285 16755 256315
rect 16885 256285 16915 256315
rect 16725 256205 16755 256235
rect 16885 256205 16915 256235
rect 16725 256125 16755 256155
rect 16885 256125 16915 256155
rect 16725 256045 16755 256075
rect 16885 256045 16915 256075
rect 16725 255965 16755 255995
rect 16885 255965 16915 255995
rect 405 255845 435 255875
rect 485 255845 515 255875
rect 565 255845 595 255875
rect 645 255845 675 255875
rect 725 255845 755 255875
rect 805 255845 835 255875
rect 885 255845 915 255875
rect 965 255845 995 255875
rect 1045 255845 1075 255875
rect 1125 255845 1155 255875
rect 1205 255845 1235 255875
rect 1285 255845 1315 255875
rect 1365 255845 1395 255875
rect 1445 255845 1475 255875
rect 1525 255845 1555 255875
rect 1605 255845 1635 255875
rect 1685 255845 1715 255875
rect 1765 255845 1795 255875
rect 1845 255845 1875 255875
rect 1925 255845 1955 255875
rect 2005 255845 2035 255875
rect 2085 255845 2115 255875
rect 2165 255845 2195 255875
rect 2245 255845 2275 255875
rect 2325 255845 2355 255875
rect 2405 255845 2435 255875
rect 2485 255845 2515 255875
rect 2565 255845 2595 255875
rect 2645 255845 2675 255875
rect 2725 255845 2755 255875
rect 3045 255845 3075 255875
rect 3125 255845 3155 255875
rect 3205 255845 3235 255875
rect 3285 255845 3315 255875
rect 3365 255845 3395 255875
rect 3445 255845 3475 255875
rect 3525 255845 3555 255875
rect 3605 255845 3635 255875
rect 3685 255845 3715 255875
rect 3765 255845 3795 255875
rect 3845 255845 3875 255875
rect 3925 255845 3955 255875
rect 4005 255845 4035 255875
rect 4085 255845 4115 255875
rect 4165 255845 4195 255875
rect 4245 255845 4275 255875
rect 4325 255845 4355 255875
rect 4405 255845 4435 255875
rect 4485 255845 4515 255875
rect 4565 255845 4595 255875
rect 4645 255845 4675 255875
rect 4725 255845 4755 255875
rect 4805 255845 4835 255875
rect 4885 255845 4915 255875
rect 4965 255845 4995 255875
rect 5045 255845 5075 255875
rect 5125 255845 5155 255875
rect 5205 255845 5235 255875
rect 5285 255845 5315 255875
rect 5365 255845 5395 255875
rect 5445 255845 5475 255875
rect 5525 255845 5555 255875
rect 5605 255845 5635 255875
rect 5685 255845 5715 255875
rect 5765 255845 5795 255875
rect 5845 255845 5875 255875
rect 5925 255845 5955 255875
rect 6005 255845 6035 255875
rect 6085 255845 6115 255875
rect 6165 255845 6195 255875
rect 6245 255845 6275 255875
rect 6325 255845 6355 255875
rect 6405 255845 6435 255875
rect 6485 255845 6515 255875
rect 6565 255845 6595 255875
rect 6645 255845 6675 255875
rect 6725 255845 6755 255875
rect 6805 255845 6835 255875
rect 6885 255845 6915 255875
rect 6965 255845 6995 255875
rect 7045 255845 7075 255875
rect 7125 255845 7155 255875
rect 7205 255845 7235 255875
rect 7285 255845 7315 255875
rect 7365 255845 7395 255875
rect 7445 255845 7475 255875
rect 7525 255845 7555 255875
rect 7605 255845 7635 255875
rect 7685 255845 7715 255875
rect 7765 255845 7795 255875
rect 7845 255845 7875 255875
rect 7925 255845 7955 255875
rect 8005 255845 8035 255875
rect 8085 255845 8115 255875
rect 8165 255845 8195 255875
rect 8245 255845 8275 255875
rect 8325 255845 8355 255875
rect 8405 255845 8435 255875
rect 8485 255845 8515 255875
rect 8565 255845 8595 255875
rect 8645 255845 8675 255875
rect 8725 255845 8755 255875
rect 8805 255845 8835 255875
rect 8885 255845 8915 255875
rect 8965 255845 8995 255875
rect 9045 255845 9075 255875
rect 9125 255845 9155 255875
rect 9205 255845 9235 255875
rect 9285 255845 9315 255875
rect 9365 255845 9395 255875
rect 9445 255845 9475 255875
rect 9525 255845 9555 255875
rect 9605 255845 9635 255875
rect 9685 255845 9715 255875
rect 9765 255845 9795 255875
rect 9845 255845 9875 255875
rect 9925 255845 9955 255875
rect 10005 255845 10035 255875
rect 10085 255845 10115 255875
rect 10165 255845 10195 255875
rect 10245 255845 10275 255875
rect 10325 255845 10355 255875
rect 10405 255845 10435 255875
rect 10485 255845 10515 255875
rect 10565 255845 10595 255875
rect 10645 255845 10675 255875
rect 10725 255845 10755 255875
rect 10805 255845 10835 255875
rect 10885 255845 10915 255875
rect 10965 255845 10995 255875
rect 11045 255845 11075 255875
rect 11125 255845 11155 255875
rect 11205 255845 11235 255875
rect 11285 255845 11315 255875
rect 11365 255845 11395 255875
rect 11445 255845 11475 255875
rect 11525 255845 11555 255875
rect 11605 255845 11635 255875
rect 11685 255845 11715 255875
rect 11765 255845 11795 255875
rect 11845 255845 11875 255875
rect 11925 255845 11955 255875
rect 12005 255845 12035 255875
rect 12085 255845 12115 255875
rect 12165 255845 12195 255875
rect 12245 255845 12275 255875
rect 12325 255845 12355 255875
rect 12405 255845 12435 255875
rect 12485 255845 12515 255875
rect 12565 255845 12595 255875
rect 12645 255845 12675 255875
rect 12725 255845 12755 255875
rect 12805 255845 12835 255875
rect 12885 255845 12915 255875
rect 12965 255845 12995 255875
rect 13045 255845 13075 255875
rect 13125 255845 13155 255875
rect 13205 255845 13235 255875
rect 13285 255845 13315 255875
rect 13365 255845 13395 255875
rect 13445 255845 13475 255875
rect 13525 255845 13555 255875
rect 13605 255845 13635 255875
rect 13685 255845 13715 255875
rect 13765 255845 13795 255875
rect 13845 255845 13875 255875
rect 13925 255845 13955 255875
rect 14005 255845 14035 255875
rect 14085 255845 14115 255875
rect 14165 255845 14195 255875
rect 14245 255845 14275 255875
rect 14325 255845 14355 255875
rect 14405 255845 14435 255875
rect 14485 255845 14515 255875
rect 14565 255845 14595 255875
rect 14645 255845 14675 255875
rect 14725 255845 14755 255875
rect 14805 255845 14835 255875
rect 14885 255845 14915 255875
rect 14965 255845 14995 255875
rect 15045 255845 15075 255875
rect 15125 255845 15155 255875
rect 15205 255845 15235 255875
rect 15285 255845 15315 255875
rect 15365 255845 15395 255875
rect 15445 255845 15475 255875
rect 15525 255845 15555 255875
rect 15605 255845 15635 255875
rect 15685 255845 15715 255875
rect 15765 255845 15795 255875
rect 15845 255845 15875 255875
rect 15925 255845 15955 255875
rect 16005 255845 16035 255875
rect 16085 255845 16115 255875
rect 16165 255845 16195 255875
rect 16245 255845 16275 255875
rect 16325 255845 16355 255875
rect 16405 255845 16435 255875
rect 16485 255845 16515 255875
rect 16565 255845 16595 255875
rect 16645 255845 16675 255875
rect 16725 255845 16755 255875
rect 16885 255845 16915 255875
rect 325 255765 355 255795
rect 16805 255765 16835 255795
rect 405 255685 435 255715
rect 485 255685 515 255715
rect 565 255685 595 255715
rect 645 255685 675 255715
rect 725 255685 755 255715
rect 805 255685 835 255715
rect 885 255685 915 255715
rect 965 255685 995 255715
rect 1045 255685 1075 255715
rect 1125 255685 1155 255715
rect 1205 255685 1235 255715
rect 1285 255685 1315 255715
rect 1365 255685 1395 255715
rect 1445 255685 1475 255715
rect 1525 255685 1555 255715
rect 1605 255685 1635 255715
rect 1685 255685 1715 255715
rect 1765 255685 1795 255715
rect 1845 255685 1875 255715
rect 1925 255685 1955 255715
rect 2005 255685 2035 255715
rect 2085 255685 2115 255715
rect 2165 255685 2195 255715
rect 2245 255685 2275 255715
rect 2325 255685 2355 255715
rect 2405 255685 2435 255715
rect 2485 255685 2515 255715
rect 2565 255685 2595 255715
rect 2645 255685 2675 255715
rect 2725 255685 2755 255715
rect 3045 255685 3075 255715
rect 3125 255685 3155 255715
rect 3205 255685 3235 255715
rect 3285 255685 3315 255715
rect 3365 255685 3395 255715
rect 3445 255685 3475 255715
rect 3525 255685 3555 255715
rect 3605 255685 3635 255715
rect 3685 255685 3715 255715
rect 3765 255685 3795 255715
rect 3845 255685 3875 255715
rect 3925 255685 3955 255715
rect 4005 255685 4035 255715
rect 4085 255685 4115 255715
rect 4165 255685 4195 255715
rect 4245 255685 4275 255715
rect 4325 255685 4355 255715
rect 4405 255685 4435 255715
rect 4485 255685 4515 255715
rect 4565 255685 4595 255715
rect 4645 255685 4675 255715
rect 4725 255685 4755 255715
rect 4805 255685 4835 255715
rect 4885 255685 4915 255715
rect 4965 255685 4995 255715
rect 5045 255685 5075 255715
rect 5125 255685 5155 255715
rect 5205 255685 5235 255715
rect 5285 255685 5315 255715
rect 5365 255685 5395 255715
rect 5445 255685 5475 255715
rect 5525 255685 5555 255715
rect 5605 255685 5635 255715
rect 5685 255685 5715 255715
rect 5765 255685 5795 255715
rect 5845 255685 5875 255715
rect 5925 255685 5955 255715
rect 6005 255685 6035 255715
rect 6085 255685 6115 255715
rect 6165 255685 6195 255715
rect 6245 255685 6275 255715
rect 6325 255685 6355 255715
rect 6405 255685 6435 255715
rect 6485 255685 6515 255715
rect 6565 255685 6595 255715
rect 6645 255685 6675 255715
rect 6725 255685 6755 255715
rect 6805 255685 6835 255715
rect 6885 255685 6915 255715
rect 6965 255685 6995 255715
rect 7045 255685 7075 255715
rect 7125 255685 7155 255715
rect 7205 255685 7235 255715
rect 7285 255685 7315 255715
rect 7365 255685 7395 255715
rect 7445 255685 7475 255715
rect 7525 255685 7555 255715
rect 7605 255685 7635 255715
rect 7685 255685 7715 255715
rect 7765 255685 7795 255715
rect 7845 255685 7875 255715
rect 7925 255685 7955 255715
rect 8005 255685 8035 255715
rect 8085 255685 8115 255715
rect 8165 255685 8195 255715
rect 8245 255685 8275 255715
rect 8325 255685 8355 255715
rect 8405 255685 8435 255715
rect 8485 255685 8515 255715
rect 8565 255685 8595 255715
rect 8645 255685 8675 255715
rect 8725 255685 8755 255715
rect 8805 255685 8835 255715
rect 8885 255685 8915 255715
rect 8965 255685 8995 255715
rect 9045 255685 9075 255715
rect 9125 255685 9155 255715
rect 9205 255685 9235 255715
rect 9285 255685 9315 255715
rect 9365 255685 9395 255715
rect 9445 255685 9475 255715
rect 9525 255685 9555 255715
rect 9605 255685 9635 255715
rect 9685 255685 9715 255715
rect 9765 255685 9795 255715
rect 9845 255685 9875 255715
rect 9925 255685 9955 255715
rect 10005 255685 10035 255715
rect 10085 255685 10115 255715
rect 10165 255685 10195 255715
rect 10245 255685 10275 255715
rect 10325 255685 10355 255715
rect 10405 255685 10435 255715
rect 10485 255685 10515 255715
rect 10565 255685 10595 255715
rect 10645 255685 10675 255715
rect 10725 255685 10755 255715
rect 10805 255685 10835 255715
rect 10885 255685 10915 255715
rect 10965 255685 10995 255715
rect 11045 255685 11075 255715
rect 11125 255685 11155 255715
rect 11205 255685 11235 255715
rect 11285 255685 11315 255715
rect 11365 255685 11395 255715
rect 11445 255685 11475 255715
rect 11525 255685 11555 255715
rect 11605 255685 11635 255715
rect 11685 255685 11715 255715
rect 11765 255685 11795 255715
rect 11845 255685 11875 255715
rect 11925 255685 11955 255715
rect 12005 255685 12035 255715
rect 12085 255685 12115 255715
rect 12165 255685 12195 255715
rect 12245 255685 12275 255715
rect 12325 255685 12355 255715
rect 12405 255685 12435 255715
rect 12485 255685 12515 255715
rect 12565 255685 12595 255715
rect 12645 255685 12675 255715
rect 12725 255685 12755 255715
rect 12805 255685 12835 255715
rect 12885 255685 12915 255715
rect 12965 255685 12995 255715
rect 13045 255685 13075 255715
rect 13125 255685 13155 255715
rect 13205 255685 13235 255715
rect 13285 255685 13315 255715
rect 13365 255685 13395 255715
rect 13445 255685 13475 255715
rect 13525 255685 13555 255715
rect 13605 255685 13635 255715
rect 13685 255685 13715 255715
rect 13765 255685 13795 255715
rect 13845 255685 13875 255715
rect 13925 255685 13955 255715
rect 14005 255685 14035 255715
rect 14085 255685 14115 255715
rect 14165 255685 14195 255715
rect 14245 255685 14275 255715
rect 14325 255685 14355 255715
rect 14405 255685 14435 255715
rect 14485 255685 14515 255715
rect 14565 255685 14595 255715
rect 14645 255685 14675 255715
rect 14725 255685 14755 255715
rect 14805 255685 14835 255715
rect 14885 255685 14915 255715
rect 14965 255685 14995 255715
rect 15045 255685 15075 255715
rect 15125 255685 15155 255715
rect 15205 255685 15235 255715
rect 15285 255685 15315 255715
rect 15365 255685 15395 255715
rect 15445 255685 15475 255715
rect 15525 255685 15555 255715
rect 15605 255685 15635 255715
rect 15685 255685 15715 255715
rect 15765 255685 15795 255715
rect 15845 255685 15875 255715
rect 15925 255685 15955 255715
rect 16005 255685 16035 255715
rect 16085 255685 16115 255715
rect 16165 255685 16195 255715
rect 16245 255685 16275 255715
rect 16325 255685 16355 255715
rect 16405 255685 16435 255715
rect 16485 255685 16515 255715
rect 16565 255685 16595 255715
rect 16645 255685 16675 255715
rect 16725 255685 16755 255715
rect 16885 255685 16915 255715
<< metal3 >>
rect 8097 351400 10597 352400
rect 8097 351200 10600 351400
rect 8097 351150 10597 351200
rect 34097 351150 36597 352400
rect 60097 351150 62597 352400
rect 82797 351150 85297 352400
rect 85447 351150 86547 352400
rect 86697 351150 87797 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 111297 351150 112397 352400
rect 112547 351150 113647 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 162147 351150 163247 352400
rect 163397 351150 164497 352400
rect 164647 351150 167147 352400
rect 206697 351150 209197 352400
rect 232697 351150 235197 352400
rect 255297 351170 257697 352400
rect 260297 351400 262697 352400
rect 271860 351816 271900 351820
rect 271860 351784 271864 351816
rect 271896 351784 271900 351816
rect 271860 351656 271900 351784
rect 272020 351816 272060 351820
rect 272020 351784 272024 351816
rect 272056 351784 272060 351816
rect 271860 351624 271864 351656
rect 271896 351624 271900 351656
rect 271860 351576 271900 351624
rect 271860 351544 271864 351576
rect 271896 351544 271900 351576
rect 271860 351496 271900 351544
rect 271860 351464 271864 351496
rect 271896 351464 271900 351496
rect 271860 351416 271900 351464
rect 260297 351200 262800 351400
rect 271860 351384 271864 351416
rect 271896 351384 271900 351416
rect 271860 351336 271900 351384
rect 271860 351304 271864 351336
rect 271896 351304 271900 351336
rect 271860 351256 271900 351304
rect 271860 351224 271864 351256
rect 271896 351224 271900 351256
rect 260297 351170 262697 351200
rect 271860 351176 271900 351224
rect 271860 351144 271864 351176
rect 271896 351144 271900 351176
rect 271860 351096 271900 351144
rect 271860 351064 271864 351096
rect 271896 351064 271900 351096
rect 271860 351016 271900 351064
rect 271860 350984 271864 351016
rect 271896 350984 271900 351016
rect 271860 350936 271900 350984
rect 271860 350904 271864 350936
rect 271896 350904 271900 350936
rect 271860 350856 271900 350904
rect 271860 350824 271864 350856
rect 271896 350824 271900 350856
rect 271860 350776 271900 350824
rect 271860 350744 271864 350776
rect 271896 350744 271900 350776
rect 271860 350696 271900 350744
rect 271860 350664 271864 350696
rect 271896 350664 271900 350696
rect 271860 350616 271900 350664
rect 271860 350584 271864 350616
rect 271896 350584 271900 350616
rect 271860 350536 271900 350584
rect 271860 350504 271864 350536
rect 271896 350504 271900 350536
rect 271860 350456 271900 350504
rect 271860 350424 271864 350456
rect 271896 350424 271900 350456
rect 258900 350200 271500 350400
rect -400 340400 850 342621
rect -400 340200 14400 340400
rect -400 340121 850 340200
rect -400 321921 830 324321
rect -400 317800 830 319321
rect -400 317790 1200 317800
rect -400 317610 1010 317790
rect 1190 317610 1200 317790
rect -400 317600 1200 317610
rect -400 316921 830 317600
rect 3200 287160 3280 287200
rect 3240 287120 3280 287160
rect -400 280600 830 282121
rect -400 280400 840 280600
rect -400 279721 830 280400
rect -400 275500 830 277121
rect 14200 275800 14400 340200
rect 16200 317790 16400 317800
rect 16200 317610 16210 317790
rect 16390 317610 16400 317790
rect 14220 275700 14300 275800
rect -400 275300 850 275500
rect -400 275200 830 275300
rect -400 275160 1200 275200
rect -400 275040 1040 275160
rect 1160 275040 1200 275160
rect -400 275000 1200 275040
rect 2400 275000 2600 275200
rect 13520 275195 13560 275200
rect 13520 275005 13525 275195
rect 13555 275005 13560 275195
rect -400 274721 830 275000
rect 13520 274880 13560 275005
rect 13680 275195 13720 275200
rect 13680 275005 13685 275195
rect 13715 275005 13720 275195
rect 13680 274920 13720 275005
rect 13840 275195 13880 275200
rect 13840 275005 13845 275195
rect 13875 275005 13880 275195
rect 13840 274920 13880 275005
rect 14000 275195 14040 275200
rect 14000 275005 14005 275195
rect 14035 275005 14040 275195
rect 14000 274920 14040 275005
rect 14160 275195 14200 275200
rect 14160 275005 14165 275195
rect 14195 275005 14200 275195
rect 14160 274920 14200 275005
rect 14240 274920 14280 275700
rect 14320 275195 14360 275200
rect 14320 275005 14325 275195
rect 14355 275005 14360 275195
rect 14320 274920 14360 275005
rect 16200 274790 16400 317610
rect 16200 274610 16210 274790
rect 16390 274610 16400 274790
rect 16200 274600 16400 274610
rect 16720 275476 16760 275480
rect 16720 275444 16724 275476
rect 16756 275444 16760 275476
rect 16720 275316 16760 275444
rect 16880 275476 16920 275480
rect 16880 275444 16884 275476
rect 16916 275444 16920 275476
rect 16720 275284 16724 275316
rect 16756 275284 16760 275316
rect 16720 274956 16760 275284
rect 16720 274924 16724 274956
rect 16756 274924 16760 274956
rect 16720 274876 16760 274924
rect 16720 274844 16724 274876
rect 16756 274844 16760 274876
rect 16720 274795 16760 274844
rect 16720 274765 16725 274795
rect 16755 274765 16760 274795
rect 16720 274715 16760 274765
rect 16720 274685 16725 274715
rect 16755 274685 16760 274715
rect 16720 274635 16760 274685
rect 16720 274605 16725 274635
rect 16755 274605 16760 274635
rect 16720 274556 16760 274605
rect 16720 274524 16724 274556
rect 16756 274524 16760 274556
rect 16720 274476 16760 274524
rect 16720 274444 16724 274476
rect 16756 274444 16760 274476
rect 16720 274396 16760 274444
rect 16720 274364 16724 274396
rect 16756 274364 16760 274396
rect 16720 274316 16760 274364
rect 16720 274284 16724 274316
rect 16756 274284 16760 274316
rect 16720 274236 16760 274284
rect 16720 274204 16724 274236
rect 16756 274204 16760 274236
rect 16720 274156 16760 274204
rect 16720 274124 16724 274156
rect 16756 274124 16760 274156
rect 16720 274076 16760 274124
rect 16720 274044 16724 274076
rect 16756 274044 16760 274076
rect 16720 273996 16760 274044
rect 16720 273964 16724 273996
rect 16756 273964 16760 273996
rect 16720 273916 16760 273964
rect 16720 273884 16724 273916
rect 16756 273884 16760 273916
rect 16720 273836 16760 273884
rect 16720 273804 16724 273836
rect 16756 273804 16760 273836
rect 16720 273756 16760 273804
rect 16720 273724 16724 273756
rect 16756 273724 16760 273756
rect 16720 273676 16760 273724
rect 16720 273644 16724 273676
rect 16756 273644 16760 273676
rect 16720 273596 16760 273644
rect 16720 273564 16724 273596
rect 16756 273564 16760 273596
rect 16720 273516 16760 273564
rect 16720 273484 16724 273516
rect 16756 273484 16760 273516
rect 16720 273436 16760 273484
rect 16720 273404 16724 273436
rect 16756 273404 16760 273436
rect 16720 273356 16760 273404
rect 16720 273324 16724 273356
rect 16756 273324 16760 273356
rect 16720 273276 16760 273324
rect 16720 273244 16724 273276
rect 16756 273244 16760 273276
rect 16720 273196 16760 273244
rect 16720 273164 16724 273196
rect 16756 273164 16760 273196
rect 16720 273116 16760 273164
rect 16720 273084 16724 273116
rect 16756 273084 16760 273116
rect 16720 273036 16760 273084
rect 16720 273004 16724 273036
rect 16756 273004 16760 273036
rect 16720 272956 16760 273004
rect 16720 272924 16724 272956
rect 16756 272924 16760 272956
rect 16720 272876 16760 272924
rect 16720 272844 16724 272876
rect 16756 272844 16760 272876
rect 16720 272796 16760 272844
rect 16720 272764 16724 272796
rect 16756 272764 16760 272796
rect 16720 272716 16760 272764
rect 16720 272684 16724 272716
rect 16756 272684 16760 272716
rect 16720 272636 16760 272684
rect 16720 272604 16724 272636
rect 16756 272604 16760 272636
rect 16720 272556 16760 272604
rect 16720 272524 16724 272556
rect 16756 272524 16760 272556
rect 16720 272476 16760 272524
rect 16720 272444 16724 272476
rect 16756 272444 16760 272476
rect 16720 272396 16760 272444
rect 16720 272364 16724 272396
rect 16756 272364 16760 272396
rect 16720 272316 16760 272364
rect 16720 272284 16724 272316
rect 16756 272284 16760 272316
rect 16720 272236 16760 272284
rect 16720 272204 16724 272236
rect 16756 272204 16760 272236
rect 16720 272156 16760 272204
rect 16720 272124 16724 272156
rect 16756 272124 16760 272156
rect 16720 272076 16760 272124
rect 16720 272044 16724 272076
rect 16756 272044 16760 272076
rect 16720 271996 16760 272044
rect 16720 271964 16724 271996
rect 16756 271964 16760 271996
rect 16720 271916 16760 271964
rect 16720 271884 16724 271916
rect 16756 271884 16760 271916
rect 16720 271836 16760 271884
rect 16720 271804 16724 271836
rect 16756 271804 16760 271836
rect 16720 271756 16760 271804
rect 16720 271724 16724 271756
rect 16756 271724 16760 271756
rect 16720 271676 16760 271724
rect 16720 271644 16724 271676
rect 16756 271644 16760 271676
rect 16720 271596 16760 271644
rect 16720 271564 16724 271596
rect 16756 271564 16760 271596
rect 16720 271516 16760 271564
rect 16720 271484 16724 271516
rect 16756 271484 16760 271516
rect 16720 271436 16760 271484
rect 16720 271404 16724 271436
rect 16756 271404 16760 271436
rect 16720 271356 16760 271404
rect 16720 271324 16724 271356
rect 16756 271324 16760 271356
rect 16720 271276 16760 271324
rect 16720 271244 16724 271276
rect 16756 271244 16760 271276
rect 16720 271196 16760 271244
rect 16720 271164 16724 271196
rect 16756 271164 16760 271196
rect 16720 271116 16760 271164
rect 16720 271084 16724 271116
rect 16756 271084 16760 271116
rect 16720 271036 16760 271084
rect 16720 271004 16724 271036
rect 16756 271004 16760 271036
rect 16720 270956 16760 271004
rect 16720 270924 16724 270956
rect 16756 270924 16760 270956
rect 16720 270876 16760 270924
rect 16720 270844 16724 270876
rect 16756 270844 16760 270876
rect 16720 270796 16760 270844
rect 16720 270764 16724 270796
rect 16756 270764 16760 270796
rect 16720 270716 16760 270764
rect 16720 270684 16724 270716
rect 16756 270684 16760 270716
rect 16720 270636 16760 270684
rect 16720 270604 16724 270636
rect 16756 270604 16760 270636
rect 16720 270556 16760 270604
rect 16720 270524 16724 270556
rect 16756 270524 16760 270556
rect 16720 270476 16760 270524
rect 16720 270444 16724 270476
rect 16756 270444 16760 270476
rect 16720 270396 16760 270444
rect 16720 270364 16724 270396
rect 16756 270364 16760 270396
rect 16720 270316 16760 270364
rect 16720 270284 16724 270316
rect 16756 270284 16760 270316
rect 16720 270236 16760 270284
rect 16720 270204 16724 270236
rect 16756 270204 16760 270236
rect 16720 270156 16760 270204
rect 16720 270124 16724 270156
rect 16756 270124 16760 270156
rect 16720 270076 16760 270124
rect 16720 270044 16724 270076
rect 16756 270044 16760 270076
rect 16720 269996 16760 270044
rect 16720 269964 16724 269996
rect 16756 269964 16760 269996
rect 16720 269916 16760 269964
rect 16720 269884 16724 269916
rect 16756 269884 16760 269916
rect 16720 269836 16760 269884
rect 16720 269804 16724 269836
rect 16756 269804 16760 269836
rect 16720 269756 16760 269804
rect 16720 269724 16724 269756
rect 16756 269724 16760 269756
rect 16720 269676 16760 269724
rect 16720 269644 16724 269676
rect 16756 269644 16760 269676
rect 16720 269596 16760 269644
rect 16720 269564 16724 269596
rect 16756 269564 16760 269596
rect 16720 269516 16760 269564
rect 16720 269484 16724 269516
rect 16756 269484 16760 269516
rect 16720 269436 16760 269484
rect 16720 269404 16724 269436
rect 16756 269404 16760 269436
rect 16720 269356 16760 269404
rect 16720 269324 16724 269356
rect 16756 269324 16760 269356
rect 16720 269276 16760 269324
rect 16720 269244 16724 269276
rect 16756 269244 16760 269276
rect 16720 269196 16760 269244
rect 16720 269164 16724 269196
rect 16756 269164 16760 269196
rect 16720 269116 16760 269164
rect 16720 269084 16724 269116
rect 16756 269084 16760 269116
rect 16720 269036 16760 269084
rect 16720 269004 16724 269036
rect 16756 269004 16760 269036
rect 16720 268956 16760 269004
rect 16720 268924 16724 268956
rect 16756 268924 16760 268956
rect 16720 268876 16760 268924
rect 16720 268844 16724 268876
rect 16756 268844 16760 268876
rect 16720 268796 16760 268844
rect 16720 268764 16724 268796
rect 16756 268764 16760 268796
rect 16720 268716 16760 268764
rect 16720 268684 16724 268716
rect 16756 268684 16760 268716
rect 16720 268636 16760 268684
rect 16720 268604 16724 268636
rect 16756 268604 16760 268636
rect 16720 268556 16760 268604
rect 16720 268524 16724 268556
rect 16756 268524 16760 268556
rect 16720 268476 16760 268524
rect 16720 268444 16724 268476
rect 16756 268444 16760 268476
rect 16720 268396 16760 268444
rect 16720 268364 16724 268396
rect 16756 268364 16760 268396
rect 16720 268316 16760 268364
rect 16720 268284 16724 268316
rect 16756 268284 16760 268316
rect 16720 268236 16760 268284
rect 16720 268204 16724 268236
rect 16756 268204 16760 268236
rect 16720 268156 16760 268204
rect 16720 268124 16724 268156
rect 16756 268124 16760 268156
rect 16720 268076 16760 268124
rect 16720 268044 16724 268076
rect 16756 268044 16760 268076
rect 16720 267996 16760 268044
rect 16720 267964 16724 267996
rect 16756 267964 16760 267996
rect 16720 267916 16760 267964
rect 16720 267884 16724 267916
rect 16756 267884 16760 267916
rect 16720 267836 16760 267884
rect 16720 267804 16724 267836
rect 16756 267804 16760 267836
rect 16720 267756 16760 267804
rect 16720 267724 16724 267756
rect 16756 267724 16760 267756
rect 16720 267676 16760 267724
rect 16720 267644 16724 267676
rect 16756 267644 16760 267676
rect 16720 267596 16760 267644
rect 16720 267564 16724 267596
rect 16756 267564 16760 267596
rect 16720 267516 16760 267564
rect 16720 267484 16724 267516
rect 16756 267484 16760 267516
rect 16720 267436 16760 267484
rect 16720 267404 16724 267436
rect 16756 267404 16760 267436
rect 16720 267356 16760 267404
rect 16720 267324 16724 267356
rect 16756 267324 16760 267356
rect 16720 267276 16760 267324
rect 16720 267244 16724 267276
rect 16756 267244 16760 267276
rect 16720 267196 16760 267244
rect 16720 267164 16724 267196
rect 16756 267164 16760 267196
rect 16720 267116 16760 267164
rect 16720 267084 16724 267116
rect 16756 267084 16760 267116
rect 16720 267036 16760 267084
rect 16720 267004 16724 267036
rect 16756 267004 16760 267036
rect 16720 266956 16760 267004
rect 16720 266924 16724 266956
rect 16756 266924 16760 266956
rect 16720 266876 16760 266924
rect 16720 266844 16724 266876
rect 16756 266844 16760 266876
rect 16720 266796 16760 266844
rect 16720 266764 16724 266796
rect 16756 266764 16760 266796
rect 16720 266716 16760 266764
rect 16720 266684 16724 266716
rect 16756 266684 16760 266716
rect 16720 266636 16760 266684
rect 16720 266604 16724 266636
rect 16756 266604 16760 266636
rect 16720 266556 16760 266604
rect 16720 266524 16724 266556
rect 16756 266524 16760 266556
rect 16720 266476 16760 266524
rect 16720 266444 16724 266476
rect 16756 266444 16760 266476
rect 16720 266396 16760 266444
rect 16720 266364 16724 266396
rect 16756 266364 16760 266396
rect 16720 266316 16760 266364
rect 16720 266284 16724 266316
rect 16756 266284 16760 266316
rect 16720 266236 16760 266284
rect 16720 266204 16724 266236
rect 16756 266204 16760 266236
rect 16720 266156 16760 266204
rect 16720 266124 16724 266156
rect 16756 266124 16760 266156
rect 16720 266076 16760 266124
rect 16720 266044 16724 266076
rect 16756 266044 16760 266076
rect 16720 265996 16760 266044
rect 16720 265964 16724 265996
rect 16756 265964 16760 265996
rect 16720 265916 16760 265964
rect 16720 265884 16724 265916
rect 16756 265884 16760 265916
rect 16720 265836 16760 265884
rect 16720 265804 16724 265836
rect 16756 265804 16760 265836
rect 16720 265756 16760 265804
rect 16720 265724 16724 265756
rect 16756 265724 16760 265756
rect 16720 265676 16760 265724
rect 16720 265644 16724 265676
rect 16756 265644 16760 265676
rect 16720 265596 16760 265644
rect 16720 265564 16724 265596
rect 16756 265564 16760 265596
rect 16720 265516 16760 265564
rect 16720 265484 16724 265516
rect 16756 265484 16760 265516
rect 16720 265436 16760 265484
rect 16720 265404 16724 265436
rect 16756 265404 16760 265436
rect 16720 265356 16760 265404
rect 16720 265324 16724 265356
rect 16756 265324 16760 265356
rect 16720 265276 16760 265324
rect 16720 265244 16724 265276
rect 16756 265244 16760 265276
rect 16720 265196 16760 265244
rect 16720 265164 16724 265196
rect 16756 265164 16760 265196
rect 16720 265116 16760 265164
rect 16720 265084 16724 265116
rect 16756 265084 16760 265116
rect 16720 265036 16760 265084
rect 16720 265004 16724 265036
rect 16756 265004 16760 265036
rect 16720 264956 16760 265004
rect 16720 264924 16724 264956
rect 16756 264924 16760 264956
rect 16720 264876 16760 264924
rect 16720 264844 16724 264876
rect 16756 264844 16760 264876
rect 16720 264796 16760 264844
rect 16720 264764 16724 264796
rect 16756 264764 16760 264796
rect 16720 264716 16760 264764
rect 16720 264684 16724 264716
rect 16756 264684 16760 264716
rect 16720 264636 16760 264684
rect 16720 264604 16724 264636
rect 16756 264604 16760 264636
rect 16720 264556 16760 264604
rect 16720 264524 16724 264556
rect 16756 264524 16760 264556
rect 16720 264476 16760 264524
rect 16720 264444 16724 264476
rect 16756 264444 16760 264476
rect 16720 264396 16760 264444
rect 16720 264364 16724 264396
rect 16756 264364 16760 264396
rect 16720 264316 16760 264364
rect 16720 264284 16724 264316
rect 16756 264284 16760 264316
rect 16720 264236 16760 264284
rect 16720 264204 16724 264236
rect 16756 264204 16760 264236
rect 16720 264156 16760 264204
rect 16720 264124 16724 264156
rect 16756 264124 16760 264156
rect 16720 264076 16760 264124
rect 16720 264044 16724 264076
rect 16756 264044 16760 264076
rect 16720 263996 16760 264044
rect 16720 263964 16724 263996
rect 16756 263964 16760 263996
rect 16720 263916 16760 263964
rect 16720 263884 16724 263916
rect 16756 263884 16760 263916
rect 16720 263836 16760 263884
rect 16720 263804 16724 263836
rect 16756 263804 16760 263836
rect 16720 263756 16760 263804
rect 16720 263724 16724 263756
rect 16756 263724 16760 263756
rect 16720 263676 16760 263724
rect 16720 263644 16724 263676
rect 16756 263644 16760 263676
rect 16720 263596 16760 263644
rect 16720 263564 16724 263596
rect 16756 263564 16760 263596
rect 16720 263516 16760 263564
rect 16720 263484 16724 263516
rect 16756 263484 16760 263516
rect 16720 263436 16760 263484
rect 16720 263404 16724 263436
rect 16756 263404 16760 263436
rect 2800 263360 2840 263400
rect 2960 263360 3000 263400
rect 3120 263360 3160 263400
rect 3280 263360 3320 263400
rect 3440 263360 3480 263400
rect 2800 263320 3480 263360
rect 16720 263356 16760 263404
rect 16720 263324 16724 263356
rect 16756 263324 16760 263356
rect 400 255876 440 255880
rect 400 255844 404 255876
rect 436 255844 440 255876
rect 200 255821 320 255840
rect -400 255800 320 255821
rect -400 255795 360 255800
rect -400 255765 325 255795
rect 355 255765 360 255795
rect 200 255760 360 255765
rect 400 255796 440 255844
rect 400 255764 404 255796
rect 436 255764 440 255796
rect 200 255720 320 255760
rect 400 255716 440 255764
rect 400 255684 404 255716
rect 436 255684 440 255716
rect 400 255680 440 255684
rect 480 255876 520 255880
rect 480 255844 484 255876
rect 516 255844 520 255876
rect 480 255796 520 255844
rect 480 255764 484 255796
rect 516 255764 520 255796
rect 480 255716 520 255764
rect 480 255684 484 255716
rect 516 255684 520 255716
rect 480 255680 520 255684
rect 560 255876 600 255880
rect 560 255844 564 255876
rect 596 255844 600 255876
rect 560 255796 600 255844
rect 560 255764 564 255796
rect 596 255764 600 255796
rect 560 255716 600 255764
rect 560 255684 564 255716
rect 596 255684 600 255716
rect 560 255680 600 255684
rect 640 255876 680 255880
rect 640 255844 644 255876
rect 676 255844 680 255876
rect 640 255796 680 255844
rect 640 255764 644 255796
rect 676 255764 680 255796
rect 640 255716 680 255764
rect 640 255684 644 255716
rect 676 255684 680 255716
rect 640 255680 680 255684
rect 720 255876 760 255880
rect 720 255844 724 255876
rect 756 255844 760 255876
rect 720 255796 760 255844
rect 720 255764 724 255796
rect 756 255764 760 255796
rect 720 255716 760 255764
rect 720 255684 724 255716
rect 756 255684 760 255716
rect 720 255680 760 255684
rect 800 255876 840 255880
rect 800 255844 804 255876
rect 836 255844 840 255876
rect 800 255796 840 255844
rect 800 255764 804 255796
rect 836 255764 840 255796
rect 800 255716 840 255764
rect 800 255684 804 255716
rect 836 255684 840 255716
rect 800 255680 840 255684
rect 880 255876 920 255880
rect 880 255844 884 255876
rect 916 255844 920 255876
rect 880 255796 920 255844
rect 880 255764 884 255796
rect 916 255764 920 255796
rect 880 255716 920 255764
rect 880 255684 884 255716
rect 916 255684 920 255716
rect 880 255680 920 255684
rect 960 255876 1000 255880
rect 960 255844 964 255876
rect 996 255844 1000 255876
rect 960 255796 1000 255844
rect 960 255764 964 255796
rect 996 255764 1000 255796
rect 960 255716 1000 255764
rect 960 255684 964 255716
rect 996 255684 1000 255716
rect 960 255680 1000 255684
rect 1040 255876 1080 255880
rect 1040 255844 1044 255876
rect 1076 255844 1080 255876
rect 1040 255796 1080 255844
rect 1040 255764 1044 255796
rect 1076 255764 1080 255796
rect 1040 255716 1080 255764
rect 1040 255684 1044 255716
rect 1076 255684 1080 255716
rect 1040 255680 1080 255684
rect 1120 255876 1160 255880
rect 1120 255844 1124 255876
rect 1156 255844 1160 255876
rect 1120 255796 1160 255844
rect 1120 255764 1124 255796
rect 1156 255764 1160 255796
rect 1120 255716 1160 255764
rect 1120 255684 1124 255716
rect 1156 255684 1160 255716
rect 1120 255680 1160 255684
rect 1200 255876 1240 255880
rect 1200 255844 1204 255876
rect 1236 255844 1240 255876
rect 1200 255796 1240 255844
rect 1200 255764 1204 255796
rect 1236 255764 1240 255796
rect 1200 255716 1240 255764
rect 1200 255684 1204 255716
rect 1236 255684 1240 255716
rect 1200 255680 1240 255684
rect 1280 255876 1320 255880
rect 1280 255844 1284 255876
rect 1316 255844 1320 255876
rect 1280 255796 1320 255844
rect 1280 255764 1284 255796
rect 1316 255764 1320 255796
rect 1280 255716 1320 255764
rect 1280 255684 1284 255716
rect 1316 255684 1320 255716
rect 1280 255680 1320 255684
rect 1360 255876 1400 255880
rect 1360 255844 1364 255876
rect 1396 255844 1400 255876
rect 1360 255796 1400 255844
rect 1360 255764 1364 255796
rect 1396 255764 1400 255796
rect 1360 255716 1400 255764
rect 1360 255684 1364 255716
rect 1396 255684 1400 255716
rect 1360 255680 1400 255684
rect 1440 255876 1480 255880
rect 1440 255844 1444 255876
rect 1476 255844 1480 255876
rect 1440 255796 1480 255844
rect 1440 255764 1444 255796
rect 1476 255764 1480 255796
rect 1440 255716 1480 255764
rect 1440 255684 1444 255716
rect 1476 255684 1480 255716
rect 1440 255680 1480 255684
rect 1520 255876 1560 255880
rect 1520 255844 1524 255876
rect 1556 255844 1560 255876
rect 1520 255796 1560 255844
rect 1520 255764 1524 255796
rect 1556 255764 1560 255796
rect 1520 255716 1560 255764
rect 1520 255684 1524 255716
rect 1556 255684 1560 255716
rect 1520 255680 1560 255684
rect 1600 255876 1640 255880
rect 1600 255844 1604 255876
rect 1636 255844 1640 255876
rect 1600 255796 1640 255844
rect 1600 255764 1604 255796
rect 1636 255764 1640 255796
rect 1600 255716 1640 255764
rect 1600 255684 1604 255716
rect 1636 255684 1640 255716
rect 1600 255680 1640 255684
rect 1680 255876 1720 255880
rect 1680 255844 1684 255876
rect 1716 255844 1720 255876
rect 1680 255796 1720 255844
rect 1680 255764 1684 255796
rect 1716 255764 1720 255796
rect 1680 255716 1720 255764
rect 1680 255684 1684 255716
rect 1716 255684 1720 255716
rect 1680 255680 1720 255684
rect 1760 255876 1800 255880
rect 1760 255844 1764 255876
rect 1796 255844 1800 255876
rect 1760 255796 1800 255844
rect 1760 255764 1764 255796
rect 1796 255764 1800 255796
rect 1760 255716 1800 255764
rect 1760 255684 1764 255716
rect 1796 255684 1800 255716
rect 1760 255680 1800 255684
rect 1840 255876 1880 255880
rect 1840 255844 1844 255876
rect 1876 255844 1880 255876
rect 1840 255796 1880 255844
rect 1840 255764 1844 255796
rect 1876 255764 1880 255796
rect 1840 255716 1880 255764
rect 1840 255684 1844 255716
rect 1876 255684 1880 255716
rect 1840 255680 1880 255684
rect 1920 255876 1960 255880
rect 1920 255844 1924 255876
rect 1956 255844 1960 255876
rect 1920 255796 1960 255844
rect 1920 255764 1924 255796
rect 1956 255764 1960 255796
rect 1920 255716 1960 255764
rect 1920 255684 1924 255716
rect 1956 255684 1960 255716
rect 1920 255680 1960 255684
rect 2000 255876 2040 255880
rect 2000 255844 2004 255876
rect 2036 255844 2040 255876
rect 2000 255796 2040 255844
rect 2000 255764 2004 255796
rect 2036 255764 2040 255796
rect 2000 255716 2040 255764
rect 2000 255684 2004 255716
rect 2036 255684 2040 255716
rect 2000 255680 2040 255684
rect 2080 255876 2120 255880
rect 2080 255844 2084 255876
rect 2116 255844 2120 255876
rect 2080 255796 2120 255844
rect 2080 255764 2084 255796
rect 2116 255764 2120 255796
rect 2080 255716 2120 255764
rect 2080 255684 2084 255716
rect 2116 255684 2120 255716
rect 2080 255680 2120 255684
rect 2160 255876 2200 255880
rect 2160 255844 2164 255876
rect 2196 255844 2200 255876
rect 2160 255796 2200 255844
rect 2160 255764 2164 255796
rect 2196 255764 2200 255796
rect 2160 255716 2200 255764
rect 2160 255684 2164 255716
rect 2196 255684 2200 255716
rect 2160 255680 2200 255684
rect 2240 255876 2280 255880
rect 2240 255844 2244 255876
rect 2276 255844 2280 255876
rect 2240 255796 2280 255844
rect 2240 255764 2244 255796
rect 2276 255764 2280 255796
rect 2240 255716 2280 255764
rect 2240 255684 2244 255716
rect 2276 255684 2280 255716
rect 2240 255680 2280 255684
rect 2320 255876 2360 255880
rect 2320 255844 2324 255876
rect 2356 255844 2360 255876
rect 2320 255796 2360 255844
rect 2320 255764 2324 255796
rect 2356 255764 2360 255796
rect 2320 255716 2360 255764
rect 2320 255684 2324 255716
rect 2356 255684 2360 255716
rect 2320 255680 2360 255684
rect 2400 255876 2440 255880
rect 2400 255844 2404 255876
rect 2436 255844 2440 255876
rect 2400 255796 2440 255844
rect 2400 255764 2404 255796
rect 2436 255764 2440 255796
rect 2400 255716 2440 255764
rect 2400 255684 2404 255716
rect 2436 255684 2440 255716
rect 2400 255680 2440 255684
rect 2480 255876 2520 255880
rect 2480 255844 2484 255876
rect 2516 255844 2520 255876
rect 2480 255796 2520 255844
rect 2480 255764 2484 255796
rect 2516 255764 2520 255796
rect 2480 255716 2520 255764
rect 2480 255684 2484 255716
rect 2516 255684 2520 255716
rect 2480 255680 2520 255684
rect 2560 255876 2600 255880
rect 2560 255844 2564 255876
rect 2596 255844 2600 255876
rect 2560 255796 2600 255844
rect 2560 255764 2564 255796
rect 2596 255764 2600 255796
rect 2560 255716 2600 255764
rect 2560 255684 2564 255716
rect 2596 255684 2600 255716
rect 2560 255680 2600 255684
rect 2640 255876 2680 255880
rect 2640 255844 2644 255876
rect 2676 255844 2680 255876
rect 2640 255796 2680 255844
rect 2640 255764 2644 255796
rect 2676 255764 2680 255796
rect 2640 255716 2680 255764
rect 2640 255684 2644 255716
rect 2676 255684 2680 255716
rect 2640 255680 2680 255684
rect 2720 255876 2760 255880
rect 2720 255844 2724 255876
rect 2756 255844 2760 255876
rect 2720 255796 2760 255844
rect 2720 255764 2724 255796
rect 2756 255764 2760 255796
rect 2720 255716 2760 255764
rect 2720 255684 2724 255716
rect 2756 255684 2760 255716
rect 2720 255680 2760 255684
rect -400 255174 240 255230
rect -400 254583 240 254639
rect -400 253992 240 254048
rect -400 253401 240 253457
rect -400 252810 240 252866
rect -400 234154 240 234210
rect -400 233563 240 233619
rect -400 232972 240 233028
rect -400 232381 240 232437
rect -400 231790 240 231846
rect -400 231199 240 231255
rect -400 212543 240 212599
rect -400 211952 240 212008
rect -400 211361 240 211417
rect -400 210770 240 210826
rect -400 210179 240 210235
rect -400 209588 240 209644
rect -400 190932 240 190988
rect -400 190341 240 190397
rect -400 189750 240 189806
rect -400 189159 240 189215
rect -400 188568 240 188624
rect -400 187977 240 188033
rect -400 169321 240 169377
rect -400 168730 240 168786
rect -400 168139 240 168195
rect -400 167548 240 167604
rect -400 166957 240 167013
rect -400 166366 240 166422
rect -400 147710 240 147766
rect -400 147119 240 147175
rect -400 146528 240 146584
rect -400 145937 240 145993
rect -400 145346 240 145402
rect -400 144755 240 144811
rect -400 126199 240 126255
rect -400 125608 240 125664
rect -400 125017 240 125073
rect -400 124426 240 124482
rect -400 123835 240 123891
rect -400 123244 240 123300
rect -400 109800 830 109844
rect 2800 109800 3000 263320
rect 16720 263276 16760 263324
rect 16720 263244 16724 263276
rect 16756 263244 16760 263276
rect 16720 263196 16760 263244
rect 16720 263164 16724 263196
rect 16756 263164 16760 263196
rect 16720 263116 16760 263164
rect 16720 263084 16724 263116
rect 16756 263084 16760 263116
rect 16720 263036 16760 263084
rect 16720 263004 16724 263036
rect 16756 263004 16760 263036
rect 16720 262956 16760 263004
rect 16720 262924 16724 262956
rect 16756 262924 16760 262956
rect 16720 262876 16760 262924
rect 16720 262844 16724 262876
rect 16756 262844 16760 262876
rect 16720 262796 16760 262844
rect 16720 262764 16724 262796
rect 16756 262764 16760 262796
rect 16720 262716 16760 262764
rect 16720 262684 16724 262716
rect 16756 262684 16760 262716
rect 16720 262636 16760 262684
rect 16720 262604 16724 262636
rect 16756 262604 16760 262636
rect 16720 262556 16760 262604
rect 16720 262524 16724 262556
rect 16756 262524 16760 262556
rect 16720 262476 16760 262524
rect 16720 262444 16724 262476
rect 16756 262444 16760 262476
rect 16720 262396 16760 262444
rect 16720 262364 16724 262396
rect 16756 262364 16760 262396
rect 16720 262316 16760 262364
rect 16720 262284 16724 262316
rect 16756 262284 16760 262316
rect 16720 262236 16760 262284
rect 16720 262204 16724 262236
rect 16756 262204 16760 262236
rect 16720 262156 16760 262204
rect 16720 262124 16724 262156
rect 16756 262124 16760 262156
rect 16720 262076 16760 262124
rect 16720 262044 16724 262076
rect 16756 262044 16760 262076
rect 16720 261996 16760 262044
rect 16720 261964 16724 261996
rect 16756 261964 16760 261996
rect 16720 261916 16760 261964
rect 16720 261884 16724 261916
rect 16756 261884 16760 261916
rect 16720 261836 16760 261884
rect 16720 261804 16724 261836
rect 16756 261804 16760 261836
rect 16720 261756 16760 261804
rect 16720 261724 16724 261756
rect 16756 261724 16760 261756
rect 16720 261676 16760 261724
rect 16720 261644 16724 261676
rect 16756 261644 16760 261676
rect 16720 261596 16760 261644
rect 16720 261564 16724 261596
rect 16756 261564 16760 261596
rect 16720 261516 16760 261564
rect 16720 261484 16724 261516
rect 16756 261484 16760 261516
rect 16720 261436 16760 261484
rect 16720 261404 16724 261436
rect 16756 261404 16760 261436
rect 16720 261356 16760 261404
rect 16720 261324 16724 261356
rect 16756 261324 16760 261356
rect 16720 261276 16760 261324
rect 16720 261244 16724 261276
rect 16756 261244 16760 261276
rect 16720 261196 16760 261244
rect 16720 261164 16724 261196
rect 16756 261164 16760 261196
rect 16720 261116 16760 261164
rect 16720 261084 16724 261116
rect 16756 261084 16760 261116
rect 16720 261036 16760 261084
rect 16720 261004 16724 261036
rect 16756 261004 16760 261036
rect 16720 260956 16760 261004
rect 16720 260924 16724 260956
rect 16756 260924 16760 260956
rect 16720 260876 16760 260924
rect 16720 260844 16724 260876
rect 16756 260844 16760 260876
rect 16720 260796 16760 260844
rect 16720 260764 16724 260796
rect 16756 260764 16760 260796
rect 16720 260716 16760 260764
rect 16720 260684 16724 260716
rect 16756 260684 16760 260716
rect 16720 260636 16760 260684
rect 16720 260604 16724 260636
rect 16756 260604 16760 260636
rect 16720 260556 16760 260604
rect 16720 260524 16724 260556
rect 16756 260524 16760 260556
rect 16720 260476 16760 260524
rect 16720 260444 16724 260476
rect 16756 260444 16760 260476
rect 16720 260396 16760 260444
rect 16720 260364 16724 260396
rect 16756 260364 16760 260396
rect 16720 260316 16760 260364
rect 16720 260284 16724 260316
rect 16756 260284 16760 260316
rect 16720 260236 16760 260284
rect 16720 260204 16724 260236
rect 16756 260204 16760 260236
rect 16720 260156 16760 260204
rect 16720 260124 16724 260156
rect 16756 260124 16760 260156
rect 16720 260076 16760 260124
rect 16720 260044 16724 260076
rect 16756 260044 16760 260076
rect 16720 259996 16760 260044
rect 16720 259964 16724 259996
rect 16756 259964 16760 259996
rect 16720 259916 16760 259964
rect 16720 259884 16724 259916
rect 16756 259884 16760 259916
rect 16720 259836 16760 259884
rect 16720 259804 16724 259836
rect 16756 259804 16760 259836
rect 16720 259756 16760 259804
rect 16720 259724 16724 259756
rect 16756 259724 16760 259756
rect 16720 259676 16760 259724
rect 16720 259644 16724 259676
rect 16756 259644 16760 259676
rect 16720 259596 16760 259644
rect 16720 259564 16724 259596
rect 16756 259564 16760 259596
rect 16720 259516 16760 259564
rect 16720 259484 16724 259516
rect 16756 259484 16760 259516
rect 16720 259436 16760 259484
rect 16720 259404 16724 259436
rect 16756 259404 16760 259436
rect 16720 259356 16760 259404
rect 16720 259324 16724 259356
rect 16756 259324 16760 259356
rect 16720 259276 16760 259324
rect 16720 259244 16724 259276
rect 16756 259244 16760 259276
rect 16720 259196 16760 259244
rect 16720 259164 16724 259196
rect 16756 259164 16760 259196
rect 16720 259116 16760 259164
rect 16720 259084 16724 259116
rect 16756 259084 16760 259116
rect 16720 259036 16760 259084
rect 16720 259004 16724 259036
rect 16756 259004 16760 259036
rect 16720 258956 16760 259004
rect 16720 258924 16724 258956
rect 16756 258924 16760 258956
rect 16720 258876 16760 258924
rect 16720 258844 16724 258876
rect 16756 258844 16760 258876
rect 16720 258796 16760 258844
rect 16720 258764 16724 258796
rect 16756 258764 16760 258796
rect 16720 258716 16760 258764
rect 16720 258684 16724 258716
rect 16756 258684 16760 258716
rect 16720 258636 16760 258684
rect 16720 258604 16724 258636
rect 16756 258604 16760 258636
rect 16720 258556 16760 258604
rect 16720 258524 16724 258556
rect 16756 258524 16760 258556
rect 16720 258476 16760 258524
rect 16720 258444 16724 258476
rect 16756 258444 16760 258476
rect 16720 258396 16760 258444
rect 16720 258364 16724 258396
rect 16756 258364 16760 258396
rect 16720 258316 16760 258364
rect 16720 258284 16724 258316
rect 16756 258284 16760 258316
rect 16720 258236 16760 258284
rect 16720 258204 16724 258236
rect 16756 258204 16760 258236
rect 16720 258156 16760 258204
rect 16720 258124 16724 258156
rect 16756 258124 16760 258156
rect 16720 258076 16760 258124
rect 16720 258044 16724 258076
rect 16756 258044 16760 258076
rect 16720 257996 16760 258044
rect 16720 257964 16724 257996
rect 16756 257964 16760 257996
rect 16720 257916 16760 257964
rect 16720 257884 16724 257916
rect 16756 257884 16760 257916
rect 16720 257836 16760 257884
rect 16720 257804 16724 257836
rect 16756 257804 16760 257836
rect 16720 257756 16760 257804
rect 16720 257724 16724 257756
rect 16756 257724 16760 257756
rect 16720 257676 16760 257724
rect 16720 257644 16724 257676
rect 16756 257644 16760 257676
rect 16720 257596 16760 257644
rect 16720 257564 16724 257596
rect 16756 257564 16760 257596
rect 16720 257516 16760 257564
rect 16720 257484 16724 257516
rect 16756 257484 16760 257516
rect 16720 257436 16760 257484
rect 16720 257404 16724 257436
rect 16756 257404 16760 257436
rect 16720 257356 16760 257404
rect 16720 257324 16724 257356
rect 16756 257324 16760 257356
rect 16720 257276 16760 257324
rect 16720 257244 16724 257276
rect 16756 257244 16760 257276
rect 16720 257196 16760 257244
rect 16720 257164 16724 257196
rect 16756 257164 16760 257196
rect 16720 257116 16760 257164
rect 16720 257084 16724 257116
rect 16756 257084 16760 257116
rect 16720 257036 16760 257084
rect 16720 257004 16724 257036
rect 16756 257004 16760 257036
rect 16720 256956 16760 257004
rect 16720 256924 16724 256956
rect 16756 256924 16760 256956
rect 16720 256876 16760 256924
rect 16720 256844 16724 256876
rect 16756 256844 16760 256876
rect 16720 256796 16760 256844
rect 16720 256764 16724 256796
rect 16756 256764 16760 256796
rect 16720 256716 16760 256764
rect 16720 256684 16724 256716
rect 16756 256684 16760 256716
rect 16720 256636 16760 256684
rect 16720 256604 16724 256636
rect 16756 256604 16760 256636
rect 16720 256556 16760 256604
rect 16720 256524 16724 256556
rect 16756 256524 16760 256556
rect 16720 256476 16760 256524
rect 16720 256444 16724 256476
rect 16756 256444 16760 256476
rect 16720 256396 16760 256444
rect 16720 256364 16724 256396
rect 16756 256364 16760 256396
rect 16720 256316 16760 256364
rect 16720 256284 16724 256316
rect 16756 256284 16760 256316
rect 16720 256236 16760 256284
rect 16720 256204 16724 256236
rect 16756 256204 16760 256236
rect 16720 256156 16760 256204
rect 16720 256124 16724 256156
rect 16756 256124 16760 256156
rect 16720 256076 16760 256124
rect 16720 256044 16724 256076
rect 16756 256044 16760 256076
rect 16720 255996 16760 256044
rect 16720 255964 16724 255996
rect 16756 255964 16760 255996
rect 3040 255876 3080 255880
rect 3040 255844 3044 255876
rect 3076 255844 3080 255876
rect 3040 255796 3080 255844
rect 3040 255764 3044 255796
rect 3076 255764 3080 255796
rect 3040 255716 3080 255764
rect 3040 255684 3044 255716
rect 3076 255684 3080 255716
rect 3040 255680 3080 255684
rect 3120 255876 3160 255880
rect 3120 255844 3124 255876
rect 3156 255844 3160 255876
rect 3120 255796 3160 255844
rect 3120 255764 3124 255796
rect 3156 255764 3160 255796
rect 3120 255716 3160 255764
rect 3120 255684 3124 255716
rect 3156 255684 3160 255716
rect 3120 255680 3160 255684
rect 3200 255876 3240 255880
rect 3200 255844 3204 255876
rect 3236 255844 3240 255876
rect 3200 255796 3240 255844
rect 3200 255764 3204 255796
rect 3236 255764 3240 255796
rect 3200 255716 3240 255764
rect 3200 255684 3204 255716
rect 3236 255684 3240 255716
rect 3200 255680 3240 255684
rect 3280 255876 3320 255880
rect 3280 255844 3284 255876
rect 3316 255844 3320 255876
rect 3280 255796 3320 255844
rect 3280 255764 3284 255796
rect 3316 255764 3320 255796
rect 3280 255716 3320 255764
rect 3280 255684 3284 255716
rect 3316 255684 3320 255716
rect 3280 255680 3320 255684
rect 3360 255876 3400 255880
rect 3360 255844 3364 255876
rect 3396 255844 3400 255876
rect 3360 255796 3400 255844
rect 3360 255764 3364 255796
rect 3396 255764 3400 255796
rect 3360 255716 3400 255764
rect 3360 255684 3364 255716
rect 3396 255684 3400 255716
rect 3360 255680 3400 255684
rect 3440 255876 3480 255880
rect 3440 255844 3444 255876
rect 3476 255844 3480 255876
rect 3440 255796 3480 255844
rect 3440 255764 3444 255796
rect 3476 255764 3480 255796
rect 3440 255716 3480 255764
rect 3440 255684 3444 255716
rect 3476 255684 3480 255716
rect 3440 255680 3480 255684
rect 3520 255876 3560 255880
rect 3520 255844 3524 255876
rect 3556 255844 3560 255876
rect 3520 255796 3560 255844
rect 3520 255764 3524 255796
rect 3556 255764 3560 255796
rect 3520 255716 3560 255764
rect 3520 255684 3524 255716
rect 3556 255684 3560 255716
rect 3520 255680 3560 255684
rect 3600 255876 3640 255880
rect 3600 255844 3604 255876
rect 3636 255844 3640 255876
rect 3600 255796 3640 255844
rect 3600 255764 3604 255796
rect 3636 255764 3640 255796
rect 3600 255716 3640 255764
rect 3600 255684 3604 255716
rect 3636 255684 3640 255716
rect 3600 255680 3640 255684
rect 3680 255876 3720 255880
rect 3680 255844 3684 255876
rect 3716 255844 3720 255876
rect 3680 255796 3720 255844
rect 3680 255764 3684 255796
rect 3716 255764 3720 255796
rect 3680 255716 3720 255764
rect 3680 255684 3684 255716
rect 3716 255684 3720 255716
rect 3680 255680 3720 255684
rect 3760 255876 3800 255880
rect 3760 255844 3764 255876
rect 3796 255844 3800 255876
rect 3760 255796 3800 255844
rect 3760 255764 3764 255796
rect 3796 255764 3800 255796
rect 3760 255716 3800 255764
rect 3760 255684 3764 255716
rect 3796 255684 3800 255716
rect 3760 255680 3800 255684
rect 3840 255876 3880 255880
rect 3840 255844 3844 255876
rect 3876 255844 3880 255876
rect 3840 255796 3880 255844
rect 3840 255764 3844 255796
rect 3876 255764 3880 255796
rect 3840 255716 3880 255764
rect 3840 255684 3844 255716
rect 3876 255684 3880 255716
rect 3840 255680 3880 255684
rect 3920 255876 3960 255880
rect 3920 255844 3924 255876
rect 3956 255844 3960 255876
rect 3920 255796 3960 255844
rect 3920 255764 3924 255796
rect 3956 255764 3960 255796
rect 3920 255716 3960 255764
rect 3920 255684 3924 255716
rect 3956 255684 3960 255716
rect 3920 255680 3960 255684
rect 4000 255876 4040 255880
rect 4000 255844 4004 255876
rect 4036 255844 4040 255876
rect 4000 255796 4040 255844
rect 4000 255764 4004 255796
rect 4036 255764 4040 255796
rect 4000 255716 4040 255764
rect 4000 255684 4004 255716
rect 4036 255684 4040 255716
rect 4000 255680 4040 255684
rect 4080 255876 4120 255880
rect 4080 255844 4084 255876
rect 4116 255844 4120 255876
rect 4080 255796 4120 255844
rect 4080 255764 4084 255796
rect 4116 255764 4120 255796
rect 4080 255716 4120 255764
rect 4080 255684 4084 255716
rect 4116 255684 4120 255716
rect 4080 255680 4120 255684
rect 4160 255876 4200 255880
rect 4160 255844 4164 255876
rect 4196 255844 4200 255876
rect 4160 255796 4200 255844
rect 4160 255764 4164 255796
rect 4196 255764 4200 255796
rect 4160 255716 4200 255764
rect 4160 255684 4164 255716
rect 4196 255684 4200 255716
rect 4160 255680 4200 255684
rect 4240 255876 4280 255880
rect 4240 255844 4244 255876
rect 4276 255844 4280 255876
rect 4240 255796 4280 255844
rect 4240 255764 4244 255796
rect 4276 255764 4280 255796
rect 4240 255716 4280 255764
rect 4240 255684 4244 255716
rect 4276 255684 4280 255716
rect 4240 255680 4280 255684
rect 4320 255876 4360 255880
rect 4320 255844 4324 255876
rect 4356 255844 4360 255876
rect 4320 255796 4360 255844
rect 4320 255764 4324 255796
rect 4356 255764 4360 255796
rect 4320 255716 4360 255764
rect 4320 255684 4324 255716
rect 4356 255684 4360 255716
rect 4320 255680 4360 255684
rect 4400 255876 4440 255880
rect 4400 255844 4404 255876
rect 4436 255844 4440 255876
rect 4400 255796 4440 255844
rect 4400 255764 4404 255796
rect 4436 255764 4440 255796
rect 4400 255716 4440 255764
rect 4400 255684 4404 255716
rect 4436 255684 4440 255716
rect 4400 255680 4440 255684
rect 4480 255876 4520 255880
rect 4480 255844 4484 255876
rect 4516 255844 4520 255876
rect 4480 255796 4520 255844
rect 4480 255764 4484 255796
rect 4516 255764 4520 255796
rect 4480 255716 4520 255764
rect 4480 255684 4484 255716
rect 4516 255684 4520 255716
rect 4480 255680 4520 255684
rect 4560 255876 4600 255880
rect 4560 255844 4564 255876
rect 4596 255844 4600 255876
rect 4560 255796 4600 255844
rect 4560 255764 4564 255796
rect 4596 255764 4600 255796
rect 4560 255716 4600 255764
rect 4560 255684 4564 255716
rect 4596 255684 4600 255716
rect 4560 255680 4600 255684
rect 4640 255876 4680 255880
rect 4640 255844 4644 255876
rect 4676 255844 4680 255876
rect 4640 255796 4680 255844
rect 4640 255764 4644 255796
rect 4676 255764 4680 255796
rect 4640 255716 4680 255764
rect 4640 255684 4644 255716
rect 4676 255684 4680 255716
rect 4640 255680 4680 255684
rect 4720 255876 4760 255880
rect 4720 255844 4724 255876
rect 4756 255844 4760 255876
rect 4720 255796 4760 255844
rect 4720 255764 4724 255796
rect 4756 255764 4760 255796
rect 4720 255716 4760 255764
rect 4720 255684 4724 255716
rect 4756 255684 4760 255716
rect 4720 255680 4760 255684
rect 4800 255876 4840 255880
rect 4800 255844 4804 255876
rect 4836 255844 4840 255876
rect 4800 255796 4840 255844
rect 4800 255764 4804 255796
rect 4836 255764 4840 255796
rect 4800 255716 4840 255764
rect 4800 255684 4804 255716
rect 4836 255684 4840 255716
rect 4800 255680 4840 255684
rect 4880 255876 4920 255880
rect 4880 255844 4884 255876
rect 4916 255844 4920 255876
rect 4880 255796 4920 255844
rect 4880 255764 4884 255796
rect 4916 255764 4920 255796
rect 4880 255716 4920 255764
rect 4880 255684 4884 255716
rect 4916 255684 4920 255716
rect 4880 255680 4920 255684
rect 4960 255876 5000 255880
rect 4960 255844 4964 255876
rect 4996 255844 5000 255876
rect 4960 255796 5000 255844
rect 4960 255764 4964 255796
rect 4996 255764 5000 255796
rect 4960 255716 5000 255764
rect 4960 255684 4964 255716
rect 4996 255684 5000 255716
rect 4960 255680 5000 255684
rect 5040 255876 5080 255880
rect 5040 255844 5044 255876
rect 5076 255844 5080 255876
rect 5040 255796 5080 255844
rect 5040 255764 5044 255796
rect 5076 255764 5080 255796
rect 5040 255716 5080 255764
rect 5040 255684 5044 255716
rect 5076 255684 5080 255716
rect 5040 255680 5080 255684
rect 5120 255876 5160 255880
rect 5120 255844 5124 255876
rect 5156 255844 5160 255876
rect 5120 255796 5160 255844
rect 5120 255764 5124 255796
rect 5156 255764 5160 255796
rect 5120 255716 5160 255764
rect 5120 255684 5124 255716
rect 5156 255684 5160 255716
rect 5120 255680 5160 255684
rect 5200 255876 5240 255880
rect 5200 255844 5204 255876
rect 5236 255844 5240 255876
rect 5200 255796 5240 255844
rect 5200 255764 5204 255796
rect 5236 255764 5240 255796
rect 5200 255716 5240 255764
rect 5200 255684 5204 255716
rect 5236 255684 5240 255716
rect 5200 255680 5240 255684
rect 5280 255876 5320 255880
rect 5280 255844 5284 255876
rect 5316 255844 5320 255876
rect 5280 255796 5320 255844
rect 5280 255764 5284 255796
rect 5316 255764 5320 255796
rect 5280 255716 5320 255764
rect 5280 255684 5284 255716
rect 5316 255684 5320 255716
rect 5280 255680 5320 255684
rect 5360 255876 5400 255880
rect 5360 255844 5364 255876
rect 5396 255844 5400 255876
rect 5360 255796 5400 255844
rect 5360 255764 5364 255796
rect 5396 255764 5400 255796
rect 5360 255716 5400 255764
rect 5360 255684 5364 255716
rect 5396 255684 5400 255716
rect 5360 255680 5400 255684
rect 5440 255876 5480 255880
rect 5440 255844 5444 255876
rect 5476 255844 5480 255876
rect 5440 255796 5480 255844
rect 5440 255764 5444 255796
rect 5476 255764 5480 255796
rect 5440 255716 5480 255764
rect 5440 255684 5444 255716
rect 5476 255684 5480 255716
rect 5440 255680 5480 255684
rect 5520 255876 5560 255880
rect 5520 255844 5524 255876
rect 5556 255844 5560 255876
rect 5520 255796 5560 255844
rect 5520 255764 5524 255796
rect 5556 255764 5560 255796
rect 5520 255716 5560 255764
rect 5520 255684 5524 255716
rect 5556 255684 5560 255716
rect 5520 255680 5560 255684
rect 5600 255876 5640 255880
rect 5600 255844 5604 255876
rect 5636 255844 5640 255876
rect 5600 255796 5640 255844
rect 5600 255764 5604 255796
rect 5636 255764 5640 255796
rect 5600 255716 5640 255764
rect 5600 255684 5604 255716
rect 5636 255684 5640 255716
rect 5600 255680 5640 255684
rect 5680 255876 5720 255880
rect 5680 255844 5684 255876
rect 5716 255844 5720 255876
rect 5680 255796 5720 255844
rect 5680 255764 5684 255796
rect 5716 255764 5720 255796
rect 5680 255716 5720 255764
rect 5680 255684 5684 255716
rect 5716 255684 5720 255716
rect 5680 255680 5720 255684
rect 5760 255876 5800 255880
rect 5760 255844 5764 255876
rect 5796 255844 5800 255876
rect 5760 255796 5800 255844
rect 5760 255764 5764 255796
rect 5796 255764 5800 255796
rect 5760 255716 5800 255764
rect 5760 255684 5764 255716
rect 5796 255684 5800 255716
rect 5760 255680 5800 255684
rect 5840 255876 5880 255880
rect 5840 255844 5844 255876
rect 5876 255844 5880 255876
rect 5840 255796 5880 255844
rect 5840 255764 5844 255796
rect 5876 255764 5880 255796
rect 5840 255716 5880 255764
rect 5840 255684 5844 255716
rect 5876 255684 5880 255716
rect 5840 255680 5880 255684
rect 5920 255876 5960 255880
rect 5920 255844 5924 255876
rect 5956 255844 5960 255876
rect 5920 255796 5960 255844
rect 5920 255764 5924 255796
rect 5956 255764 5960 255796
rect 5920 255716 5960 255764
rect 5920 255684 5924 255716
rect 5956 255684 5960 255716
rect 5920 255680 5960 255684
rect 6000 255876 6040 255880
rect 6000 255844 6004 255876
rect 6036 255844 6040 255876
rect 6000 255796 6040 255844
rect 6000 255764 6004 255796
rect 6036 255764 6040 255796
rect 6000 255716 6040 255764
rect 6000 255684 6004 255716
rect 6036 255684 6040 255716
rect 6000 255680 6040 255684
rect 6080 255876 6120 255880
rect 6080 255844 6084 255876
rect 6116 255844 6120 255876
rect 6080 255796 6120 255844
rect 6080 255764 6084 255796
rect 6116 255764 6120 255796
rect 6080 255716 6120 255764
rect 6080 255684 6084 255716
rect 6116 255684 6120 255716
rect 6080 255680 6120 255684
rect 6160 255876 6200 255880
rect 6160 255844 6164 255876
rect 6196 255844 6200 255876
rect 6160 255796 6200 255844
rect 6160 255764 6164 255796
rect 6196 255764 6200 255796
rect 6160 255716 6200 255764
rect 6160 255684 6164 255716
rect 6196 255684 6200 255716
rect 6160 255680 6200 255684
rect 6240 255876 6280 255880
rect 6240 255844 6244 255876
rect 6276 255844 6280 255876
rect 6240 255796 6280 255844
rect 6240 255764 6244 255796
rect 6276 255764 6280 255796
rect 6240 255716 6280 255764
rect 6240 255684 6244 255716
rect 6276 255684 6280 255716
rect 6240 255680 6280 255684
rect 6320 255876 6360 255880
rect 6320 255844 6324 255876
rect 6356 255844 6360 255876
rect 6320 255796 6360 255844
rect 6320 255764 6324 255796
rect 6356 255764 6360 255796
rect 6320 255716 6360 255764
rect 6320 255684 6324 255716
rect 6356 255684 6360 255716
rect 6320 255680 6360 255684
rect 6400 255876 6440 255880
rect 6400 255844 6404 255876
rect 6436 255844 6440 255876
rect 6400 255796 6440 255844
rect 6400 255764 6404 255796
rect 6436 255764 6440 255796
rect 6400 255716 6440 255764
rect 6400 255684 6404 255716
rect 6436 255684 6440 255716
rect 6400 255680 6440 255684
rect 6480 255876 6520 255880
rect 6480 255844 6484 255876
rect 6516 255844 6520 255876
rect 6480 255796 6520 255844
rect 6480 255764 6484 255796
rect 6516 255764 6520 255796
rect 6480 255716 6520 255764
rect 6480 255684 6484 255716
rect 6516 255684 6520 255716
rect 6480 255680 6520 255684
rect 6560 255876 6600 255880
rect 6560 255844 6564 255876
rect 6596 255844 6600 255876
rect 6560 255796 6600 255844
rect 6560 255764 6564 255796
rect 6596 255764 6600 255796
rect 6560 255716 6600 255764
rect 6560 255684 6564 255716
rect 6596 255684 6600 255716
rect 6560 255680 6600 255684
rect 6640 255876 6680 255880
rect 6640 255844 6644 255876
rect 6676 255844 6680 255876
rect 6640 255796 6680 255844
rect 6640 255764 6644 255796
rect 6676 255764 6680 255796
rect 6640 255716 6680 255764
rect 6640 255684 6644 255716
rect 6676 255684 6680 255716
rect 6640 255680 6680 255684
rect 6720 255876 6760 255880
rect 6720 255844 6724 255876
rect 6756 255844 6760 255876
rect 6720 255796 6760 255844
rect 6720 255764 6724 255796
rect 6756 255764 6760 255796
rect 6720 255716 6760 255764
rect 6720 255684 6724 255716
rect 6756 255684 6760 255716
rect 6720 255680 6760 255684
rect 6800 255876 6840 255880
rect 6800 255844 6804 255876
rect 6836 255844 6840 255876
rect 6800 255796 6840 255844
rect 6800 255764 6804 255796
rect 6836 255764 6840 255796
rect 6800 255716 6840 255764
rect 6800 255684 6804 255716
rect 6836 255684 6840 255716
rect 6800 255680 6840 255684
rect 6880 255876 6920 255880
rect 6880 255844 6884 255876
rect 6916 255844 6920 255876
rect 6880 255796 6920 255844
rect 6880 255764 6884 255796
rect 6916 255764 6920 255796
rect 6880 255716 6920 255764
rect 6880 255684 6884 255716
rect 6916 255684 6920 255716
rect 6880 255680 6920 255684
rect 6960 255876 7000 255880
rect 6960 255844 6964 255876
rect 6996 255844 7000 255876
rect 6960 255796 7000 255844
rect 6960 255764 6964 255796
rect 6996 255764 7000 255796
rect 6960 255716 7000 255764
rect 6960 255684 6964 255716
rect 6996 255684 7000 255716
rect 6960 255680 7000 255684
rect 7040 255876 7080 255880
rect 7040 255844 7044 255876
rect 7076 255844 7080 255876
rect 7040 255796 7080 255844
rect 7040 255764 7044 255796
rect 7076 255764 7080 255796
rect 7040 255716 7080 255764
rect 7040 255684 7044 255716
rect 7076 255684 7080 255716
rect 7040 255680 7080 255684
rect 7120 255876 7160 255880
rect 7120 255844 7124 255876
rect 7156 255844 7160 255876
rect 7120 255796 7160 255844
rect 7120 255764 7124 255796
rect 7156 255764 7160 255796
rect 7120 255716 7160 255764
rect 7120 255684 7124 255716
rect 7156 255684 7160 255716
rect 7120 255680 7160 255684
rect 7200 255876 7240 255880
rect 7200 255844 7204 255876
rect 7236 255844 7240 255876
rect 7200 255796 7240 255844
rect 7200 255764 7204 255796
rect 7236 255764 7240 255796
rect 7200 255716 7240 255764
rect 7200 255684 7204 255716
rect 7236 255684 7240 255716
rect 7200 255680 7240 255684
rect 7280 255876 7320 255880
rect 7280 255844 7284 255876
rect 7316 255844 7320 255876
rect 7280 255796 7320 255844
rect 7280 255764 7284 255796
rect 7316 255764 7320 255796
rect 7280 255716 7320 255764
rect 7280 255684 7284 255716
rect 7316 255684 7320 255716
rect 7280 255680 7320 255684
rect 7360 255876 7400 255880
rect 7360 255844 7364 255876
rect 7396 255844 7400 255876
rect 7360 255796 7400 255844
rect 7360 255764 7364 255796
rect 7396 255764 7400 255796
rect 7360 255716 7400 255764
rect 7360 255684 7364 255716
rect 7396 255684 7400 255716
rect 7360 255680 7400 255684
rect 7440 255876 7480 255880
rect 7440 255844 7444 255876
rect 7476 255844 7480 255876
rect 7440 255796 7480 255844
rect 7440 255764 7444 255796
rect 7476 255764 7480 255796
rect 7440 255716 7480 255764
rect 7440 255684 7444 255716
rect 7476 255684 7480 255716
rect 7440 255680 7480 255684
rect 7520 255876 7560 255880
rect 7520 255844 7524 255876
rect 7556 255844 7560 255876
rect 7520 255796 7560 255844
rect 7520 255764 7524 255796
rect 7556 255764 7560 255796
rect 7520 255716 7560 255764
rect 7520 255684 7524 255716
rect 7556 255684 7560 255716
rect 7520 255680 7560 255684
rect 7600 255876 7640 255880
rect 7600 255844 7604 255876
rect 7636 255844 7640 255876
rect 7600 255796 7640 255844
rect 7600 255764 7604 255796
rect 7636 255764 7640 255796
rect 7600 255716 7640 255764
rect 7600 255684 7604 255716
rect 7636 255684 7640 255716
rect 7600 255680 7640 255684
rect 7680 255876 7720 255880
rect 7680 255844 7684 255876
rect 7716 255844 7720 255876
rect 7680 255796 7720 255844
rect 7680 255764 7684 255796
rect 7716 255764 7720 255796
rect 7680 255716 7720 255764
rect 7680 255684 7684 255716
rect 7716 255684 7720 255716
rect 7680 255680 7720 255684
rect 7760 255876 7800 255880
rect 7760 255844 7764 255876
rect 7796 255844 7800 255876
rect 7760 255796 7800 255844
rect 7760 255764 7764 255796
rect 7796 255764 7800 255796
rect 7760 255716 7800 255764
rect 7760 255684 7764 255716
rect 7796 255684 7800 255716
rect 7760 255680 7800 255684
rect 7840 255876 7880 255880
rect 7840 255844 7844 255876
rect 7876 255844 7880 255876
rect 7840 255796 7880 255844
rect 7840 255764 7844 255796
rect 7876 255764 7880 255796
rect 7840 255716 7880 255764
rect 7840 255684 7844 255716
rect 7876 255684 7880 255716
rect 7840 255680 7880 255684
rect 7920 255876 7960 255880
rect 7920 255844 7924 255876
rect 7956 255844 7960 255876
rect 7920 255796 7960 255844
rect 7920 255764 7924 255796
rect 7956 255764 7960 255796
rect 7920 255716 7960 255764
rect 7920 255684 7924 255716
rect 7956 255684 7960 255716
rect 7920 255680 7960 255684
rect 8000 255876 8040 255880
rect 8000 255844 8004 255876
rect 8036 255844 8040 255876
rect 8000 255796 8040 255844
rect 8000 255764 8004 255796
rect 8036 255764 8040 255796
rect 8000 255716 8040 255764
rect 8000 255684 8004 255716
rect 8036 255684 8040 255716
rect 8000 255680 8040 255684
rect 8080 255876 8120 255880
rect 8080 255844 8084 255876
rect 8116 255844 8120 255876
rect 8080 255796 8120 255844
rect 8080 255764 8084 255796
rect 8116 255764 8120 255796
rect 8080 255716 8120 255764
rect 8080 255684 8084 255716
rect 8116 255684 8120 255716
rect 8080 255680 8120 255684
rect 8160 255876 8200 255880
rect 8160 255844 8164 255876
rect 8196 255844 8200 255876
rect 8160 255796 8200 255844
rect 8160 255764 8164 255796
rect 8196 255764 8200 255796
rect 8160 255716 8200 255764
rect 8160 255684 8164 255716
rect 8196 255684 8200 255716
rect 8160 255680 8200 255684
rect 8240 255876 8280 255880
rect 8240 255844 8244 255876
rect 8276 255844 8280 255876
rect 8240 255796 8280 255844
rect 8240 255764 8244 255796
rect 8276 255764 8280 255796
rect 8240 255716 8280 255764
rect 8240 255684 8244 255716
rect 8276 255684 8280 255716
rect 8240 255680 8280 255684
rect 8320 255876 8360 255880
rect 8320 255844 8324 255876
rect 8356 255844 8360 255876
rect 8320 255796 8360 255844
rect 8320 255764 8324 255796
rect 8356 255764 8360 255796
rect 8320 255716 8360 255764
rect 8320 255684 8324 255716
rect 8356 255684 8360 255716
rect 8320 255680 8360 255684
rect 8400 255876 8440 255880
rect 8400 255844 8404 255876
rect 8436 255844 8440 255876
rect 8400 255796 8440 255844
rect 8400 255764 8404 255796
rect 8436 255764 8440 255796
rect 8400 255716 8440 255764
rect 8400 255684 8404 255716
rect 8436 255684 8440 255716
rect 8400 255680 8440 255684
rect 8480 255876 8520 255880
rect 8480 255844 8484 255876
rect 8516 255844 8520 255876
rect 8480 255796 8520 255844
rect 8480 255764 8484 255796
rect 8516 255764 8520 255796
rect 8480 255716 8520 255764
rect 8480 255684 8484 255716
rect 8516 255684 8520 255716
rect 8480 255680 8520 255684
rect 8560 255876 8600 255880
rect 8560 255844 8564 255876
rect 8596 255844 8600 255876
rect 8560 255796 8600 255844
rect 8560 255764 8564 255796
rect 8596 255764 8600 255796
rect 8560 255716 8600 255764
rect 8560 255684 8564 255716
rect 8596 255684 8600 255716
rect 8560 255680 8600 255684
rect 8640 255876 8680 255880
rect 8640 255844 8644 255876
rect 8676 255844 8680 255876
rect 8640 255796 8680 255844
rect 8640 255764 8644 255796
rect 8676 255764 8680 255796
rect 8640 255716 8680 255764
rect 8640 255684 8644 255716
rect 8676 255684 8680 255716
rect 8640 255680 8680 255684
rect 8720 255876 8760 255880
rect 8720 255844 8724 255876
rect 8756 255844 8760 255876
rect 8720 255796 8760 255844
rect 8720 255764 8724 255796
rect 8756 255764 8760 255796
rect 8720 255716 8760 255764
rect 8720 255684 8724 255716
rect 8756 255684 8760 255716
rect 8720 255680 8760 255684
rect 8800 255876 8840 255880
rect 8800 255844 8804 255876
rect 8836 255844 8840 255876
rect 8800 255796 8840 255844
rect 8800 255764 8804 255796
rect 8836 255764 8840 255796
rect 8800 255716 8840 255764
rect 8800 255684 8804 255716
rect 8836 255684 8840 255716
rect 8800 255680 8840 255684
rect 8880 255876 8920 255880
rect 8880 255844 8884 255876
rect 8916 255844 8920 255876
rect 8880 255796 8920 255844
rect 8880 255764 8884 255796
rect 8916 255764 8920 255796
rect 8880 255716 8920 255764
rect 8880 255684 8884 255716
rect 8916 255684 8920 255716
rect 8880 255680 8920 255684
rect 8960 255876 9000 255880
rect 8960 255844 8964 255876
rect 8996 255844 9000 255876
rect 8960 255796 9000 255844
rect 8960 255764 8964 255796
rect 8996 255764 9000 255796
rect 8960 255716 9000 255764
rect 8960 255684 8964 255716
rect 8996 255684 9000 255716
rect 8960 255680 9000 255684
rect 9040 255876 9080 255880
rect 9040 255844 9044 255876
rect 9076 255844 9080 255876
rect 9040 255796 9080 255844
rect 9040 255764 9044 255796
rect 9076 255764 9080 255796
rect 9040 255716 9080 255764
rect 9040 255684 9044 255716
rect 9076 255684 9080 255716
rect 9040 255680 9080 255684
rect 9120 255876 9160 255880
rect 9120 255844 9124 255876
rect 9156 255844 9160 255876
rect 9120 255796 9160 255844
rect 9120 255764 9124 255796
rect 9156 255764 9160 255796
rect 9120 255716 9160 255764
rect 9120 255684 9124 255716
rect 9156 255684 9160 255716
rect 9120 255680 9160 255684
rect 9200 255876 9240 255880
rect 9200 255844 9204 255876
rect 9236 255844 9240 255876
rect 9200 255796 9240 255844
rect 9200 255764 9204 255796
rect 9236 255764 9240 255796
rect 9200 255716 9240 255764
rect 9200 255684 9204 255716
rect 9236 255684 9240 255716
rect 9200 255680 9240 255684
rect 9280 255876 9320 255880
rect 9280 255844 9284 255876
rect 9316 255844 9320 255876
rect 9280 255796 9320 255844
rect 9280 255764 9284 255796
rect 9316 255764 9320 255796
rect 9280 255716 9320 255764
rect 9280 255684 9284 255716
rect 9316 255684 9320 255716
rect 9280 255680 9320 255684
rect 9360 255876 9400 255880
rect 9360 255844 9364 255876
rect 9396 255844 9400 255876
rect 9360 255796 9400 255844
rect 9360 255764 9364 255796
rect 9396 255764 9400 255796
rect 9360 255716 9400 255764
rect 9360 255684 9364 255716
rect 9396 255684 9400 255716
rect 9360 255680 9400 255684
rect 9440 255876 9480 255880
rect 9440 255844 9444 255876
rect 9476 255844 9480 255876
rect 9440 255796 9480 255844
rect 9440 255764 9444 255796
rect 9476 255764 9480 255796
rect 9440 255716 9480 255764
rect 9440 255684 9444 255716
rect 9476 255684 9480 255716
rect 9440 255680 9480 255684
rect 9520 255876 9560 255880
rect 9520 255844 9524 255876
rect 9556 255844 9560 255876
rect 9520 255796 9560 255844
rect 9520 255764 9524 255796
rect 9556 255764 9560 255796
rect 9520 255716 9560 255764
rect 9520 255684 9524 255716
rect 9556 255684 9560 255716
rect 9520 255680 9560 255684
rect 9600 255876 9640 255880
rect 9600 255844 9604 255876
rect 9636 255844 9640 255876
rect 9600 255796 9640 255844
rect 9600 255764 9604 255796
rect 9636 255764 9640 255796
rect 9600 255716 9640 255764
rect 9600 255684 9604 255716
rect 9636 255684 9640 255716
rect 9600 255680 9640 255684
rect 9680 255876 9720 255880
rect 9680 255844 9684 255876
rect 9716 255844 9720 255876
rect 9680 255796 9720 255844
rect 9680 255764 9684 255796
rect 9716 255764 9720 255796
rect 9680 255716 9720 255764
rect 9680 255684 9684 255716
rect 9716 255684 9720 255716
rect 9680 255680 9720 255684
rect 9760 255876 9800 255880
rect 9760 255844 9764 255876
rect 9796 255844 9800 255876
rect 9760 255796 9800 255844
rect 9760 255764 9764 255796
rect 9796 255764 9800 255796
rect 9760 255716 9800 255764
rect 9760 255684 9764 255716
rect 9796 255684 9800 255716
rect 9760 255680 9800 255684
rect 9840 255876 9880 255880
rect 9840 255844 9844 255876
rect 9876 255844 9880 255876
rect 9840 255796 9880 255844
rect 9840 255764 9844 255796
rect 9876 255764 9880 255796
rect 9840 255716 9880 255764
rect 9840 255684 9844 255716
rect 9876 255684 9880 255716
rect 9840 255680 9880 255684
rect 9920 255876 9960 255880
rect 9920 255844 9924 255876
rect 9956 255844 9960 255876
rect 9920 255796 9960 255844
rect 9920 255764 9924 255796
rect 9956 255764 9960 255796
rect 9920 255716 9960 255764
rect 9920 255684 9924 255716
rect 9956 255684 9960 255716
rect 9920 255680 9960 255684
rect 10000 255876 10040 255880
rect 10000 255844 10004 255876
rect 10036 255844 10040 255876
rect 10000 255796 10040 255844
rect 10000 255764 10004 255796
rect 10036 255764 10040 255796
rect 10000 255716 10040 255764
rect 10000 255684 10004 255716
rect 10036 255684 10040 255716
rect 10000 255680 10040 255684
rect 10080 255876 10120 255880
rect 10080 255844 10084 255876
rect 10116 255844 10120 255876
rect 10080 255796 10120 255844
rect 10080 255764 10084 255796
rect 10116 255764 10120 255796
rect 10080 255716 10120 255764
rect 10080 255684 10084 255716
rect 10116 255684 10120 255716
rect 10080 255680 10120 255684
rect 10160 255876 10200 255880
rect 10160 255844 10164 255876
rect 10196 255844 10200 255876
rect 10160 255796 10200 255844
rect 10160 255764 10164 255796
rect 10196 255764 10200 255796
rect 10160 255716 10200 255764
rect 10160 255684 10164 255716
rect 10196 255684 10200 255716
rect 10160 255680 10200 255684
rect 10240 255876 10280 255880
rect 10240 255844 10244 255876
rect 10276 255844 10280 255876
rect 10240 255796 10280 255844
rect 10240 255764 10244 255796
rect 10276 255764 10280 255796
rect 10240 255716 10280 255764
rect 10240 255684 10244 255716
rect 10276 255684 10280 255716
rect 10240 255680 10280 255684
rect 10320 255876 10360 255880
rect 10320 255844 10324 255876
rect 10356 255844 10360 255876
rect 10320 255796 10360 255844
rect 10320 255764 10324 255796
rect 10356 255764 10360 255796
rect 10320 255716 10360 255764
rect 10320 255684 10324 255716
rect 10356 255684 10360 255716
rect 10320 255680 10360 255684
rect 10400 255876 10440 255880
rect 10400 255844 10404 255876
rect 10436 255844 10440 255876
rect 10400 255796 10440 255844
rect 10400 255764 10404 255796
rect 10436 255764 10440 255796
rect 10400 255716 10440 255764
rect 10400 255684 10404 255716
rect 10436 255684 10440 255716
rect 10400 255680 10440 255684
rect 10480 255876 10520 255880
rect 10480 255844 10484 255876
rect 10516 255844 10520 255876
rect 10480 255796 10520 255844
rect 10480 255764 10484 255796
rect 10516 255764 10520 255796
rect 10480 255716 10520 255764
rect 10480 255684 10484 255716
rect 10516 255684 10520 255716
rect 10480 255680 10520 255684
rect 10560 255876 10600 255880
rect 10560 255844 10564 255876
rect 10596 255844 10600 255876
rect 10560 255796 10600 255844
rect 10560 255764 10564 255796
rect 10596 255764 10600 255796
rect 10560 255716 10600 255764
rect 10560 255684 10564 255716
rect 10596 255684 10600 255716
rect 10560 255680 10600 255684
rect 10640 255876 10680 255880
rect 10640 255844 10644 255876
rect 10676 255844 10680 255876
rect 10640 255796 10680 255844
rect 10640 255764 10644 255796
rect 10676 255764 10680 255796
rect 10640 255716 10680 255764
rect 10640 255684 10644 255716
rect 10676 255684 10680 255716
rect 10640 255680 10680 255684
rect 10720 255876 10760 255880
rect 10720 255844 10724 255876
rect 10756 255844 10760 255876
rect 10720 255796 10760 255844
rect 10720 255764 10724 255796
rect 10756 255764 10760 255796
rect 10720 255716 10760 255764
rect 10720 255684 10724 255716
rect 10756 255684 10760 255716
rect 10720 255680 10760 255684
rect 10800 255876 10840 255880
rect 10800 255844 10804 255876
rect 10836 255844 10840 255876
rect 10800 255796 10840 255844
rect 10800 255764 10804 255796
rect 10836 255764 10840 255796
rect 10800 255716 10840 255764
rect 10800 255684 10804 255716
rect 10836 255684 10840 255716
rect 10800 255680 10840 255684
rect 10880 255876 10920 255880
rect 10880 255844 10884 255876
rect 10916 255844 10920 255876
rect 10880 255796 10920 255844
rect 10880 255764 10884 255796
rect 10916 255764 10920 255796
rect 10880 255716 10920 255764
rect 10880 255684 10884 255716
rect 10916 255684 10920 255716
rect 10880 255680 10920 255684
rect 10960 255876 11000 255880
rect 10960 255844 10964 255876
rect 10996 255844 11000 255876
rect 10960 255796 11000 255844
rect 10960 255764 10964 255796
rect 10996 255764 11000 255796
rect 10960 255716 11000 255764
rect 10960 255684 10964 255716
rect 10996 255684 11000 255716
rect 10960 255680 11000 255684
rect 11040 255876 11080 255880
rect 11040 255844 11044 255876
rect 11076 255844 11080 255876
rect 11040 255796 11080 255844
rect 11040 255764 11044 255796
rect 11076 255764 11080 255796
rect 11040 255716 11080 255764
rect 11040 255684 11044 255716
rect 11076 255684 11080 255716
rect 11040 255680 11080 255684
rect 11120 255876 11160 255880
rect 11120 255844 11124 255876
rect 11156 255844 11160 255876
rect 11120 255796 11160 255844
rect 11120 255764 11124 255796
rect 11156 255764 11160 255796
rect 11120 255716 11160 255764
rect 11120 255684 11124 255716
rect 11156 255684 11160 255716
rect 11120 255680 11160 255684
rect 11200 255876 11240 255880
rect 11200 255844 11204 255876
rect 11236 255844 11240 255876
rect 11200 255796 11240 255844
rect 11200 255764 11204 255796
rect 11236 255764 11240 255796
rect 11200 255716 11240 255764
rect 11200 255684 11204 255716
rect 11236 255684 11240 255716
rect 11200 255680 11240 255684
rect 11280 255876 11320 255880
rect 11280 255844 11284 255876
rect 11316 255844 11320 255876
rect 11280 255796 11320 255844
rect 11280 255764 11284 255796
rect 11316 255764 11320 255796
rect 11280 255716 11320 255764
rect 11280 255684 11284 255716
rect 11316 255684 11320 255716
rect 11280 255680 11320 255684
rect 11360 255876 11400 255880
rect 11360 255844 11364 255876
rect 11396 255844 11400 255876
rect 11360 255796 11400 255844
rect 11360 255764 11364 255796
rect 11396 255764 11400 255796
rect 11360 255716 11400 255764
rect 11360 255684 11364 255716
rect 11396 255684 11400 255716
rect 11360 255680 11400 255684
rect 11440 255876 11480 255880
rect 11440 255844 11444 255876
rect 11476 255844 11480 255876
rect 11440 255796 11480 255844
rect 11440 255764 11444 255796
rect 11476 255764 11480 255796
rect 11440 255716 11480 255764
rect 11440 255684 11444 255716
rect 11476 255684 11480 255716
rect 11440 255680 11480 255684
rect 11520 255876 11560 255880
rect 11520 255844 11524 255876
rect 11556 255844 11560 255876
rect 11520 255796 11560 255844
rect 11520 255764 11524 255796
rect 11556 255764 11560 255796
rect 11520 255716 11560 255764
rect 11520 255684 11524 255716
rect 11556 255684 11560 255716
rect 11520 255680 11560 255684
rect 11600 255876 11640 255880
rect 11600 255844 11604 255876
rect 11636 255844 11640 255876
rect 11600 255796 11640 255844
rect 11600 255764 11604 255796
rect 11636 255764 11640 255796
rect 11600 255716 11640 255764
rect 11600 255684 11604 255716
rect 11636 255684 11640 255716
rect 11600 255680 11640 255684
rect 11680 255876 11720 255880
rect 11680 255844 11684 255876
rect 11716 255844 11720 255876
rect 11680 255796 11720 255844
rect 11680 255764 11684 255796
rect 11716 255764 11720 255796
rect 11680 255716 11720 255764
rect 11680 255684 11684 255716
rect 11716 255684 11720 255716
rect 11680 255680 11720 255684
rect 11760 255876 11800 255880
rect 11760 255844 11764 255876
rect 11796 255844 11800 255876
rect 11760 255796 11800 255844
rect 11760 255764 11764 255796
rect 11796 255764 11800 255796
rect 11760 255716 11800 255764
rect 11760 255684 11764 255716
rect 11796 255684 11800 255716
rect 11760 255680 11800 255684
rect 11840 255876 11880 255880
rect 11840 255844 11844 255876
rect 11876 255844 11880 255876
rect 11840 255796 11880 255844
rect 11840 255764 11844 255796
rect 11876 255764 11880 255796
rect 11840 255716 11880 255764
rect 11840 255684 11844 255716
rect 11876 255684 11880 255716
rect 11840 255680 11880 255684
rect 11920 255876 11960 255880
rect 11920 255844 11924 255876
rect 11956 255844 11960 255876
rect 11920 255796 11960 255844
rect 11920 255764 11924 255796
rect 11956 255764 11960 255796
rect 11920 255716 11960 255764
rect 11920 255684 11924 255716
rect 11956 255684 11960 255716
rect 11920 255680 11960 255684
rect 12000 255876 12040 255880
rect 12000 255844 12004 255876
rect 12036 255844 12040 255876
rect 12000 255796 12040 255844
rect 12000 255764 12004 255796
rect 12036 255764 12040 255796
rect 12000 255716 12040 255764
rect 12000 255684 12004 255716
rect 12036 255684 12040 255716
rect 12000 255680 12040 255684
rect 12080 255876 12120 255880
rect 12080 255844 12084 255876
rect 12116 255844 12120 255876
rect 12080 255796 12120 255844
rect 12080 255764 12084 255796
rect 12116 255764 12120 255796
rect 12080 255716 12120 255764
rect 12080 255684 12084 255716
rect 12116 255684 12120 255716
rect 12080 255680 12120 255684
rect 12160 255876 12200 255880
rect 12160 255844 12164 255876
rect 12196 255844 12200 255876
rect 12160 255796 12200 255844
rect 12160 255764 12164 255796
rect 12196 255764 12200 255796
rect 12160 255716 12200 255764
rect 12160 255684 12164 255716
rect 12196 255684 12200 255716
rect 12160 255680 12200 255684
rect 12240 255876 12280 255880
rect 12240 255844 12244 255876
rect 12276 255844 12280 255876
rect 12240 255796 12280 255844
rect 12240 255764 12244 255796
rect 12276 255764 12280 255796
rect 12240 255716 12280 255764
rect 12240 255684 12244 255716
rect 12276 255684 12280 255716
rect 12240 255680 12280 255684
rect 12320 255876 12360 255880
rect 12320 255844 12324 255876
rect 12356 255844 12360 255876
rect 12320 255796 12360 255844
rect 12320 255764 12324 255796
rect 12356 255764 12360 255796
rect 12320 255716 12360 255764
rect 12320 255684 12324 255716
rect 12356 255684 12360 255716
rect 12320 255680 12360 255684
rect 12400 255876 12440 255880
rect 12400 255844 12404 255876
rect 12436 255844 12440 255876
rect 12400 255796 12440 255844
rect 12400 255764 12404 255796
rect 12436 255764 12440 255796
rect 12400 255716 12440 255764
rect 12400 255684 12404 255716
rect 12436 255684 12440 255716
rect 12400 255680 12440 255684
rect 12480 255876 12520 255880
rect 12480 255844 12484 255876
rect 12516 255844 12520 255876
rect 12480 255796 12520 255844
rect 12480 255764 12484 255796
rect 12516 255764 12520 255796
rect 12480 255716 12520 255764
rect 12480 255684 12484 255716
rect 12516 255684 12520 255716
rect 12480 255680 12520 255684
rect 12560 255876 12600 255880
rect 12560 255844 12564 255876
rect 12596 255844 12600 255876
rect 12560 255796 12600 255844
rect 12560 255764 12564 255796
rect 12596 255764 12600 255796
rect 12560 255716 12600 255764
rect 12560 255684 12564 255716
rect 12596 255684 12600 255716
rect 12560 255680 12600 255684
rect 12640 255876 12680 255880
rect 12640 255844 12644 255876
rect 12676 255844 12680 255876
rect 12640 255796 12680 255844
rect 12640 255764 12644 255796
rect 12676 255764 12680 255796
rect 12640 255716 12680 255764
rect 12640 255684 12644 255716
rect 12676 255684 12680 255716
rect 12640 255680 12680 255684
rect 12720 255876 12760 255880
rect 12720 255844 12724 255876
rect 12756 255844 12760 255876
rect 12720 255796 12760 255844
rect 12720 255764 12724 255796
rect 12756 255764 12760 255796
rect 12720 255716 12760 255764
rect 12720 255684 12724 255716
rect 12756 255684 12760 255716
rect 12720 255680 12760 255684
rect 12800 255876 12840 255880
rect 12800 255844 12804 255876
rect 12836 255844 12840 255876
rect 12800 255796 12840 255844
rect 12800 255764 12804 255796
rect 12836 255764 12840 255796
rect 12800 255716 12840 255764
rect 12800 255684 12804 255716
rect 12836 255684 12840 255716
rect 12800 255680 12840 255684
rect 12880 255876 12920 255880
rect 12880 255844 12884 255876
rect 12916 255844 12920 255876
rect 12880 255796 12920 255844
rect 12880 255764 12884 255796
rect 12916 255764 12920 255796
rect 12880 255716 12920 255764
rect 12880 255684 12884 255716
rect 12916 255684 12920 255716
rect 12880 255680 12920 255684
rect 12960 255876 13000 255880
rect 12960 255844 12964 255876
rect 12996 255844 13000 255876
rect 12960 255796 13000 255844
rect 12960 255764 12964 255796
rect 12996 255764 13000 255796
rect 12960 255716 13000 255764
rect 12960 255684 12964 255716
rect 12996 255684 13000 255716
rect 12960 255680 13000 255684
rect 13040 255876 13080 255880
rect 13040 255844 13044 255876
rect 13076 255844 13080 255876
rect 13040 255796 13080 255844
rect 13040 255764 13044 255796
rect 13076 255764 13080 255796
rect 13040 255716 13080 255764
rect 13040 255684 13044 255716
rect 13076 255684 13080 255716
rect 13040 255680 13080 255684
rect 13120 255876 13160 255880
rect 13120 255844 13124 255876
rect 13156 255844 13160 255876
rect 13120 255796 13160 255844
rect 13120 255764 13124 255796
rect 13156 255764 13160 255796
rect 13120 255716 13160 255764
rect 13120 255684 13124 255716
rect 13156 255684 13160 255716
rect 13120 255680 13160 255684
rect 13200 255876 13240 255880
rect 13200 255844 13204 255876
rect 13236 255844 13240 255876
rect 13200 255796 13240 255844
rect 13200 255764 13204 255796
rect 13236 255764 13240 255796
rect 13200 255716 13240 255764
rect 13200 255684 13204 255716
rect 13236 255684 13240 255716
rect 13200 255680 13240 255684
rect 13280 255876 13320 255880
rect 13280 255844 13284 255876
rect 13316 255844 13320 255876
rect 13280 255796 13320 255844
rect 13280 255764 13284 255796
rect 13316 255764 13320 255796
rect 13280 255716 13320 255764
rect 13280 255684 13284 255716
rect 13316 255684 13320 255716
rect 13280 255680 13320 255684
rect 13360 255876 13400 255880
rect 13360 255844 13364 255876
rect 13396 255844 13400 255876
rect 13360 255796 13400 255844
rect 13360 255764 13364 255796
rect 13396 255764 13400 255796
rect 13360 255716 13400 255764
rect 13360 255684 13364 255716
rect 13396 255684 13400 255716
rect 13360 255680 13400 255684
rect 13440 255876 13480 255880
rect 13440 255844 13444 255876
rect 13476 255844 13480 255876
rect 13440 255796 13480 255844
rect 13440 255764 13444 255796
rect 13476 255764 13480 255796
rect 13440 255716 13480 255764
rect 13440 255684 13444 255716
rect 13476 255684 13480 255716
rect 13440 255680 13480 255684
rect 13520 255876 13560 255880
rect 13520 255844 13524 255876
rect 13556 255844 13560 255876
rect 13520 255796 13560 255844
rect 13520 255764 13524 255796
rect 13556 255764 13560 255796
rect 13520 255716 13560 255764
rect 13520 255684 13524 255716
rect 13556 255684 13560 255716
rect 13520 255680 13560 255684
rect 13600 255876 13640 255880
rect 13600 255844 13604 255876
rect 13636 255844 13640 255876
rect 13600 255796 13640 255844
rect 13600 255764 13604 255796
rect 13636 255764 13640 255796
rect 13600 255716 13640 255764
rect 13600 255684 13604 255716
rect 13636 255684 13640 255716
rect 13600 255680 13640 255684
rect 13680 255876 13720 255880
rect 13680 255844 13684 255876
rect 13716 255844 13720 255876
rect 13680 255796 13720 255844
rect 13680 255764 13684 255796
rect 13716 255764 13720 255796
rect 13680 255716 13720 255764
rect 13680 255684 13684 255716
rect 13716 255684 13720 255716
rect 13680 255680 13720 255684
rect 13760 255876 13800 255880
rect 13760 255844 13764 255876
rect 13796 255844 13800 255876
rect 13760 255796 13800 255844
rect 13760 255764 13764 255796
rect 13796 255764 13800 255796
rect 13760 255716 13800 255764
rect 13760 255684 13764 255716
rect 13796 255684 13800 255716
rect 13760 255680 13800 255684
rect 13840 255876 13880 255880
rect 13840 255844 13844 255876
rect 13876 255844 13880 255876
rect 13840 255796 13880 255844
rect 13840 255764 13844 255796
rect 13876 255764 13880 255796
rect 13840 255716 13880 255764
rect 13840 255684 13844 255716
rect 13876 255684 13880 255716
rect 13840 255680 13880 255684
rect 13920 255876 13960 255880
rect 13920 255844 13924 255876
rect 13956 255844 13960 255876
rect 13920 255796 13960 255844
rect 13920 255764 13924 255796
rect 13956 255764 13960 255796
rect 13920 255716 13960 255764
rect 13920 255684 13924 255716
rect 13956 255684 13960 255716
rect 13920 255680 13960 255684
rect 14000 255876 14040 255880
rect 14000 255844 14004 255876
rect 14036 255844 14040 255876
rect 14000 255796 14040 255844
rect 14000 255764 14004 255796
rect 14036 255764 14040 255796
rect 14000 255716 14040 255764
rect 14000 255684 14004 255716
rect 14036 255684 14040 255716
rect 14000 255680 14040 255684
rect 14080 255876 14120 255880
rect 14080 255844 14084 255876
rect 14116 255844 14120 255876
rect 14080 255796 14120 255844
rect 14080 255764 14084 255796
rect 14116 255764 14120 255796
rect 14080 255716 14120 255764
rect 14080 255684 14084 255716
rect 14116 255684 14120 255716
rect 14080 255680 14120 255684
rect 14160 255876 14200 255880
rect 14160 255844 14164 255876
rect 14196 255844 14200 255876
rect 14160 255796 14200 255844
rect 14160 255764 14164 255796
rect 14196 255764 14200 255796
rect 14160 255716 14200 255764
rect 14160 255684 14164 255716
rect 14196 255684 14200 255716
rect 14160 255680 14200 255684
rect 14240 255876 14280 255880
rect 14240 255844 14244 255876
rect 14276 255844 14280 255876
rect 14240 255796 14280 255844
rect 14240 255764 14244 255796
rect 14276 255764 14280 255796
rect 14240 255716 14280 255764
rect 14240 255684 14244 255716
rect 14276 255684 14280 255716
rect 14240 255680 14280 255684
rect 14320 255876 14360 255880
rect 14320 255844 14324 255876
rect 14356 255844 14360 255876
rect 14320 255796 14360 255844
rect 14320 255764 14324 255796
rect 14356 255764 14360 255796
rect 14320 255716 14360 255764
rect 14320 255684 14324 255716
rect 14356 255684 14360 255716
rect 14320 255680 14360 255684
rect 14400 255876 14440 255880
rect 14400 255844 14404 255876
rect 14436 255844 14440 255876
rect 14400 255796 14440 255844
rect 14400 255764 14404 255796
rect 14436 255764 14440 255796
rect 14400 255716 14440 255764
rect 14400 255684 14404 255716
rect 14436 255684 14440 255716
rect 14400 255680 14440 255684
rect 14480 255876 14520 255880
rect 14480 255844 14484 255876
rect 14516 255844 14520 255876
rect 14480 255796 14520 255844
rect 14480 255764 14484 255796
rect 14516 255764 14520 255796
rect 14480 255716 14520 255764
rect 14480 255684 14484 255716
rect 14516 255684 14520 255716
rect 14480 255680 14520 255684
rect 14560 255876 14600 255880
rect 14560 255844 14564 255876
rect 14596 255844 14600 255876
rect 14560 255796 14600 255844
rect 14560 255764 14564 255796
rect 14596 255764 14600 255796
rect 14560 255716 14600 255764
rect 14560 255684 14564 255716
rect 14596 255684 14600 255716
rect 14560 255680 14600 255684
rect 14640 255876 14680 255880
rect 14640 255844 14644 255876
rect 14676 255844 14680 255876
rect 14640 255796 14680 255844
rect 14640 255764 14644 255796
rect 14676 255764 14680 255796
rect 14640 255716 14680 255764
rect 14640 255684 14644 255716
rect 14676 255684 14680 255716
rect 14640 255680 14680 255684
rect 14720 255876 14760 255880
rect 14720 255844 14724 255876
rect 14756 255844 14760 255876
rect 14720 255796 14760 255844
rect 14720 255764 14724 255796
rect 14756 255764 14760 255796
rect 14720 255716 14760 255764
rect 14720 255684 14724 255716
rect 14756 255684 14760 255716
rect 14720 255680 14760 255684
rect 14800 255876 14840 255880
rect 14800 255844 14804 255876
rect 14836 255844 14840 255876
rect 14800 255796 14840 255844
rect 14800 255764 14804 255796
rect 14836 255764 14840 255796
rect 14800 255716 14840 255764
rect 14800 255684 14804 255716
rect 14836 255684 14840 255716
rect 14800 255680 14840 255684
rect 14880 255876 14920 255880
rect 14880 255844 14884 255876
rect 14916 255844 14920 255876
rect 14880 255796 14920 255844
rect 14880 255764 14884 255796
rect 14916 255764 14920 255796
rect 14880 255716 14920 255764
rect 14880 255684 14884 255716
rect 14916 255684 14920 255716
rect 14880 255680 14920 255684
rect 14960 255876 15000 255880
rect 14960 255844 14964 255876
rect 14996 255844 15000 255876
rect 14960 255796 15000 255844
rect 14960 255764 14964 255796
rect 14996 255764 15000 255796
rect 14960 255716 15000 255764
rect 14960 255684 14964 255716
rect 14996 255684 15000 255716
rect 14960 255680 15000 255684
rect 15040 255876 15080 255880
rect 15040 255844 15044 255876
rect 15076 255844 15080 255876
rect 15040 255796 15080 255844
rect 15040 255764 15044 255796
rect 15076 255764 15080 255796
rect 15040 255716 15080 255764
rect 15040 255684 15044 255716
rect 15076 255684 15080 255716
rect 15040 255680 15080 255684
rect 15120 255876 15160 255880
rect 15120 255844 15124 255876
rect 15156 255844 15160 255876
rect 15120 255796 15160 255844
rect 15120 255764 15124 255796
rect 15156 255764 15160 255796
rect 15120 255716 15160 255764
rect 15120 255684 15124 255716
rect 15156 255684 15160 255716
rect 15120 255680 15160 255684
rect 15200 255876 15240 255880
rect 15200 255844 15204 255876
rect 15236 255844 15240 255876
rect 15200 255796 15240 255844
rect 15200 255764 15204 255796
rect 15236 255764 15240 255796
rect 15200 255716 15240 255764
rect 15200 255684 15204 255716
rect 15236 255684 15240 255716
rect 15200 255680 15240 255684
rect 15280 255876 15320 255880
rect 15280 255844 15284 255876
rect 15316 255844 15320 255876
rect 15280 255796 15320 255844
rect 15280 255764 15284 255796
rect 15316 255764 15320 255796
rect 15280 255716 15320 255764
rect 15280 255684 15284 255716
rect 15316 255684 15320 255716
rect 15280 255680 15320 255684
rect 15360 255876 15400 255880
rect 15360 255844 15364 255876
rect 15396 255844 15400 255876
rect 15360 255796 15400 255844
rect 15360 255764 15364 255796
rect 15396 255764 15400 255796
rect 15360 255716 15400 255764
rect 15360 255684 15364 255716
rect 15396 255684 15400 255716
rect 15360 255680 15400 255684
rect 15440 255876 15480 255880
rect 15440 255844 15444 255876
rect 15476 255844 15480 255876
rect 15440 255796 15480 255844
rect 15440 255764 15444 255796
rect 15476 255764 15480 255796
rect 15440 255716 15480 255764
rect 15440 255684 15444 255716
rect 15476 255684 15480 255716
rect 15440 255680 15480 255684
rect 15520 255876 15560 255880
rect 15520 255844 15524 255876
rect 15556 255844 15560 255876
rect 15520 255796 15560 255844
rect 15520 255764 15524 255796
rect 15556 255764 15560 255796
rect 15520 255716 15560 255764
rect 15520 255684 15524 255716
rect 15556 255684 15560 255716
rect 15520 255680 15560 255684
rect 15600 255876 15640 255880
rect 15600 255844 15604 255876
rect 15636 255844 15640 255876
rect 15600 255796 15640 255844
rect 15600 255764 15604 255796
rect 15636 255764 15640 255796
rect 15600 255716 15640 255764
rect 15600 255684 15604 255716
rect 15636 255684 15640 255716
rect 15600 255680 15640 255684
rect 15680 255876 15720 255880
rect 15680 255844 15684 255876
rect 15716 255844 15720 255876
rect 15680 255796 15720 255844
rect 15680 255764 15684 255796
rect 15716 255764 15720 255796
rect 15680 255716 15720 255764
rect 15680 255684 15684 255716
rect 15716 255684 15720 255716
rect 15680 255680 15720 255684
rect 15760 255876 15800 255880
rect 15760 255844 15764 255876
rect 15796 255844 15800 255876
rect 15760 255796 15800 255844
rect 15760 255764 15764 255796
rect 15796 255764 15800 255796
rect 15760 255716 15800 255764
rect 15760 255684 15764 255716
rect 15796 255684 15800 255716
rect 15760 255680 15800 255684
rect 15840 255876 15880 255880
rect 15840 255844 15844 255876
rect 15876 255844 15880 255876
rect 15840 255796 15880 255844
rect 15840 255764 15844 255796
rect 15876 255764 15880 255796
rect 15840 255716 15880 255764
rect 15840 255684 15844 255716
rect 15876 255684 15880 255716
rect 15840 255680 15880 255684
rect 15920 255876 15960 255880
rect 15920 255844 15924 255876
rect 15956 255844 15960 255876
rect 15920 255796 15960 255844
rect 15920 255764 15924 255796
rect 15956 255764 15960 255796
rect 15920 255716 15960 255764
rect 15920 255684 15924 255716
rect 15956 255684 15960 255716
rect 15920 255680 15960 255684
rect 16000 255876 16040 255880
rect 16000 255844 16004 255876
rect 16036 255844 16040 255876
rect 16000 255796 16040 255844
rect 16000 255764 16004 255796
rect 16036 255764 16040 255796
rect 16000 255716 16040 255764
rect 16000 255684 16004 255716
rect 16036 255684 16040 255716
rect 16000 255680 16040 255684
rect 16080 255876 16120 255880
rect 16080 255844 16084 255876
rect 16116 255844 16120 255876
rect 16080 255796 16120 255844
rect 16080 255764 16084 255796
rect 16116 255764 16120 255796
rect 16080 255716 16120 255764
rect 16080 255684 16084 255716
rect 16116 255684 16120 255716
rect 16080 255680 16120 255684
rect 16160 255876 16200 255880
rect 16160 255844 16164 255876
rect 16196 255844 16200 255876
rect 16160 255796 16200 255844
rect 16160 255764 16164 255796
rect 16196 255764 16200 255796
rect 16160 255716 16200 255764
rect 16160 255684 16164 255716
rect 16196 255684 16200 255716
rect 16160 255680 16200 255684
rect 16240 255876 16280 255880
rect 16240 255844 16244 255876
rect 16276 255844 16280 255876
rect 16240 255796 16280 255844
rect 16240 255764 16244 255796
rect 16276 255764 16280 255796
rect 16240 255716 16280 255764
rect 16240 255684 16244 255716
rect 16276 255684 16280 255716
rect 16240 255680 16280 255684
rect 16320 255876 16360 255880
rect 16320 255844 16324 255876
rect 16356 255844 16360 255876
rect 16320 255796 16360 255844
rect 16320 255764 16324 255796
rect 16356 255764 16360 255796
rect 16320 255716 16360 255764
rect 16320 255684 16324 255716
rect 16356 255684 16360 255716
rect 16320 255680 16360 255684
rect 16400 255876 16440 255880
rect 16400 255844 16404 255876
rect 16436 255844 16440 255876
rect 16400 255796 16440 255844
rect 16400 255764 16404 255796
rect 16436 255764 16440 255796
rect 16400 255716 16440 255764
rect 16400 255684 16404 255716
rect 16436 255684 16440 255716
rect 16400 255680 16440 255684
rect 16480 255876 16520 255880
rect 16480 255844 16484 255876
rect 16516 255844 16520 255876
rect 16480 255796 16520 255844
rect 16480 255764 16484 255796
rect 16516 255764 16520 255796
rect 16480 255716 16520 255764
rect 16480 255684 16484 255716
rect 16516 255684 16520 255716
rect 16480 255680 16520 255684
rect 16560 255876 16600 255880
rect 16560 255844 16564 255876
rect 16596 255844 16600 255876
rect 16560 255796 16600 255844
rect 16560 255764 16564 255796
rect 16596 255764 16600 255796
rect 16560 255716 16600 255764
rect 16560 255684 16564 255716
rect 16596 255684 16600 255716
rect 16560 255680 16600 255684
rect 16640 255876 16680 255880
rect 16640 255844 16644 255876
rect 16676 255844 16680 255876
rect 16640 255796 16680 255844
rect 16640 255764 16644 255796
rect 16676 255764 16680 255796
rect 16640 255716 16680 255764
rect 16640 255684 16644 255716
rect 16676 255684 16680 255716
rect 16640 255680 16680 255684
rect 16720 255876 16760 255964
rect 16720 255844 16724 255876
rect 16756 255844 16760 255876
rect 16720 255796 16760 255844
rect 16720 255764 16724 255796
rect 16756 255764 16760 255796
rect 16720 255716 16760 255764
rect 16800 275395 16840 275400
rect 16800 275365 16805 275395
rect 16835 275365 16840 275395
rect 16800 255795 16840 275365
rect 16800 255765 16805 255795
rect 16835 255765 16840 255795
rect 16800 255760 16840 255765
rect 16880 275396 16920 275444
rect 16880 275364 16884 275396
rect 16916 275364 16920 275396
rect 16880 275316 16920 275364
rect 16880 275284 16884 275316
rect 16916 275284 16920 275316
rect 16880 274956 16920 275284
rect 16960 275476 17000 275480
rect 16960 275444 16964 275476
rect 16996 275444 17000 275476
rect 16960 275396 17000 275444
rect 16960 275364 16964 275396
rect 16996 275364 17000 275396
rect 16960 275316 17000 275364
rect 16960 275284 16964 275316
rect 16996 275284 17000 275316
rect 16960 275280 17000 275284
rect 17040 275476 17080 275480
rect 17040 275444 17044 275476
rect 17076 275444 17080 275476
rect 17040 275396 17080 275444
rect 17040 275364 17044 275396
rect 17076 275364 17080 275396
rect 17040 275316 17080 275364
rect 17120 275476 17160 275480
rect 17120 275444 17124 275476
rect 17156 275444 17160 275476
rect 17120 275395 17160 275444
rect 17120 275365 17125 275395
rect 17155 275365 17160 275395
rect 17120 275360 17160 275365
rect 17200 275476 17240 275480
rect 17200 275444 17204 275476
rect 17236 275444 17240 275476
rect 17040 275284 17044 275316
rect 17076 275284 17080 275316
rect 17040 275280 17080 275284
rect 17200 275316 17240 275444
rect 17200 275284 17204 275316
rect 17236 275284 17240 275316
rect 17200 275280 17240 275284
rect 16880 274924 16884 274956
rect 16916 274924 16920 274956
rect 16880 274876 16920 274924
rect 27920 275195 27960 275440
rect 27920 275005 27925 275195
rect 27955 275005 27960 275195
rect 27920 274880 27960 275005
rect 28080 275195 28120 275440
rect 28080 275005 28085 275195
rect 28115 275005 28120 275195
rect 28080 274920 28120 275005
rect 28240 275195 28280 275440
rect 28240 275005 28245 275195
rect 28275 275005 28280 275195
rect 28240 274920 28280 275005
rect 28400 275356 28440 275440
rect 28400 275324 28404 275356
rect 28436 275324 28440 275356
rect 28400 275276 28440 275324
rect 28400 275244 28404 275276
rect 28436 275244 28440 275276
rect 28400 275195 28440 275244
rect 28400 275005 28405 275195
rect 28435 275005 28440 275195
rect 28400 274920 28440 275005
rect 28480 274920 28520 275400
rect 28560 275356 28600 275440
rect 28560 275324 28564 275356
rect 28596 275324 28600 275356
rect 28560 275276 28600 275324
rect 28560 275244 28564 275276
rect 28596 275244 28600 275276
rect 28560 275195 28600 275244
rect 28560 275005 28565 275195
rect 28595 275005 28600 275195
rect 28560 274920 28600 275005
rect 28640 274920 28680 275400
rect 28720 275356 28760 275440
rect 28720 275324 28724 275356
rect 28756 275324 28760 275356
rect 28720 275276 28760 275324
rect 28720 275244 28724 275276
rect 28756 275244 28760 275276
rect 28720 275195 28760 275244
rect 28720 275005 28725 275195
rect 28755 275005 28760 275195
rect 28720 274920 28760 275005
rect 258900 275190 259100 350200
rect 271300 350100 271500 350200
rect 271860 350376 271900 350424
rect 271860 350344 271864 350376
rect 271896 350344 271900 350376
rect 271860 350296 271900 350344
rect 271860 350264 271864 350296
rect 271896 350264 271900 350296
rect 271860 350216 271900 350264
rect 271860 350184 271864 350216
rect 271896 350184 271900 350216
rect 271860 350136 271900 350184
rect 271860 350104 271864 350136
rect 271896 350104 271900 350136
rect 271220 350060 271580 350100
rect 271220 349980 271260 350060
rect 271380 350020 271420 350060
rect 271540 350020 271580 350060
rect 271860 350056 271900 350104
rect 271860 350024 271864 350056
rect 271896 350024 271900 350056
rect 271860 350020 271900 350024
rect 271940 351735 271980 351740
rect 271940 351705 271945 351735
rect 271975 351705 271980 351735
rect 271940 349980 271980 351705
rect 272020 351736 272060 351784
rect 272020 351704 272024 351736
rect 272056 351704 272060 351736
rect 272020 351656 272060 351704
rect 272020 351624 272024 351656
rect 272056 351624 272060 351656
rect 272020 351576 272060 351624
rect 272100 351816 272140 351820
rect 272100 351784 272104 351816
rect 272136 351784 272140 351816
rect 272100 351736 272140 351784
rect 272100 351704 272104 351736
rect 272136 351704 272140 351736
rect 272100 351656 272140 351704
rect 272100 351624 272104 351656
rect 272136 351624 272140 351656
rect 272100 351620 272140 351624
rect 272180 351816 272220 351820
rect 272180 351784 272184 351816
rect 272216 351784 272220 351816
rect 272180 351736 272220 351784
rect 272180 351704 272184 351736
rect 272216 351704 272220 351736
rect 272180 351656 272220 351704
rect 272180 351624 272184 351656
rect 272216 351624 272220 351656
rect 272180 351620 272220 351624
rect 272260 351816 272300 351820
rect 272260 351784 272264 351816
rect 272296 351784 272300 351816
rect 272260 351736 272300 351784
rect 272260 351704 272264 351736
rect 272296 351704 272300 351736
rect 272260 351656 272300 351704
rect 272260 351624 272264 351656
rect 272296 351624 272300 351656
rect 272260 351620 272300 351624
rect 272340 351816 272380 351820
rect 272340 351784 272344 351816
rect 272376 351784 272380 351816
rect 272340 351736 272380 351784
rect 272340 351704 272344 351736
rect 272376 351704 272380 351736
rect 272340 351656 272380 351704
rect 272340 351624 272344 351656
rect 272376 351624 272380 351656
rect 272340 351620 272380 351624
rect 272420 351816 272460 351820
rect 272420 351784 272424 351816
rect 272456 351784 272460 351816
rect 272420 351736 272460 351784
rect 272420 351704 272424 351736
rect 272456 351704 272460 351736
rect 272420 351656 272460 351704
rect 272420 351624 272424 351656
rect 272456 351624 272460 351656
rect 272420 351620 272460 351624
rect 272500 351816 272540 351820
rect 272500 351784 272504 351816
rect 272536 351784 272540 351816
rect 272500 351736 272540 351784
rect 272500 351704 272504 351736
rect 272536 351704 272540 351736
rect 272500 351656 272540 351704
rect 272500 351624 272504 351656
rect 272536 351624 272540 351656
rect 272500 351620 272540 351624
rect 272580 351816 272620 351820
rect 272580 351784 272584 351816
rect 272616 351784 272620 351816
rect 272580 351736 272620 351784
rect 272580 351704 272584 351736
rect 272616 351704 272620 351736
rect 272580 351656 272620 351704
rect 272580 351624 272584 351656
rect 272616 351624 272620 351656
rect 272580 351620 272620 351624
rect 272660 351816 272700 351820
rect 272660 351784 272664 351816
rect 272696 351784 272700 351816
rect 272660 351736 272700 351784
rect 272660 351704 272664 351736
rect 272696 351704 272700 351736
rect 272660 351656 272700 351704
rect 272660 351624 272664 351656
rect 272696 351624 272700 351656
rect 272660 351620 272700 351624
rect 272740 351816 272780 351820
rect 272740 351784 272744 351816
rect 272776 351784 272780 351816
rect 272740 351736 272780 351784
rect 272740 351704 272744 351736
rect 272776 351704 272780 351736
rect 272740 351656 272780 351704
rect 272740 351624 272744 351656
rect 272776 351624 272780 351656
rect 272740 351620 272780 351624
rect 272820 351816 272860 351820
rect 272820 351784 272824 351816
rect 272856 351784 272860 351816
rect 272820 351736 272860 351784
rect 272820 351704 272824 351736
rect 272856 351704 272860 351736
rect 272820 351656 272860 351704
rect 272820 351624 272824 351656
rect 272856 351624 272860 351656
rect 272820 351620 272860 351624
rect 272900 351816 272940 351820
rect 272900 351784 272904 351816
rect 272936 351784 272940 351816
rect 272900 351736 272940 351784
rect 272900 351704 272904 351736
rect 272936 351704 272940 351736
rect 272900 351656 272940 351704
rect 272900 351624 272904 351656
rect 272936 351624 272940 351656
rect 272900 351620 272940 351624
rect 272980 351816 273020 351820
rect 272980 351784 272984 351816
rect 273016 351784 273020 351816
rect 272980 351736 273020 351784
rect 272980 351704 272984 351736
rect 273016 351704 273020 351736
rect 272980 351656 273020 351704
rect 272980 351624 272984 351656
rect 273016 351624 273020 351656
rect 272980 351620 273020 351624
rect 273060 351816 273100 351820
rect 273060 351784 273064 351816
rect 273096 351784 273100 351816
rect 273060 351736 273100 351784
rect 273060 351704 273064 351736
rect 273096 351704 273100 351736
rect 273060 351656 273100 351704
rect 273060 351624 273064 351656
rect 273096 351624 273100 351656
rect 273060 351620 273100 351624
rect 273140 351816 273180 351820
rect 273140 351784 273144 351816
rect 273176 351784 273180 351816
rect 273140 351736 273180 351784
rect 273140 351704 273144 351736
rect 273176 351704 273180 351736
rect 273140 351656 273180 351704
rect 273140 351624 273144 351656
rect 273176 351624 273180 351656
rect 273140 351620 273180 351624
rect 273220 351816 273260 351820
rect 273220 351784 273224 351816
rect 273256 351784 273260 351816
rect 273220 351736 273260 351784
rect 273220 351704 273224 351736
rect 273256 351704 273260 351736
rect 273220 351656 273260 351704
rect 273220 351624 273224 351656
rect 273256 351624 273260 351656
rect 273220 351620 273260 351624
rect 273300 351816 273340 351820
rect 273300 351784 273304 351816
rect 273336 351784 273340 351816
rect 273300 351736 273340 351784
rect 273300 351704 273304 351736
rect 273336 351704 273340 351736
rect 273300 351656 273340 351704
rect 273300 351624 273304 351656
rect 273336 351624 273340 351656
rect 273300 351620 273340 351624
rect 273380 351816 273420 351820
rect 273380 351784 273384 351816
rect 273416 351784 273420 351816
rect 273380 351736 273420 351784
rect 273380 351704 273384 351736
rect 273416 351704 273420 351736
rect 273380 351656 273420 351704
rect 273380 351624 273384 351656
rect 273416 351624 273420 351656
rect 273380 351620 273420 351624
rect 273460 351816 273500 351820
rect 273460 351784 273464 351816
rect 273496 351784 273500 351816
rect 273460 351736 273500 351784
rect 273460 351704 273464 351736
rect 273496 351704 273500 351736
rect 273460 351656 273500 351704
rect 273460 351624 273464 351656
rect 273496 351624 273500 351656
rect 273460 351620 273500 351624
rect 273540 351816 273580 351820
rect 273540 351784 273544 351816
rect 273576 351784 273580 351816
rect 273540 351736 273580 351784
rect 273540 351704 273544 351736
rect 273576 351704 273580 351736
rect 273540 351656 273580 351704
rect 273540 351624 273544 351656
rect 273576 351624 273580 351656
rect 273540 351620 273580 351624
rect 273620 351816 273660 351820
rect 273620 351784 273624 351816
rect 273656 351784 273660 351816
rect 273620 351736 273660 351784
rect 273620 351704 273624 351736
rect 273656 351704 273660 351736
rect 273620 351656 273660 351704
rect 273620 351624 273624 351656
rect 273656 351624 273660 351656
rect 273620 351620 273660 351624
rect 273700 351816 273740 351820
rect 273700 351784 273704 351816
rect 273736 351784 273740 351816
rect 273700 351736 273740 351784
rect 273700 351704 273704 351736
rect 273736 351704 273740 351736
rect 273700 351656 273740 351704
rect 273700 351624 273704 351656
rect 273736 351624 273740 351656
rect 273700 351620 273740 351624
rect 273780 351816 273820 351820
rect 273780 351784 273784 351816
rect 273816 351784 273820 351816
rect 273780 351736 273820 351784
rect 273780 351704 273784 351736
rect 273816 351704 273820 351736
rect 273780 351656 273820 351704
rect 273780 351624 273784 351656
rect 273816 351624 273820 351656
rect 273780 351620 273820 351624
rect 273860 351816 273900 351820
rect 273860 351784 273864 351816
rect 273896 351784 273900 351816
rect 273860 351736 273900 351784
rect 273860 351704 273864 351736
rect 273896 351704 273900 351736
rect 273860 351656 273900 351704
rect 273860 351624 273864 351656
rect 273896 351624 273900 351656
rect 273860 351620 273900 351624
rect 273940 351816 273980 351820
rect 273940 351784 273944 351816
rect 273976 351784 273980 351816
rect 273940 351736 273980 351784
rect 273940 351704 273944 351736
rect 273976 351704 273980 351736
rect 273940 351656 273980 351704
rect 273940 351624 273944 351656
rect 273976 351624 273980 351656
rect 273940 351620 273980 351624
rect 274020 351816 274060 351820
rect 274020 351784 274024 351816
rect 274056 351784 274060 351816
rect 274020 351736 274060 351784
rect 274020 351704 274024 351736
rect 274056 351704 274060 351736
rect 274020 351656 274060 351704
rect 274020 351624 274024 351656
rect 274056 351624 274060 351656
rect 274020 351620 274060 351624
rect 274100 351816 274140 351820
rect 274100 351784 274104 351816
rect 274136 351784 274140 351816
rect 274100 351736 274140 351784
rect 274100 351704 274104 351736
rect 274136 351704 274140 351736
rect 274100 351656 274140 351704
rect 274100 351624 274104 351656
rect 274136 351624 274140 351656
rect 274100 351620 274140 351624
rect 274180 351816 274220 351820
rect 274180 351784 274184 351816
rect 274216 351784 274220 351816
rect 274180 351736 274220 351784
rect 274180 351704 274184 351736
rect 274216 351704 274220 351736
rect 274180 351656 274220 351704
rect 274180 351624 274184 351656
rect 274216 351624 274220 351656
rect 274180 351620 274220 351624
rect 274260 351816 274300 351820
rect 274260 351784 274264 351816
rect 274296 351784 274300 351816
rect 274260 351736 274300 351784
rect 274260 351704 274264 351736
rect 274296 351704 274300 351736
rect 274260 351656 274300 351704
rect 274260 351624 274264 351656
rect 274296 351624 274300 351656
rect 274260 351620 274300 351624
rect 274340 351816 274380 351820
rect 274340 351784 274344 351816
rect 274376 351784 274380 351816
rect 274340 351736 274380 351784
rect 274340 351704 274344 351736
rect 274376 351704 274380 351736
rect 274340 351656 274380 351704
rect 274340 351624 274344 351656
rect 274376 351624 274380 351656
rect 274340 351620 274380 351624
rect 274420 351816 274460 351820
rect 274420 351784 274424 351816
rect 274456 351784 274460 351816
rect 274420 351736 274460 351784
rect 274420 351704 274424 351736
rect 274456 351704 274460 351736
rect 274420 351656 274460 351704
rect 274420 351624 274424 351656
rect 274456 351624 274460 351656
rect 274420 351620 274460 351624
rect 274500 351816 274540 351820
rect 274500 351784 274504 351816
rect 274536 351784 274540 351816
rect 274500 351736 274540 351784
rect 274500 351704 274504 351736
rect 274536 351704 274540 351736
rect 274500 351656 274540 351704
rect 274500 351624 274504 351656
rect 274536 351624 274540 351656
rect 274500 351620 274540 351624
rect 274580 351816 274620 351820
rect 274580 351784 274584 351816
rect 274616 351784 274620 351816
rect 274580 351736 274620 351784
rect 274580 351704 274584 351736
rect 274616 351704 274620 351736
rect 274580 351656 274620 351704
rect 274580 351624 274584 351656
rect 274616 351624 274620 351656
rect 274580 351620 274620 351624
rect 274660 351816 274700 351820
rect 274660 351784 274664 351816
rect 274696 351784 274700 351816
rect 274660 351736 274700 351784
rect 274660 351704 274664 351736
rect 274696 351704 274700 351736
rect 274660 351656 274700 351704
rect 274660 351624 274664 351656
rect 274696 351624 274700 351656
rect 274660 351620 274700 351624
rect 274740 351816 274780 351820
rect 274740 351784 274744 351816
rect 274776 351784 274780 351816
rect 274740 351736 274780 351784
rect 274740 351704 274744 351736
rect 274776 351704 274780 351736
rect 274740 351656 274780 351704
rect 274740 351624 274744 351656
rect 274776 351624 274780 351656
rect 274740 351620 274780 351624
rect 274820 351816 274860 351820
rect 274820 351784 274824 351816
rect 274856 351784 274860 351816
rect 274820 351736 274860 351784
rect 274820 351704 274824 351736
rect 274856 351704 274860 351736
rect 274820 351656 274860 351704
rect 274820 351624 274824 351656
rect 274856 351624 274860 351656
rect 274820 351620 274860 351624
rect 274900 351816 274940 351820
rect 274900 351784 274904 351816
rect 274936 351784 274940 351816
rect 274900 351736 274940 351784
rect 274900 351704 274904 351736
rect 274936 351704 274940 351736
rect 274900 351656 274940 351704
rect 274900 351624 274904 351656
rect 274936 351624 274940 351656
rect 274900 351620 274940 351624
rect 274980 351816 275020 351820
rect 274980 351784 274984 351816
rect 275016 351784 275020 351816
rect 274980 351736 275020 351784
rect 274980 351704 274984 351736
rect 275016 351704 275020 351736
rect 274980 351656 275020 351704
rect 274980 351624 274984 351656
rect 275016 351624 275020 351656
rect 274980 351620 275020 351624
rect 275060 351816 275100 351820
rect 275060 351784 275064 351816
rect 275096 351784 275100 351816
rect 275060 351736 275100 351784
rect 275060 351704 275064 351736
rect 275096 351704 275100 351736
rect 275060 351656 275100 351704
rect 275060 351624 275064 351656
rect 275096 351624 275100 351656
rect 275060 351620 275100 351624
rect 275140 351816 275180 351820
rect 275140 351784 275144 351816
rect 275176 351784 275180 351816
rect 275140 351736 275180 351784
rect 275140 351704 275144 351736
rect 275176 351704 275180 351736
rect 275140 351656 275180 351704
rect 275140 351624 275144 351656
rect 275176 351624 275180 351656
rect 275140 351620 275180 351624
rect 275220 351816 275260 351820
rect 275220 351784 275224 351816
rect 275256 351784 275260 351816
rect 275220 351736 275260 351784
rect 275220 351704 275224 351736
rect 275256 351704 275260 351736
rect 275220 351656 275260 351704
rect 275220 351624 275224 351656
rect 275256 351624 275260 351656
rect 275220 351620 275260 351624
rect 275300 351816 275340 351820
rect 275300 351784 275304 351816
rect 275336 351784 275340 351816
rect 275300 351736 275340 351784
rect 275300 351704 275304 351736
rect 275336 351704 275340 351736
rect 275300 351656 275340 351704
rect 275300 351624 275304 351656
rect 275336 351624 275340 351656
rect 275300 351620 275340 351624
rect 275380 351816 275420 351820
rect 275380 351784 275384 351816
rect 275416 351784 275420 351816
rect 275380 351736 275420 351784
rect 275380 351704 275384 351736
rect 275416 351704 275420 351736
rect 275380 351656 275420 351704
rect 275380 351624 275384 351656
rect 275416 351624 275420 351656
rect 275380 351620 275420 351624
rect 275460 351816 275500 351820
rect 275460 351784 275464 351816
rect 275496 351784 275500 351816
rect 275460 351736 275500 351784
rect 275460 351704 275464 351736
rect 275496 351704 275500 351736
rect 275460 351656 275500 351704
rect 275460 351624 275464 351656
rect 275496 351624 275500 351656
rect 275460 351620 275500 351624
rect 275540 351816 275580 351820
rect 275540 351784 275544 351816
rect 275576 351784 275580 351816
rect 275540 351736 275580 351784
rect 275540 351704 275544 351736
rect 275576 351704 275580 351736
rect 275540 351656 275580 351704
rect 275540 351624 275544 351656
rect 275576 351624 275580 351656
rect 275540 351620 275580 351624
rect 275620 351816 275660 351820
rect 275620 351784 275624 351816
rect 275656 351784 275660 351816
rect 275620 351736 275660 351784
rect 275620 351704 275624 351736
rect 275656 351704 275660 351736
rect 275620 351656 275660 351704
rect 275620 351624 275624 351656
rect 275656 351624 275660 351656
rect 275620 351620 275660 351624
rect 275700 351816 275740 351820
rect 275700 351784 275704 351816
rect 275736 351784 275740 351816
rect 275700 351736 275740 351784
rect 275700 351704 275704 351736
rect 275736 351704 275740 351736
rect 275700 351656 275740 351704
rect 275700 351624 275704 351656
rect 275736 351624 275740 351656
rect 275700 351620 275740 351624
rect 275780 351816 275820 351820
rect 275780 351784 275784 351816
rect 275816 351784 275820 351816
rect 275780 351736 275820 351784
rect 275780 351704 275784 351736
rect 275816 351704 275820 351736
rect 275780 351656 275820 351704
rect 275780 351624 275784 351656
rect 275816 351624 275820 351656
rect 275780 351620 275820 351624
rect 275860 351816 275900 351820
rect 275860 351784 275864 351816
rect 275896 351784 275900 351816
rect 275860 351736 275900 351784
rect 275860 351704 275864 351736
rect 275896 351704 275900 351736
rect 275860 351656 275900 351704
rect 275860 351624 275864 351656
rect 275896 351624 275900 351656
rect 275860 351620 275900 351624
rect 275940 351816 275980 351820
rect 275940 351784 275944 351816
rect 275976 351784 275980 351816
rect 275940 351736 275980 351784
rect 275940 351704 275944 351736
rect 275976 351704 275980 351736
rect 275940 351656 275980 351704
rect 275940 351624 275944 351656
rect 275976 351624 275980 351656
rect 275940 351620 275980 351624
rect 276020 351816 276060 351820
rect 276020 351784 276024 351816
rect 276056 351784 276060 351816
rect 276020 351736 276060 351784
rect 276020 351704 276024 351736
rect 276056 351704 276060 351736
rect 276020 351656 276060 351704
rect 276020 351624 276024 351656
rect 276056 351624 276060 351656
rect 276020 351620 276060 351624
rect 276100 351816 276140 351820
rect 276100 351784 276104 351816
rect 276136 351784 276140 351816
rect 276100 351736 276140 351784
rect 276100 351704 276104 351736
rect 276136 351704 276140 351736
rect 276100 351656 276140 351704
rect 276100 351624 276104 351656
rect 276136 351624 276140 351656
rect 276100 351620 276140 351624
rect 276180 351816 276220 351820
rect 276180 351784 276184 351816
rect 276216 351784 276220 351816
rect 276180 351736 276220 351784
rect 276180 351704 276184 351736
rect 276216 351704 276220 351736
rect 276180 351656 276220 351704
rect 276180 351624 276184 351656
rect 276216 351624 276220 351656
rect 276180 351620 276220 351624
rect 276260 351816 276300 351820
rect 276260 351784 276264 351816
rect 276296 351784 276300 351816
rect 276260 351736 276300 351784
rect 276260 351704 276264 351736
rect 276296 351704 276300 351736
rect 276260 351656 276300 351704
rect 276260 351624 276264 351656
rect 276296 351624 276300 351656
rect 276260 351620 276300 351624
rect 276340 351816 276380 351820
rect 276340 351784 276344 351816
rect 276376 351784 276380 351816
rect 276340 351736 276380 351784
rect 276340 351704 276344 351736
rect 276376 351704 276380 351736
rect 276340 351656 276380 351704
rect 276340 351624 276344 351656
rect 276376 351624 276380 351656
rect 276340 351620 276380 351624
rect 276420 351816 276460 351820
rect 276420 351784 276424 351816
rect 276456 351784 276460 351816
rect 276420 351736 276460 351784
rect 276420 351704 276424 351736
rect 276456 351704 276460 351736
rect 276420 351656 276460 351704
rect 276420 351624 276424 351656
rect 276456 351624 276460 351656
rect 276420 351620 276460 351624
rect 276500 351816 276540 351820
rect 276500 351784 276504 351816
rect 276536 351784 276540 351816
rect 276500 351736 276540 351784
rect 276500 351704 276504 351736
rect 276536 351704 276540 351736
rect 276500 351656 276540 351704
rect 276500 351624 276504 351656
rect 276536 351624 276540 351656
rect 276500 351620 276540 351624
rect 276580 351816 276620 351820
rect 276580 351784 276584 351816
rect 276616 351784 276620 351816
rect 276580 351736 276620 351784
rect 276580 351704 276584 351736
rect 276616 351704 276620 351736
rect 276580 351656 276620 351704
rect 276580 351624 276584 351656
rect 276616 351624 276620 351656
rect 276580 351620 276620 351624
rect 276660 351816 276700 351820
rect 276660 351784 276664 351816
rect 276696 351784 276700 351816
rect 276660 351736 276700 351784
rect 276660 351704 276664 351736
rect 276696 351704 276700 351736
rect 276660 351656 276700 351704
rect 276660 351624 276664 351656
rect 276696 351624 276700 351656
rect 276660 351620 276700 351624
rect 276740 351816 276780 351820
rect 276740 351784 276744 351816
rect 276776 351784 276780 351816
rect 276740 351736 276780 351784
rect 276740 351704 276744 351736
rect 276776 351704 276780 351736
rect 276740 351656 276780 351704
rect 276740 351624 276744 351656
rect 276776 351624 276780 351656
rect 276740 351620 276780 351624
rect 276820 351816 276860 351820
rect 276820 351784 276824 351816
rect 276856 351784 276860 351816
rect 276820 351736 276860 351784
rect 276820 351704 276824 351736
rect 276856 351704 276860 351736
rect 276820 351656 276860 351704
rect 276820 351624 276824 351656
rect 276856 351624 276860 351656
rect 276820 351620 276860 351624
rect 276900 351816 276940 351820
rect 276900 351784 276904 351816
rect 276936 351784 276940 351816
rect 276900 351736 276940 351784
rect 276900 351704 276904 351736
rect 276936 351704 276940 351736
rect 276900 351656 276940 351704
rect 276900 351624 276904 351656
rect 276936 351624 276940 351656
rect 276900 351620 276940 351624
rect 276980 351816 277020 351820
rect 276980 351784 276984 351816
rect 277016 351784 277020 351816
rect 276980 351736 277020 351784
rect 276980 351704 276984 351736
rect 277016 351704 277020 351736
rect 276980 351656 277020 351704
rect 276980 351624 276984 351656
rect 277016 351624 277020 351656
rect 276980 351620 277020 351624
rect 277060 351816 277100 351820
rect 277060 351784 277064 351816
rect 277096 351784 277100 351816
rect 277060 351736 277100 351784
rect 277060 351704 277064 351736
rect 277096 351704 277100 351736
rect 277060 351656 277100 351704
rect 277060 351624 277064 351656
rect 277096 351624 277100 351656
rect 277060 351620 277100 351624
rect 277140 351816 277180 351820
rect 277140 351784 277144 351816
rect 277176 351784 277180 351816
rect 277140 351736 277180 351784
rect 277140 351704 277144 351736
rect 277176 351704 277180 351736
rect 277140 351656 277180 351704
rect 277140 351624 277144 351656
rect 277176 351624 277180 351656
rect 277140 351620 277180 351624
rect 277220 351816 277260 351820
rect 277220 351784 277224 351816
rect 277256 351784 277260 351816
rect 277220 351736 277260 351784
rect 277220 351704 277224 351736
rect 277256 351704 277260 351736
rect 277220 351656 277260 351704
rect 277220 351624 277224 351656
rect 277256 351624 277260 351656
rect 277220 351620 277260 351624
rect 277300 351816 277340 351820
rect 277300 351784 277304 351816
rect 277336 351784 277340 351816
rect 277300 351736 277340 351784
rect 277300 351704 277304 351736
rect 277336 351704 277340 351736
rect 277300 351656 277340 351704
rect 277300 351624 277304 351656
rect 277336 351624 277340 351656
rect 277300 351620 277340 351624
rect 277380 351816 277420 351820
rect 277380 351784 277384 351816
rect 277416 351784 277420 351816
rect 277380 351736 277420 351784
rect 277380 351704 277384 351736
rect 277416 351704 277420 351736
rect 277380 351656 277420 351704
rect 277380 351624 277384 351656
rect 277416 351624 277420 351656
rect 277380 351620 277420 351624
rect 277460 351816 277500 351820
rect 277460 351784 277464 351816
rect 277496 351784 277500 351816
rect 277460 351736 277500 351784
rect 277460 351704 277464 351736
rect 277496 351704 277500 351736
rect 277460 351656 277500 351704
rect 277460 351624 277464 351656
rect 277496 351624 277500 351656
rect 277460 351620 277500 351624
rect 277540 351816 277580 351820
rect 277540 351784 277544 351816
rect 277576 351784 277580 351816
rect 277540 351736 277580 351784
rect 277540 351704 277544 351736
rect 277576 351704 277580 351736
rect 277540 351656 277580 351704
rect 277540 351624 277544 351656
rect 277576 351624 277580 351656
rect 277540 351620 277580 351624
rect 277620 351816 277660 351820
rect 277620 351784 277624 351816
rect 277656 351784 277660 351816
rect 277620 351736 277660 351784
rect 277620 351704 277624 351736
rect 277656 351704 277660 351736
rect 277620 351656 277660 351704
rect 277620 351624 277624 351656
rect 277656 351624 277660 351656
rect 277620 351620 277660 351624
rect 277700 351816 277740 351820
rect 277700 351784 277704 351816
rect 277736 351784 277740 351816
rect 277700 351736 277740 351784
rect 277700 351704 277704 351736
rect 277736 351704 277740 351736
rect 277700 351656 277740 351704
rect 277700 351624 277704 351656
rect 277736 351624 277740 351656
rect 277700 351620 277740 351624
rect 277780 351816 277820 351820
rect 277780 351784 277784 351816
rect 277816 351784 277820 351816
rect 277780 351736 277820 351784
rect 277780 351704 277784 351736
rect 277816 351704 277820 351736
rect 277780 351656 277820 351704
rect 277780 351624 277784 351656
rect 277816 351624 277820 351656
rect 277780 351620 277820 351624
rect 277860 351816 277900 351820
rect 277860 351784 277864 351816
rect 277896 351784 277900 351816
rect 277860 351736 277900 351784
rect 277860 351704 277864 351736
rect 277896 351704 277900 351736
rect 277860 351656 277900 351704
rect 277860 351624 277864 351656
rect 277896 351624 277900 351656
rect 277860 351620 277900 351624
rect 277940 351816 277980 351820
rect 277940 351784 277944 351816
rect 277976 351784 277980 351816
rect 277940 351736 277980 351784
rect 277940 351704 277944 351736
rect 277976 351704 277980 351736
rect 277940 351656 277980 351704
rect 277940 351624 277944 351656
rect 277976 351624 277980 351656
rect 277940 351620 277980 351624
rect 278020 351816 278060 351820
rect 278020 351784 278024 351816
rect 278056 351784 278060 351816
rect 278020 351736 278060 351784
rect 278020 351704 278024 351736
rect 278056 351704 278060 351736
rect 278020 351656 278060 351704
rect 278020 351624 278024 351656
rect 278056 351624 278060 351656
rect 278020 351620 278060 351624
rect 278100 351816 278140 351820
rect 278100 351784 278104 351816
rect 278136 351784 278140 351816
rect 278100 351736 278140 351784
rect 278100 351704 278104 351736
rect 278136 351704 278140 351736
rect 278100 351656 278140 351704
rect 278100 351624 278104 351656
rect 278136 351624 278140 351656
rect 278100 351620 278140 351624
rect 278180 351816 278220 351820
rect 278180 351784 278184 351816
rect 278216 351784 278220 351816
rect 278180 351736 278220 351784
rect 278180 351704 278184 351736
rect 278216 351704 278220 351736
rect 278180 351656 278220 351704
rect 278180 351624 278184 351656
rect 278216 351624 278220 351656
rect 278180 351620 278220 351624
rect 278260 351816 278300 351820
rect 278260 351784 278264 351816
rect 278296 351784 278300 351816
rect 278260 351736 278300 351784
rect 278260 351704 278264 351736
rect 278296 351704 278300 351736
rect 278260 351656 278300 351704
rect 278260 351624 278264 351656
rect 278296 351624 278300 351656
rect 278260 351620 278300 351624
rect 278340 351816 278380 351820
rect 278340 351784 278344 351816
rect 278376 351784 278380 351816
rect 278340 351736 278380 351784
rect 278340 351704 278344 351736
rect 278376 351704 278380 351736
rect 278340 351656 278380 351704
rect 278340 351624 278344 351656
rect 278376 351624 278380 351656
rect 278340 351620 278380 351624
rect 278420 351816 278460 351820
rect 278420 351784 278424 351816
rect 278456 351784 278460 351816
rect 278420 351736 278460 351784
rect 278420 351704 278424 351736
rect 278456 351704 278460 351736
rect 278420 351656 278460 351704
rect 278420 351624 278424 351656
rect 278456 351624 278460 351656
rect 278420 351620 278460 351624
rect 278500 351816 278540 351820
rect 278500 351784 278504 351816
rect 278536 351784 278540 351816
rect 278500 351736 278540 351784
rect 278500 351704 278504 351736
rect 278536 351704 278540 351736
rect 278500 351656 278540 351704
rect 278500 351624 278504 351656
rect 278536 351624 278540 351656
rect 278500 351620 278540 351624
rect 278580 351816 278620 351820
rect 278580 351784 278584 351816
rect 278616 351784 278620 351816
rect 278580 351736 278620 351784
rect 278580 351704 278584 351736
rect 278616 351704 278620 351736
rect 278580 351656 278620 351704
rect 278580 351624 278584 351656
rect 278616 351624 278620 351656
rect 278580 351620 278620 351624
rect 278660 351816 278700 351820
rect 278660 351784 278664 351816
rect 278696 351784 278700 351816
rect 278660 351736 278700 351784
rect 278660 351704 278664 351736
rect 278696 351704 278700 351736
rect 278660 351656 278700 351704
rect 278660 351624 278664 351656
rect 278696 351624 278700 351656
rect 278660 351620 278700 351624
rect 278740 351816 278780 351820
rect 278740 351784 278744 351816
rect 278776 351784 278780 351816
rect 278740 351736 278780 351784
rect 278740 351704 278744 351736
rect 278776 351704 278780 351736
rect 278740 351656 278780 351704
rect 278740 351624 278744 351656
rect 278776 351624 278780 351656
rect 278740 351620 278780 351624
rect 278820 351816 278860 351820
rect 278820 351784 278824 351816
rect 278856 351784 278860 351816
rect 278820 351736 278860 351784
rect 278820 351704 278824 351736
rect 278856 351704 278860 351736
rect 278820 351656 278860 351704
rect 278820 351624 278824 351656
rect 278856 351624 278860 351656
rect 278820 351620 278860 351624
rect 278900 351816 278940 351820
rect 278900 351784 278904 351816
rect 278936 351784 278940 351816
rect 278900 351736 278940 351784
rect 278900 351704 278904 351736
rect 278936 351704 278940 351736
rect 278900 351656 278940 351704
rect 278900 351624 278904 351656
rect 278936 351624 278940 351656
rect 278900 351620 278940 351624
rect 278980 351816 279020 351820
rect 278980 351784 278984 351816
rect 279016 351784 279020 351816
rect 278980 351736 279020 351784
rect 278980 351704 278984 351736
rect 279016 351704 279020 351736
rect 278980 351656 279020 351704
rect 278980 351624 278984 351656
rect 279016 351624 279020 351656
rect 278980 351620 279020 351624
rect 279060 351816 279100 351820
rect 279060 351784 279064 351816
rect 279096 351784 279100 351816
rect 279060 351736 279100 351784
rect 279060 351704 279064 351736
rect 279096 351704 279100 351736
rect 279060 351656 279100 351704
rect 279060 351624 279064 351656
rect 279096 351624 279100 351656
rect 279060 351620 279100 351624
rect 279140 351816 279180 351820
rect 279140 351784 279144 351816
rect 279176 351784 279180 351816
rect 279140 351736 279180 351784
rect 279140 351704 279144 351736
rect 279176 351704 279180 351736
rect 279140 351656 279180 351704
rect 279140 351624 279144 351656
rect 279176 351624 279180 351656
rect 279140 351620 279180 351624
rect 279220 351816 279260 351820
rect 279220 351784 279224 351816
rect 279256 351784 279260 351816
rect 279220 351736 279260 351784
rect 279220 351704 279224 351736
rect 279256 351704 279260 351736
rect 279220 351656 279260 351704
rect 279220 351624 279224 351656
rect 279256 351624 279260 351656
rect 279220 351620 279260 351624
rect 279300 351816 279340 351820
rect 279300 351784 279304 351816
rect 279336 351784 279340 351816
rect 279300 351736 279340 351784
rect 279300 351704 279304 351736
rect 279336 351704 279340 351736
rect 279300 351656 279340 351704
rect 279300 351624 279304 351656
rect 279336 351624 279340 351656
rect 279300 351620 279340 351624
rect 279380 351816 279420 351820
rect 279380 351784 279384 351816
rect 279416 351784 279420 351816
rect 279380 351736 279420 351784
rect 279380 351704 279384 351736
rect 279416 351704 279420 351736
rect 279380 351656 279420 351704
rect 279380 351624 279384 351656
rect 279416 351624 279420 351656
rect 279380 351620 279420 351624
rect 279460 351816 279500 351820
rect 279460 351784 279464 351816
rect 279496 351784 279500 351816
rect 279460 351736 279500 351784
rect 279460 351704 279464 351736
rect 279496 351704 279500 351736
rect 279460 351656 279500 351704
rect 279460 351624 279464 351656
rect 279496 351624 279500 351656
rect 279460 351620 279500 351624
rect 279540 351816 279580 351820
rect 279540 351784 279544 351816
rect 279576 351784 279580 351816
rect 279540 351736 279580 351784
rect 279540 351704 279544 351736
rect 279576 351704 279580 351736
rect 279540 351656 279580 351704
rect 279540 351624 279544 351656
rect 279576 351624 279580 351656
rect 279540 351620 279580 351624
rect 279620 351816 279660 351820
rect 279620 351784 279624 351816
rect 279656 351784 279660 351816
rect 279620 351736 279660 351784
rect 279620 351704 279624 351736
rect 279656 351704 279660 351736
rect 279620 351656 279660 351704
rect 279620 351624 279624 351656
rect 279656 351624 279660 351656
rect 279620 351620 279660 351624
rect 279700 351816 279740 351820
rect 279700 351784 279704 351816
rect 279736 351784 279740 351816
rect 279700 351736 279740 351784
rect 279700 351704 279704 351736
rect 279736 351704 279740 351736
rect 279700 351656 279740 351704
rect 279700 351624 279704 351656
rect 279736 351624 279740 351656
rect 279700 351620 279740 351624
rect 279780 351816 279820 351820
rect 279780 351784 279784 351816
rect 279816 351784 279820 351816
rect 279780 351736 279820 351784
rect 279780 351704 279784 351736
rect 279816 351704 279820 351736
rect 279780 351656 279820 351704
rect 279780 351624 279784 351656
rect 279816 351624 279820 351656
rect 279780 351620 279820 351624
rect 279860 351816 279900 351820
rect 279860 351784 279864 351816
rect 279896 351784 279900 351816
rect 279860 351736 279900 351784
rect 279860 351704 279864 351736
rect 279896 351704 279900 351736
rect 279860 351656 279900 351704
rect 279860 351624 279864 351656
rect 279896 351624 279900 351656
rect 279860 351620 279900 351624
rect 279940 351816 279980 351820
rect 279940 351784 279944 351816
rect 279976 351784 279980 351816
rect 279940 351736 279980 351784
rect 279940 351704 279944 351736
rect 279976 351704 279980 351736
rect 279940 351656 279980 351704
rect 279940 351624 279944 351656
rect 279976 351624 279980 351656
rect 279940 351620 279980 351624
rect 280020 351816 280060 351820
rect 280020 351784 280024 351816
rect 280056 351784 280060 351816
rect 280020 351736 280060 351784
rect 280020 351704 280024 351736
rect 280056 351704 280060 351736
rect 280020 351656 280060 351704
rect 280020 351624 280024 351656
rect 280056 351624 280060 351656
rect 280020 351620 280060 351624
rect 280100 351816 280140 351820
rect 280100 351784 280104 351816
rect 280136 351784 280140 351816
rect 280100 351736 280140 351784
rect 280100 351704 280104 351736
rect 280136 351704 280140 351736
rect 280100 351656 280140 351704
rect 280100 351624 280104 351656
rect 280136 351624 280140 351656
rect 280100 351620 280140 351624
rect 280180 351816 280220 351820
rect 280180 351784 280184 351816
rect 280216 351784 280220 351816
rect 280180 351736 280220 351784
rect 280180 351704 280184 351736
rect 280216 351704 280220 351736
rect 280180 351656 280220 351704
rect 280180 351624 280184 351656
rect 280216 351624 280220 351656
rect 280180 351620 280220 351624
rect 280260 351816 280300 351820
rect 280260 351784 280264 351816
rect 280296 351784 280300 351816
rect 280260 351736 280300 351784
rect 280260 351704 280264 351736
rect 280296 351704 280300 351736
rect 280260 351656 280300 351704
rect 280260 351624 280264 351656
rect 280296 351624 280300 351656
rect 280260 351620 280300 351624
rect 280340 351816 280380 351820
rect 280340 351784 280344 351816
rect 280376 351784 280380 351816
rect 280340 351736 280380 351784
rect 280340 351704 280344 351736
rect 280376 351704 280380 351736
rect 280340 351656 280380 351704
rect 280340 351624 280344 351656
rect 280376 351624 280380 351656
rect 280340 351620 280380 351624
rect 280420 351816 280460 351820
rect 280420 351784 280424 351816
rect 280456 351784 280460 351816
rect 280420 351736 280460 351784
rect 280420 351704 280424 351736
rect 280456 351704 280460 351736
rect 280420 351656 280460 351704
rect 280420 351624 280424 351656
rect 280456 351624 280460 351656
rect 280420 351620 280460 351624
rect 280500 351816 280540 351820
rect 280500 351784 280504 351816
rect 280536 351784 280540 351816
rect 280500 351736 280540 351784
rect 280500 351704 280504 351736
rect 280536 351704 280540 351736
rect 280500 351656 280540 351704
rect 280500 351624 280504 351656
rect 280536 351624 280540 351656
rect 280500 351620 280540 351624
rect 280580 351816 280620 351820
rect 280580 351784 280584 351816
rect 280616 351784 280620 351816
rect 280580 351736 280620 351784
rect 280580 351704 280584 351736
rect 280616 351704 280620 351736
rect 280580 351656 280620 351704
rect 280580 351624 280584 351656
rect 280616 351624 280620 351656
rect 280580 351620 280620 351624
rect 280660 351816 280700 351820
rect 280660 351784 280664 351816
rect 280696 351784 280700 351816
rect 280660 351736 280700 351784
rect 280660 351704 280664 351736
rect 280696 351704 280700 351736
rect 280660 351656 280700 351704
rect 280660 351624 280664 351656
rect 280696 351624 280700 351656
rect 280660 351620 280700 351624
rect 280740 351816 280780 351820
rect 280740 351784 280744 351816
rect 280776 351784 280780 351816
rect 280740 351736 280780 351784
rect 280740 351704 280744 351736
rect 280776 351704 280780 351736
rect 280740 351656 280780 351704
rect 280740 351624 280744 351656
rect 280776 351624 280780 351656
rect 280740 351620 280780 351624
rect 280820 351816 280860 351820
rect 280820 351784 280824 351816
rect 280856 351784 280860 351816
rect 280820 351736 280860 351784
rect 280820 351704 280824 351736
rect 280856 351704 280860 351736
rect 280820 351656 280860 351704
rect 280820 351624 280824 351656
rect 280856 351624 280860 351656
rect 280820 351620 280860 351624
rect 280900 351816 280940 351820
rect 280900 351784 280904 351816
rect 280936 351784 280940 351816
rect 280900 351736 280940 351784
rect 280900 351704 280904 351736
rect 280936 351704 280940 351736
rect 280900 351656 280940 351704
rect 280900 351624 280904 351656
rect 280936 351624 280940 351656
rect 280900 351620 280940 351624
rect 280980 351816 281020 351820
rect 280980 351784 280984 351816
rect 281016 351784 281020 351816
rect 280980 351736 281020 351784
rect 280980 351704 280984 351736
rect 281016 351704 281020 351736
rect 280980 351656 281020 351704
rect 280980 351624 280984 351656
rect 281016 351624 281020 351656
rect 280980 351620 281020 351624
rect 281060 351816 281100 351820
rect 281060 351784 281064 351816
rect 281096 351784 281100 351816
rect 281060 351736 281100 351784
rect 281060 351704 281064 351736
rect 281096 351704 281100 351736
rect 281060 351656 281100 351704
rect 281060 351624 281064 351656
rect 281096 351624 281100 351656
rect 281060 351620 281100 351624
rect 281140 351816 281180 351820
rect 281140 351784 281144 351816
rect 281176 351784 281180 351816
rect 281140 351736 281180 351784
rect 281140 351704 281144 351736
rect 281176 351704 281180 351736
rect 281140 351656 281180 351704
rect 281140 351624 281144 351656
rect 281176 351624 281180 351656
rect 281140 351620 281180 351624
rect 281220 351816 281260 351820
rect 281220 351784 281224 351816
rect 281256 351784 281260 351816
rect 281220 351736 281260 351784
rect 281220 351704 281224 351736
rect 281256 351704 281260 351736
rect 281220 351656 281260 351704
rect 281220 351624 281224 351656
rect 281256 351624 281260 351656
rect 281220 351620 281260 351624
rect 281300 351816 281340 351820
rect 281300 351784 281304 351816
rect 281336 351784 281340 351816
rect 281300 351736 281340 351784
rect 281300 351704 281304 351736
rect 281336 351704 281340 351736
rect 281300 351656 281340 351704
rect 281300 351624 281304 351656
rect 281336 351624 281340 351656
rect 281300 351620 281340 351624
rect 281380 351816 281420 351820
rect 281380 351784 281384 351816
rect 281416 351784 281420 351816
rect 281380 351736 281420 351784
rect 281380 351704 281384 351736
rect 281416 351704 281420 351736
rect 281380 351656 281420 351704
rect 281380 351624 281384 351656
rect 281416 351624 281420 351656
rect 281380 351620 281420 351624
rect 281460 351816 281500 351820
rect 281460 351784 281464 351816
rect 281496 351784 281500 351816
rect 281460 351736 281500 351784
rect 281460 351704 281464 351736
rect 281496 351704 281500 351736
rect 281460 351656 281500 351704
rect 281460 351624 281464 351656
rect 281496 351624 281500 351656
rect 281460 351620 281500 351624
rect 281540 351816 281580 351820
rect 281540 351784 281544 351816
rect 281576 351784 281580 351816
rect 281540 351736 281580 351784
rect 281540 351704 281544 351736
rect 281576 351704 281580 351736
rect 281540 351656 281580 351704
rect 281540 351624 281544 351656
rect 281576 351624 281580 351656
rect 281540 351620 281580 351624
rect 281620 351816 281660 351820
rect 281620 351784 281624 351816
rect 281656 351784 281660 351816
rect 281620 351736 281660 351784
rect 281620 351704 281624 351736
rect 281656 351704 281660 351736
rect 281620 351656 281660 351704
rect 281620 351624 281624 351656
rect 281656 351624 281660 351656
rect 281620 351620 281660 351624
rect 281700 351816 281740 351820
rect 281700 351784 281704 351816
rect 281736 351784 281740 351816
rect 281700 351736 281740 351784
rect 281700 351704 281704 351736
rect 281736 351704 281740 351736
rect 281700 351656 281740 351704
rect 281700 351624 281704 351656
rect 281736 351624 281740 351656
rect 281700 351620 281740 351624
rect 281780 351816 281820 351820
rect 281780 351784 281784 351816
rect 281816 351784 281820 351816
rect 281780 351736 281820 351784
rect 281780 351704 281784 351736
rect 281816 351704 281820 351736
rect 281780 351656 281820 351704
rect 281780 351624 281784 351656
rect 281816 351624 281820 351656
rect 281780 351620 281820 351624
rect 281860 351816 281900 351820
rect 281860 351784 281864 351816
rect 281896 351784 281900 351816
rect 281860 351736 281900 351784
rect 281860 351704 281864 351736
rect 281896 351704 281900 351736
rect 281860 351656 281900 351704
rect 281860 351624 281864 351656
rect 281896 351624 281900 351656
rect 281860 351620 281900 351624
rect 281940 351816 281980 351820
rect 281940 351784 281944 351816
rect 281976 351784 281980 351816
rect 281940 351736 281980 351784
rect 281940 351704 281944 351736
rect 281976 351704 281980 351736
rect 281940 351656 281980 351704
rect 281940 351624 281944 351656
rect 281976 351624 281980 351656
rect 281940 351620 281980 351624
rect 282020 351816 282060 351820
rect 282020 351784 282024 351816
rect 282056 351784 282060 351816
rect 282020 351736 282060 351784
rect 282020 351704 282024 351736
rect 282056 351704 282060 351736
rect 282020 351656 282060 351704
rect 282020 351624 282024 351656
rect 282056 351624 282060 351656
rect 282020 351620 282060 351624
rect 282100 351816 282140 351820
rect 282100 351784 282104 351816
rect 282136 351784 282140 351816
rect 282100 351736 282140 351784
rect 282100 351704 282104 351736
rect 282136 351704 282140 351736
rect 282100 351656 282140 351704
rect 282100 351624 282104 351656
rect 282136 351624 282140 351656
rect 282100 351620 282140 351624
rect 282180 351816 282220 351820
rect 282180 351784 282184 351816
rect 282216 351784 282220 351816
rect 282180 351736 282220 351784
rect 282180 351704 282184 351736
rect 282216 351704 282220 351736
rect 282180 351656 282220 351704
rect 282180 351624 282184 351656
rect 282216 351624 282220 351656
rect 282180 351620 282220 351624
rect 282260 351816 282300 351820
rect 282260 351784 282264 351816
rect 282296 351784 282300 351816
rect 282260 351736 282300 351784
rect 282260 351704 282264 351736
rect 282296 351704 282300 351736
rect 282260 351656 282300 351704
rect 282260 351624 282264 351656
rect 282296 351624 282300 351656
rect 282260 351620 282300 351624
rect 282340 351816 282380 351820
rect 282340 351784 282344 351816
rect 282376 351784 282380 351816
rect 282340 351736 282380 351784
rect 282340 351704 282344 351736
rect 282376 351704 282380 351736
rect 282340 351656 282380 351704
rect 282340 351624 282344 351656
rect 282376 351624 282380 351656
rect 282340 351620 282380 351624
rect 282420 351816 282460 351820
rect 282420 351784 282424 351816
rect 282456 351784 282460 351816
rect 282420 351736 282460 351784
rect 282420 351704 282424 351736
rect 282456 351704 282460 351736
rect 282420 351656 282460 351704
rect 282420 351624 282424 351656
rect 282456 351624 282460 351656
rect 282420 351620 282460 351624
rect 282500 351816 282540 351820
rect 282500 351784 282504 351816
rect 282536 351784 282540 351816
rect 282500 351736 282540 351784
rect 282500 351704 282504 351736
rect 282536 351704 282540 351736
rect 282500 351656 282540 351704
rect 282500 351624 282504 351656
rect 282536 351624 282540 351656
rect 282500 351620 282540 351624
rect 282580 351816 282620 351820
rect 282580 351784 282584 351816
rect 282616 351784 282620 351816
rect 282580 351736 282620 351784
rect 282580 351704 282584 351736
rect 282616 351704 282620 351736
rect 282580 351656 282620 351704
rect 282580 351624 282584 351656
rect 282616 351624 282620 351656
rect 282580 351620 282620 351624
rect 282660 351816 282700 351820
rect 282660 351784 282664 351816
rect 282696 351784 282700 351816
rect 282660 351736 282700 351784
rect 282660 351704 282664 351736
rect 282696 351704 282700 351736
rect 282660 351656 282700 351704
rect 282660 351624 282664 351656
rect 282696 351624 282700 351656
rect 282660 351620 282700 351624
rect 282740 351816 282780 351820
rect 282740 351784 282744 351816
rect 282776 351784 282780 351816
rect 282740 351736 282780 351784
rect 282740 351704 282744 351736
rect 282776 351704 282780 351736
rect 282740 351656 282780 351704
rect 282740 351624 282744 351656
rect 282776 351624 282780 351656
rect 282740 351620 282780 351624
rect 282820 351816 282860 351820
rect 282820 351784 282824 351816
rect 282856 351784 282860 351816
rect 282820 351736 282860 351784
rect 282820 351704 282824 351736
rect 282856 351704 282860 351736
rect 282820 351656 282860 351704
rect 282820 351624 282824 351656
rect 282856 351624 282860 351656
rect 282820 351620 282860 351624
rect 282900 351816 282940 351820
rect 282900 351784 282904 351816
rect 282936 351784 282940 351816
rect 282900 351736 282940 351784
rect 282900 351704 282904 351736
rect 282936 351704 282940 351736
rect 282900 351656 282940 351704
rect 282900 351624 282904 351656
rect 282936 351624 282940 351656
rect 282900 351620 282940 351624
rect 282980 351816 283020 351820
rect 282980 351784 282984 351816
rect 283016 351784 283020 351816
rect 282980 351736 283020 351784
rect 282980 351704 282984 351736
rect 283016 351704 283020 351736
rect 282980 351656 283020 351704
rect 282980 351624 282984 351656
rect 283016 351624 283020 351656
rect 282980 351620 283020 351624
rect 283060 351816 283100 351820
rect 283060 351784 283064 351816
rect 283096 351784 283100 351816
rect 283060 351736 283100 351784
rect 283060 351704 283064 351736
rect 283096 351704 283100 351736
rect 283060 351656 283100 351704
rect 283060 351624 283064 351656
rect 283096 351624 283100 351656
rect 283060 351620 283100 351624
rect 283140 351816 283180 351820
rect 283140 351784 283144 351816
rect 283176 351784 283180 351816
rect 283140 351736 283180 351784
rect 283297 351740 285797 352400
rect 283140 351704 283144 351736
rect 283176 351704 283180 351736
rect 283140 351656 283180 351704
rect 283220 351735 285797 351740
rect 283220 351705 283225 351735
rect 283255 351705 285797 351735
rect 283220 351700 285797 351705
rect 283140 351624 283144 351656
rect 283176 351624 283180 351656
rect 283140 351620 283180 351624
rect 272020 351544 272024 351576
rect 272056 351544 272060 351576
rect 272020 351496 272060 351544
rect 272020 351464 272024 351496
rect 272056 351464 272060 351496
rect 272020 351416 272060 351464
rect 272020 351384 272024 351416
rect 272056 351384 272060 351416
rect 272020 351336 272060 351384
rect 272020 351304 272024 351336
rect 272056 351304 272060 351336
rect 272020 351256 272060 351304
rect 272020 351224 272024 351256
rect 272056 351224 272060 351256
rect 272020 351176 272060 351224
rect 272020 351144 272024 351176
rect 272056 351144 272060 351176
rect 283297 351150 285797 351700
rect 272020 351096 272060 351144
rect 272020 351064 272024 351096
rect 272056 351064 272060 351096
rect 272020 351016 272060 351064
rect 272020 350984 272024 351016
rect 272056 350984 272060 351016
rect 272020 350936 272060 350984
rect 272020 350904 272024 350936
rect 272056 350904 272060 350936
rect 272020 350856 272060 350904
rect 272020 350824 272024 350856
rect 272056 350824 272060 350856
rect 272020 350776 272060 350824
rect 272020 350744 272024 350776
rect 272056 350744 272060 350776
rect 272020 350696 272060 350744
rect 272020 350664 272024 350696
rect 272056 350664 272060 350696
rect 272020 350616 272060 350664
rect 272020 350584 272024 350616
rect 272056 350584 272060 350616
rect 272020 350536 272060 350584
rect 272020 350504 272024 350536
rect 272056 350504 272060 350536
rect 272020 350456 272060 350504
rect 272020 350424 272024 350456
rect 272056 350424 272060 350456
rect 272020 350376 272060 350424
rect 272020 350344 272024 350376
rect 272056 350344 272060 350376
rect 272020 350296 272060 350344
rect 272020 350264 272024 350296
rect 272056 350264 272060 350296
rect 272020 350216 272060 350264
rect 272020 350184 272024 350216
rect 272056 350184 272060 350216
rect 272020 350136 272060 350184
rect 272020 350104 272024 350136
rect 272056 350104 272060 350136
rect 272020 350056 272060 350104
rect 272020 350024 272024 350056
rect 272056 350024 272060 350056
rect 272020 350020 272060 350024
rect 291150 338992 292400 341492
rect 260500 338460 260540 338500
rect 260660 338460 260700 338500
rect 260820 338460 260860 338500
rect 260500 338420 260860 338460
rect 260600 277400 260800 338420
rect 291170 319892 292400 322292
rect 291170 314892 292400 317292
rect 291760 294736 292400 294792
rect 291760 294145 292400 294201
rect 291760 293554 292400 293610
rect 291760 292963 292400 293019
rect 291760 292372 292400 292428
rect 291760 291781 292400 291837
rect 291170 277400 292400 277681
rect 260600 277200 292400 277400
rect 291170 275281 292400 277200
rect 258900 275010 258910 275190
rect 259090 275010 259100 275190
rect 258900 275000 259100 275010
rect 16880 274844 16884 274876
rect 16916 274844 16920 274876
rect 16880 274795 16920 274844
rect 16880 274765 16885 274795
rect 16915 274765 16920 274795
rect 16880 274715 16920 274765
rect 16880 274685 16885 274715
rect 16915 274685 16920 274715
rect 16880 274635 16920 274685
rect 16880 274605 16885 274635
rect 16915 274605 16920 274635
rect 16880 274556 16920 274605
rect 16880 274524 16884 274556
rect 16916 274524 16920 274556
rect 16880 274476 16920 274524
rect 16880 274444 16884 274476
rect 16916 274444 16920 274476
rect 16880 274396 16920 274444
rect 16880 274364 16884 274396
rect 16916 274364 16920 274396
rect 16880 274316 16920 274364
rect 16880 274284 16884 274316
rect 16916 274284 16920 274316
rect 16880 274236 16920 274284
rect 16880 274204 16884 274236
rect 16916 274204 16920 274236
rect 16880 274156 16920 274204
rect 16880 274124 16884 274156
rect 16916 274124 16920 274156
rect 16880 274076 16920 274124
rect 16880 274044 16884 274076
rect 16916 274044 16920 274076
rect 16880 273996 16920 274044
rect 16880 273964 16884 273996
rect 16916 273964 16920 273996
rect 16880 273916 16920 273964
rect 16880 273884 16884 273916
rect 16916 273884 16920 273916
rect 16880 273836 16920 273884
rect 16880 273804 16884 273836
rect 16916 273804 16920 273836
rect 16880 273756 16920 273804
rect 16880 273724 16884 273756
rect 16916 273724 16920 273756
rect 16880 273676 16920 273724
rect 16880 273644 16884 273676
rect 16916 273644 16920 273676
rect 16880 273596 16920 273644
rect 16880 273564 16884 273596
rect 16916 273564 16920 273596
rect 16880 273516 16920 273564
rect 16880 273484 16884 273516
rect 16916 273484 16920 273516
rect 16880 273436 16920 273484
rect 16880 273404 16884 273436
rect 16916 273404 16920 273436
rect 16880 273356 16920 273404
rect 16880 273324 16884 273356
rect 16916 273324 16920 273356
rect 16880 273276 16920 273324
rect 16880 273244 16884 273276
rect 16916 273244 16920 273276
rect 16880 273196 16920 273244
rect 16880 273164 16884 273196
rect 16916 273164 16920 273196
rect 16880 273116 16920 273164
rect 16880 273084 16884 273116
rect 16916 273084 16920 273116
rect 16880 273036 16920 273084
rect 16880 273004 16884 273036
rect 16916 273004 16920 273036
rect 16880 272956 16920 273004
rect 16880 272924 16884 272956
rect 16916 272924 16920 272956
rect 16880 272876 16920 272924
rect 16880 272844 16884 272876
rect 16916 272844 16920 272876
rect 16880 272796 16920 272844
rect 16880 272764 16884 272796
rect 16916 272764 16920 272796
rect 16880 272716 16920 272764
rect 16880 272684 16884 272716
rect 16916 272684 16920 272716
rect 16880 272636 16920 272684
rect 16880 272604 16884 272636
rect 16916 272604 16920 272636
rect 16880 272556 16920 272604
rect 16880 272524 16884 272556
rect 16916 272524 16920 272556
rect 16880 272476 16920 272524
rect 16880 272444 16884 272476
rect 16916 272444 16920 272476
rect 16880 272396 16920 272444
rect 16880 272364 16884 272396
rect 16916 272364 16920 272396
rect 16880 272316 16920 272364
rect 16880 272284 16884 272316
rect 16916 272284 16920 272316
rect 16880 272236 16920 272284
rect 16880 272204 16884 272236
rect 16916 272204 16920 272236
rect 16880 272156 16920 272204
rect 16880 272124 16884 272156
rect 16916 272124 16920 272156
rect 16880 272076 16920 272124
rect 16880 272044 16884 272076
rect 16916 272044 16920 272076
rect 16880 271996 16920 272044
rect 16880 271964 16884 271996
rect 16916 271964 16920 271996
rect 16880 271916 16920 271964
rect 16880 271884 16884 271916
rect 16916 271884 16920 271916
rect 16880 271836 16920 271884
rect 16880 271804 16884 271836
rect 16916 271804 16920 271836
rect 16880 271756 16920 271804
rect 16880 271724 16884 271756
rect 16916 271724 16920 271756
rect 16880 271676 16920 271724
rect 16880 271644 16884 271676
rect 16916 271644 16920 271676
rect 16880 271596 16920 271644
rect 16880 271564 16884 271596
rect 16916 271564 16920 271596
rect 16880 271516 16920 271564
rect 16880 271484 16884 271516
rect 16916 271484 16920 271516
rect 16880 271436 16920 271484
rect 16880 271404 16884 271436
rect 16916 271404 16920 271436
rect 16880 271356 16920 271404
rect 16880 271324 16884 271356
rect 16916 271324 16920 271356
rect 16880 271276 16920 271324
rect 16880 271244 16884 271276
rect 16916 271244 16920 271276
rect 16880 271196 16920 271244
rect 16880 271164 16884 271196
rect 16916 271164 16920 271196
rect 16880 271116 16920 271164
rect 16880 271084 16884 271116
rect 16916 271084 16920 271116
rect 16880 271036 16920 271084
rect 16880 271004 16884 271036
rect 16916 271004 16920 271036
rect 16880 270956 16920 271004
rect 16880 270924 16884 270956
rect 16916 270924 16920 270956
rect 16880 270876 16920 270924
rect 16880 270844 16884 270876
rect 16916 270844 16920 270876
rect 16880 270796 16920 270844
rect 16880 270764 16884 270796
rect 16916 270764 16920 270796
rect 16880 270716 16920 270764
rect 16880 270684 16884 270716
rect 16916 270684 16920 270716
rect 16880 270636 16920 270684
rect 16880 270604 16884 270636
rect 16916 270604 16920 270636
rect 16880 270556 16920 270604
rect 16880 270524 16884 270556
rect 16916 270524 16920 270556
rect 16880 270476 16920 270524
rect 16880 270444 16884 270476
rect 16916 270444 16920 270476
rect 16880 270396 16920 270444
rect 16880 270364 16884 270396
rect 16916 270364 16920 270396
rect 16880 270316 16920 270364
rect 16880 270284 16884 270316
rect 16916 270284 16920 270316
rect 16880 270236 16920 270284
rect 291170 270281 292400 272681
rect 16880 270204 16884 270236
rect 16916 270204 16920 270236
rect 16880 270156 16920 270204
rect 16880 270124 16884 270156
rect 16916 270124 16920 270156
rect 16880 270076 16920 270124
rect 16880 270044 16884 270076
rect 16916 270044 16920 270076
rect 16880 269996 16920 270044
rect 16880 269964 16884 269996
rect 16916 269964 16920 269996
rect 16880 269916 16920 269964
rect 16880 269884 16884 269916
rect 16916 269884 16920 269916
rect 16880 269836 16920 269884
rect 16880 269804 16884 269836
rect 16916 269804 16920 269836
rect 16880 269756 16920 269804
rect 16880 269724 16884 269756
rect 16916 269724 16920 269756
rect 16880 269676 16920 269724
rect 16880 269644 16884 269676
rect 16916 269644 16920 269676
rect 16880 269596 16920 269644
rect 16880 269564 16884 269596
rect 16916 269564 16920 269596
rect 16880 269516 16920 269564
rect 16880 269484 16884 269516
rect 16916 269484 16920 269516
rect 16880 269436 16920 269484
rect 16880 269404 16884 269436
rect 16916 269404 16920 269436
rect 16880 269356 16920 269404
rect 16880 269324 16884 269356
rect 16916 269324 16920 269356
rect 16880 269276 16920 269324
rect 16880 269244 16884 269276
rect 16916 269244 16920 269276
rect 16880 269196 16920 269244
rect 16880 269164 16884 269196
rect 16916 269164 16920 269196
rect 16880 269116 16920 269164
rect 16880 269084 16884 269116
rect 16916 269084 16920 269116
rect 16880 269036 16920 269084
rect 16880 269004 16884 269036
rect 16916 269004 16920 269036
rect 16880 268956 16920 269004
rect 16880 268924 16884 268956
rect 16916 268924 16920 268956
rect 16880 268876 16920 268924
rect 16880 268844 16884 268876
rect 16916 268844 16920 268876
rect 16880 268796 16920 268844
rect 16880 268764 16884 268796
rect 16916 268764 16920 268796
rect 16880 268716 16920 268764
rect 16880 268684 16884 268716
rect 16916 268684 16920 268716
rect 16880 268636 16920 268684
rect 16880 268604 16884 268636
rect 16916 268604 16920 268636
rect 16880 268556 16920 268604
rect 16880 268524 16884 268556
rect 16916 268524 16920 268556
rect 16880 268476 16920 268524
rect 16880 268444 16884 268476
rect 16916 268444 16920 268476
rect 16880 268396 16920 268444
rect 16880 268364 16884 268396
rect 16916 268364 16920 268396
rect 16880 268316 16920 268364
rect 16880 268284 16884 268316
rect 16916 268284 16920 268316
rect 16880 268236 16920 268284
rect 16880 268204 16884 268236
rect 16916 268204 16920 268236
rect 16880 268156 16920 268204
rect 16880 268124 16884 268156
rect 16916 268124 16920 268156
rect 16880 268076 16920 268124
rect 16880 268044 16884 268076
rect 16916 268044 16920 268076
rect 16880 267996 16920 268044
rect 16880 267964 16884 267996
rect 16916 267964 16920 267996
rect 16880 267916 16920 267964
rect 16880 267884 16884 267916
rect 16916 267884 16920 267916
rect 16880 267836 16920 267884
rect 16880 267804 16884 267836
rect 16916 267804 16920 267836
rect 16880 267756 16920 267804
rect 16880 267724 16884 267756
rect 16916 267724 16920 267756
rect 16880 267676 16920 267724
rect 16880 267644 16884 267676
rect 16916 267644 16920 267676
rect 16880 267596 16920 267644
rect 16880 267564 16884 267596
rect 16916 267564 16920 267596
rect 16880 267516 16920 267564
rect 16880 267484 16884 267516
rect 16916 267484 16920 267516
rect 16880 267436 16920 267484
rect 16880 267404 16884 267436
rect 16916 267404 16920 267436
rect 16880 267356 16920 267404
rect 16880 267324 16884 267356
rect 16916 267324 16920 267356
rect 16880 267276 16920 267324
rect 16880 267244 16884 267276
rect 16916 267244 16920 267276
rect 16880 267196 16920 267244
rect 16880 267164 16884 267196
rect 16916 267164 16920 267196
rect 16880 267116 16920 267164
rect 16880 267084 16884 267116
rect 16916 267084 16920 267116
rect 16880 267036 16920 267084
rect 16880 267004 16884 267036
rect 16916 267004 16920 267036
rect 16880 266956 16920 267004
rect 16880 266924 16884 266956
rect 16916 266924 16920 266956
rect 16880 266876 16920 266924
rect 16880 266844 16884 266876
rect 16916 266844 16920 266876
rect 16880 266796 16920 266844
rect 16880 266764 16884 266796
rect 16916 266764 16920 266796
rect 16880 266716 16920 266764
rect 16880 266684 16884 266716
rect 16916 266684 16920 266716
rect 16880 266636 16920 266684
rect 16880 266604 16884 266636
rect 16916 266604 16920 266636
rect 16880 266556 16920 266604
rect 16880 266524 16884 266556
rect 16916 266524 16920 266556
rect 16880 266476 16920 266524
rect 16880 266444 16884 266476
rect 16916 266444 16920 266476
rect 16880 266396 16920 266444
rect 16880 266364 16884 266396
rect 16916 266364 16920 266396
rect 16880 266316 16920 266364
rect 16880 266284 16884 266316
rect 16916 266284 16920 266316
rect 16880 266236 16920 266284
rect 16880 266204 16884 266236
rect 16916 266204 16920 266236
rect 16880 266156 16920 266204
rect 16880 266124 16884 266156
rect 16916 266124 16920 266156
rect 16880 266076 16920 266124
rect 16880 266044 16884 266076
rect 16916 266044 16920 266076
rect 16880 265996 16920 266044
rect 16880 265964 16884 265996
rect 16916 265964 16920 265996
rect 16880 265916 16920 265964
rect 16880 265884 16884 265916
rect 16916 265884 16920 265916
rect 16880 265836 16920 265884
rect 16880 265804 16884 265836
rect 16916 265804 16920 265836
rect 16880 265756 16920 265804
rect 16880 265724 16884 265756
rect 16916 265724 16920 265756
rect 16880 265676 16920 265724
rect 16880 265644 16884 265676
rect 16916 265644 16920 265676
rect 16880 265596 16920 265644
rect 16880 265564 16884 265596
rect 16916 265564 16920 265596
rect 16880 265516 16920 265564
rect 16880 265484 16884 265516
rect 16916 265484 16920 265516
rect 16880 265436 16920 265484
rect 16880 265404 16884 265436
rect 16916 265404 16920 265436
rect 16880 265356 16920 265404
rect 16880 265324 16884 265356
rect 16916 265324 16920 265356
rect 16880 265276 16920 265324
rect 16880 265244 16884 265276
rect 16916 265244 16920 265276
rect 16880 265196 16920 265244
rect 16880 265164 16884 265196
rect 16916 265164 16920 265196
rect 16880 265116 16920 265164
rect 16880 265084 16884 265116
rect 16916 265084 16920 265116
rect 16880 265036 16920 265084
rect 16880 265004 16884 265036
rect 16916 265004 16920 265036
rect 16880 264956 16920 265004
rect 16880 264924 16884 264956
rect 16916 264924 16920 264956
rect 16880 264876 16920 264924
rect 16880 264844 16884 264876
rect 16916 264844 16920 264876
rect 16880 264796 16920 264844
rect 16880 264764 16884 264796
rect 16916 264764 16920 264796
rect 16880 264716 16920 264764
rect 16880 264684 16884 264716
rect 16916 264684 16920 264716
rect 16880 264636 16920 264684
rect 16880 264604 16884 264636
rect 16916 264604 16920 264636
rect 16880 264556 16920 264604
rect 16880 264524 16884 264556
rect 16916 264524 16920 264556
rect 16880 264476 16920 264524
rect 16880 264444 16884 264476
rect 16916 264444 16920 264476
rect 16880 264396 16920 264444
rect 16880 264364 16884 264396
rect 16916 264364 16920 264396
rect 16880 264316 16920 264364
rect 16880 264284 16884 264316
rect 16916 264284 16920 264316
rect 16880 264236 16920 264284
rect 16880 264204 16884 264236
rect 16916 264204 16920 264236
rect 16880 264156 16920 264204
rect 16880 264124 16884 264156
rect 16916 264124 16920 264156
rect 16880 264076 16920 264124
rect 16880 264044 16884 264076
rect 16916 264044 16920 264076
rect 16880 263996 16920 264044
rect 16880 263964 16884 263996
rect 16916 263964 16920 263996
rect 16880 263916 16920 263964
rect 16880 263884 16884 263916
rect 16916 263884 16920 263916
rect 16880 263836 16920 263884
rect 16880 263804 16884 263836
rect 16916 263804 16920 263836
rect 16880 263756 16920 263804
rect 16880 263724 16884 263756
rect 16916 263724 16920 263756
rect 16880 263676 16920 263724
rect 16880 263644 16884 263676
rect 16916 263644 16920 263676
rect 16880 263596 16920 263644
rect 16880 263564 16884 263596
rect 16916 263564 16920 263596
rect 16880 263516 16920 263564
rect 16880 263484 16884 263516
rect 16916 263484 16920 263516
rect 16880 263436 16920 263484
rect 16880 263404 16884 263436
rect 16916 263404 16920 263436
rect 16880 263356 16920 263404
rect 16880 263324 16884 263356
rect 16916 263324 16920 263356
rect 16880 263276 16920 263324
rect 16880 263244 16884 263276
rect 16916 263244 16920 263276
rect 16880 263196 16920 263244
rect 16880 263164 16884 263196
rect 16916 263164 16920 263196
rect 16880 263116 16920 263164
rect 16880 263084 16884 263116
rect 16916 263084 16920 263116
rect 16880 263036 16920 263084
rect 16880 263004 16884 263036
rect 16916 263004 16920 263036
rect 16880 262956 16920 263004
rect 16880 262924 16884 262956
rect 16916 262924 16920 262956
rect 16880 262876 16920 262924
rect 16880 262844 16884 262876
rect 16916 262844 16920 262876
rect 16880 262796 16920 262844
rect 16880 262764 16884 262796
rect 16916 262764 16920 262796
rect 16880 262716 16920 262764
rect 16880 262684 16884 262716
rect 16916 262684 16920 262716
rect 16880 262636 16920 262684
rect 16880 262604 16884 262636
rect 16916 262604 16920 262636
rect 16880 262556 16920 262604
rect 16880 262524 16884 262556
rect 16916 262524 16920 262556
rect 16880 262476 16920 262524
rect 16880 262444 16884 262476
rect 16916 262444 16920 262476
rect 16880 262396 16920 262444
rect 16880 262364 16884 262396
rect 16916 262364 16920 262396
rect 16880 262316 16920 262364
rect 16880 262284 16884 262316
rect 16916 262284 16920 262316
rect 16880 262236 16920 262284
rect 16880 262204 16884 262236
rect 16916 262204 16920 262236
rect 16880 262156 16920 262204
rect 16880 262124 16884 262156
rect 16916 262124 16920 262156
rect 16880 262076 16920 262124
rect 16880 262044 16884 262076
rect 16916 262044 16920 262076
rect 16880 261996 16920 262044
rect 16880 261964 16884 261996
rect 16916 261964 16920 261996
rect 16880 261916 16920 261964
rect 16880 261884 16884 261916
rect 16916 261884 16920 261916
rect 16880 261836 16920 261884
rect 16880 261804 16884 261836
rect 16916 261804 16920 261836
rect 16880 261756 16920 261804
rect 16880 261724 16884 261756
rect 16916 261724 16920 261756
rect 16880 261676 16920 261724
rect 16880 261644 16884 261676
rect 16916 261644 16920 261676
rect 16880 261596 16920 261644
rect 16880 261564 16884 261596
rect 16916 261564 16920 261596
rect 16880 261516 16920 261564
rect 16880 261484 16884 261516
rect 16916 261484 16920 261516
rect 16880 261436 16920 261484
rect 16880 261404 16884 261436
rect 16916 261404 16920 261436
rect 16880 261356 16920 261404
rect 16880 261324 16884 261356
rect 16916 261324 16920 261356
rect 16880 261276 16920 261324
rect 16880 261244 16884 261276
rect 16916 261244 16920 261276
rect 16880 261196 16920 261244
rect 16880 261164 16884 261196
rect 16916 261164 16920 261196
rect 16880 261116 16920 261164
rect 16880 261084 16884 261116
rect 16916 261084 16920 261116
rect 16880 261036 16920 261084
rect 16880 261004 16884 261036
rect 16916 261004 16920 261036
rect 16880 260956 16920 261004
rect 16880 260924 16884 260956
rect 16916 260924 16920 260956
rect 16880 260876 16920 260924
rect 16880 260844 16884 260876
rect 16916 260844 16920 260876
rect 16880 260796 16920 260844
rect 16880 260764 16884 260796
rect 16916 260764 16920 260796
rect 16880 260716 16920 260764
rect 16880 260684 16884 260716
rect 16916 260684 16920 260716
rect 16880 260636 16920 260684
rect 16880 260604 16884 260636
rect 16916 260604 16920 260636
rect 16880 260556 16920 260604
rect 16880 260524 16884 260556
rect 16916 260524 16920 260556
rect 16880 260476 16920 260524
rect 16880 260444 16884 260476
rect 16916 260444 16920 260476
rect 16880 260396 16920 260444
rect 16880 260364 16884 260396
rect 16916 260364 16920 260396
rect 16880 260316 16920 260364
rect 16880 260284 16884 260316
rect 16916 260284 16920 260316
rect 16880 260236 16920 260284
rect 16880 260204 16884 260236
rect 16916 260204 16920 260236
rect 16880 260156 16920 260204
rect 16880 260124 16884 260156
rect 16916 260124 16920 260156
rect 16880 260076 16920 260124
rect 16880 260044 16884 260076
rect 16916 260044 16920 260076
rect 16880 259996 16920 260044
rect 16880 259964 16884 259996
rect 16916 259964 16920 259996
rect 16880 259916 16920 259964
rect 16880 259884 16884 259916
rect 16916 259884 16920 259916
rect 16880 259836 16920 259884
rect 16880 259804 16884 259836
rect 16916 259804 16920 259836
rect 16880 259756 16920 259804
rect 16880 259724 16884 259756
rect 16916 259724 16920 259756
rect 16880 259676 16920 259724
rect 16880 259644 16884 259676
rect 16916 259644 16920 259676
rect 16880 259596 16920 259644
rect 16880 259564 16884 259596
rect 16916 259564 16920 259596
rect 16880 259516 16920 259564
rect 16880 259484 16884 259516
rect 16916 259484 16920 259516
rect 16880 259436 16920 259484
rect 16880 259404 16884 259436
rect 16916 259404 16920 259436
rect 16880 259356 16920 259404
rect 16880 259324 16884 259356
rect 16916 259324 16920 259356
rect 16880 259276 16920 259324
rect 16880 259244 16884 259276
rect 16916 259244 16920 259276
rect 16880 259196 16920 259244
rect 16880 259164 16884 259196
rect 16916 259164 16920 259196
rect 16880 259116 16920 259164
rect 16880 259084 16884 259116
rect 16916 259084 16920 259116
rect 16880 259036 16920 259084
rect 16880 259004 16884 259036
rect 16916 259004 16920 259036
rect 16880 258956 16920 259004
rect 16880 258924 16884 258956
rect 16916 258924 16920 258956
rect 16880 258876 16920 258924
rect 16880 258844 16884 258876
rect 16916 258844 16920 258876
rect 16880 258796 16920 258844
rect 16880 258764 16884 258796
rect 16916 258764 16920 258796
rect 16880 258716 16920 258764
rect 16880 258684 16884 258716
rect 16916 258684 16920 258716
rect 16880 258636 16920 258684
rect 16880 258604 16884 258636
rect 16916 258604 16920 258636
rect 16880 258556 16920 258604
rect 16880 258524 16884 258556
rect 16916 258524 16920 258556
rect 16880 258476 16920 258524
rect 16880 258444 16884 258476
rect 16916 258444 16920 258476
rect 16880 258396 16920 258444
rect 16880 258364 16884 258396
rect 16916 258364 16920 258396
rect 16880 258316 16920 258364
rect 16880 258284 16884 258316
rect 16916 258284 16920 258316
rect 16880 258236 16920 258284
rect 16880 258204 16884 258236
rect 16916 258204 16920 258236
rect 16880 258156 16920 258204
rect 16880 258124 16884 258156
rect 16916 258124 16920 258156
rect 16880 258076 16920 258124
rect 16880 258044 16884 258076
rect 16916 258044 16920 258076
rect 16880 257996 16920 258044
rect 16880 257964 16884 257996
rect 16916 257964 16920 257996
rect 16880 257916 16920 257964
rect 16880 257884 16884 257916
rect 16916 257884 16920 257916
rect 16880 257836 16920 257884
rect 16880 257804 16884 257836
rect 16916 257804 16920 257836
rect 16880 257756 16920 257804
rect 16880 257724 16884 257756
rect 16916 257724 16920 257756
rect 16880 257676 16920 257724
rect 16880 257644 16884 257676
rect 16916 257644 16920 257676
rect 16880 257596 16920 257644
rect 16880 257564 16884 257596
rect 16916 257564 16920 257596
rect 16880 257516 16920 257564
rect 16880 257484 16884 257516
rect 16916 257484 16920 257516
rect 16880 257436 16920 257484
rect 16880 257404 16884 257436
rect 16916 257404 16920 257436
rect 16880 257356 16920 257404
rect 16880 257324 16884 257356
rect 16916 257324 16920 257356
rect 16880 257276 16920 257324
rect 16880 257244 16884 257276
rect 16916 257244 16920 257276
rect 16880 257196 16920 257244
rect 16880 257164 16884 257196
rect 16916 257164 16920 257196
rect 16880 257116 16920 257164
rect 16880 257084 16884 257116
rect 16916 257084 16920 257116
rect 16880 257036 16920 257084
rect 16880 257004 16884 257036
rect 16916 257004 16920 257036
rect 16880 256956 16920 257004
rect 16880 256924 16884 256956
rect 16916 256924 16920 256956
rect 16880 256876 16920 256924
rect 16880 256844 16884 256876
rect 16916 256844 16920 256876
rect 16880 256796 16920 256844
rect 16880 256764 16884 256796
rect 16916 256764 16920 256796
rect 16880 256716 16920 256764
rect 16880 256684 16884 256716
rect 16916 256684 16920 256716
rect 16880 256636 16920 256684
rect 16880 256604 16884 256636
rect 16916 256604 16920 256636
rect 16880 256556 16920 256604
rect 16880 256524 16884 256556
rect 16916 256524 16920 256556
rect 16880 256476 16920 256524
rect 16880 256444 16884 256476
rect 16916 256444 16920 256476
rect 16880 256396 16920 256444
rect 16880 256364 16884 256396
rect 16916 256364 16920 256396
rect 16880 256316 16920 256364
rect 16880 256284 16884 256316
rect 16916 256284 16920 256316
rect 16880 256236 16920 256284
rect 16880 256204 16884 256236
rect 16916 256204 16920 256236
rect 16880 256156 16920 256204
rect 16880 256124 16884 256156
rect 16916 256124 16920 256156
rect 16880 256076 16920 256124
rect 16880 256044 16884 256076
rect 16916 256044 16920 256076
rect 16880 255996 16920 256044
rect 16880 255964 16884 255996
rect 16916 255964 16920 255996
rect 16880 255876 16920 255964
rect 16880 255844 16884 255876
rect 16916 255844 16920 255876
rect 16720 255684 16724 255716
rect 16756 255684 16760 255716
rect 16720 255680 16760 255684
rect 16880 255716 16920 255844
rect 16880 255684 16884 255716
rect 16916 255684 16920 255716
rect 16880 255680 16920 255684
rect 291760 250025 292400 250081
rect 291760 249434 292400 249490
rect 291760 248843 292400 248899
rect 291760 248252 292400 248308
rect 291760 247661 292400 247717
rect 291760 247070 292400 247126
rect 291760 227814 292400 227870
rect 291760 227223 292400 227279
rect 291760 226632 292400 226688
rect 291760 226041 292400 226097
rect 291760 225450 292400 225506
rect 291760 224859 292400 224915
rect 291760 205603 292400 205659
rect 291760 205012 292400 205068
rect 291760 204421 292400 204477
rect 291760 203830 292400 203886
rect 291760 203239 292400 203295
rect 291760 202648 292400 202704
rect 291760 182392 292400 182448
rect 291760 181801 292400 181857
rect 291760 181210 292400 181266
rect 291760 180619 292400 180675
rect 291760 180028 292400 180084
rect 291760 179437 292400 179493
rect 291760 159781 292400 159837
rect 291760 159190 292400 159246
rect 291760 158599 292400 158655
rect 291760 158008 292400 158064
rect 291760 157417 292400 157473
rect 291760 156826 292400 156882
rect 291760 137570 292400 137626
rect 291760 136979 292400 137035
rect 291760 136388 292400 136444
rect 291760 135797 292400 135853
rect 291760 135206 292400 135262
rect 291760 134615 292400 134671
rect 291170 117615 292400 120015
rect 291170 112615 292400 115015
rect -400 109600 3000 109800
rect -400 107444 830 109600
rect -400 102444 830 104844
rect 291170 95715 292400 98115
rect 291170 90715 292400 93115
rect -400 86444 830 88844
rect -400 81444 830 83844
rect 291170 73415 292400 75815
rect 291170 68415 292400 70815
rect -400 62388 240 62444
rect -400 61797 240 61853
rect -400 61206 240 61262
rect -400 60615 240 60671
rect -400 60024 240 60080
rect -400 59433 240 59489
rect 291760 47559 292400 47615
rect 291760 46968 292400 47024
rect 291760 46377 292400 46433
rect 291760 45786 292400 45842
rect -400 40777 240 40833
rect -400 40186 240 40242
rect -400 39595 240 39651
rect -400 39004 240 39060
rect -400 38413 240 38469
rect -400 37822 240 37878
rect 291760 25230 292400 25286
rect 291760 24639 292400 24695
rect 291760 24048 292400 24104
rect 291760 23457 292400 23513
rect -400 19166 240 19222
rect -400 18575 240 18631
rect -400 17984 240 18040
rect -400 17393 240 17449
rect -400 16802 240 16858
rect -400 16211 240 16267
rect 291760 12001 292400 12057
rect 291760 11410 292400 11466
rect 291760 10819 292400 10875
rect 291760 10228 292400 10284
rect 291760 9637 292400 9693
rect 291760 9046 292400 9102
rect -400 8455 240 8511
rect 291760 8455 292400 8511
rect -400 7864 240 7920
rect 291760 7864 292400 7920
rect -400 7273 240 7329
rect 291760 7273 292400 7329
rect -400 6682 240 6738
rect 291760 6682 292400 6738
rect -400 6091 240 6147
rect 291760 6091 292400 6147
rect -400 5500 240 5556
rect 291760 5500 292400 5556
rect -400 4909 240 4965
rect 291760 4909 292400 4965
rect -400 4318 240 4374
rect 291760 4318 292400 4374
rect -400 3727 240 3783
rect 291760 3727 292400 3783
rect -400 3136 240 3192
rect 291760 3136 292400 3192
rect -400 2545 240 2601
rect 291760 2545 292400 2601
rect -400 1954 240 2010
rect 291760 1954 292400 2010
rect -400 1363 240 1419
rect 291760 1363 292400 1419
rect -400 772 240 828
rect 291760 772 292400 828
<< via3 >>
rect 271864 351815 271896 351816
rect 271864 351785 271865 351815
rect 271865 351785 271895 351815
rect 271895 351785 271896 351815
rect 271864 351784 271896 351785
rect 272024 351815 272056 351816
rect 272024 351785 272025 351815
rect 272025 351785 272055 351815
rect 272055 351785 272056 351815
rect 272024 351784 272056 351785
rect 271864 351655 271896 351656
rect 271864 351625 271865 351655
rect 271865 351625 271895 351655
rect 271895 351625 271896 351655
rect 271864 351624 271896 351625
rect 271864 351575 271896 351576
rect 271864 351545 271865 351575
rect 271865 351545 271895 351575
rect 271895 351545 271896 351575
rect 271864 351544 271896 351545
rect 271864 351495 271896 351496
rect 271864 351465 271865 351495
rect 271865 351465 271895 351495
rect 271895 351465 271896 351495
rect 271864 351464 271896 351465
rect 271864 351415 271896 351416
rect 271864 351385 271865 351415
rect 271865 351385 271895 351415
rect 271895 351385 271896 351415
rect 271864 351384 271896 351385
rect 271864 351335 271896 351336
rect 271864 351305 271865 351335
rect 271865 351305 271895 351335
rect 271895 351305 271896 351335
rect 271864 351304 271896 351305
rect 271864 351255 271896 351256
rect 271864 351225 271865 351255
rect 271865 351225 271895 351255
rect 271895 351225 271896 351255
rect 271864 351224 271896 351225
rect 271864 351175 271896 351176
rect 271864 351145 271865 351175
rect 271865 351145 271895 351175
rect 271895 351145 271896 351175
rect 271864 351144 271896 351145
rect 271864 351095 271896 351096
rect 271864 351065 271865 351095
rect 271865 351065 271895 351095
rect 271895 351065 271896 351095
rect 271864 351064 271896 351065
rect 271864 351015 271896 351016
rect 271864 350985 271865 351015
rect 271865 350985 271895 351015
rect 271895 350985 271896 351015
rect 271864 350984 271896 350985
rect 271864 350935 271896 350936
rect 271864 350905 271865 350935
rect 271865 350905 271895 350935
rect 271895 350905 271896 350935
rect 271864 350904 271896 350905
rect 271864 350855 271896 350856
rect 271864 350825 271865 350855
rect 271865 350825 271895 350855
rect 271895 350825 271896 350855
rect 271864 350824 271896 350825
rect 271864 350775 271896 350776
rect 271864 350745 271865 350775
rect 271865 350745 271895 350775
rect 271895 350745 271896 350775
rect 271864 350744 271896 350745
rect 271864 350695 271896 350696
rect 271864 350665 271865 350695
rect 271865 350665 271895 350695
rect 271895 350665 271896 350695
rect 271864 350664 271896 350665
rect 271864 350615 271896 350616
rect 271864 350585 271865 350615
rect 271865 350585 271895 350615
rect 271895 350585 271896 350615
rect 271864 350584 271896 350585
rect 271864 350535 271896 350536
rect 271864 350505 271865 350535
rect 271865 350505 271895 350535
rect 271895 350505 271896 350535
rect 271864 350504 271896 350505
rect 271864 350455 271896 350456
rect 271864 350425 271865 350455
rect 271865 350425 271895 350455
rect 271895 350425 271896 350455
rect 271864 350424 271896 350425
rect 1010 317610 1190 317790
rect 16210 317610 16390 317790
rect 1040 275040 1160 275160
rect 16210 274610 16390 274790
rect 16724 275475 16756 275476
rect 16724 275445 16725 275475
rect 16725 275445 16755 275475
rect 16755 275445 16756 275475
rect 16724 275444 16756 275445
rect 16884 275475 16916 275476
rect 16884 275445 16885 275475
rect 16885 275445 16915 275475
rect 16915 275445 16916 275475
rect 16884 275444 16916 275445
rect 16724 275315 16756 275316
rect 16724 275285 16725 275315
rect 16725 275285 16755 275315
rect 16755 275285 16756 275315
rect 16724 275284 16756 275285
rect 16724 274955 16756 274956
rect 16724 274925 16725 274955
rect 16725 274925 16755 274955
rect 16755 274925 16756 274955
rect 16724 274924 16756 274925
rect 16724 274875 16756 274876
rect 16724 274845 16725 274875
rect 16725 274845 16755 274875
rect 16755 274845 16756 274875
rect 16724 274844 16756 274845
rect 16724 274555 16756 274556
rect 16724 274525 16725 274555
rect 16725 274525 16755 274555
rect 16755 274525 16756 274555
rect 16724 274524 16756 274525
rect 16724 274475 16756 274476
rect 16724 274445 16725 274475
rect 16725 274445 16755 274475
rect 16755 274445 16756 274475
rect 16724 274444 16756 274445
rect 16724 274395 16756 274396
rect 16724 274365 16725 274395
rect 16725 274365 16755 274395
rect 16755 274365 16756 274395
rect 16724 274364 16756 274365
rect 16724 274315 16756 274316
rect 16724 274285 16725 274315
rect 16725 274285 16755 274315
rect 16755 274285 16756 274315
rect 16724 274284 16756 274285
rect 16724 274235 16756 274236
rect 16724 274205 16725 274235
rect 16725 274205 16755 274235
rect 16755 274205 16756 274235
rect 16724 274204 16756 274205
rect 16724 274155 16756 274156
rect 16724 274125 16725 274155
rect 16725 274125 16755 274155
rect 16755 274125 16756 274155
rect 16724 274124 16756 274125
rect 16724 274075 16756 274076
rect 16724 274045 16725 274075
rect 16725 274045 16755 274075
rect 16755 274045 16756 274075
rect 16724 274044 16756 274045
rect 16724 273995 16756 273996
rect 16724 273965 16725 273995
rect 16725 273965 16755 273995
rect 16755 273965 16756 273995
rect 16724 273964 16756 273965
rect 16724 273915 16756 273916
rect 16724 273885 16725 273915
rect 16725 273885 16755 273915
rect 16755 273885 16756 273915
rect 16724 273884 16756 273885
rect 16724 273835 16756 273836
rect 16724 273805 16725 273835
rect 16725 273805 16755 273835
rect 16755 273805 16756 273835
rect 16724 273804 16756 273805
rect 16724 273755 16756 273756
rect 16724 273725 16725 273755
rect 16725 273725 16755 273755
rect 16755 273725 16756 273755
rect 16724 273724 16756 273725
rect 16724 273675 16756 273676
rect 16724 273645 16725 273675
rect 16725 273645 16755 273675
rect 16755 273645 16756 273675
rect 16724 273644 16756 273645
rect 16724 273595 16756 273596
rect 16724 273565 16725 273595
rect 16725 273565 16755 273595
rect 16755 273565 16756 273595
rect 16724 273564 16756 273565
rect 16724 273515 16756 273516
rect 16724 273485 16725 273515
rect 16725 273485 16755 273515
rect 16755 273485 16756 273515
rect 16724 273484 16756 273485
rect 16724 273435 16756 273436
rect 16724 273405 16725 273435
rect 16725 273405 16755 273435
rect 16755 273405 16756 273435
rect 16724 273404 16756 273405
rect 16724 273355 16756 273356
rect 16724 273325 16725 273355
rect 16725 273325 16755 273355
rect 16755 273325 16756 273355
rect 16724 273324 16756 273325
rect 16724 273275 16756 273276
rect 16724 273245 16725 273275
rect 16725 273245 16755 273275
rect 16755 273245 16756 273275
rect 16724 273244 16756 273245
rect 16724 273195 16756 273196
rect 16724 273165 16725 273195
rect 16725 273165 16755 273195
rect 16755 273165 16756 273195
rect 16724 273164 16756 273165
rect 16724 273115 16756 273116
rect 16724 273085 16725 273115
rect 16725 273085 16755 273115
rect 16755 273085 16756 273115
rect 16724 273084 16756 273085
rect 16724 273035 16756 273036
rect 16724 273005 16725 273035
rect 16725 273005 16755 273035
rect 16755 273005 16756 273035
rect 16724 273004 16756 273005
rect 16724 272955 16756 272956
rect 16724 272925 16725 272955
rect 16725 272925 16755 272955
rect 16755 272925 16756 272955
rect 16724 272924 16756 272925
rect 16724 272875 16756 272876
rect 16724 272845 16725 272875
rect 16725 272845 16755 272875
rect 16755 272845 16756 272875
rect 16724 272844 16756 272845
rect 16724 272795 16756 272796
rect 16724 272765 16725 272795
rect 16725 272765 16755 272795
rect 16755 272765 16756 272795
rect 16724 272764 16756 272765
rect 16724 272715 16756 272716
rect 16724 272685 16725 272715
rect 16725 272685 16755 272715
rect 16755 272685 16756 272715
rect 16724 272684 16756 272685
rect 16724 272635 16756 272636
rect 16724 272605 16725 272635
rect 16725 272605 16755 272635
rect 16755 272605 16756 272635
rect 16724 272604 16756 272605
rect 16724 272555 16756 272556
rect 16724 272525 16725 272555
rect 16725 272525 16755 272555
rect 16755 272525 16756 272555
rect 16724 272524 16756 272525
rect 16724 272475 16756 272476
rect 16724 272445 16725 272475
rect 16725 272445 16755 272475
rect 16755 272445 16756 272475
rect 16724 272444 16756 272445
rect 16724 272395 16756 272396
rect 16724 272365 16725 272395
rect 16725 272365 16755 272395
rect 16755 272365 16756 272395
rect 16724 272364 16756 272365
rect 16724 272315 16756 272316
rect 16724 272285 16725 272315
rect 16725 272285 16755 272315
rect 16755 272285 16756 272315
rect 16724 272284 16756 272285
rect 16724 272235 16756 272236
rect 16724 272205 16725 272235
rect 16725 272205 16755 272235
rect 16755 272205 16756 272235
rect 16724 272204 16756 272205
rect 16724 272155 16756 272156
rect 16724 272125 16725 272155
rect 16725 272125 16755 272155
rect 16755 272125 16756 272155
rect 16724 272124 16756 272125
rect 16724 272075 16756 272076
rect 16724 272045 16725 272075
rect 16725 272045 16755 272075
rect 16755 272045 16756 272075
rect 16724 272044 16756 272045
rect 16724 271995 16756 271996
rect 16724 271965 16725 271995
rect 16725 271965 16755 271995
rect 16755 271965 16756 271995
rect 16724 271964 16756 271965
rect 16724 271915 16756 271916
rect 16724 271885 16725 271915
rect 16725 271885 16755 271915
rect 16755 271885 16756 271915
rect 16724 271884 16756 271885
rect 16724 271835 16756 271836
rect 16724 271805 16725 271835
rect 16725 271805 16755 271835
rect 16755 271805 16756 271835
rect 16724 271804 16756 271805
rect 16724 271755 16756 271756
rect 16724 271725 16725 271755
rect 16725 271725 16755 271755
rect 16755 271725 16756 271755
rect 16724 271724 16756 271725
rect 16724 271675 16756 271676
rect 16724 271645 16725 271675
rect 16725 271645 16755 271675
rect 16755 271645 16756 271675
rect 16724 271644 16756 271645
rect 16724 271595 16756 271596
rect 16724 271565 16725 271595
rect 16725 271565 16755 271595
rect 16755 271565 16756 271595
rect 16724 271564 16756 271565
rect 16724 271515 16756 271516
rect 16724 271485 16725 271515
rect 16725 271485 16755 271515
rect 16755 271485 16756 271515
rect 16724 271484 16756 271485
rect 16724 271435 16756 271436
rect 16724 271405 16725 271435
rect 16725 271405 16755 271435
rect 16755 271405 16756 271435
rect 16724 271404 16756 271405
rect 16724 271355 16756 271356
rect 16724 271325 16725 271355
rect 16725 271325 16755 271355
rect 16755 271325 16756 271355
rect 16724 271324 16756 271325
rect 16724 271275 16756 271276
rect 16724 271245 16725 271275
rect 16725 271245 16755 271275
rect 16755 271245 16756 271275
rect 16724 271244 16756 271245
rect 16724 271195 16756 271196
rect 16724 271165 16725 271195
rect 16725 271165 16755 271195
rect 16755 271165 16756 271195
rect 16724 271164 16756 271165
rect 16724 271115 16756 271116
rect 16724 271085 16725 271115
rect 16725 271085 16755 271115
rect 16755 271085 16756 271115
rect 16724 271084 16756 271085
rect 16724 271035 16756 271036
rect 16724 271005 16725 271035
rect 16725 271005 16755 271035
rect 16755 271005 16756 271035
rect 16724 271004 16756 271005
rect 16724 270955 16756 270956
rect 16724 270925 16725 270955
rect 16725 270925 16755 270955
rect 16755 270925 16756 270955
rect 16724 270924 16756 270925
rect 16724 270875 16756 270876
rect 16724 270845 16725 270875
rect 16725 270845 16755 270875
rect 16755 270845 16756 270875
rect 16724 270844 16756 270845
rect 16724 270795 16756 270796
rect 16724 270765 16725 270795
rect 16725 270765 16755 270795
rect 16755 270765 16756 270795
rect 16724 270764 16756 270765
rect 16724 270715 16756 270716
rect 16724 270685 16725 270715
rect 16725 270685 16755 270715
rect 16755 270685 16756 270715
rect 16724 270684 16756 270685
rect 16724 270635 16756 270636
rect 16724 270605 16725 270635
rect 16725 270605 16755 270635
rect 16755 270605 16756 270635
rect 16724 270604 16756 270605
rect 16724 270555 16756 270556
rect 16724 270525 16725 270555
rect 16725 270525 16755 270555
rect 16755 270525 16756 270555
rect 16724 270524 16756 270525
rect 16724 270475 16756 270476
rect 16724 270445 16725 270475
rect 16725 270445 16755 270475
rect 16755 270445 16756 270475
rect 16724 270444 16756 270445
rect 16724 270395 16756 270396
rect 16724 270365 16725 270395
rect 16725 270365 16755 270395
rect 16755 270365 16756 270395
rect 16724 270364 16756 270365
rect 16724 270315 16756 270316
rect 16724 270285 16725 270315
rect 16725 270285 16755 270315
rect 16755 270285 16756 270315
rect 16724 270284 16756 270285
rect 16724 270235 16756 270236
rect 16724 270205 16725 270235
rect 16725 270205 16755 270235
rect 16755 270205 16756 270235
rect 16724 270204 16756 270205
rect 16724 270155 16756 270156
rect 16724 270125 16725 270155
rect 16725 270125 16755 270155
rect 16755 270125 16756 270155
rect 16724 270124 16756 270125
rect 16724 270075 16756 270076
rect 16724 270045 16725 270075
rect 16725 270045 16755 270075
rect 16755 270045 16756 270075
rect 16724 270044 16756 270045
rect 16724 269995 16756 269996
rect 16724 269965 16725 269995
rect 16725 269965 16755 269995
rect 16755 269965 16756 269995
rect 16724 269964 16756 269965
rect 16724 269915 16756 269916
rect 16724 269885 16725 269915
rect 16725 269885 16755 269915
rect 16755 269885 16756 269915
rect 16724 269884 16756 269885
rect 16724 269835 16756 269836
rect 16724 269805 16725 269835
rect 16725 269805 16755 269835
rect 16755 269805 16756 269835
rect 16724 269804 16756 269805
rect 16724 269755 16756 269756
rect 16724 269725 16725 269755
rect 16725 269725 16755 269755
rect 16755 269725 16756 269755
rect 16724 269724 16756 269725
rect 16724 269675 16756 269676
rect 16724 269645 16725 269675
rect 16725 269645 16755 269675
rect 16755 269645 16756 269675
rect 16724 269644 16756 269645
rect 16724 269595 16756 269596
rect 16724 269565 16725 269595
rect 16725 269565 16755 269595
rect 16755 269565 16756 269595
rect 16724 269564 16756 269565
rect 16724 269515 16756 269516
rect 16724 269485 16725 269515
rect 16725 269485 16755 269515
rect 16755 269485 16756 269515
rect 16724 269484 16756 269485
rect 16724 269435 16756 269436
rect 16724 269405 16725 269435
rect 16725 269405 16755 269435
rect 16755 269405 16756 269435
rect 16724 269404 16756 269405
rect 16724 269355 16756 269356
rect 16724 269325 16725 269355
rect 16725 269325 16755 269355
rect 16755 269325 16756 269355
rect 16724 269324 16756 269325
rect 16724 269275 16756 269276
rect 16724 269245 16725 269275
rect 16725 269245 16755 269275
rect 16755 269245 16756 269275
rect 16724 269244 16756 269245
rect 16724 269195 16756 269196
rect 16724 269165 16725 269195
rect 16725 269165 16755 269195
rect 16755 269165 16756 269195
rect 16724 269164 16756 269165
rect 16724 269115 16756 269116
rect 16724 269085 16725 269115
rect 16725 269085 16755 269115
rect 16755 269085 16756 269115
rect 16724 269084 16756 269085
rect 16724 269035 16756 269036
rect 16724 269005 16725 269035
rect 16725 269005 16755 269035
rect 16755 269005 16756 269035
rect 16724 269004 16756 269005
rect 16724 268955 16756 268956
rect 16724 268925 16725 268955
rect 16725 268925 16755 268955
rect 16755 268925 16756 268955
rect 16724 268924 16756 268925
rect 16724 268875 16756 268876
rect 16724 268845 16725 268875
rect 16725 268845 16755 268875
rect 16755 268845 16756 268875
rect 16724 268844 16756 268845
rect 16724 268795 16756 268796
rect 16724 268765 16725 268795
rect 16725 268765 16755 268795
rect 16755 268765 16756 268795
rect 16724 268764 16756 268765
rect 16724 268715 16756 268716
rect 16724 268685 16725 268715
rect 16725 268685 16755 268715
rect 16755 268685 16756 268715
rect 16724 268684 16756 268685
rect 16724 268635 16756 268636
rect 16724 268605 16725 268635
rect 16725 268605 16755 268635
rect 16755 268605 16756 268635
rect 16724 268604 16756 268605
rect 16724 268555 16756 268556
rect 16724 268525 16725 268555
rect 16725 268525 16755 268555
rect 16755 268525 16756 268555
rect 16724 268524 16756 268525
rect 16724 268475 16756 268476
rect 16724 268445 16725 268475
rect 16725 268445 16755 268475
rect 16755 268445 16756 268475
rect 16724 268444 16756 268445
rect 16724 268395 16756 268396
rect 16724 268365 16725 268395
rect 16725 268365 16755 268395
rect 16755 268365 16756 268395
rect 16724 268364 16756 268365
rect 16724 268315 16756 268316
rect 16724 268285 16725 268315
rect 16725 268285 16755 268315
rect 16755 268285 16756 268315
rect 16724 268284 16756 268285
rect 16724 268235 16756 268236
rect 16724 268205 16725 268235
rect 16725 268205 16755 268235
rect 16755 268205 16756 268235
rect 16724 268204 16756 268205
rect 16724 268155 16756 268156
rect 16724 268125 16725 268155
rect 16725 268125 16755 268155
rect 16755 268125 16756 268155
rect 16724 268124 16756 268125
rect 16724 268075 16756 268076
rect 16724 268045 16725 268075
rect 16725 268045 16755 268075
rect 16755 268045 16756 268075
rect 16724 268044 16756 268045
rect 16724 267995 16756 267996
rect 16724 267965 16725 267995
rect 16725 267965 16755 267995
rect 16755 267965 16756 267995
rect 16724 267964 16756 267965
rect 16724 267915 16756 267916
rect 16724 267885 16725 267915
rect 16725 267885 16755 267915
rect 16755 267885 16756 267915
rect 16724 267884 16756 267885
rect 16724 267835 16756 267836
rect 16724 267805 16725 267835
rect 16725 267805 16755 267835
rect 16755 267805 16756 267835
rect 16724 267804 16756 267805
rect 16724 267755 16756 267756
rect 16724 267725 16725 267755
rect 16725 267725 16755 267755
rect 16755 267725 16756 267755
rect 16724 267724 16756 267725
rect 16724 267675 16756 267676
rect 16724 267645 16725 267675
rect 16725 267645 16755 267675
rect 16755 267645 16756 267675
rect 16724 267644 16756 267645
rect 16724 267595 16756 267596
rect 16724 267565 16725 267595
rect 16725 267565 16755 267595
rect 16755 267565 16756 267595
rect 16724 267564 16756 267565
rect 16724 267515 16756 267516
rect 16724 267485 16725 267515
rect 16725 267485 16755 267515
rect 16755 267485 16756 267515
rect 16724 267484 16756 267485
rect 16724 267435 16756 267436
rect 16724 267405 16725 267435
rect 16725 267405 16755 267435
rect 16755 267405 16756 267435
rect 16724 267404 16756 267405
rect 16724 267355 16756 267356
rect 16724 267325 16725 267355
rect 16725 267325 16755 267355
rect 16755 267325 16756 267355
rect 16724 267324 16756 267325
rect 16724 267275 16756 267276
rect 16724 267245 16725 267275
rect 16725 267245 16755 267275
rect 16755 267245 16756 267275
rect 16724 267244 16756 267245
rect 16724 267195 16756 267196
rect 16724 267165 16725 267195
rect 16725 267165 16755 267195
rect 16755 267165 16756 267195
rect 16724 267164 16756 267165
rect 16724 267115 16756 267116
rect 16724 267085 16725 267115
rect 16725 267085 16755 267115
rect 16755 267085 16756 267115
rect 16724 267084 16756 267085
rect 16724 267035 16756 267036
rect 16724 267005 16725 267035
rect 16725 267005 16755 267035
rect 16755 267005 16756 267035
rect 16724 267004 16756 267005
rect 16724 266955 16756 266956
rect 16724 266925 16725 266955
rect 16725 266925 16755 266955
rect 16755 266925 16756 266955
rect 16724 266924 16756 266925
rect 16724 266875 16756 266876
rect 16724 266845 16725 266875
rect 16725 266845 16755 266875
rect 16755 266845 16756 266875
rect 16724 266844 16756 266845
rect 16724 266795 16756 266796
rect 16724 266765 16725 266795
rect 16725 266765 16755 266795
rect 16755 266765 16756 266795
rect 16724 266764 16756 266765
rect 16724 266715 16756 266716
rect 16724 266685 16725 266715
rect 16725 266685 16755 266715
rect 16755 266685 16756 266715
rect 16724 266684 16756 266685
rect 16724 266635 16756 266636
rect 16724 266605 16725 266635
rect 16725 266605 16755 266635
rect 16755 266605 16756 266635
rect 16724 266604 16756 266605
rect 16724 266555 16756 266556
rect 16724 266525 16725 266555
rect 16725 266525 16755 266555
rect 16755 266525 16756 266555
rect 16724 266524 16756 266525
rect 16724 266475 16756 266476
rect 16724 266445 16725 266475
rect 16725 266445 16755 266475
rect 16755 266445 16756 266475
rect 16724 266444 16756 266445
rect 16724 266395 16756 266396
rect 16724 266365 16725 266395
rect 16725 266365 16755 266395
rect 16755 266365 16756 266395
rect 16724 266364 16756 266365
rect 16724 266315 16756 266316
rect 16724 266285 16725 266315
rect 16725 266285 16755 266315
rect 16755 266285 16756 266315
rect 16724 266284 16756 266285
rect 16724 266235 16756 266236
rect 16724 266205 16725 266235
rect 16725 266205 16755 266235
rect 16755 266205 16756 266235
rect 16724 266204 16756 266205
rect 16724 266155 16756 266156
rect 16724 266125 16725 266155
rect 16725 266125 16755 266155
rect 16755 266125 16756 266155
rect 16724 266124 16756 266125
rect 16724 266075 16756 266076
rect 16724 266045 16725 266075
rect 16725 266045 16755 266075
rect 16755 266045 16756 266075
rect 16724 266044 16756 266045
rect 16724 265995 16756 265996
rect 16724 265965 16725 265995
rect 16725 265965 16755 265995
rect 16755 265965 16756 265995
rect 16724 265964 16756 265965
rect 16724 265915 16756 265916
rect 16724 265885 16725 265915
rect 16725 265885 16755 265915
rect 16755 265885 16756 265915
rect 16724 265884 16756 265885
rect 16724 265835 16756 265836
rect 16724 265805 16725 265835
rect 16725 265805 16755 265835
rect 16755 265805 16756 265835
rect 16724 265804 16756 265805
rect 16724 265755 16756 265756
rect 16724 265725 16725 265755
rect 16725 265725 16755 265755
rect 16755 265725 16756 265755
rect 16724 265724 16756 265725
rect 16724 265675 16756 265676
rect 16724 265645 16725 265675
rect 16725 265645 16755 265675
rect 16755 265645 16756 265675
rect 16724 265644 16756 265645
rect 16724 265595 16756 265596
rect 16724 265565 16725 265595
rect 16725 265565 16755 265595
rect 16755 265565 16756 265595
rect 16724 265564 16756 265565
rect 16724 265515 16756 265516
rect 16724 265485 16725 265515
rect 16725 265485 16755 265515
rect 16755 265485 16756 265515
rect 16724 265484 16756 265485
rect 16724 265435 16756 265436
rect 16724 265405 16725 265435
rect 16725 265405 16755 265435
rect 16755 265405 16756 265435
rect 16724 265404 16756 265405
rect 16724 265355 16756 265356
rect 16724 265325 16725 265355
rect 16725 265325 16755 265355
rect 16755 265325 16756 265355
rect 16724 265324 16756 265325
rect 16724 265275 16756 265276
rect 16724 265245 16725 265275
rect 16725 265245 16755 265275
rect 16755 265245 16756 265275
rect 16724 265244 16756 265245
rect 16724 265195 16756 265196
rect 16724 265165 16725 265195
rect 16725 265165 16755 265195
rect 16755 265165 16756 265195
rect 16724 265164 16756 265165
rect 16724 265115 16756 265116
rect 16724 265085 16725 265115
rect 16725 265085 16755 265115
rect 16755 265085 16756 265115
rect 16724 265084 16756 265085
rect 16724 265035 16756 265036
rect 16724 265005 16725 265035
rect 16725 265005 16755 265035
rect 16755 265005 16756 265035
rect 16724 265004 16756 265005
rect 16724 264955 16756 264956
rect 16724 264925 16725 264955
rect 16725 264925 16755 264955
rect 16755 264925 16756 264955
rect 16724 264924 16756 264925
rect 16724 264875 16756 264876
rect 16724 264845 16725 264875
rect 16725 264845 16755 264875
rect 16755 264845 16756 264875
rect 16724 264844 16756 264845
rect 16724 264795 16756 264796
rect 16724 264765 16725 264795
rect 16725 264765 16755 264795
rect 16755 264765 16756 264795
rect 16724 264764 16756 264765
rect 16724 264715 16756 264716
rect 16724 264685 16725 264715
rect 16725 264685 16755 264715
rect 16755 264685 16756 264715
rect 16724 264684 16756 264685
rect 16724 264635 16756 264636
rect 16724 264605 16725 264635
rect 16725 264605 16755 264635
rect 16755 264605 16756 264635
rect 16724 264604 16756 264605
rect 16724 264555 16756 264556
rect 16724 264525 16725 264555
rect 16725 264525 16755 264555
rect 16755 264525 16756 264555
rect 16724 264524 16756 264525
rect 16724 264475 16756 264476
rect 16724 264445 16725 264475
rect 16725 264445 16755 264475
rect 16755 264445 16756 264475
rect 16724 264444 16756 264445
rect 16724 264395 16756 264396
rect 16724 264365 16725 264395
rect 16725 264365 16755 264395
rect 16755 264365 16756 264395
rect 16724 264364 16756 264365
rect 16724 264315 16756 264316
rect 16724 264285 16725 264315
rect 16725 264285 16755 264315
rect 16755 264285 16756 264315
rect 16724 264284 16756 264285
rect 16724 264235 16756 264236
rect 16724 264205 16725 264235
rect 16725 264205 16755 264235
rect 16755 264205 16756 264235
rect 16724 264204 16756 264205
rect 16724 264155 16756 264156
rect 16724 264125 16725 264155
rect 16725 264125 16755 264155
rect 16755 264125 16756 264155
rect 16724 264124 16756 264125
rect 16724 264075 16756 264076
rect 16724 264045 16725 264075
rect 16725 264045 16755 264075
rect 16755 264045 16756 264075
rect 16724 264044 16756 264045
rect 16724 263995 16756 263996
rect 16724 263965 16725 263995
rect 16725 263965 16755 263995
rect 16755 263965 16756 263995
rect 16724 263964 16756 263965
rect 16724 263915 16756 263916
rect 16724 263885 16725 263915
rect 16725 263885 16755 263915
rect 16755 263885 16756 263915
rect 16724 263884 16756 263885
rect 16724 263835 16756 263836
rect 16724 263805 16725 263835
rect 16725 263805 16755 263835
rect 16755 263805 16756 263835
rect 16724 263804 16756 263805
rect 16724 263755 16756 263756
rect 16724 263725 16725 263755
rect 16725 263725 16755 263755
rect 16755 263725 16756 263755
rect 16724 263724 16756 263725
rect 16724 263675 16756 263676
rect 16724 263645 16725 263675
rect 16725 263645 16755 263675
rect 16755 263645 16756 263675
rect 16724 263644 16756 263645
rect 16724 263595 16756 263596
rect 16724 263565 16725 263595
rect 16725 263565 16755 263595
rect 16755 263565 16756 263595
rect 16724 263564 16756 263565
rect 16724 263515 16756 263516
rect 16724 263485 16725 263515
rect 16725 263485 16755 263515
rect 16755 263485 16756 263515
rect 16724 263484 16756 263485
rect 16724 263435 16756 263436
rect 16724 263405 16725 263435
rect 16725 263405 16755 263435
rect 16755 263405 16756 263435
rect 16724 263404 16756 263405
rect 16724 263355 16756 263356
rect 16724 263325 16725 263355
rect 16725 263325 16755 263355
rect 16755 263325 16756 263355
rect 16724 263324 16756 263325
rect 404 255875 436 255876
rect 404 255845 405 255875
rect 405 255845 435 255875
rect 435 255845 436 255875
rect 404 255844 436 255845
rect 404 255764 436 255796
rect 404 255715 436 255716
rect 404 255685 405 255715
rect 405 255685 435 255715
rect 435 255685 436 255715
rect 404 255684 436 255685
rect 484 255875 516 255876
rect 484 255845 485 255875
rect 485 255845 515 255875
rect 515 255845 516 255875
rect 484 255844 516 255845
rect 484 255764 516 255796
rect 484 255715 516 255716
rect 484 255685 485 255715
rect 485 255685 515 255715
rect 515 255685 516 255715
rect 484 255684 516 255685
rect 564 255875 596 255876
rect 564 255845 565 255875
rect 565 255845 595 255875
rect 595 255845 596 255875
rect 564 255844 596 255845
rect 564 255764 596 255796
rect 564 255715 596 255716
rect 564 255685 565 255715
rect 565 255685 595 255715
rect 595 255685 596 255715
rect 564 255684 596 255685
rect 644 255875 676 255876
rect 644 255845 645 255875
rect 645 255845 675 255875
rect 675 255845 676 255875
rect 644 255844 676 255845
rect 644 255764 676 255796
rect 644 255715 676 255716
rect 644 255685 645 255715
rect 645 255685 675 255715
rect 675 255685 676 255715
rect 644 255684 676 255685
rect 724 255875 756 255876
rect 724 255845 725 255875
rect 725 255845 755 255875
rect 755 255845 756 255875
rect 724 255844 756 255845
rect 724 255764 756 255796
rect 724 255715 756 255716
rect 724 255685 725 255715
rect 725 255685 755 255715
rect 755 255685 756 255715
rect 724 255684 756 255685
rect 804 255875 836 255876
rect 804 255845 805 255875
rect 805 255845 835 255875
rect 835 255845 836 255875
rect 804 255844 836 255845
rect 804 255764 836 255796
rect 804 255715 836 255716
rect 804 255685 805 255715
rect 805 255685 835 255715
rect 835 255685 836 255715
rect 804 255684 836 255685
rect 884 255875 916 255876
rect 884 255845 885 255875
rect 885 255845 915 255875
rect 915 255845 916 255875
rect 884 255844 916 255845
rect 884 255764 916 255796
rect 884 255715 916 255716
rect 884 255685 885 255715
rect 885 255685 915 255715
rect 915 255685 916 255715
rect 884 255684 916 255685
rect 964 255875 996 255876
rect 964 255845 965 255875
rect 965 255845 995 255875
rect 995 255845 996 255875
rect 964 255844 996 255845
rect 964 255764 996 255796
rect 964 255715 996 255716
rect 964 255685 965 255715
rect 965 255685 995 255715
rect 995 255685 996 255715
rect 964 255684 996 255685
rect 1044 255875 1076 255876
rect 1044 255845 1045 255875
rect 1045 255845 1075 255875
rect 1075 255845 1076 255875
rect 1044 255844 1076 255845
rect 1044 255764 1076 255796
rect 1044 255715 1076 255716
rect 1044 255685 1045 255715
rect 1045 255685 1075 255715
rect 1075 255685 1076 255715
rect 1044 255684 1076 255685
rect 1124 255875 1156 255876
rect 1124 255845 1125 255875
rect 1125 255845 1155 255875
rect 1155 255845 1156 255875
rect 1124 255844 1156 255845
rect 1124 255764 1156 255796
rect 1124 255715 1156 255716
rect 1124 255685 1125 255715
rect 1125 255685 1155 255715
rect 1155 255685 1156 255715
rect 1124 255684 1156 255685
rect 1204 255875 1236 255876
rect 1204 255845 1205 255875
rect 1205 255845 1235 255875
rect 1235 255845 1236 255875
rect 1204 255844 1236 255845
rect 1204 255764 1236 255796
rect 1204 255715 1236 255716
rect 1204 255685 1205 255715
rect 1205 255685 1235 255715
rect 1235 255685 1236 255715
rect 1204 255684 1236 255685
rect 1284 255875 1316 255876
rect 1284 255845 1285 255875
rect 1285 255845 1315 255875
rect 1315 255845 1316 255875
rect 1284 255844 1316 255845
rect 1284 255764 1316 255796
rect 1284 255715 1316 255716
rect 1284 255685 1285 255715
rect 1285 255685 1315 255715
rect 1315 255685 1316 255715
rect 1284 255684 1316 255685
rect 1364 255875 1396 255876
rect 1364 255845 1365 255875
rect 1365 255845 1395 255875
rect 1395 255845 1396 255875
rect 1364 255844 1396 255845
rect 1364 255764 1396 255796
rect 1364 255715 1396 255716
rect 1364 255685 1365 255715
rect 1365 255685 1395 255715
rect 1395 255685 1396 255715
rect 1364 255684 1396 255685
rect 1444 255875 1476 255876
rect 1444 255845 1445 255875
rect 1445 255845 1475 255875
rect 1475 255845 1476 255875
rect 1444 255844 1476 255845
rect 1444 255764 1476 255796
rect 1444 255715 1476 255716
rect 1444 255685 1445 255715
rect 1445 255685 1475 255715
rect 1475 255685 1476 255715
rect 1444 255684 1476 255685
rect 1524 255875 1556 255876
rect 1524 255845 1525 255875
rect 1525 255845 1555 255875
rect 1555 255845 1556 255875
rect 1524 255844 1556 255845
rect 1524 255764 1556 255796
rect 1524 255715 1556 255716
rect 1524 255685 1525 255715
rect 1525 255685 1555 255715
rect 1555 255685 1556 255715
rect 1524 255684 1556 255685
rect 1604 255875 1636 255876
rect 1604 255845 1605 255875
rect 1605 255845 1635 255875
rect 1635 255845 1636 255875
rect 1604 255844 1636 255845
rect 1604 255764 1636 255796
rect 1604 255715 1636 255716
rect 1604 255685 1605 255715
rect 1605 255685 1635 255715
rect 1635 255685 1636 255715
rect 1604 255684 1636 255685
rect 1684 255875 1716 255876
rect 1684 255845 1685 255875
rect 1685 255845 1715 255875
rect 1715 255845 1716 255875
rect 1684 255844 1716 255845
rect 1684 255764 1716 255796
rect 1684 255715 1716 255716
rect 1684 255685 1685 255715
rect 1685 255685 1715 255715
rect 1715 255685 1716 255715
rect 1684 255684 1716 255685
rect 1764 255875 1796 255876
rect 1764 255845 1765 255875
rect 1765 255845 1795 255875
rect 1795 255845 1796 255875
rect 1764 255844 1796 255845
rect 1764 255764 1796 255796
rect 1764 255715 1796 255716
rect 1764 255685 1765 255715
rect 1765 255685 1795 255715
rect 1795 255685 1796 255715
rect 1764 255684 1796 255685
rect 1844 255875 1876 255876
rect 1844 255845 1845 255875
rect 1845 255845 1875 255875
rect 1875 255845 1876 255875
rect 1844 255844 1876 255845
rect 1844 255764 1876 255796
rect 1844 255715 1876 255716
rect 1844 255685 1845 255715
rect 1845 255685 1875 255715
rect 1875 255685 1876 255715
rect 1844 255684 1876 255685
rect 1924 255875 1956 255876
rect 1924 255845 1925 255875
rect 1925 255845 1955 255875
rect 1955 255845 1956 255875
rect 1924 255844 1956 255845
rect 1924 255764 1956 255796
rect 1924 255715 1956 255716
rect 1924 255685 1925 255715
rect 1925 255685 1955 255715
rect 1955 255685 1956 255715
rect 1924 255684 1956 255685
rect 2004 255875 2036 255876
rect 2004 255845 2005 255875
rect 2005 255845 2035 255875
rect 2035 255845 2036 255875
rect 2004 255844 2036 255845
rect 2004 255764 2036 255796
rect 2004 255715 2036 255716
rect 2004 255685 2005 255715
rect 2005 255685 2035 255715
rect 2035 255685 2036 255715
rect 2004 255684 2036 255685
rect 2084 255875 2116 255876
rect 2084 255845 2085 255875
rect 2085 255845 2115 255875
rect 2115 255845 2116 255875
rect 2084 255844 2116 255845
rect 2084 255764 2116 255796
rect 2084 255715 2116 255716
rect 2084 255685 2085 255715
rect 2085 255685 2115 255715
rect 2115 255685 2116 255715
rect 2084 255684 2116 255685
rect 2164 255875 2196 255876
rect 2164 255845 2165 255875
rect 2165 255845 2195 255875
rect 2195 255845 2196 255875
rect 2164 255844 2196 255845
rect 2164 255764 2196 255796
rect 2164 255715 2196 255716
rect 2164 255685 2165 255715
rect 2165 255685 2195 255715
rect 2195 255685 2196 255715
rect 2164 255684 2196 255685
rect 2244 255875 2276 255876
rect 2244 255845 2245 255875
rect 2245 255845 2275 255875
rect 2275 255845 2276 255875
rect 2244 255844 2276 255845
rect 2244 255764 2276 255796
rect 2244 255715 2276 255716
rect 2244 255685 2245 255715
rect 2245 255685 2275 255715
rect 2275 255685 2276 255715
rect 2244 255684 2276 255685
rect 2324 255875 2356 255876
rect 2324 255845 2325 255875
rect 2325 255845 2355 255875
rect 2355 255845 2356 255875
rect 2324 255844 2356 255845
rect 2324 255764 2356 255796
rect 2324 255715 2356 255716
rect 2324 255685 2325 255715
rect 2325 255685 2355 255715
rect 2355 255685 2356 255715
rect 2324 255684 2356 255685
rect 2404 255875 2436 255876
rect 2404 255845 2405 255875
rect 2405 255845 2435 255875
rect 2435 255845 2436 255875
rect 2404 255844 2436 255845
rect 2404 255764 2436 255796
rect 2404 255715 2436 255716
rect 2404 255685 2405 255715
rect 2405 255685 2435 255715
rect 2435 255685 2436 255715
rect 2404 255684 2436 255685
rect 2484 255875 2516 255876
rect 2484 255845 2485 255875
rect 2485 255845 2515 255875
rect 2515 255845 2516 255875
rect 2484 255844 2516 255845
rect 2484 255764 2516 255796
rect 2484 255715 2516 255716
rect 2484 255685 2485 255715
rect 2485 255685 2515 255715
rect 2515 255685 2516 255715
rect 2484 255684 2516 255685
rect 2564 255875 2596 255876
rect 2564 255845 2565 255875
rect 2565 255845 2595 255875
rect 2595 255845 2596 255875
rect 2564 255844 2596 255845
rect 2564 255764 2596 255796
rect 2564 255715 2596 255716
rect 2564 255685 2565 255715
rect 2565 255685 2595 255715
rect 2595 255685 2596 255715
rect 2564 255684 2596 255685
rect 2644 255875 2676 255876
rect 2644 255845 2645 255875
rect 2645 255845 2675 255875
rect 2675 255845 2676 255875
rect 2644 255844 2676 255845
rect 2644 255764 2676 255796
rect 2644 255715 2676 255716
rect 2644 255685 2645 255715
rect 2645 255685 2675 255715
rect 2675 255685 2676 255715
rect 2644 255684 2676 255685
rect 2724 255875 2756 255876
rect 2724 255845 2725 255875
rect 2725 255845 2755 255875
rect 2755 255845 2756 255875
rect 2724 255844 2756 255845
rect 2724 255764 2756 255796
rect 2724 255715 2756 255716
rect 2724 255685 2725 255715
rect 2725 255685 2755 255715
rect 2755 255685 2756 255715
rect 2724 255684 2756 255685
rect 16724 263275 16756 263276
rect 16724 263245 16725 263275
rect 16725 263245 16755 263275
rect 16755 263245 16756 263275
rect 16724 263244 16756 263245
rect 16724 263195 16756 263196
rect 16724 263165 16725 263195
rect 16725 263165 16755 263195
rect 16755 263165 16756 263195
rect 16724 263164 16756 263165
rect 16724 263115 16756 263116
rect 16724 263085 16725 263115
rect 16725 263085 16755 263115
rect 16755 263085 16756 263115
rect 16724 263084 16756 263085
rect 16724 263035 16756 263036
rect 16724 263005 16725 263035
rect 16725 263005 16755 263035
rect 16755 263005 16756 263035
rect 16724 263004 16756 263005
rect 16724 262955 16756 262956
rect 16724 262925 16725 262955
rect 16725 262925 16755 262955
rect 16755 262925 16756 262955
rect 16724 262924 16756 262925
rect 16724 262875 16756 262876
rect 16724 262845 16725 262875
rect 16725 262845 16755 262875
rect 16755 262845 16756 262875
rect 16724 262844 16756 262845
rect 16724 262795 16756 262796
rect 16724 262765 16725 262795
rect 16725 262765 16755 262795
rect 16755 262765 16756 262795
rect 16724 262764 16756 262765
rect 16724 262715 16756 262716
rect 16724 262685 16725 262715
rect 16725 262685 16755 262715
rect 16755 262685 16756 262715
rect 16724 262684 16756 262685
rect 16724 262635 16756 262636
rect 16724 262605 16725 262635
rect 16725 262605 16755 262635
rect 16755 262605 16756 262635
rect 16724 262604 16756 262605
rect 16724 262555 16756 262556
rect 16724 262525 16725 262555
rect 16725 262525 16755 262555
rect 16755 262525 16756 262555
rect 16724 262524 16756 262525
rect 16724 262475 16756 262476
rect 16724 262445 16725 262475
rect 16725 262445 16755 262475
rect 16755 262445 16756 262475
rect 16724 262444 16756 262445
rect 16724 262395 16756 262396
rect 16724 262365 16725 262395
rect 16725 262365 16755 262395
rect 16755 262365 16756 262395
rect 16724 262364 16756 262365
rect 16724 262315 16756 262316
rect 16724 262285 16725 262315
rect 16725 262285 16755 262315
rect 16755 262285 16756 262315
rect 16724 262284 16756 262285
rect 16724 262235 16756 262236
rect 16724 262205 16725 262235
rect 16725 262205 16755 262235
rect 16755 262205 16756 262235
rect 16724 262204 16756 262205
rect 16724 262155 16756 262156
rect 16724 262125 16725 262155
rect 16725 262125 16755 262155
rect 16755 262125 16756 262155
rect 16724 262124 16756 262125
rect 16724 262075 16756 262076
rect 16724 262045 16725 262075
rect 16725 262045 16755 262075
rect 16755 262045 16756 262075
rect 16724 262044 16756 262045
rect 16724 261995 16756 261996
rect 16724 261965 16725 261995
rect 16725 261965 16755 261995
rect 16755 261965 16756 261995
rect 16724 261964 16756 261965
rect 16724 261915 16756 261916
rect 16724 261885 16725 261915
rect 16725 261885 16755 261915
rect 16755 261885 16756 261915
rect 16724 261884 16756 261885
rect 16724 261835 16756 261836
rect 16724 261805 16725 261835
rect 16725 261805 16755 261835
rect 16755 261805 16756 261835
rect 16724 261804 16756 261805
rect 16724 261755 16756 261756
rect 16724 261725 16725 261755
rect 16725 261725 16755 261755
rect 16755 261725 16756 261755
rect 16724 261724 16756 261725
rect 16724 261675 16756 261676
rect 16724 261645 16725 261675
rect 16725 261645 16755 261675
rect 16755 261645 16756 261675
rect 16724 261644 16756 261645
rect 16724 261595 16756 261596
rect 16724 261565 16725 261595
rect 16725 261565 16755 261595
rect 16755 261565 16756 261595
rect 16724 261564 16756 261565
rect 16724 261515 16756 261516
rect 16724 261485 16725 261515
rect 16725 261485 16755 261515
rect 16755 261485 16756 261515
rect 16724 261484 16756 261485
rect 16724 261435 16756 261436
rect 16724 261405 16725 261435
rect 16725 261405 16755 261435
rect 16755 261405 16756 261435
rect 16724 261404 16756 261405
rect 16724 261355 16756 261356
rect 16724 261325 16725 261355
rect 16725 261325 16755 261355
rect 16755 261325 16756 261355
rect 16724 261324 16756 261325
rect 16724 261275 16756 261276
rect 16724 261245 16725 261275
rect 16725 261245 16755 261275
rect 16755 261245 16756 261275
rect 16724 261244 16756 261245
rect 16724 261195 16756 261196
rect 16724 261165 16725 261195
rect 16725 261165 16755 261195
rect 16755 261165 16756 261195
rect 16724 261164 16756 261165
rect 16724 261115 16756 261116
rect 16724 261085 16725 261115
rect 16725 261085 16755 261115
rect 16755 261085 16756 261115
rect 16724 261084 16756 261085
rect 16724 261035 16756 261036
rect 16724 261005 16725 261035
rect 16725 261005 16755 261035
rect 16755 261005 16756 261035
rect 16724 261004 16756 261005
rect 16724 260955 16756 260956
rect 16724 260925 16725 260955
rect 16725 260925 16755 260955
rect 16755 260925 16756 260955
rect 16724 260924 16756 260925
rect 16724 260875 16756 260876
rect 16724 260845 16725 260875
rect 16725 260845 16755 260875
rect 16755 260845 16756 260875
rect 16724 260844 16756 260845
rect 16724 260795 16756 260796
rect 16724 260765 16725 260795
rect 16725 260765 16755 260795
rect 16755 260765 16756 260795
rect 16724 260764 16756 260765
rect 16724 260715 16756 260716
rect 16724 260685 16725 260715
rect 16725 260685 16755 260715
rect 16755 260685 16756 260715
rect 16724 260684 16756 260685
rect 16724 260635 16756 260636
rect 16724 260605 16725 260635
rect 16725 260605 16755 260635
rect 16755 260605 16756 260635
rect 16724 260604 16756 260605
rect 16724 260555 16756 260556
rect 16724 260525 16725 260555
rect 16725 260525 16755 260555
rect 16755 260525 16756 260555
rect 16724 260524 16756 260525
rect 16724 260475 16756 260476
rect 16724 260445 16725 260475
rect 16725 260445 16755 260475
rect 16755 260445 16756 260475
rect 16724 260444 16756 260445
rect 16724 260395 16756 260396
rect 16724 260365 16725 260395
rect 16725 260365 16755 260395
rect 16755 260365 16756 260395
rect 16724 260364 16756 260365
rect 16724 260315 16756 260316
rect 16724 260285 16725 260315
rect 16725 260285 16755 260315
rect 16755 260285 16756 260315
rect 16724 260284 16756 260285
rect 16724 260235 16756 260236
rect 16724 260205 16725 260235
rect 16725 260205 16755 260235
rect 16755 260205 16756 260235
rect 16724 260204 16756 260205
rect 16724 260155 16756 260156
rect 16724 260125 16725 260155
rect 16725 260125 16755 260155
rect 16755 260125 16756 260155
rect 16724 260124 16756 260125
rect 16724 260075 16756 260076
rect 16724 260045 16725 260075
rect 16725 260045 16755 260075
rect 16755 260045 16756 260075
rect 16724 260044 16756 260045
rect 16724 259995 16756 259996
rect 16724 259965 16725 259995
rect 16725 259965 16755 259995
rect 16755 259965 16756 259995
rect 16724 259964 16756 259965
rect 16724 259915 16756 259916
rect 16724 259885 16725 259915
rect 16725 259885 16755 259915
rect 16755 259885 16756 259915
rect 16724 259884 16756 259885
rect 16724 259835 16756 259836
rect 16724 259805 16725 259835
rect 16725 259805 16755 259835
rect 16755 259805 16756 259835
rect 16724 259804 16756 259805
rect 16724 259755 16756 259756
rect 16724 259725 16725 259755
rect 16725 259725 16755 259755
rect 16755 259725 16756 259755
rect 16724 259724 16756 259725
rect 16724 259675 16756 259676
rect 16724 259645 16725 259675
rect 16725 259645 16755 259675
rect 16755 259645 16756 259675
rect 16724 259644 16756 259645
rect 16724 259595 16756 259596
rect 16724 259565 16725 259595
rect 16725 259565 16755 259595
rect 16755 259565 16756 259595
rect 16724 259564 16756 259565
rect 16724 259515 16756 259516
rect 16724 259485 16725 259515
rect 16725 259485 16755 259515
rect 16755 259485 16756 259515
rect 16724 259484 16756 259485
rect 16724 259435 16756 259436
rect 16724 259405 16725 259435
rect 16725 259405 16755 259435
rect 16755 259405 16756 259435
rect 16724 259404 16756 259405
rect 16724 259355 16756 259356
rect 16724 259325 16725 259355
rect 16725 259325 16755 259355
rect 16755 259325 16756 259355
rect 16724 259324 16756 259325
rect 16724 259275 16756 259276
rect 16724 259245 16725 259275
rect 16725 259245 16755 259275
rect 16755 259245 16756 259275
rect 16724 259244 16756 259245
rect 16724 259195 16756 259196
rect 16724 259165 16725 259195
rect 16725 259165 16755 259195
rect 16755 259165 16756 259195
rect 16724 259164 16756 259165
rect 16724 259115 16756 259116
rect 16724 259085 16725 259115
rect 16725 259085 16755 259115
rect 16755 259085 16756 259115
rect 16724 259084 16756 259085
rect 16724 259035 16756 259036
rect 16724 259005 16725 259035
rect 16725 259005 16755 259035
rect 16755 259005 16756 259035
rect 16724 259004 16756 259005
rect 16724 258955 16756 258956
rect 16724 258925 16725 258955
rect 16725 258925 16755 258955
rect 16755 258925 16756 258955
rect 16724 258924 16756 258925
rect 16724 258875 16756 258876
rect 16724 258845 16725 258875
rect 16725 258845 16755 258875
rect 16755 258845 16756 258875
rect 16724 258844 16756 258845
rect 16724 258795 16756 258796
rect 16724 258765 16725 258795
rect 16725 258765 16755 258795
rect 16755 258765 16756 258795
rect 16724 258764 16756 258765
rect 16724 258715 16756 258716
rect 16724 258685 16725 258715
rect 16725 258685 16755 258715
rect 16755 258685 16756 258715
rect 16724 258684 16756 258685
rect 16724 258635 16756 258636
rect 16724 258605 16725 258635
rect 16725 258605 16755 258635
rect 16755 258605 16756 258635
rect 16724 258604 16756 258605
rect 16724 258555 16756 258556
rect 16724 258525 16725 258555
rect 16725 258525 16755 258555
rect 16755 258525 16756 258555
rect 16724 258524 16756 258525
rect 16724 258475 16756 258476
rect 16724 258445 16725 258475
rect 16725 258445 16755 258475
rect 16755 258445 16756 258475
rect 16724 258444 16756 258445
rect 16724 258395 16756 258396
rect 16724 258365 16725 258395
rect 16725 258365 16755 258395
rect 16755 258365 16756 258395
rect 16724 258364 16756 258365
rect 16724 258315 16756 258316
rect 16724 258285 16725 258315
rect 16725 258285 16755 258315
rect 16755 258285 16756 258315
rect 16724 258284 16756 258285
rect 16724 258235 16756 258236
rect 16724 258205 16725 258235
rect 16725 258205 16755 258235
rect 16755 258205 16756 258235
rect 16724 258204 16756 258205
rect 16724 258155 16756 258156
rect 16724 258125 16725 258155
rect 16725 258125 16755 258155
rect 16755 258125 16756 258155
rect 16724 258124 16756 258125
rect 16724 258075 16756 258076
rect 16724 258045 16725 258075
rect 16725 258045 16755 258075
rect 16755 258045 16756 258075
rect 16724 258044 16756 258045
rect 16724 257995 16756 257996
rect 16724 257965 16725 257995
rect 16725 257965 16755 257995
rect 16755 257965 16756 257995
rect 16724 257964 16756 257965
rect 16724 257915 16756 257916
rect 16724 257885 16725 257915
rect 16725 257885 16755 257915
rect 16755 257885 16756 257915
rect 16724 257884 16756 257885
rect 16724 257835 16756 257836
rect 16724 257805 16725 257835
rect 16725 257805 16755 257835
rect 16755 257805 16756 257835
rect 16724 257804 16756 257805
rect 16724 257755 16756 257756
rect 16724 257725 16725 257755
rect 16725 257725 16755 257755
rect 16755 257725 16756 257755
rect 16724 257724 16756 257725
rect 16724 257675 16756 257676
rect 16724 257645 16725 257675
rect 16725 257645 16755 257675
rect 16755 257645 16756 257675
rect 16724 257644 16756 257645
rect 16724 257595 16756 257596
rect 16724 257565 16725 257595
rect 16725 257565 16755 257595
rect 16755 257565 16756 257595
rect 16724 257564 16756 257565
rect 16724 257515 16756 257516
rect 16724 257485 16725 257515
rect 16725 257485 16755 257515
rect 16755 257485 16756 257515
rect 16724 257484 16756 257485
rect 16724 257435 16756 257436
rect 16724 257405 16725 257435
rect 16725 257405 16755 257435
rect 16755 257405 16756 257435
rect 16724 257404 16756 257405
rect 16724 257355 16756 257356
rect 16724 257325 16725 257355
rect 16725 257325 16755 257355
rect 16755 257325 16756 257355
rect 16724 257324 16756 257325
rect 16724 257275 16756 257276
rect 16724 257245 16725 257275
rect 16725 257245 16755 257275
rect 16755 257245 16756 257275
rect 16724 257244 16756 257245
rect 16724 257195 16756 257196
rect 16724 257165 16725 257195
rect 16725 257165 16755 257195
rect 16755 257165 16756 257195
rect 16724 257164 16756 257165
rect 16724 257115 16756 257116
rect 16724 257085 16725 257115
rect 16725 257085 16755 257115
rect 16755 257085 16756 257115
rect 16724 257084 16756 257085
rect 16724 257035 16756 257036
rect 16724 257005 16725 257035
rect 16725 257005 16755 257035
rect 16755 257005 16756 257035
rect 16724 257004 16756 257005
rect 16724 256955 16756 256956
rect 16724 256925 16725 256955
rect 16725 256925 16755 256955
rect 16755 256925 16756 256955
rect 16724 256924 16756 256925
rect 16724 256875 16756 256876
rect 16724 256845 16725 256875
rect 16725 256845 16755 256875
rect 16755 256845 16756 256875
rect 16724 256844 16756 256845
rect 16724 256795 16756 256796
rect 16724 256765 16725 256795
rect 16725 256765 16755 256795
rect 16755 256765 16756 256795
rect 16724 256764 16756 256765
rect 16724 256715 16756 256716
rect 16724 256685 16725 256715
rect 16725 256685 16755 256715
rect 16755 256685 16756 256715
rect 16724 256684 16756 256685
rect 16724 256635 16756 256636
rect 16724 256605 16725 256635
rect 16725 256605 16755 256635
rect 16755 256605 16756 256635
rect 16724 256604 16756 256605
rect 16724 256555 16756 256556
rect 16724 256525 16725 256555
rect 16725 256525 16755 256555
rect 16755 256525 16756 256555
rect 16724 256524 16756 256525
rect 16724 256475 16756 256476
rect 16724 256445 16725 256475
rect 16725 256445 16755 256475
rect 16755 256445 16756 256475
rect 16724 256444 16756 256445
rect 16724 256395 16756 256396
rect 16724 256365 16725 256395
rect 16725 256365 16755 256395
rect 16755 256365 16756 256395
rect 16724 256364 16756 256365
rect 16724 256315 16756 256316
rect 16724 256285 16725 256315
rect 16725 256285 16755 256315
rect 16755 256285 16756 256315
rect 16724 256284 16756 256285
rect 16724 256235 16756 256236
rect 16724 256205 16725 256235
rect 16725 256205 16755 256235
rect 16755 256205 16756 256235
rect 16724 256204 16756 256205
rect 16724 256155 16756 256156
rect 16724 256125 16725 256155
rect 16725 256125 16755 256155
rect 16755 256125 16756 256155
rect 16724 256124 16756 256125
rect 16724 256075 16756 256076
rect 16724 256045 16725 256075
rect 16725 256045 16755 256075
rect 16755 256045 16756 256075
rect 16724 256044 16756 256045
rect 16724 255995 16756 255996
rect 16724 255965 16725 255995
rect 16725 255965 16755 255995
rect 16755 255965 16756 255995
rect 16724 255964 16756 255965
rect 3044 255875 3076 255876
rect 3044 255845 3045 255875
rect 3045 255845 3075 255875
rect 3075 255845 3076 255875
rect 3044 255844 3076 255845
rect 3044 255764 3076 255796
rect 3044 255715 3076 255716
rect 3044 255685 3045 255715
rect 3045 255685 3075 255715
rect 3075 255685 3076 255715
rect 3044 255684 3076 255685
rect 3124 255875 3156 255876
rect 3124 255845 3125 255875
rect 3125 255845 3155 255875
rect 3155 255845 3156 255875
rect 3124 255844 3156 255845
rect 3124 255764 3156 255796
rect 3124 255715 3156 255716
rect 3124 255685 3125 255715
rect 3125 255685 3155 255715
rect 3155 255685 3156 255715
rect 3124 255684 3156 255685
rect 3204 255875 3236 255876
rect 3204 255845 3205 255875
rect 3205 255845 3235 255875
rect 3235 255845 3236 255875
rect 3204 255844 3236 255845
rect 3204 255764 3236 255796
rect 3204 255715 3236 255716
rect 3204 255685 3205 255715
rect 3205 255685 3235 255715
rect 3235 255685 3236 255715
rect 3204 255684 3236 255685
rect 3284 255875 3316 255876
rect 3284 255845 3285 255875
rect 3285 255845 3315 255875
rect 3315 255845 3316 255875
rect 3284 255844 3316 255845
rect 3284 255764 3316 255796
rect 3284 255715 3316 255716
rect 3284 255685 3285 255715
rect 3285 255685 3315 255715
rect 3315 255685 3316 255715
rect 3284 255684 3316 255685
rect 3364 255875 3396 255876
rect 3364 255845 3365 255875
rect 3365 255845 3395 255875
rect 3395 255845 3396 255875
rect 3364 255844 3396 255845
rect 3364 255764 3396 255796
rect 3364 255715 3396 255716
rect 3364 255685 3365 255715
rect 3365 255685 3395 255715
rect 3395 255685 3396 255715
rect 3364 255684 3396 255685
rect 3444 255875 3476 255876
rect 3444 255845 3445 255875
rect 3445 255845 3475 255875
rect 3475 255845 3476 255875
rect 3444 255844 3476 255845
rect 3444 255764 3476 255796
rect 3444 255715 3476 255716
rect 3444 255685 3445 255715
rect 3445 255685 3475 255715
rect 3475 255685 3476 255715
rect 3444 255684 3476 255685
rect 3524 255875 3556 255876
rect 3524 255845 3525 255875
rect 3525 255845 3555 255875
rect 3555 255845 3556 255875
rect 3524 255844 3556 255845
rect 3524 255764 3556 255796
rect 3524 255715 3556 255716
rect 3524 255685 3525 255715
rect 3525 255685 3555 255715
rect 3555 255685 3556 255715
rect 3524 255684 3556 255685
rect 3604 255875 3636 255876
rect 3604 255845 3605 255875
rect 3605 255845 3635 255875
rect 3635 255845 3636 255875
rect 3604 255844 3636 255845
rect 3604 255764 3636 255796
rect 3604 255715 3636 255716
rect 3604 255685 3605 255715
rect 3605 255685 3635 255715
rect 3635 255685 3636 255715
rect 3604 255684 3636 255685
rect 3684 255875 3716 255876
rect 3684 255845 3685 255875
rect 3685 255845 3715 255875
rect 3715 255845 3716 255875
rect 3684 255844 3716 255845
rect 3684 255764 3716 255796
rect 3684 255715 3716 255716
rect 3684 255685 3685 255715
rect 3685 255685 3715 255715
rect 3715 255685 3716 255715
rect 3684 255684 3716 255685
rect 3764 255875 3796 255876
rect 3764 255845 3765 255875
rect 3765 255845 3795 255875
rect 3795 255845 3796 255875
rect 3764 255844 3796 255845
rect 3764 255764 3796 255796
rect 3764 255715 3796 255716
rect 3764 255685 3765 255715
rect 3765 255685 3795 255715
rect 3795 255685 3796 255715
rect 3764 255684 3796 255685
rect 3844 255875 3876 255876
rect 3844 255845 3845 255875
rect 3845 255845 3875 255875
rect 3875 255845 3876 255875
rect 3844 255844 3876 255845
rect 3844 255764 3876 255796
rect 3844 255715 3876 255716
rect 3844 255685 3845 255715
rect 3845 255685 3875 255715
rect 3875 255685 3876 255715
rect 3844 255684 3876 255685
rect 3924 255875 3956 255876
rect 3924 255845 3925 255875
rect 3925 255845 3955 255875
rect 3955 255845 3956 255875
rect 3924 255844 3956 255845
rect 3924 255764 3956 255796
rect 3924 255715 3956 255716
rect 3924 255685 3925 255715
rect 3925 255685 3955 255715
rect 3955 255685 3956 255715
rect 3924 255684 3956 255685
rect 4004 255875 4036 255876
rect 4004 255845 4005 255875
rect 4005 255845 4035 255875
rect 4035 255845 4036 255875
rect 4004 255844 4036 255845
rect 4004 255764 4036 255796
rect 4004 255715 4036 255716
rect 4004 255685 4005 255715
rect 4005 255685 4035 255715
rect 4035 255685 4036 255715
rect 4004 255684 4036 255685
rect 4084 255875 4116 255876
rect 4084 255845 4085 255875
rect 4085 255845 4115 255875
rect 4115 255845 4116 255875
rect 4084 255844 4116 255845
rect 4084 255764 4116 255796
rect 4084 255715 4116 255716
rect 4084 255685 4085 255715
rect 4085 255685 4115 255715
rect 4115 255685 4116 255715
rect 4084 255684 4116 255685
rect 4164 255875 4196 255876
rect 4164 255845 4165 255875
rect 4165 255845 4195 255875
rect 4195 255845 4196 255875
rect 4164 255844 4196 255845
rect 4164 255764 4196 255796
rect 4164 255715 4196 255716
rect 4164 255685 4165 255715
rect 4165 255685 4195 255715
rect 4195 255685 4196 255715
rect 4164 255684 4196 255685
rect 4244 255875 4276 255876
rect 4244 255845 4245 255875
rect 4245 255845 4275 255875
rect 4275 255845 4276 255875
rect 4244 255844 4276 255845
rect 4244 255764 4276 255796
rect 4244 255715 4276 255716
rect 4244 255685 4245 255715
rect 4245 255685 4275 255715
rect 4275 255685 4276 255715
rect 4244 255684 4276 255685
rect 4324 255875 4356 255876
rect 4324 255845 4325 255875
rect 4325 255845 4355 255875
rect 4355 255845 4356 255875
rect 4324 255844 4356 255845
rect 4324 255764 4356 255796
rect 4324 255715 4356 255716
rect 4324 255685 4325 255715
rect 4325 255685 4355 255715
rect 4355 255685 4356 255715
rect 4324 255684 4356 255685
rect 4404 255875 4436 255876
rect 4404 255845 4405 255875
rect 4405 255845 4435 255875
rect 4435 255845 4436 255875
rect 4404 255844 4436 255845
rect 4404 255764 4436 255796
rect 4404 255715 4436 255716
rect 4404 255685 4405 255715
rect 4405 255685 4435 255715
rect 4435 255685 4436 255715
rect 4404 255684 4436 255685
rect 4484 255875 4516 255876
rect 4484 255845 4485 255875
rect 4485 255845 4515 255875
rect 4515 255845 4516 255875
rect 4484 255844 4516 255845
rect 4484 255764 4516 255796
rect 4484 255715 4516 255716
rect 4484 255685 4485 255715
rect 4485 255685 4515 255715
rect 4515 255685 4516 255715
rect 4484 255684 4516 255685
rect 4564 255875 4596 255876
rect 4564 255845 4565 255875
rect 4565 255845 4595 255875
rect 4595 255845 4596 255875
rect 4564 255844 4596 255845
rect 4564 255764 4596 255796
rect 4564 255715 4596 255716
rect 4564 255685 4565 255715
rect 4565 255685 4595 255715
rect 4595 255685 4596 255715
rect 4564 255684 4596 255685
rect 4644 255875 4676 255876
rect 4644 255845 4645 255875
rect 4645 255845 4675 255875
rect 4675 255845 4676 255875
rect 4644 255844 4676 255845
rect 4644 255764 4676 255796
rect 4644 255715 4676 255716
rect 4644 255685 4645 255715
rect 4645 255685 4675 255715
rect 4675 255685 4676 255715
rect 4644 255684 4676 255685
rect 4724 255875 4756 255876
rect 4724 255845 4725 255875
rect 4725 255845 4755 255875
rect 4755 255845 4756 255875
rect 4724 255844 4756 255845
rect 4724 255764 4756 255796
rect 4724 255715 4756 255716
rect 4724 255685 4725 255715
rect 4725 255685 4755 255715
rect 4755 255685 4756 255715
rect 4724 255684 4756 255685
rect 4804 255875 4836 255876
rect 4804 255845 4805 255875
rect 4805 255845 4835 255875
rect 4835 255845 4836 255875
rect 4804 255844 4836 255845
rect 4804 255764 4836 255796
rect 4804 255715 4836 255716
rect 4804 255685 4805 255715
rect 4805 255685 4835 255715
rect 4835 255685 4836 255715
rect 4804 255684 4836 255685
rect 4884 255875 4916 255876
rect 4884 255845 4885 255875
rect 4885 255845 4915 255875
rect 4915 255845 4916 255875
rect 4884 255844 4916 255845
rect 4884 255764 4916 255796
rect 4884 255715 4916 255716
rect 4884 255685 4885 255715
rect 4885 255685 4915 255715
rect 4915 255685 4916 255715
rect 4884 255684 4916 255685
rect 4964 255875 4996 255876
rect 4964 255845 4965 255875
rect 4965 255845 4995 255875
rect 4995 255845 4996 255875
rect 4964 255844 4996 255845
rect 4964 255764 4996 255796
rect 4964 255715 4996 255716
rect 4964 255685 4965 255715
rect 4965 255685 4995 255715
rect 4995 255685 4996 255715
rect 4964 255684 4996 255685
rect 5044 255875 5076 255876
rect 5044 255845 5045 255875
rect 5045 255845 5075 255875
rect 5075 255845 5076 255875
rect 5044 255844 5076 255845
rect 5044 255764 5076 255796
rect 5044 255715 5076 255716
rect 5044 255685 5045 255715
rect 5045 255685 5075 255715
rect 5075 255685 5076 255715
rect 5044 255684 5076 255685
rect 5124 255875 5156 255876
rect 5124 255845 5125 255875
rect 5125 255845 5155 255875
rect 5155 255845 5156 255875
rect 5124 255844 5156 255845
rect 5124 255764 5156 255796
rect 5124 255715 5156 255716
rect 5124 255685 5125 255715
rect 5125 255685 5155 255715
rect 5155 255685 5156 255715
rect 5124 255684 5156 255685
rect 5204 255875 5236 255876
rect 5204 255845 5205 255875
rect 5205 255845 5235 255875
rect 5235 255845 5236 255875
rect 5204 255844 5236 255845
rect 5204 255764 5236 255796
rect 5204 255715 5236 255716
rect 5204 255685 5205 255715
rect 5205 255685 5235 255715
rect 5235 255685 5236 255715
rect 5204 255684 5236 255685
rect 5284 255875 5316 255876
rect 5284 255845 5285 255875
rect 5285 255845 5315 255875
rect 5315 255845 5316 255875
rect 5284 255844 5316 255845
rect 5284 255764 5316 255796
rect 5284 255715 5316 255716
rect 5284 255685 5285 255715
rect 5285 255685 5315 255715
rect 5315 255685 5316 255715
rect 5284 255684 5316 255685
rect 5364 255875 5396 255876
rect 5364 255845 5365 255875
rect 5365 255845 5395 255875
rect 5395 255845 5396 255875
rect 5364 255844 5396 255845
rect 5364 255764 5396 255796
rect 5364 255715 5396 255716
rect 5364 255685 5365 255715
rect 5365 255685 5395 255715
rect 5395 255685 5396 255715
rect 5364 255684 5396 255685
rect 5444 255875 5476 255876
rect 5444 255845 5445 255875
rect 5445 255845 5475 255875
rect 5475 255845 5476 255875
rect 5444 255844 5476 255845
rect 5444 255764 5476 255796
rect 5444 255715 5476 255716
rect 5444 255685 5445 255715
rect 5445 255685 5475 255715
rect 5475 255685 5476 255715
rect 5444 255684 5476 255685
rect 5524 255875 5556 255876
rect 5524 255845 5525 255875
rect 5525 255845 5555 255875
rect 5555 255845 5556 255875
rect 5524 255844 5556 255845
rect 5524 255764 5556 255796
rect 5524 255715 5556 255716
rect 5524 255685 5525 255715
rect 5525 255685 5555 255715
rect 5555 255685 5556 255715
rect 5524 255684 5556 255685
rect 5604 255875 5636 255876
rect 5604 255845 5605 255875
rect 5605 255845 5635 255875
rect 5635 255845 5636 255875
rect 5604 255844 5636 255845
rect 5604 255764 5636 255796
rect 5604 255715 5636 255716
rect 5604 255685 5605 255715
rect 5605 255685 5635 255715
rect 5635 255685 5636 255715
rect 5604 255684 5636 255685
rect 5684 255875 5716 255876
rect 5684 255845 5685 255875
rect 5685 255845 5715 255875
rect 5715 255845 5716 255875
rect 5684 255844 5716 255845
rect 5684 255764 5716 255796
rect 5684 255715 5716 255716
rect 5684 255685 5685 255715
rect 5685 255685 5715 255715
rect 5715 255685 5716 255715
rect 5684 255684 5716 255685
rect 5764 255875 5796 255876
rect 5764 255845 5765 255875
rect 5765 255845 5795 255875
rect 5795 255845 5796 255875
rect 5764 255844 5796 255845
rect 5764 255764 5796 255796
rect 5764 255715 5796 255716
rect 5764 255685 5765 255715
rect 5765 255685 5795 255715
rect 5795 255685 5796 255715
rect 5764 255684 5796 255685
rect 5844 255875 5876 255876
rect 5844 255845 5845 255875
rect 5845 255845 5875 255875
rect 5875 255845 5876 255875
rect 5844 255844 5876 255845
rect 5844 255764 5876 255796
rect 5844 255715 5876 255716
rect 5844 255685 5845 255715
rect 5845 255685 5875 255715
rect 5875 255685 5876 255715
rect 5844 255684 5876 255685
rect 5924 255875 5956 255876
rect 5924 255845 5925 255875
rect 5925 255845 5955 255875
rect 5955 255845 5956 255875
rect 5924 255844 5956 255845
rect 5924 255764 5956 255796
rect 5924 255715 5956 255716
rect 5924 255685 5925 255715
rect 5925 255685 5955 255715
rect 5955 255685 5956 255715
rect 5924 255684 5956 255685
rect 6004 255875 6036 255876
rect 6004 255845 6005 255875
rect 6005 255845 6035 255875
rect 6035 255845 6036 255875
rect 6004 255844 6036 255845
rect 6004 255764 6036 255796
rect 6004 255715 6036 255716
rect 6004 255685 6005 255715
rect 6005 255685 6035 255715
rect 6035 255685 6036 255715
rect 6004 255684 6036 255685
rect 6084 255875 6116 255876
rect 6084 255845 6085 255875
rect 6085 255845 6115 255875
rect 6115 255845 6116 255875
rect 6084 255844 6116 255845
rect 6084 255764 6116 255796
rect 6084 255715 6116 255716
rect 6084 255685 6085 255715
rect 6085 255685 6115 255715
rect 6115 255685 6116 255715
rect 6084 255684 6116 255685
rect 6164 255875 6196 255876
rect 6164 255845 6165 255875
rect 6165 255845 6195 255875
rect 6195 255845 6196 255875
rect 6164 255844 6196 255845
rect 6164 255764 6196 255796
rect 6164 255715 6196 255716
rect 6164 255685 6165 255715
rect 6165 255685 6195 255715
rect 6195 255685 6196 255715
rect 6164 255684 6196 255685
rect 6244 255875 6276 255876
rect 6244 255845 6245 255875
rect 6245 255845 6275 255875
rect 6275 255845 6276 255875
rect 6244 255844 6276 255845
rect 6244 255764 6276 255796
rect 6244 255715 6276 255716
rect 6244 255685 6245 255715
rect 6245 255685 6275 255715
rect 6275 255685 6276 255715
rect 6244 255684 6276 255685
rect 6324 255875 6356 255876
rect 6324 255845 6325 255875
rect 6325 255845 6355 255875
rect 6355 255845 6356 255875
rect 6324 255844 6356 255845
rect 6324 255764 6356 255796
rect 6324 255715 6356 255716
rect 6324 255685 6325 255715
rect 6325 255685 6355 255715
rect 6355 255685 6356 255715
rect 6324 255684 6356 255685
rect 6404 255875 6436 255876
rect 6404 255845 6405 255875
rect 6405 255845 6435 255875
rect 6435 255845 6436 255875
rect 6404 255844 6436 255845
rect 6404 255764 6436 255796
rect 6404 255715 6436 255716
rect 6404 255685 6405 255715
rect 6405 255685 6435 255715
rect 6435 255685 6436 255715
rect 6404 255684 6436 255685
rect 6484 255875 6516 255876
rect 6484 255845 6485 255875
rect 6485 255845 6515 255875
rect 6515 255845 6516 255875
rect 6484 255844 6516 255845
rect 6484 255764 6516 255796
rect 6484 255715 6516 255716
rect 6484 255685 6485 255715
rect 6485 255685 6515 255715
rect 6515 255685 6516 255715
rect 6484 255684 6516 255685
rect 6564 255875 6596 255876
rect 6564 255845 6565 255875
rect 6565 255845 6595 255875
rect 6595 255845 6596 255875
rect 6564 255844 6596 255845
rect 6564 255764 6596 255796
rect 6564 255715 6596 255716
rect 6564 255685 6565 255715
rect 6565 255685 6595 255715
rect 6595 255685 6596 255715
rect 6564 255684 6596 255685
rect 6644 255875 6676 255876
rect 6644 255845 6645 255875
rect 6645 255845 6675 255875
rect 6675 255845 6676 255875
rect 6644 255844 6676 255845
rect 6644 255764 6676 255796
rect 6644 255715 6676 255716
rect 6644 255685 6645 255715
rect 6645 255685 6675 255715
rect 6675 255685 6676 255715
rect 6644 255684 6676 255685
rect 6724 255875 6756 255876
rect 6724 255845 6725 255875
rect 6725 255845 6755 255875
rect 6755 255845 6756 255875
rect 6724 255844 6756 255845
rect 6724 255764 6756 255796
rect 6724 255715 6756 255716
rect 6724 255685 6725 255715
rect 6725 255685 6755 255715
rect 6755 255685 6756 255715
rect 6724 255684 6756 255685
rect 6804 255875 6836 255876
rect 6804 255845 6805 255875
rect 6805 255845 6835 255875
rect 6835 255845 6836 255875
rect 6804 255844 6836 255845
rect 6804 255764 6836 255796
rect 6804 255715 6836 255716
rect 6804 255685 6805 255715
rect 6805 255685 6835 255715
rect 6835 255685 6836 255715
rect 6804 255684 6836 255685
rect 6884 255875 6916 255876
rect 6884 255845 6885 255875
rect 6885 255845 6915 255875
rect 6915 255845 6916 255875
rect 6884 255844 6916 255845
rect 6884 255764 6916 255796
rect 6884 255715 6916 255716
rect 6884 255685 6885 255715
rect 6885 255685 6915 255715
rect 6915 255685 6916 255715
rect 6884 255684 6916 255685
rect 6964 255875 6996 255876
rect 6964 255845 6965 255875
rect 6965 255845 6995 255875
rect 6995 255845 6996 255875
rect 6964 255844 6996 255845
rect 6964 255764 6996 255796
rect 6964 255715 6996 255716
rect 6964 255685 6965 255715
rect 6965 255685 6995 255715
rect 6995 255685 6996 255715
rect 6964 255684 6996 255685
rect 7044 255875 7076 255876
rect 7044 255845 7045 255875
rect 7045 255845 7075 255875
rect 7075 255845 7076 255875
rect 7044 255844 7076 255845
rect 7044 255764 7076 255796
rect 7044 255715 7076 255716
rect 7044 255685 7045 255715
rect 7045 255685 7075 255715
rect 7075 255685 7076 255715
rect 7044 255684 7076 255685
rect 7124 255875 7156 255876
rect 7124 255845 7125 255875
rect 7125 255845 7155 255875
rect 7155 255845 7156 255875
rect 7124 255844 7156 255845
rect 7124 255764 7156 255796
rect 7124 255715 7156 255716
rect 7124 255685 7125 255715
rect 7125 255685 7155 255715
rect 7155 255685 7156 255715
rect 7124 255684 7156 255685
rect 7204 255875 7236 255876
rect 7204 255845 7205 255875
rect 7205 255845 7235 255875
rect 7235 255845 7236 255875
rect 7204 255844 7236 255845
rect 7204 255764 7236 255796
rect 7204 255715 7236 255716
rect 7204 255685 7205 255715
rect 7205 255685 7235 255715
rect 7235 255685 7236 255715
rect 7204 255684 7236 255685
rect 7284 255875 7316 255876
rect 7284 255845 7285 255875
rect 7285 255845 7315 255875
rect 7315 255845 7316 255875
rect 7284 255844 7316 255845
rect 7284 255764 7316 255796
rect 7284 255715 7316 255716
rect 7284 255685 7285 255715
rect 7285 255685 7315 255715
rect 7315 255685 7316 255715
rect 7284 255684 7316 255685
rect 7364 255875 7396 255876
rect 7364 255845 7365 255875
rect 7365 255845 7395 255875
rect 7395 255845 7396 255875
rect 7364 255844 7396 255845
rect 7364 255764 7396 255796
rect 7364 255715 7396 255716
rect 7364 255685 7365 255715
rect 7365 255685 7395 255715
rect 7395 255685 7396 255715
rect 7364 255684 7396 255685
rect 7444 255875 7476 255876
rect 7444 255845 7445 255875
rect 7445 255845 7475 255875
rect 7475 255845 7476 255875
rect 7444 255844 7476 255845
rect 7444 255764 7476 255796
rect 7444 255715 7476 255716
rect 7444 255685 7445 255715
rect 7445 255685 7475 255715
rect 7475 255685 7476 255715
rect 7444 255684 7476 255685
rect 7524 255875 7556 255876
rect 7524 255845 7525 255875
rect 7525 255845 7555 255875
rect 7555 255845 7556 255875
rect 7524 255844 7556 255845
rect 7524 255764 7556 255796
rect 7524 255715 7556 255716
rect 7524 255685 7525 255715
rect 7525 255685 7555 255715
rect 7555 255685 7556 255715
rect 7524 255684 7556 255685
rect 7604 255875 7636 255876
rect 7604 255845 7605 255875
rect 7605 255845 7635 255875
rect 7635 255845 7636 255875
rect 7604 255844 7636 255845
rect 7604 255764 7636 255796
rect 7604 255715 7636 255716
rect 7604 255685 7605 255715
rect 7605 255685 7635 255715
rect 7635 255685 7636 255715
rect 7604 255684 7636 255685
rect 7684 255875 7716 255876
rect 7684 255845 7685 255875
rect 7685 255845 7715 255875
rect 7715 255845 7716 255875
rect 7684 255844 7716 255845
rect 7684 255764 7716 255796
rect 7684 255715 7716 255716
rect 7684 255685 7685 255715
rect 7685 255685 7715 255715
rect 7715 255685 7716 255715
rect 7684 255684 7716 255685
rect 7764 255875 7796 255876
rect 7764 255845 7765 255875
rect 7765 255845 7795 255875
rect 7795 255845 7796 255875
rect 7764 255844 7796 255845
rect 7764 255764 7796 255796
rect 7764 255715 7796 255716
rect 7764 255685 7765 255715
rect 7765 255685 7795 255715
rect 7795 255685 7796 255715
rect 7764 255684 7796 255685
rect 7844 255875 7876 255876
rect 7844 255845 7845 255875
rect 7845 255845 7875 255875
rect 7875 255845 7876 255875
rect 7844 255844 7876 255845
rect 7844 255764 7876 255796
rect 7844 255715 7876 255716
rect 7844 255685 7845 255715
rect 7845 255685 7875 255715
rect 7875 255685 7876 255715
rect 7844 255684 7876 255685
rect 7924 255875 7956 255876
rect 7924 255845 7925 255875
rect 7925 255845 7955 255875
rect 7955 255845 7956 255875
rect 7924 255844 7956 255845
rect 7924 255764 7956 255796
rect 7924 255715 7956 255716
rect 7924 255685 7925 255715
rect 7925 255685 7955 255715
rect 7955 255685 7956 255715
rect 7924 255684 7956 255685
rect 8004 255875 8036 255876
rect 8004 255845 8005 255875
rect 8005 255845 8035 255875
rect 8035 255845 8036 255875
rect 8004 255844 8036 255845
rect 8004 255764 8036 255796
rect 8004 255715 8036 255716
rect 8004 255685 8005 255715
rect 8005 255685 8035 255715
rect 8035 255685 8036 255715
rect 8004 255684 8036 255685
rect 8084 255875 8116 255876
rect 8084 255845 8085 255875
rect 8085 255845 8115 255875
rect 8115 255845 8116 255875
rect 8084 255844 8116 255845
rect 8084 255764 8116 255796
rect 8084 255715 8116 255716
rect 8084 255685 8085 255715
rect 8085 255685 8115 255715
rect 8115 255685 8116 255715
rect 8084 255684 8116 255685
rect 8164 255875 8196 255876
rect 8164 255845 8165 255875
rect 8165 255845 8195 255875
rect 8195 255845 8196 255875
rect 8164 255844 8196 255845
rect 8164 255764 8196 255796
rect 8164 255715 8196 255716
rect 8164 255685 8165 255715
rect 8165 255685 8195 255715
rect 8195 255685 8196 255715
rect 8164 255684 8196 255685
rect 8244 255875 8276 255876
rect 8244 255845 8245 255875
rect 8245 255845 8275 255875
rect 8275 255845 8276 255875
rect 8244 255844 8276 255845
rect 8244 255764 8276 255796
rect 8244 255715 8276 255716
rect 8244 255685 8245 255715
rect 8245 255685 8275 255715
rect 8275 255685 8276 255715
rect 8244 255684 8276 255685
rect 8324 255875 8356 255876
rect 8324 255845 8325 255875
rect 8325 255845 8355 255875
rect 8355 255845 8356 255875
rect 8324 255844 8356 255845
rect 8324 255764 8356 255796
rect 8324 255715 8356 255716
rect 8324 255685 8325 255715
rect 8325 255685 8355 255715
rect 8355 255685 8356 255715
rect 8324 255684 8356 255685
rect 8404 255875 8436 255876
rect 8404 255845 8405 255875
rect 8405 255845 8435 255875
rect 8435 255845 8436 255875
rect 8404 255844 8436 255845
rect 8404 255764 8436 255796
rect 8404 255715 8436 255716
rect 8404 255685 8405 255715
rect 8405 255685 8435 255715
rect 8435 255685 8436 255715
rect 8404 255684 8436 255685
rect 8484 255875 8516 255876
rect 8484 255845 8485 255875
rect 8485 255845 8515 255875
rect 8515 255845 8516 255875
rect 8484 255844 8516 255845
rect 8484 255764 8516 255796
rect 8484 255715 8516 255716
rect 8484 255685 8485 255715
rect 8485 255685 8515 255715
rect 8515 255685 8516 255715
rect 8484 255684 8516 255685
rect 8564 255875 8596 255876
rect 8564 255845 8565 255875
rect 8565 255845 8595 255875
rect 8595 255845 8596 255875
rect 8564 255844 8596 255845
rect 8564 255764 8596 255796
rect 8564 255715 8596 255716
rect 8564 255685 8565 255715
rect 8565 255685 8595 255715
rect 8595 255685 8596 255715
rect 8564 255684 8596 255685
rect 8644 255875 8676 255876
rect 8644 255845 8645 255875
rect 8645 255845 8675 255875
rect 8675 255845 8676 255875
rect 8644 255844 8676 255845
rect 8644 255764 8676 255796
rect 8644 255715 8676 255716
rect 8644 255685 8645 255715
rect 8645 255685 8675 255715
rect 8675 255685 8676 255715
rect 8644 255684 8676 255685
rect 8724 255875 8756 255876
rect 8724 255845 8725 255875
rect 8725 255845 8755 255875
rect 8755 255845 8756 255875
rect 8724 255844 8756 255845
rect 8724 255764 8756 255796
rect 8724 255715 8756 255716
rect 8724 255685 8725 255715
rect 8725 255685 8755 255715
rect 8755 255685 8756 255715
rect 8724 255684 8756 255685
rect 8804 255875 8836 255876
rect 8804 255845 8805 255875
rect 8805 255845 8835 255875
rect 8835 255845 8836 255875
rect 8804 255844 8836 255845
rect 8804 255764 8836 255796
rect 8804 255715 8836 255716
rect 8804 255685 8805 255715
rect 8805 255685 8835 255715
rect 8835 255685 8836 255715
rect 8804 255684 8836 255685
rect 8884 255875 8916 255876
rect 8884 255845 8885 255875
rect 8885 255845 8915 255875
rect 8915 255845 8916 255875
rect 8884 255844 8916 255845
rect 8884 255764 8916 255796
rect 8884 255715 8916 255716
rect 8884 255685 8885 255715
rect 8885 255685 8915 255715
rect 8915 255685 8916 255715
rect 8884 255684 8916 255685
rect 8964 255875 8996 255876
rect 8964 255845 8965 255875
rect 8965 255845 8995 255875
rect 8995 255845 8996 255875
rect 8964 255844 8996 255845
rect 8964 255764 8996 255796
rect 8964 255715 8996 255716
rect 8964 255685 8965 255715
rect 8965 255685 8995 255715
rect 8995 255685 8996 255715
rect 8964 255684 8996 255685
rect 9044 255875 9076 255876
rect 9044 255845 9045 255875
rect 9045 255845 9075 255875
rect 9075 255845 9076 255875
rect 9044 255844 9076 255845
rect 9044 255764 9076 255796
rect 9044 255715 9076 255716
rect 9044 255685 9045 255715
rect 9045 255685 9075 255715
rect 9075 255685 9076 255715
rect 9044 255684 9076 255685
rect 9124 255875 9156 255876
rect 9124 255845 9125 255875
rect 9125 255845 9155 255875
rect 9155 255845 9156 255875
rect 9124 255844 9156 255845
rect 9124 255764 9156 255796
rect 9124 255715 9156 255716
rect 9124 255685 9125 255715
rect 9125 255685 9155 255715
rect 9155 255685 9156 255715
rect 9124 255684 9156 255685
rect 9204 255875 9236 255876
rect 9204 255845 9205 255875
rect 9205 255845 9235 255875
rect 9235 255845 9236 255875
rect 9204 255844 9236 255845
rect 9204 255764 9236 255796
rect 9204 255715 9236 255716
rect 9204 255685 9205 255715
rect 9205 255685 9235 255715
rect 9235 255685 9236 255715
rect 9204 255684 9236 255685
rect 9284 255875 9316 255876
rect 9284 255845 9285 255875
rect 9285 255845 9315 255875
rect 9315 255845 9316 255875
rect 9284 255844 9316 255845
rect 9284 255764 9316 255796
rect 9284 255715 9316 255716
rect 9284 255685 9285 255715
rect 9285 255685 9315 255715
rect 9315 255685 9316 255715
rect 9284 255684 9316 255685
rect 9364 255875 9396 255876
rect 9364 255845 9365 255875
rect 9365 255845 9395 255875
rect 9395 255845 9396 255875
rect 9364 255844 9396 255845
rect 9364 255764 9396 255796
rect 9364 255715 9396 255716
rect 9364 255685 9365 255715
rect 9365 255685 9395 255715
rect 9395 255685 9396 255715
rect 9364 255684 9396 255685
rect 9444 255875 9476 255876
rect 9444 255845 9445 255875
rect 9445 255845 9475 255875
rect 9475 255845 9476 255875
rect 9444 255844 9476 255845
rect 9444 255764 9476 255796
rect 9444 255715 9476 255716
rect 9444 255685 9445 255715
rect 9445 255685 9475 255715
rect 9475 255685 9476 255715
rect 9444 255684 9476 255685
rect 9524 255875 9556 255876
rect 9524 255845 9525 255875
rect 9525 255845 9555 255875
rect 9555 255845 9556 255875
rect 9524 255844 9556 255845
rect 9524 255764 9556 255796
rect 9524 255715 9556 255716
rect 9524 255685 9525 255715
rect 9525 255685 9555 255715
rect 9555 255685 9556 255715
rect 9524 255684 9556 255685
rect 9604 255875 9636 255876
rect 9604 255845 9605 255875
rect 9605 255845 9635 255875
rect 9635 255845 9636 255875
rect 9604 255844 9636 255845
rect 9604 255764 9636 255796
rect 9604 255715 9636 255716
rect 9604 255685 9605 255715
rect 9605 255685 9635 255715
rect 9635 255685 9636 255715
rect 9604 255684 9636 255685
rect 9684 255875 9716 255876
rect 9684 255845 9685 255875
rect 9685 255845 9715 255875
rect 9715 255845 9716 255875
rect 9684 255844 9716 255845
rect 9684 255764 9716 255796
rect 9684 255715 9716 255716
rect 9684 255685 9685 255715
rect 9685 255685 9715 255715
rect 9715 255685 9716 255715
rect 9684 255684 9716 255685
rect 9764 255875 9796 255876
rect 9764 255845 9765 255875
rect 9765 255845 9795 255875
rect 9795 255845 9796 255875
rect 9764 255844 9796 255845
rect 9764 255764 9796 255796
rect 9764 255715 9796 255716
rect 9764 255685 9765 255715
rect 9765 255685 9795 255715
rect 9795 255685 9796 255715
rect 9764 255684 9796 255685
rect 9844 255875 9876 255876
rect 9844 255845 9845 255875
rect 9845 255845 9875 255875
rect 9875 255845 9876 255875
rect 9844 255844 9876 255845
rect 9844 255764 9876 255796
rect 9844 255715 9876 255716
rect 9844 255685 9845 255715
rect 9845 255685 9875 255715
rect 9875 255685 9876 255715
rect 9844 255684 9876 255685
rect 9924 255875 9956 255876
rect 9924 255845 9925 255875
rect 9925 255845 9955 255875
rect 9955 255845 9956 255875
rect 9924 255844 9956 255845
rect 9924 255764 9956 255796
rect 9924 255715 9956 255716
rect 9924 255685 9925 255715
rect 9925 255685 9955 255715
rect 9955 255685 9956 255715
rect 9924 255684 9956 255685
rect 10004 255875 10036 255876
rect 10004 255845 10005 255875
rect 10005 255845 10035 255875
rect 10035 255845 10036 255875
rect 10004 255844 10036 255845
rect 10004 255764 10036 255796
rect 10004 255715 10036 255716
rect 10004 255685 10005 255715
rect 10005 255685 10035 255715
rect 10035 255685 10036 255715
rect 10004 255684 10036 255685
rect 10084 255875 10116 255876
rect 10084 255845 10085 255875
rect 10085 255845 10115 255875
rect 10115 255845 10116 255875
rect 10084 255844 10116 255845
rect 10084 255764 10116 255796
rect 10084 255715 10116 255716
rect 10084 255685 10085 255715
rect 10085 255685 10115 255715
rect 10115 255685 10116 255715
rect 10084 255684 10116 255685
rect 10164 255875 10196 255876
rect 10164 255845 10165 255875
rect 10165 255845 10195 255875
rect 10195 255845 10196 255875
rect 10164 255844 10196 255845
rect 10164 255764 10196 255796
rect 10164 255715 10196 255716
rect 10164 255685 10165 255715
rect 10165 255685 10195 255715
rect 10195 255685 10196 255715
rect 10164 255684 10196 255685
rect 10244 255875 10276 255876
rect 10244 255845 10245 255875
rect 10245 255845 10275 255875
rect 10275 255845 10276 255875
rect 10244 255844 10276 255845
rect 10244 255764 10276 255796
rect 10244 255715 10276 255716
rect 10244 255685 10245 255715
rect 10245 255685 10275 255715
rect 10275 255685 10276 255715
rect 10244 255684 10276 255685
rect 10324 255875 10356 255876
rect 10324 255845 10325 255875
rect 10325 255845 10355 255875
rect 10355 255845 10356 255875
rect 10324 255844 10356 255845
rect 10324 255764 10356 255796
rect 10324 255715 10356 255716
rect 10324 255685 10325 255715
rect 10325 255685 10355 255715
rect 10355 255685 10356 255715
rect 10324 255684 10356 255685
rect 10404 255875 10436 255876
rect 10404 255845 10405 255875
rect 10405 255845 10435 255875
rect 10435 255845 10436 255875
rect 10404 255844 10436 255845
rect 10404 255764 10436 255796
rect 10404 255715 10436 255716
rect 10404 255685 10405 255715
rect 10405 255685 10435 255715
rect 10435 255685 10436 255715
rect 10404 255684 10436 255685
rect 10484 255875 10516 255876
rect 10484 255845 10485 255875
rect 10485 255845 10515 255875
rect 10515 255845 10516 255875
rect 10484 255844 10516 255845
rect 10484 255764 10516 255796
rect 10484 255715 10516 255716
rect 10484 255685 10485 255715
rect 10485 255685 10515 255715
rect 10515 255685 10516 255715
rect 10484 255684 10516 255685
rect 10564 255875 10596 255876
rect 10564 255845 10565 255875
rect 10565 255845 10595 255875
rect 10595 255845 10596 255875
rect 10564 255844 10596 255845
rect 10564 255764 10596 255796
rect 10564 255715 10596 255716
rect 10564 255685 10565 255715
rect 10565 255685 10595 255715
rect 10595 255685 10596 255715
rect 10564 255684 10596 255685
rect 10644 255875 10676 255876
rect 10644 255845 10645 255875
rect 10645 255845 10675 255875
rect 10675 255845 10676 255875
rect 10644 255844 10676 255845
rect 10644 255764 10676 255796
rect 10644 255715 10676 255716
rect 10644 255685 10645 255715
rect 10645 255685 10675 255715
rect 10675 255685 10676 255715
rect 10644 255684 10676 255685
rect 10724 255875 10756 255876
rect 10724 255845 10725 255875
rect 10725 255845 10755 255875
rect 10755 255845 10756 255875
rect 10724 255844 10756 255845
rect 10724 255764 10756 255796
rect 10724 255715 10756 255716
rect 10724 255685 10725 255715
rect 10725 255685 10755 255715
rect 10755 255685 10756 255715
rect 10724 255684 10756 255685
rect 10804 255875 10836 255876
rect 10804 255845 10805 255875
rect 10805 255845 10835 255875
rect 10835 255845 10836 255875
rect 10804 255844 10836 255845
rect 10804 255764 10836 255796
rect 10804 255715 10836 255716
rect 10804 255685 10805 255715
rect 10805 255685 10835 255715
rect 10835 255685 10836 255715
rect 10804 255684 10836 255685
rect 10884 255875 10916 255876
rect 10884 255845 10885 255875
rect 10885 255845 10915 255875
rect 10915 255845 10916 255875
rect 10884 255844 10916 255845
rect 10884 255764 10916 255796
rect 10884 255715 10916 255716
rect 10884 255685 10885 255715
rect 10885 255685 10915 255715
rect 10915 255685 10916 255715
rect 10884 255684 10916 255685
rect 10964 255875 10996 255876
rect 10964 255845 10965 255875
rect 10965 255845 10995 255875
rect 10995 255845 10996 255875
rect 10964 255844 10996 255845
rect 10964 255764 10996 255796
rect 10964 255715 10996 255716
rect 10964 255685 10965 255715
rect 10965 255685 10995 255715
rect 10995 255685 10996 255715
rect 10964 255684 10996 255685
rect 11044 255875 11076 255876
rect 11044 255845 11045 255875
rect 11045 255845 11075 255875
rect 11075 255845 11076 255875
rect 11044 255844 11076 255845
rect 11044 255764 11076 255796
rect 11044 255715 11076 255716
rect 11044 255685 11045 255715
rect 11045 255685 11075 255715
rect 11075 255685 11076 255715
rect 11044 255684 11076 255685
rect 11124 255875 11156 255876
rect 11124 255845 11125 255875
rect 11125 255845 11155 255875
rect 11155 255845 11156 255875
rect 11124 255844 11156 255845
rect 11124 255764 11156 255796
rect 11124 255715 11156 255716
rect 11124 255685 11125 255715
rect 11125 255685 11155 255715
rect 11155 255685 11156 255715
rect 11124 255684 11156 255685
rect 11204 255875 11236 255876
rect 11204 255845 11205 255875
rect 11205 255845 11235 255875
rect 11235 255845 11236 255875
rect 11204 255844 11236 255845
rect 11204 255764 11236 255796
rect 11204 255715 11236 255716
rect 11204 255685 11205 255715
rect 11205 255685 11235 255715
rect 11235 255685 11236 255715
rect 11204 255684 11236 255685
rect 11284 255875 11316 255876
rect 11284 255845 11285 255875
rect 11285 255845 11315 255875
rect 11315 255845 11316 255875
rect 11284 255844 11316 255845
rect 11284 255764 11316 255796
rect 11284 255715 11316 255716
rect 11284 255685 11285 255715
rect 11285 255685 11315 255715
rect 11315 255685 11316 255715
rect 11284 255684 11316 255685
rect 11364 255875 11396 255876
rect 11364 255845 11365 255875
rect 11365 255845 11395 255875
rect 11395 255845 11396 255875
rect 11364 255844 11396 255845
rect 11364 255764 11396 255796
rect 11364 255715 11396 255716
rect 11364 255685 11365 255715
rect 11365 255685 11395 255715
rect 11395 255685 11396 255715
rect 11364 255684 11396 255685
rect 11444 255875 11476 255876
rect 11444 255845 11445 255875
rect 11445 255845 11475 255875
rect 11475 255845 11476 255875
rect 11444 255844 11476 255845
rect 11444 255764 11476 255796
rect 11444 255715 11476 255716
rect 11444 255685 11445 255715
rect 11445 255685 11475 255715
rect 11475 255685 11476 255715
rect 11444 255684 11476 255685
rect 11524 255875 11556 255876
rect 11524 255845 11525 255875
rect 11525 255845 11555 255875
rect 11555 255845 11556 255875
rect 11524 255844 11556 255845
rect 11524 255764 11556 255796
rect 11524 255715 11556 255716
rect 11524 255685 11525 255715
rect 11525 255685 11555 255715
rect 11555 255685 11556 255715
rect 11524 255684 11556 255685
rect 11604 255875 11636 255876
rect 11604 255845 11605 255875
rect 11605 255845 11635 255875
rect 11635 255845 11636 255875
rect 11604 255844 11636 255845
rect 11604 255764 11636 255796
rect 11604 255715 11636 255716
rect 11604 255685 11605 255715
rect 11605 255685 11635 255715
rect 11635 255685 11636 255715
rect 11604 255684 11636 255685
rect 11684 255875 11716 255876
rect 11684 255845 11685 255875
rect 11685 255845 11715 255875
rect 11715 255845 11716 255875
rect 11684 255844 11716 255845
rect 11684 255764 11716 255796
rect 11684 255715 11716 255716
rect 11684 255685 11685 255715
rect 11685 255685 11715 255715
rect 11715 255685 11716 255715
rect 11684 255684 11716 255685
rect 11764 255875 11796 255876
rect 11764 255845 11765 255875
rect 11765 255845 11795 255875
rect 11795 255845 11796 255875
rect 11764 255844 11796 255845
rect 11764 255764 11796 255796
rect 11764 255715 11796 255716
rect 11764 255685 11765 255715
rect 11765 255685 11795 255715
rect 11795 255685 11796 255715
rect 11764 255684 11796 255685
rect 11844 255875 11876 255876
rect 11844 255845 11845 255875
rect 11845 255845 11875 255875
rect 11875 255845 11876 255875
rect 11844 255844 11876 255845
rect 11844 255764 11876 255796
rect 11844 255715 11876 255716
rect 11844 255685 11845 255715
rect 11845 255685 11875 255715
rect 11875 255685 11876 255715
rect 11844 255684 11876 255685
rect 11924 255875 11956 255876
rect 11924 255845 11925 255875
rect 11925 255845 11955 255875
rect 11955 255845 11956 255875
rect 11924 255844 11956 255845
rect 11924 255764 11956 255796
rect 11924 255715 11956 255716
rect 11924 255685 11925 255715
rect 11925 255685 11955 255715
rect 11955 255685 11956 255715
rect 11924 255684 11956 255685
rect 12004 255875 12036 255876
rect 12004 255845 12005 255875
rect 12005 255845 12035 255875
rect 12035 255845 12036 255875
rect 12004 255844 12036 255845
rect 12004 255764 12036 255796
rect 12004 255715 12036 255716
rect 12004 255685 12005 255715
rect 12005 255685 12035 255715
rect 12035 255685 12036 255715
rect 12004 255684 12036 255685
rect 12084 255875 12116 255876
rect 12084 255845 12085 255875
rect 12085 255845 12115 255875
rect 12115 255845 12116 255875
rect 12084 255844 12116 255845
rect 12084 255764 12116 255796
rect 12084 255715 12116 255716
rect 12084 255685 12085 255715
rect 12085 255685 12115 255715
rect 12115 255685 12116 255715
rect 12084 255684 12116 255685
rect 12164 255875 12196 255876
rect 12164 255845 12165 255875
rect 12165 255845 12195 255875
rect 12195 255845 12196 255875
rect 12164 255844 12196 255845
rect 12164 255764 12196 255796
rect 12164 255715 12196 255716
rect 12164 255685 12165 255715
rect 12165 255685 12195 255715
rect 12195 255685 12196 255715
rect 12164 255684 12196 255685
rect 12244 255875 12276 255876
rect 12244 255845 12245 255875
rect 12245 255845 12275 255875
rect 12275 255845 12276 255875
rect 12244 255844 12276 255845
rect 12244 255764 12276 255796
rect 12244 255715 12276 255716
rect 12244 255685 12245 255715
rect 12245 255685 12275 255715
rect 12275 255685 12276 255715
rect 12244 255684 12276 255685
rect 12324 255875 12356 255876
rect 12324 255845 12325 255875
rect 12325 255845 12355 255875
rect 12355 255845 12356 255875
rect 12324 255844 12356 255845
rect 12324 255764 12356 255796
rect 12324 255715 12356 255716
rect 12324 255685 12325 255715
rect 12325 255685 12355 255715
rect 12355 255685 12356 255715
rect 12324 255684 12356 255685
rect 12404 255875 12436 255876
rect 12404 255845 12405 255875
rect 12405 255845 12435 255875
rect 12435 255845 12436 255875
rect 12404 255844 12436 255845
rect 12404 255764 12436 255796
rect 12404 255715 12436 255716
rect 12404 255685 12405 255715
rect 12405 255685 12435 255715
rect 12435 255685 12436 255715
rect 12404 255684 12436 255685
rect 12484 255875 12516 255876
rect 12484 255845 12485 255875
rect 12485 255845 12515 255875
rect 12515 255845 12516 255875
rect 12484 255844 12516 255845
rect 12484 255764 12516 255796
rect 12484 255715 12516 255716
rect 12484 255685 12485 255715
rect 12485 255685 12515 255715
rect 12515 255685 12516 255715
rect 12484 255684 12516 255685
rect 12564 255875 12596 255876
rect 12564 255845 12565 255875
rect 12565 255845 12595 255875
rect 12595 255845 12596 255875
rect 12564 255844 12596 255845
rect 12564 255764 12596 255796
rect 12564 255715 12596 255716
rect 12564 255685 12565 255715
rect 12565 255685 12595 255715
rect 12595 255685 12596 255715
rect 12564 255684 12596 255685
rect 12644 255875 12676 255876
rect 12644 255845 12645 255875
rect 12645 255845 12675 255875
rect 12675 255845 12676 255875
rect 12644 255844 12676 255845
rect 12644 255764 12676 255796
rect 12644 255715 12676 255716
rect 12644 255685 12645 255715
rect 12645 255685 12675 255715
rect 12675 255685 12676 255715
rect 12644 255684 12676 255685
rect 12724 255875 12756 255876
rect 12724 255845 12725 255875
rect 12725 255845 12755 255875
rect 12755 255845 12756 255875
rect 12724 255844 12756 255845
rect 12724 255764 12756 255796
rect 12724 255715 12756 255716
rect 12724 255685 12725 255715
rect 12725 255685 12755 255715
rect 12755 255685 12756 255715
rect 12724 255684 12756 255685
rect 12804 255875 12836 255876
rect 12804 255845 12805 255875
rect 12805 255845 12835 255875
rect 12835 255845 12836 255875
rect 12804 255844 12836 255845
rect 12804 255764 12836 255796
rect 12804 255715 12836 255716
rect 12804 255685 12805 255715
rect 12805 255685 12835 255715
rect 12835 255685 12836 255715
rect 12804 255684 12836 255685
rect 12884 255875 12916 255876
rect 12884 255845 12885 255875
rect 12885 255845 12915 255875
rect 12915 255845 12916 255875
rect 12884 255844 12916 255845
rect 12884 255764 12916 255796
rect 12884 255715 12916 255716
rect 12884 255685 12885 255715
rect 12885 255685 12915 255715
rect 12915 255685 12916 255715
rect 12884 255684 12916 255685
rect 12964 255875 12996 255876
rect 12964 255845 12965 255875
rect 12965 255845 12995 255875
rect 12995 255845 12996 255875
rect 12964 255844 12996 255845
rect 12964 255764 12996 255796
rect 12964 255715 12996 255716
rect 12964 255685 12965 255715
rect 12965 255685 12995 255715
rect 12995 255685 12996 255715
rect 12964 255684 12996 255685
rect 13044 255875 13076 255876
rect 13044 255845 13045 255875
rect 13045 255845 13075 255875
rect 13075 255845 13076 255875
rect 13044 255844 13076 255845
rect 13044 255764 13076 255796
rect 13044 255715 13076 255716
rect 13044 255685 13045 255715
rect 13045 255685 13075 255715
rect 13075 255685 13076 255715
rect 13044 255684 13076 255685
rect 13124 255875 13156 255876
rect 13124 255845 13125 255875
rect 13125 255845 13155 255875
rect 13155 255845 13156 255875
rect 13124 255844 13156 255845
rect 13124 255764 13156 255796
rect 13124 255715 13156 255716
rect 13124 255685 13125 255715
rect 13125 255685 13155 255715
rect 13155 255685 13156 255715
rect 13124 255684 13156 255685
rect 13204 255875 13236 255876
rect 13204 255845 13205 255875
rect 13205 255845 13235 255875
rect 13235 255845 13236 255875
rect 13204 255844 13236 255845
rect 13204 255764 13236 255796
rect 13204 255715 13236 255716
rect 13204 255685 13205 255715
rect 13205 255685 13235 255715
rect 13235 255685 13236 255715
rect 13204 255684 13236 255685
rect 13284 255875 13316 255876
rect 13284 255845 13285 255875
rect 13285 255845 13315 255875
rect 13315 255845 13316 255875
rect 13284 255844 13316 255845
rect 13284 255764 13316 255796
rect 13284 255715 13316 255716
rect 13284 255685 13285 255715
rect 13285 255685 13315 255715
rect 13315 255685 13316 255715
rect 13284 255684 13316 255685
rect 13364 255875 13396 255876
rect 13364 255845 13365 255875
rect 13365 255845 13395 255875
rect 13395 255845 13396 255875
rect 13364 255844 13396 255845
rect 13364 255764 13396 255796
rect 13364 255715 13396 255716
rect 13364 255685 13365 255715
rect 13365 255685 13395 255715
rect 13395 255685 13396 255715
rect 13364 255684 13396 255685
rect 13444 255875 13476 255876
rect 13444 255845 13445 255875
rect 13445 255845 13475 255875
rect 13475 255845 13476 255875
rect 13444 255844 13476 255845
rect 13444 255764 13476 255796
rect 13444 255715 13476 255716
rect 13444 255685 13445 255715
rect 13445 255685 13475 255715
rect 13475 255685 13476 255715
rect 13444 255684 13476 255685
rect 13524 255875 13556 255876
rect 13524 255845 13525 255875
rect 13525 255845 13555 255875
rect 13555 255845 13556 255875
rect 13524 255844 13556 255845
rect 13524 255764 13556 255796
rect 13524 255715 13556 255716
rect 13524 255685 13525 255715
rect 13525 255685 13555 255715
rect 13555 255685 13556 255715
rect 13524 255684 13556 255685
rect 13604 255875 13636 255876
rect 13604 255845 13605 255875
rect 13605 255845 13635 255875
rect 13635 255845 13636 255875
rect 13604 255844 13636 255845
rect 13604 255764 13636 255796
rect 13604 255715 13636 255716
rect 13604 255685 13605 255715
rect 13605 255685 13635 255715
rect 13635 255685 13636 255715
rect 13604 255684 13636 255685
rect 13684 255875 13716 255876
rect 13684 255845 13685 255875
rect 13685 255845 13715 255875
rect 13715 255845 13716 255875
rect 13684 255844 13716 255845
rect 13684 255764 13716 255796
rect 13684 255715 13716 255716
rect 13684 255685 13685 255715
rect 13685 255685 13715 255715
rect 13715 255685 13716 255715
rect 13684 255684 13716 255685
rect 13764 255875 13796 255876
rect 13764 255845 13765 255875
rect 13765 255845 13795 255875
rect 13795 255845 13796 255875
rect 13764 255844 13796 255845
rect 13764 255764 13796 255796
rect 13764 255715 13796 255716
rect 13764 255685 13765 255715
rect 13765 255685 13795 255715
rect 13795 255685 13796 255715
rect 13764 255684 13796 255685
rect 13844 255875 13876 255876
rect 13844 255845 13845 255875
rect 13845 255845 13875 255875
rect 13875 255845 13876 255875
rect 13844 255844 13876 255845
rect 13844 255764 13876 255796
rect 13844 255715 13876 255716
rect 13844 255685 13845 255715
rect 13845 255685 13875 255715
rect 13875 255685 13876 255715
rect 13844 255684 13876 255685
rect 13924 255875 13956 255876
rect 13924 255845 13925 255875
rect 13925 255845 13955 255875
rect 13955 255845 13956 255875
rect 13924 255844 13956 255845
rect 13924 255764 13956 255796
rect 13924 255715 13956 255716
rect 13924 255685 13925 255715
rect 13925 255685 13955 255715
rect 13955 255685 13956 255715
rect 13924 255684 13956 255685
rect 14004 255875 14036 255876
rect 14004 255845 14005 255875
rect 14005 255845 14035 255875
rect 14035 255845 14036 255875
rect 14004 255844 14036 255845
rect 14004 255764 14036 255796
rect 14004 255715 14036 255716
rect 14004 255685 14005 255715
rect 14005 255685 14035 255715
rect 14035 255685 14036 255715
rect 14004 255684 14036 255685
rect 14084 255875 14116 255876
rect 14084 255845 14085 255875
rect 14085 255845 14115 255875
rect 14115 255845 14116 255875
rect 14084 255844 14116 255845
rect 14084 255764 14116 255796
rect 14084 255715 14116 255716
rect 14084 255685 14085 255715
rect 14085 255685 14115 255715
rect 14115 255685 14116 255715
rect 14084 255684 14116 255685
rect 14164 255875 14196 255876
rect 14164 255845 14165 255875
rect 14165 255845 14195 255875
rect 14195 255845 14196 255875
rect 14164 255844 14196 255845
rect 14164 255764 14196 255796
rect 14164 255715 14196 255716
rect 14164 255685 14165 255715
rect 14165 255685 14195 255715
rect 14195 255685 14196 255715
rect 14164 255684 14196 255685
rect 14244 255875 14276 255876
rect 14244 255845 14245 255875
rect 14245 255845 14275 255875
rect 14275 255845 14276 255875
rect 14244 255844 14276 255845
rect 14244 255764 14276 255796
rect 14244 255715 14276 255716
rect 14244 255685 14245 255715
rect 14245 255685 14275 255715
rect 14275 255685 14276 255715
rect 14244 255684 14276 255685
rect 14324 255875 14356 255876
rect 14324 255845 14325 255875
rect 14325 255845 14355 255875
rect 14355 255845 14356 255875
rect 14324 255844 14356 255845
rect 14324 255764 14356 255796
rect 14324 255715 14356 255716
rect 14324 255685 14325 255715
rect 14325 255685 14355 255715
rect 14355 255685 14356 255715
rect 14324 255684 14356 255685
rect 14404 255875 14436 255876
rect 14404 255845 14405 255875
rect 14405 255845 14435 255875
rect 14435 255845 14436 255875
rect 14404 255844 14436 255845
rect 14404 255764 14436 255796
rect 14404 255715 14436 255716
rect 14404 255685 14405 255715
rect 14405 255685 14435 255715
rect 14435 255685 14436 255715
rect 14404 255684 14436 255685
rect 14484 255875 14516 255876
rect 14484 255845 14485 255875
rect 14485 255845 14515 255875
rect 14515 255845 14516 255875
rect 14484 255844 14516 255845
rect 14484 255764 14516 255796
rect 14484 255715 14516 255716
rect 14484 255685 14485 255715
rect 14485 255685 14515 255715
rect 14515 255685 14516 255715
rect 14484 255684 14516 255685
rect 14564 255875 14596 255876
rect 14564 255845 14565 255875
rect 14565 255845 14595 255875
rect 14595 255845 14596 255875
rect 14564 255844 14596 255845
rect 14564 255764 14596 255796
rect 14564 255715 14596 255716
rect 14564 255685 14565 255715
rect 14565 255685 14595 255715
rect 14595 255685 14596 255715
rect 14564 255684 14596 255685
rect 14644 255875 14676 255876
rect 14644 255845 14645 255875
rect 14645 255845 14675 255875
rect 14675 255845 14676 255875
rect 14644 255844 14676 255845
rect 14644 255764 14676 255796
rect 14644 255715 14676 255716
rect 14644 255685 14645 255715
rect 14645 255685 14675 255715
rect 14675 255685 14676 255715
rect 14644 255684 14676 255685
rect 14724 255875 14756 255876
rect 14724 255845 14725 255875
rect 14725 255845 14755 255875
rect 14755 255845 14756 255875
rect 14724 255844 14756 255845
rect 14724 255764 14756 255796
rect 14724 255715 14756 255716
rect 14724 255685 14725 255715
rect 14725 255685 14755 255715
rect 14755 255685 14756 255715
rect 14724 255684 14756 255685
rect 14804 255875 14836 255876
rect 14804 255845 14805 255875
rect 14805 255845 14835 255875
rect 14835 255845 14836 255875
rect 14804 255844 14836 255845
rect 14804 255764 14836 255796
rect 14804 255715 14836 255716
rect 14804 255685 14805 255715
rect 14805 255685 14835 255715
rect 14835 255685 14836 255715
rect 14804 255684 14836 255685
rect 14884 255875 14916 255876
rect 14884 255845 14885 255875
rect 14885 255845 14915 255875
rect 14915 255845 14916 255875
rect 14884 255844 14916 255845
rect 14884 255764 14916 255796
rect 14884 255715 14916 255716
rect 14884 255685 14885 255715
rect 14885 255685 14915 255715
rect 14915 255685 14916 255715
rect 14884 255684 14916 255685
rect 14964 255875 14996 255876
rect 14964 255845 14965 255875
rect 14965 255845 14995 255875
rect 14995 255845 14996 255875
rect 14964 255844 14996 255845
rect 14964 255764 14996 255796
rect 14964 255715 14996 255716
rect 14964 255685 14965 255715
rect 14965 255685 14995 255715
rect 14995 255685 14996 255715
rect 14964 255684 14996 255685
rect 15044 255875 15076 255876
rect 15044 255845 15045 255875
rect 15045 255845 15075 255875
rect 15075 255845 15076 255875
rect 15044 255844 15076 255845
rect 15044 255764 15076 255796
rect 15044 255715 15076 255716
rect 15044 255685 15045 255715
rect 15045 255685 15075 255715
rect 15075 255685 15076 255715
rect 15044 255684 15076 255685
rect 15124 255875 15156 255876
rect 15124 255845 15125 255875
rect 15125 255845 15155 255875
rect 15155 255845 15156 255875
rect 15124 255844 15156 255845
rect 15124 255764 15156 255796
rect 15124 255715 15156 255716
rect 15124 255685 15125 255715
rect 15125 255685 15155 255715
rect 15155 255685 15156 255715
rect 15124 255684 15156 255685
rect 15204 255875 15236 255876
rect 15204 255845 15205 255875
rect 15205 255845 15235 255875
rect 15235 255845 15236 255875
rect 15204 255844 15236 255845
rect 15204 255764 15236 255796
rect 15204 255715 15236 255716
rect 15204 255685 15205 255715
rect 15205 255685 15235 255715
rect 15235 255685 15236 255715
rect 15204 255684 15236 255685
rect 15284 255875 15316 255876
rect 15284 255845 15285 255875
rect 15285 255845 15315 255875
rect 15315 255845 15316 255875
rect 15284 255844 15316 255845
rect 15284 255764 15316 255796
rect 15284 255715 15316 255716
rect 15284 255685 15285 255715
rect 15285 255685 15315 255715
rect 15315 255685 15316 255715
rect 15284 255684 15316 255685
rect 15364 255875 15396 255876
rect 15364 255845 15365 255875
rect 15365 255845 15395 255875
rect 15395 255845 15396 255875
rect 15364 255844 15396 255845
rect 15364 255764 15396 255796
rect 15364 255715 15396 255716
rect 15364 255685 15365 255715
rect 15365 255685 15395 255715
rect 15395 255685 15396 255715
rect 15364 255684 15396 255685
rect 15444 255875 15476 255876
rect 15444 255845 15445 255875
rect 15445 255845 15475 255875
rect 15475 255845 15476 255875
rect 15444 255844 15476 255845
rect 15444 255764 15476 255796
rect 15444 255715 15476 255716
rect 15444 255685 15445 255715
rect 15445 255685 15475 255715
rect 15475 255685 15476 255715
rect 15444 255684 15476 255685
rect 15524 255875 15556 255876
rect 15524 255845 15525 255875
rect 15525 255845 15555 255875
rect 15555 255845 15556 255875
rect 15524 255844 15556 255845
rect 15524 255764 15556 255796
rect 15524 255715 15556 255716
rect 15524 255685 15525 255715
rect 15525 255685 15555 255715
rect 15555 255685 15556 255715
rect 15524 255684 15556 255685
rect 15604 255875 15636 255876
rect 15604 255845 15605 255875
rect 15605 255845 15635 255875
rect 15635 255845 15636 255875
rect 15604 255844 15636 255845
rect 15604 255764 15636 255796
rect 15604 255715 15636 255716
rect 15604 255685 15605 255715
rect 15605 255685 15635 255715
rect 15635 255685 15636 255715
rect 15604 255684 15636 255685
rect 15684 255875 15716 255876
rect 15684 255845 15685 255875
rect 15685 255845 15715 255875
rect 15715 255845 15716 255875
rect 15684 255844 15716 255845
rect 15684 255764 15716 255796
rect 15684 255715 15716 255716
rect 15684 255685 15685 255715
rect 15685 255685 15715 255715
rect 15715 255685 15716 255715
rect 15684 255684 15716 255685
rect 15764 255875 15796 255876
rect 15764 255845 15765 255875
rect 15765 255845 15795 255875
rect 15795 255845 15796 255875
rect 15764 255844 15796 255845
rect 15764 255764 15796 255796
rect 15764 255715 15796 255716
rect 15764 255685 15765 255715
rect 15765 255685 15795 255715
rect 15795 255685 15796 255715
rect 15764 255684 15796 255685
rect 15844 255875 15876 255876
rect 15844 255845 15845 255875
rect 15845 255845 15875 255875
rect 15875 255845 15876 255875
rect 15844 255844 15876 255845
rect 15844 255764 15876 255796
rect 15844 255715 15876 255716
rect 15844 255685 15845 255715
rect 15845 255685 15875 255715
rect 15875 255685 15876 255715
rect 15844 255684 15876 255685
rect 15924 255875 15956 255876
rect 15924 255845 15925 255875
rect 15925 255845 15955 255875
rect 15955 255845 15956 255875
rect 15924 255844 15956 255845
rect 15924 255764 15956 255796
rect 15924 255715 15956 255716
rect 15924 255685 15925 255715
rect 15925 255685 15955 255715
rect 15955 255685 15956 255715
rect 15924 255684 15956 255685
rect 16004 255875 16036 255876
rect 16004 255845 16005 255875
rect 16005 255845 16035 255875
rect 16035 255845 16036 255875
rect 16004 255844 16036 255845
rect 16004 255764 16036 255796
rect 16004 255715 16036 255716
rect 16004 255685 16005 255715
rect 16005 255685 16035 255715
rect 16035 255685 16036 255715
rect 16004 255684 16036 255685
rect 16084 255875 16116 255876
rect 16084 255845 16085 255875
rect 16085 255845 16115 255875
rect 16115 255845 16116 255875
rect 16084 255844 16116 255845
rect 16084 255764 16116 255796
rect 16084 255715 16116 255716
rect 16084 255685 16085 255715
rect 16085 255685 16115 255715
rect 16115 255685 16116 255715
rect 16084 255684 16116 255685
rect 16164 255875 16196 255876
rect 16164 255845 16165 255875
rect 16165 255845 16195 255875
rect 16195 255845 16196 255875
rect 16164 255844 16196 255845
rect 16164 255764 16196 255796
rect 16164 255715 16196 255716
rect 16164 255685 16165 255715
rect 16165 255685 16195 255715
rect 16195 255685 16196 255715
rect 16164 255684 16196 255685
rect 16244 255875 16276 255876
rect 16244 255845 16245 255875
rect 16245 255845 16275 255875
rect 16275 255845 16276 255875
rect 16244 255844 16276 255845
rect 16244 255764 16276 255796
rect 16244 255715 16276 255716
rect 16244 255685 16245 255715
rect 16245 255685 16275 255715
rect 16275 255685 16276 255715
rect 16244 255684 16276 255685
rect 16324 255875 16356 255876
rect 16324 255845 16325 255875
rect 16325 255845 16355 255875
rect 16355 255845 16356 255875
rect 16324 255844 16356 255845
rect 16324 255764 16356 255796
rect 16324 255715 16356 255716
rect 16324 255685 16325 255715
rect 16325 255685 16355 255715
rect 16355 255685 16356 255715
rect 16324 255684 16356 255685
rect 16404 255875 16436 255876
rect 16404 255845 16405 255875
rect 16405 255845 16435 255875
rect 16435 255845 16436 255875
rect 16404 255844 16436 255845
rect 16404 255764 16436 255796
rect 16404 255715 16436 255716
rect 16404 255685 16405 255715
rect 16405 255685 16435 255715
rect 16435 255685 16436 255715
rect 16404 255684 16436 255685
rect 16484 255875 16516 255876
rect 16484 255845 16485 255875
rect 16485 255845 16515 255875
rect 16515 255845 16516 255875
rect 16484 255844 16516 255845
rect 16484 255764 16516 255796
rect 16484 255715 16516 255716
rect 16484 255685 16485 255715
rect 16485 255685 16515 255715
rect 16515 255685 16516 255715
rect 16484 255684 16516 255685
rect 16564 255875 16596 255876
rect 16564 255845 16565 255875
rect 16565 255845 16595 255875
rect 16595 255845 16596 255875
rect 16564 255844 16596 255845
rect 16564 255764 16596 255796
rect 16564 255715 16596 255716
rect 16564 255685 16565 255715
rect 16565 255685 16595 255715
rect 16595 255685 16596 255715
rect 16564 255684 16596 255685
rect 16644 255875 16676 255876
rect 16644 255845 16645 255875
rect 16645 255845 16675 255875
rect 16675 255845 16676 255875
rect 16644 255844 16676 255845
rect 16644 255764 16676 255796
rect 16644 255715 16676 255716
rect 16644 255685 16645 255715
rect 16645 255685 16675 255715
rect 16675 255685 16676 255715
rect 16644 255684 16676 255685
rect 16724 255875 16756 255876
rect 16724 255845 16725 255875
rect 16725 255845 16755 255875
rect 16755 255845 16756 255875
rect 16724 255844 16756 255845
rect 16724 255764 16756 255796
rect 16884 275364 16916 275396
rect 16884 275315 16916 275316
rect 16884 275285 16885 275315
rect 16885 275285 16915 275315
rect 16915 275285 16916 275315
rect 16884 275284 16916 275285
rect 16964 275475 16996 275476
rect 16964 275445 16965 275475
rect 16965 275445 16995 275475
rect 16995 275445 16996 275475
rect 16964 275444 16996 275445
rect 16964 275364 16996 275396
rect 16964 275315 16996 275316
rect 16964 275285 16965 275315
rect 16965 275285 16995 275315
rect 16995 275285 16996 275315
rect 16964 275284 16996 275285
rect 17044 275475 17076 275476
rect 17044 275445 17045 275475
rect 17045 275445 17075 275475
rect 17075 275445 17076 275475
rect 17044 275444 17076 275445
rect 17044 275364 17076 275396
rect 17124 275475 17156 275476
rect 17124 275445 17125 275475
rect 17125 275445 17155 275475
rect 17155 275445 17156 275475
rect 17124 275444 17156 275445
rect 17204 275475 17236 275476
rect 17204 275445 17205 275475
rect 17205 275445 17235 275475
rect 17235 275445 17236 275475
rect 17204 275444 17236 275445
rect 17044 275315 17076 275316
rect 17044 275285 17045 275315
rect 17045 275285 17075 275315
rect 17075 275285 17076 275315
rect 17044 275284 17076 275285
rect 17204 275315 17236 275316
rect 17204 275285 17205 275315
rect 17205 275285 17235 275315
rect 17235 275285 17236 275315
rect 17204 275284 17236 275285
rect 16884 274955 16916 274956
rect 16884 274925 16885 274955
rect 16885 274925 16915 274955
rect 16915 274925 16916 274955
rect 16884 274924 16916 274925
rect 28404 275355 28436 275356
rect 28404 275325 28405 275355
rect 28405 275325 28435 275355
rect 28435 275325 28436 275355
rect 28404 275324 28436 275325
rect 28404 275275 28436 275276
rect 28404 275245 28405 275275
rect 28405 275245 28435 275275
rect 28435 275245 28436 275275
rect 28404 275244 28436 275245
rect 28564 275355 28596 275356
rect 28564 275325 28565 275355
rect 28565 275325 28595 275355
rect 28595 275325 28596 275355
rect 28564 275324 28596 275325
rect 28564 275275 28596 275276
rect 28564 275245 28565 275275
rect 28565 275245 28595 275275
rect 28595 275245 28596 275275
rect 28564 275244 28596 275245
rect 28724 275355 28756 275356
rect 28724 275325 28725 275355
rect 28725 275325 28755 275355
rect 28755 275325 28756 275355
rect 28724 275324 28756 275325
rect 28724 275275 28756 275276
rect 28724 275245 28725 275275
rect 28725 275245 28755 275275
rect 28755 275245 28756 275275
rect 28724 275244 28756 275245
rect 271864 350375 271896 350376
rect 271864 350345 271865 350375
rect 271865 350345 271895 350375
rect 271895 350345 271896 350375
rect 271864 350344 271896 350345
rect 271864 350295 271896 350296
rect 271864 350265 271865 350295
rect 271865 350265 271895 350295
rect 271895 350265 271896 350295
rect 271864 350264 271896 350265
rect 271864 350215 271896 350216
rect 271864 350185 271865 350215
rect 271865 350185 271895 350215
rect 271895 350185 271896 350215
rect 271864 350184 271896 350185
rect 271864 350135 271896 350136
rect 271864 350105 271865 350135
rect 271865 350105 271895 350135
rect 271895 350105 271896 350135
rect 271864 350104 271896 350105
rect 271864 350055 271896 350056
rect 271864 350025 271865 350055
rect 271865 350025 271895 350055
rect 271895 350025 271896 350055
rect 271864 350024 271896 350025
rect 272024 351704 272056 351736
rect 272024 351655 272056 351656
rect 272024 351625 272025 351655
rect 272025 351625 272055 351655
rect 272055 351625 272056 351655
rect 272024 351624 272056 351625
rect 272104 351815 272136 351816
rect 272104 351785 272105 351815
rect 272105 351785 272135 351815
rect 272135 351785 272136 351815
rect 272104 351784 272136 351785
rect 272104 351704 272136 351736
rect 272104 351655 272136 351656
rect 272104 351625 272105 351655
rect 272105 351625 272135 351655
rect 272135 351625 272136 351655
rect 272104 351624 272136 351625
rect 272184 351815 272216 351816
rect 272184 351785 272185 351815
rect 272185 351785 272215 351815
rect 272215 351785 272216 351815
rect 272184 351784 272216 351785
rect 272184 351704 272216 351736
rect 272184 351655 272216 351656
rect 272184 351625 272185 351655
rect 272185 351625 272215 351655
rect 272215 351625 272216 351655
rect 272184 351624 272216 351625
rect 272264 351815 272296 351816
rect 272264 351785 272265 351815
rect 272265 351785 272295 351815
rect 272295 351785 272296 351815
rect 272264 351784 272296 351785
rect 272264 351704 272296 351736
rect 272264 351655 272296 351656
rect 272264 351625 272265 351655
rect 272265 351625 272295 351655
rect 272295 351625 272296 351655
rect 272264 351624 272296 351625
rect 272344 351815 272376 351816
rect 272344 351785 272345 351815
rect 272345 351785 272375 351815
rect 272375 351785 272376 351815
rect 272344 351784 272376 351785
rect 272344 351704 272376 351736
rect 272344 351655 272376 351656
rect 272344 351625 272345 351655
rect 272345 351625 272375 351655
rect 272375 351625 272376 351655
rect 272344 351624 272376 351625
rect 272424 351815 272456 351816
rect 272424 351785 272425 351815
rect 272425 351785 272455 351815
rect 272455 351785 272456 351815
rect 272424 351784 272456 351785
rect 272424 351704 272456 351736
rect 272424 351655 272456 351656
rect 272424 351625 272425 351655
rect 272425 351625 272455 351655
rect 272455 351625 272456 351655
rect 272424 351624 272456 351625
rect 272504 351815 272536 351816
rect 272504 351785 272505 351815
rect 272505 351785 272535 351815
rect 272535 351785 272536 351815
rect 272504 351784 272536 351785
rect 272504 351704 272536 351736
rect 272504 351655 272536 351656
rect 272504 351625 272505 351655
rect 272505 351625 272535 351655
rect 272535 351625 272536 351655
rect 272504 351624 272536 351625
rect 272584 351815 272616 351816
rect 272584 351785 272585 351815
rect 272585 351785 272615 351815
rect 272615 351785 272616 351815
rect 272584 351784 272616 351785
rect 272584 351704 272616 351736
rect 272584 351655 272616 351656
rect 272584 351625 272585 351655
rect 272585 351625 272615 351655
rect 272615 351625 272616 351655
rect 272584 351624 272616 351625
rect 272664 351815 272696 351816
rect 272664 351785 272665 351815
rect 272665 351785 272695 351815
rect 272695 351785 272696 351815
rect 272664 351784 272696 351785
rect 272664 351704 272696 351736
rect 272664 351655 272696 351656
rect 272664 351625 272665 351655
rect 272665 351625 272695 351655
rect 272695 351625 272696 351655
rect 272664 351624 272696 351625
rect 272744 351815 272776 351816
rect 272744 351785 272745 351815
rect 272745 351785 272775 351815
rect 272775 351785 272776 351815
rect 272744 351784 272776 351785
rect 272744 351704 272776 351736
rect 272744 351655 272776 351656
rect 272744 351625 272745 351655
rect 272745 351625 272775 351655
rect 272775 351625 272776 351655
rect 272744 351624 272776 351625
rect 272824 351815 272856 351816
rect 272824 351785 272825 351815
rect 272825 351785 272855 351815
rect 272855 351785 272856 351815
rect 272824 351784 272856 351785
rect 272824 351704 272856 351736
rect 272824 351655 272856 351656
rect 272824 351625 272825 351655
rect 272825 351625 272855 351655
rect 272855 351625 272856 351655
rect 272824 351624 272856 351625
rect 272904 351815 272936 351816
rect 272904 351785 272905 351815
rect 272905 351785 272935 351815
rect 272935 351785 272936 351815
rect 272904 351784 272936 351785
rect 272904 351704 272936 351736
rect 272904 351655 272936 351656
rect 272904 351625 272905 351655
rect 272905 351625 272935 351655
rect 272935 351625 272936 351655
rect 272904 351624 272936 351625
rect 272984 351815 273016 351816
rect 272984 351785 272985 351815
rect 272985 351785 273015 351815
rect 273015 351785 273016 351815
rect 272984 351784 273016 351785
rect 272984 351704 273016 351736
rect 272984 351655 273016 351656
rect 272984 351625 272985 351655
rect 272985 351625 273015 351655
rect 273015 351625 273016 351655
rect 272984 351624 273016 351625
rect 273064 351815 273096 351816
rect 273064 351785 273065 351815
rect 273065 351785 273095 351815
rect 273095 351785 273096 351815
rect 273064 351784 273096 351785
rect 273064 351704 273096 351736
rect 273064 351655 273096 351656
rect 273064 351625 273065 351655
rect 273065 351625 273095 351655
rect 273095 351625 273096 351655
rect 273064 351624 273096 351625
rect 273144 351815 273176 351816
rect 273144 351785 273145 351815
rect 273145 351785 273175 351815
rect 273175 351785 273176 351815
rect 273144 351784 273176 351785
rect 273144 351704 273176 351736
rect 273144 351655 273176 351656
rect 273144 351625 273145 351655
rect 273145 351625 273175 351655
rect 273175 351625 273176 351655
rect 273144 351624 273176 351625
rect 273224 351815 273256 351816
rect 273224 351785 273225 351815
rect 273225 351785 273255 351815
rect 273255 351785 273256 351815
rect 273224 351784 273256 351785
rect 273224 351704 273256 351736
rect 273224 351655 273256 351656
rect 273224 351625 273225 351655
rect 273225 351625 273255 351655
rect 273255 351625 273256 351655
rect 273224 351624 273256 351625
rect 273304 351815 273336 351816
rect 273304 351785 273305 351815
rect 273305 351785 273335 351815
rect 273335 351785 273336 351815
rect 273304 351784 273336 351785
rect 273304 351704 273336 351736
rect 273304 351655 273336 351656
rect 273304 351625 273305 351655
rect 273305 351625 273335 351655
rect 273335 351625 273336 351655
rect 273304 351624 273336 351625
rect 273384 351815 273416 351816
rect 273384 351785 273385 351815
rect 273385 351785 273415 351815
rect 273415 351785 273416 351815
rect 273384 351784 273416 351785
rect 273384 351704 273416 351736
rect 273384 351655 273416 351656
rect 273384 351625 273385 351655
rect 273385 351625 273415 351655
rect 273415 351625 273416 351655
rect 273384 351624 273416 351625
rect 273464 351815 273496 351816
rect 273464 351785 273465 351815
rect 273465 351785 273495 351815
rect 273495 351785 273496 351815
rect 273464 351784 273496 351785
rect 273464 351704 273496 351736
rect 273464 351655 273496 351656
rect 273464 351625 273465 351655
rect 273465 351625 273495 351655
rect 273495 351625 273496 351655
rect 273464 351624 273496 351625
rect 273544 351815 273576 351816
rect 273544 351785 273545 351815
rect 273545 351785 273575 351815
rect 273575 351785 273576 351815
rect 273544 351784 273576 351785
rect 273544 351704 273576 351736
rect 273544 351655 273576 351656
rect 273544 351625 273545 351655
rect 273545 351625 273575 351655
rect 273575 351625 273576 351655
rect 273544 351624 273576 351625
rect 273624 351815 273656 351816
rect 273624 351785 273625 351815
rect 273625 351785 273655 351815
rect 273655 351785 273656 351815
rect 273624 351784 273656 351785
rect 273624 351704 273656 351736
rect 273624 351655 273656 351656
rect 273624 351625 273625 351655
rect 273625 351625 273655 351655
rect 273655 351625 273656 351655
rect 273624 351624 273656 351625
rect 273704 351815 273736 351816
rect 273704 351785 273705 351815
rect 273705 351785 273735 351815
rect 273735 351785 273736 351815
rect 273704 351784 273736 351785
rect 273704 351704 273736 351736
rect 273704 351655 273736 351656
rect 273704 351625 273705 351655
rect 273705 351625 273735 351655
rect 273735 351625 273736 351655
rect 273704 351624 273736 351625
rect 273784 351815 273816 351816
rect 273784 351785 273785 351815
rect 273785 351785 273815 351815
rect 273815 351785 273816 351815
rect 273784 351784 273816 351785
rect 273784 351704 273816 351736
rect 273784 351655 273816 351656
rect 273784 351625 273785 351655
rect 273785 351625 273815 351655
rect 273815 351625 273816 351655
rect 273784 351624 273816 351625
rect 273864 351815 273896 351816
rect 273864 351785 273865 351815
rect 273865 351785 273895 351815
rect 273895 351785 273896 351815
rect 273864 351784 273896 351785
rect 273864 351704 273896 351736
rect 273864 351655 273896 351656
rect 273864 351625 273865 351655
rect 273865 351625 273895 351655
rect 273895 351625 273896 351655
rect 273864 351624 273896 351625
rect 273944 351815 273976 351816
rect 273944 351785 273945 351815
rect 273945 351785 273975 351815
rect 273975 351785 273976 351815
rect 273944 351784 273976 351785
rect 273944 351704 273976 351736
rect 273944 351655 273976 351656
rect 273944 351625 273945 351655
rect 273945 351625 273975 351655
rect 273975 351625 273976 351655
rect 273944 351624 273976 351625
rect 274024 351815 274056 351816
rect 274024 351785 274025 351815
rect 274025 351785 274055 351815
rect 274055 351785 274056 351815
rect 274024 351784 274056 351785
rect 274024 351704 274056 351736
rect 274024 351655 274056 351656
rect 274024 351625 274025 351655
rect 274025 351625 274055 351655
rect 274055 351625 274056 351655
rect 274024 351624 274056 351625
rect 274104 351815 274136 351816
rect 274104 351785 274105 351815
rect 274105 351785 274135 351815
rect 274135 351785 274136 351815
rect 274104 351784 274136 351785
rect 274104 351704 274136 351736
rect 274104 351655 274136 351656
rect 274104 351625 274105 351655
rect 274105 351625 274135 351655
rect 274135 351625 274136 351655
rect 274104 351624 274136 351625
rect 274184 351815 274216 351816
rect 274184 351785 274185 351815
rect 274185 351785 274215 351815
rect 274215 351785 274216 351815
rect 274184 351784 274216 351785
rect 274184 351704 274216 351736
rect 274184 351655 274216 351656
rect 274184 351625 274185 351655
rect 274185 351625 274215 351655
rect 274215 351625 274216 351655
rect 274184 351624 274216 351625
rect 274264 351815 274296 351816
rect 274264 351785 274265 351815
rect 274265 351785 274295 351815
rect 274295 351785 274296 351815
rect 274264 351784 274296 351785
rect 274264 351704 274296 351736
rect 274264 351655 274296 351656
rect 274264 351625 274265 351655
rect 274265 351625 274295 351655
rect 274295 351625 274296 351655
rect 274264 351624 274296 351625
rect 274344 351815 274376 351816
rect 274344 351785 274345 351815
rect 274345 351785 274375 351815
rect 274375 351785 274376 351815
rect 274344 351784 274376 351785
rect 274344 351704 274376 351736
rect 274344 351655 274376 351656
rect 274344 351625 274345 351655
rect 274345 351625 274375 351655
rect 274375 351625 274376 351655
rect 274344 351624 274376 351625
rect 274424 351815 274456 351816
rect 274424 351785 274425 351815
rect 274425 351785 274455 351815
rect 274455 351785 274456 351815
rect 274424 351784 274456 351785
rect 274424 351704 274456 351736
rect 274424 351655 274456 351656
rect 274424 351625 274425 351655
rect 274425 351625 274455 351655
rect 274455 351625 274456 351655
rect 274424 351624 274456 351625
rect 274504 351815 274536 351816
rect 274504 351785 274505 351815
rect 274505 351785 274535 351815
rect 274535 351785 274536 351815
rect 274504 351784 274536 351785
rect 274504 351704 274536 351736
rect 274504 351655 274536 351656
rect 274504 351625 274505 351655
rect 274505 351625 274535 351655
rect 274535 351625 274536 351655
rect 274504 351624 274536 351625
rect 274584 351815 274616 351816
rect 274584 351785 274585 351815
rect 274585 351785 274615 351815
rect 274615 351785 274616 351815
rect 274584 351784 274616 351785
rect 274584 351704 274616 351736
rect 274584 351655 274616 351656
rect 274584 351625 274585 351655
rect 274585 351625 274615 351655
rect 274615 351625 274616 351655
rect 274584 351624 274616 351625
rect 274664 351815 274696 351816
rect 274664 351785 274665 351815
rect 274665 351785 274695 351815
rect 274695 351785 274696 351815
rect 274664 351784 274696 351785
rect 274664 351704 274696 351736
rect 274664 351655 274696 351656
rect 274664 351625 274665 351655
rect 274665 351625 274695 351655
rect 274695 351625 274696 351655
rect 274664 351624 274696 351625
rect 274744 351815 274776 351816
rect 274744 351785 274745 351815
rect 274745 351785 274775 351815
rect 274775 351785 274776 351815
rect 274744 351784 274776 351785
rect 274744 351704 274776 351736
rect 274744 351655 274776 351656
rect 274744 351625 274745 351655
rect 274745 351625 274775 351655
rect 274775 351625 274776 351655
rect 274744 351624 274776 351625
rect 274824 351815 274856 351816
rect 274824 351785 274825 351815
rect 274825 351785 274855 351815
rect 274855 351785 274856 351815
rect 274824 351784 274856 351785
rect 274824 351704 274856 351736
rect 274824 351655 274856 351656
rect 274824 351625 274825 351655
rect 274825 351625 274855 351655
rect 274855 351625 274856 351655
rect 274824 351624 274856 351625
rect 274904 351815 274936 351816
rect 274904 351785 274905 351815
rect 274905 351785 274935 351815
rect 274935 351785 274936 351815
rect 274904 351784 274936 351785
rect 274904 351704 274936 351736
rect 274904 351655 274936 351656
rect 274904 351625 274905 351655
rect 274905 351625 274935 351655
rect 274935 351625 274936 351655
rect 274904 351624 274936 351625
rect 274984 351815 275016 351816
rect 274984 351785 274985 351815
rect 274985 351785 275015 351815
rect 275015 351785 275016 351815
rect 274984 351784 275016 351785
rect 274984 351704 275016 351736
rect 274984 351655 275016 351656
rect 274984 351625 274985 351655
rect 274985 351625 275015 351655
rect 275015 351625 275016 351655
rect 274984 351624 275016 351625
rect 275064 351815 275096 351816
rect 275064 351785 275065 351815
rect 275065 351785 275095 351815
rect 275095 351785 275096 351815
rect 275064 351784 275096 351785
rect 275064 351704 275096 351736
rect 275064 351655 275096 351656
rect 275064 351625 275065 351655
rect 275065 351625 275095 351655
rect 275095 351625 275096 351655
rect 275064 351624 275096 351625
rect 275144 351815 275176 351816
rect 275144 351785 275145 351815
rect 275145 351785 275175 351815
rect 275175 351785 275176 351815
rect 275144 351784 275176 351785
rect 275144 351704 275176 351736
rect 275144 351655 275176 351656
rect 275144 351625 275145 351655
rect 275145 351625 275175 351655
rect 275175 351625 275176 351655
rect 275144 351624 275176 351625
rect 275224 351815 275256 351816
rect 275224 351785 275225 351815
rect 275225 351785 275255 351815
rect 275255 351785 275256 351815
rect 275224 351784 275256 351785
rect 275224 351704 275256 351736
rect 275224 351655 275256 351656
rect 275224 351625 275225 351655
rect 275225 351625 275255 351655
rect 275255 351625 275256 351655
rect 275224 351624 275256 351625
rect 275304 351815 275336 351816
rect 275304 351785 275305 351815
rect 275305 351785 275335 351815
rect 275335 351785 275336 351815
rect 275304 351784 275336 351785
rect 275304 351704 275336 351736
rect 275304 351655 275336 351656
rect 275304 351625 275305 351655
rect 275305 351625 275335 351655
rect 275335 351625 275336 351655
rect 275304 351624 275336 351625
rect 275384 351815 275416 351816
rect 275384 351785 275385 351815
rect 275385 351785 275415 351815
rect 275415 351785 275416 351815
rect 275384 351784 275416 351785
rect 275384 351704 275416 351736
rect 275384 351655 275416 351656
rect 275384 351625 275385 351655
rect 275385 351625 275415 351655
rect 275415 351625 275416 351655
rect 275384 351624 275416 351625
rect 275464 351815 275496 351816
rect 275464 351785 275465 351815
rect 275465 351785 275495 351815
rect 275495 351785 275496 351815
rect 275464 351784 275496 351785
rect 275464 351704 275496 351736
rect 275464 351655 275496 351656
rect 275464 351625 275465 351655
rect 275465 351625 275495 351655
rect 275495 351625 275496 351655
rect 275464 351624 275496 351625
rect 275544 351815 275576 351816
rect 275544 351785 275545 351815
rect 275545 351785 275575 351815
rect 275575 351785 275576 351815
rect 275544 351784 275576 351785
rect 275544 351704 275576 351736
rect 275544 351655 275576 351656
rect 275544 351625 275545 351655
rect 275545 351625 275575 351655
rect 275575 351625 275576 351655
rect 275544 351624 275576 351625
rect 275624 351815 275656 351816
rect 275624 351785 275625 351815
rect 275625 351785 275655 351815
rect 275655 351785 275656 351815
rect 275624 351784 275656 351785
rect 275624 351704 275656 351736
rect 275624 351655 275656 351656
rect 275624 351625 275625 351655
rect 275625 351625 275655 351655
rect 275655 351625 275656 351655
rect 275624 351624 275656 351625
rect 275704 351815 275736 351816
rect 275704 351785 275705 351815
rect 275705 351785 275735 351815
rect 275735 351785 275736 351815
rect 275704 351784 275736 351785
rect 275704 351704 275736 351736
rect 275704 351655 275736 351656
rect 275704 351625 275705 351655
rect 275705 351625 275735 351655
rect 275735 351625 275736 351655
rect 275704 351624 275736 351625
rect 275784 351815 275816 351816
rect 275784 351785 275785 351815
rect 275785 351785 275815 351815
rect 275815 351785 275816 351815
rect 275784 351784 275816 351785
rect 275784 351704 275816 351736
rect 275784 351655 275816 351656
rect 275784 351625 275785 351655
rect 275785 351625 275815 351655
rect 275815 351625 275816 351655
rect 275784 351624 275816 351625
rect 275864 351815 275896 351816
rect 275864 351785 275865 351815
rect 275865 351785 275895 351815
rect 275895 351785 275896 351815
rect 275864 351784 275896 351785
rect 275864 351704 275896 351736
rect 275864 351655 275896 351656
rect 275864 351625 275865 351655
rect 275865 351625 275895 351655
rect 275895 351625 275896 351655
rect 275864 351624 275896 351625
rect 275944 351815 275976 351816
rect 275944 351785 275945 351815
rect 275945 351785 275975 351815
rect 275975 351785 275976 351815
rect 275944 351784 275976 351785
rect 275944 351704 275976 351736
rect 275944 351655 275976 351656
rect 275944 351625 275945 351655
rect 275945 351625 275975 351655
rect 275975 351625 275976 351655
rect 275944 351624 275976 351625
rect 276024 351815 276056 351816
rect 276024 351785 276025 351815
rect 276025 351785 276055 351815
rect 276055 351785 276056 351815
rect 276024 351784 276056 351785
rect 276024 351704 276056 351736
rect 276024 351655 276056 351656
rect 276024 351625 276025 351655
rect 276025 351625 276055 351655
rect 276055 351625 276056 351655
rect 276024 351624 276056 351625
rect 276104 351815 276136 351816
rect 276104 351785 276105 351815
rect 276105 351785 276135 351815
rect 276135 351785 276136 351815
rect 276104 351784 276136 351785
rect 276104 351704 276136 351736
rect 276104 351655 276136 351656
rect 276104 351625 276105 351655
rect 276105 351625 276135 351655
rect 276135 351625 276136 351655
rect 276104 351624 276136 351625
rect 276184 351815 276216 351816
rect 276184 351785 276185 351815
rect 276185 351785 276215 351815
rect 276215 351785 276216 351815
rect 276184 351784 276216 351785
rect 276184 351704 276216 351736
rect 276184 351655 276216 351656
rect 276184 351625 276185 351655
rect 276185 351625 276215 351655
rect 276215 351625 276216 351655
rect 276184 351624 276216 351625
rect 276264 351815 276296 351816
rect 276264 351785 276265 351815
rect 276265 351785 276295 351815
rect 276295 351785 276296 351815
rect 276264 351784 276296 351785
rect 276264 351704 276296 351736
rect 276264 351655 276296 351656
rect 276264 351625 276265 351655
rect 276265 351625 276295 351655
rect 276295 351625 276296 351655
rect 276264 351624 276296 351625
rect 276344 351815 276376 351816
rect 276344 351785 276345 351815
rect 276345 351785 276375 351815
rect 276375 351785 276376 351815
rect 276344 351784 276376 351785
rect 276344 351704 276376 351736
rect 276344 351655 276376 351656
rect 276344 351625 276345 351655
rect 276345 351625 276375 351655
rect 276375 351625 276376 351655
rect 276344 351624 276376 351625
rect 276424 351815 276456 351816
rect 276424 351785 276425 351815
rect 276425 351785 276455 351815
rect 276455 351785 276456 351815
rect 276424 351784 276456 351785
rect 276424 351704 276456 351736
rect 276424 351655 276456 351656
rect 276424 351625 276425 351655
rect 276425 351625 276455 351655
rect 276455 351625 276456 351655
rect 276424 351624 276456 351625
rect 276504 351815 276536 351816
rect 276504 351785 276505 351815
rect 276505 351785 276535 351815
rect 276535 351785 276536 351815
rect 276504 351784 276536 351785
rect 276504 351704 276536 351736
rect 276504 351655 276536 351656
rect 276504 351625 276505 351655
rect 276505 351625 276535 351655
rect 276535 351625 276536 351655
rect 276504 351624 276536 351625
rect 276584 351815 276616 351816
rect 276584 351785 276585 351815
rect 276585 351785 276615 351815
rect 276615 351785 276616 351815
rect 276584 351784 276616 351785
rect 276584 351704 276616 351736
rect 276584 351655 276616 351656
rect 276584 351625 276585 351655
rect 276585 351625 276615 351655
rect 276615 351625 276616 351655
rect 276584 351624 276616 351625
rect 276664 351815 276696 351816
rect 276664 351785 276665 351815
rect 276665 351785 276695 351815
rect 276695 351785 276696 351815
rect 276664 351784 276696 351785
rect 276664 351704 276696 351736
rect 276664 351655 276696 351656
rect 276664 351625 276665 351655
rect 276665 351625 276695 351655
rect 276695 351625 276696 351655
rect 276664 351624 276696 351625
rect 276744 351815 276776 351816
rect 276744 351785 276745 351815
rect 276745 351785 276775 351815
rect 276775 351785 276776 351815
rect 276744 351784 276776 351785
rect 276744 351704 276776 351736
rect 276744 351655 276776 351656
rect 276744 351625 276745 351655
rect 276745 351625 276775 351655
rect 276775 351625 276776 351655
rect 276744 351624 276776 351625
rect 276824 351815 276856 351816
rect 276824 351785 276825 351815
rect 276825 351785 276855 351815
rect 276855 351785 276856 351815
rect 276824 351784 276856 351785
rect 276824 351704 276856 351736
rect 276824 351655 276856 351656
rect 276824 351625 276825 351655
rect 276825 351625 276855 351655
rect 276855 351625 276856 351655
rect 276824 351624 276856 351625
rect 276904 351815 276936 351816
rect 276904 351785 276905 351815
rect 276905 351785 276935 351815
rect 276935 351785 276936 351815
rect 276904 351784 276936 351785
rect 276904 351704 276936 351736
rect 276904 351655 276936 351656
rect 276904 351625 276905 351655
rect 276905 351625 276935 351655
rect 276935 351625 276936 351655
rect 276904 351624 276936 351625
rect 276984 351815 277016 351816
rect 276984 351785 276985 351815
rect 276985 351785 277015 351815
rect 277015 351785 277016 351815
rect 276984 351784 277016 351785
rect 276984 351704 277016 351736
rect 276984 351655 277016 351656
rect 276984 351625 276985 351655
rect 276985 351625 277015 351655
rect 277015 351625 277016 351655
rect 276984 351624 277016 351625
rect 277064 351815 277096 351816
rect 277064 351785 277065 351815
rect 277065 351785 277095 351815
rect 277095 351785 277096 351815
rect 277064 351784 277096 351785
rect 277064 351704 277096 351736
rect 277064 351655 277096 351656
rect 277064 351625 277065 351655
rect 277065 351625 277095 351655
rect 277095 351625 277096 351655
rect 277064 351624 277096 351625
rect 277144 351815 277176 351816
rect 277144 351785 277145 351815
rect 277145 351785 277175 351815
rect 277175 351785 277176 351815
rect 277144 351784 277176 351785
rect 277144 351704 277176 351736
rect 277144 351655 277176 351656
rect 277144 351625 277145 351655
rect 277145 351625 277175 351655
rect 277175 351625 277176 351655
rect 277144 351624 277176 351625
rect 277224 351815 277256 351816
rect 277224 351785 277225 351815
rect 277225 351785 277255 351815
rect 277255 351785 277256 351815
rect 277224 351784 277256 351785
rect 277224 351704 277256 351736
rect 277224 351655 277256 351656
rect 277224 351625 277225 351655
rect 277225 351625 277255 351655
rect 277255 351625 277256 351655
rect 277224 351624 277256 351625
rect 277304 351815 277336 351816
rect 277304 351785 277305 351815
rect 277305 351785 277335 351815
rect 277335 351785 277336 351815
rect 277304 351784 277336 351785
rect 277304 351704 277336 351736
rect 277304 351655 277336 351656
rect 277304 351625 277305 351655
rect 277305 351625 277335 351655
rect 277335 351625 277336 351655
rect 277304 351624 277336 351625
rect 277384 351815 277416 351816
rect 277384 351785 277385 351815
rect 277385 351785 277415 351815
rect 277415 351785 277416 351815
rect 277384 351784 277416 351785
rect 277384 351704 277416 351736
rect 277384 351655 277416 351656
rect 277384 351625 277385 351655
rect 277385 351625 277415 351655
rect 277415 351625 277416 351655
rect 277384 351624 277416 351625
rect 277464 351815 277496 351816
rect 277464 351785 277465 351815
rect 277465 351785 277495 351815
rect 277495 351785 277496 351815
rect 277464 351784 277496 351785
rect 277464 351704 277496 351736
rect 277464 351655 277496 351656
rect 277464 351625 277465 351655
rect 277465 351625 277495 351655
rect 277495 351625 277496 351655
rect 277464 351624 277496 351625
rect 277544 351815 277576 351816
rect 277544 351785 277545 351815
rect 277545 351785 277575 351815
rect 277575 351785 277576 351815
rect 277544 351784 277576 351785
rect 277544 351704 277576 351736
rect 277544 351655 277576 351656
rect 277544 351625 277545 351655
rect 277545 351625 277575 351655
rect 277575 351625 277576 351655
rect 277544 351624 277576 351625
rect 277624 351815 277656 351816
rect 277624 351785 277625 351815
rect 277625 351785 277655 351815
rect 277655 351785 277656 351815
rect 277624 351784 277656 351785
rect 277624 351704 277656 351736
rect 277624 351655 277656 351656
rect 277624 351625 277625 351655
rect 277625 351625 277655 351655
rect 277655 351625 277656 351655
rect 277624 351624 277656 351625
rect 277704 351815 277736 351816
rect 277704 351785 277705 351815
rect 277705 351785 277735 351815
rect 277735 351785 277736 351815
rect 277704 351784 277736 351785
rect 277704 351704 277736 351736
rect 277704 351655 277736 351656
rect 277704 351625 277705 351655
rect 277705 351625 277735 351655
rect 277735 351625 277736 351655
rect 277704 351624 277736 351625
rect 277784 351815 277816 351816
rect 277784 351785 277785 351815
rect 277785 351785 277815 351815
rect 277815 351785 277816 351815
rect 277784 351784 277816 351785
rect 277784 351704 277816 351736
rect 277784 351655 277816 351656
rect 277784 351625 277785 351655
rect 277785 351625 277815 351655
rect 277815 351625 277816 351655
rect 277784 351624 277816 351625
rect 277864 351815 277896 351816
rect 277864 351785 277865 351815
rect 277865 351785 277895 351815
rect 277895 351785 277896 351815
rect 277864 351784 277896 351785
rect 277864 351704 277896 351736
rect 277864 351655 277896 351656
rect 277864 351625 277865 351655
rect 277865 351625 277895 351655
rect 277895 351625 277896 351655
rect 277864 351624 277896 351625
rect 277944 351815 277976 351816
rect 277944 351785 277945 351815
rect 277945 351785 277975 351815
rect 277975 351785 277976 351815
rect 277944 351784 277976 351785
rect 277944 351704 277976 351736
rect 277944 351655 277976 351656
rect 277944 351625 277945 351655
rect 277945 351625 277975 351655
rect 277975 351625 277976 351655
rect 277944 351624 277976 351625
rect 278024 351815 278056 351816
rect 278024 351785 278025 351815
rect 278025 351785 278055 351815
rect 278055 351785 278056 351815
rect 278024 351784 278056 351785
rect 278024 351704 278056 351736
rect 278024 351655 278056 351656
rect 278024 351625 278025 351655
rect 278025 351625 278055 351655
rect 278055 351625 278056 351655
rect 278024 351624 278056 351625
rect 278104 351815 278136 351816
rect 278104 351785 278105 351815
rect 278105 351785 278135 351815
rect 278135 351785 278136 351815
rect 278104 351784 278136 351785
rect 278104 351704 278136 351736
rect 278104 351655 278136 351656
rect 278104 351625 278105 351655
rect 278105 351625 278135 351655
rect 278135 351625 278136 351655
rect 278104 351624 278136 351625
rect 278184 351815 278216 351816
rect 278184 351785 278185 351815
rect 278185 351785 278215 351815
rect 278215 351785 278216 351815
rect 278184 351784 278216 351785
rect 278184 351704 278216 351736
rect 278184 351655 278216 351656
rect 278184 351625 278185 351655
rect 278185 351625 278215 351655
rect 278215 351625 278216 351655
rect 278184 351624 278216 351625
rect 278264 351815 278296 351816
rect 278264 351785 278265 351815
rect 278265 351785 278295 351815
rect 278295 351785 278296 351815
rect 278264 351784 278296 351785
rect 278264 351704 278296 351736
rect 278264 351655 278296 351656
rect 278264 351625 278265 351655
rect 278265 351625 278295 351655
rect 278295 351625 278296 351655
rect 278264 351624 278296 351625
rect 278344 351815 278376 351816
rect 278344 351785 278345 351815
rect 278345 351785 278375 351815
rect 278375 351785 278376 351815
rect 278344 351784 278376 351785
rect 278344 351704 278376 351736
rect 278344 351655 278376 351656
rect 278344 351625 278345 351655
rect 278345 351625 278375 351655
rect 278375 351625 278376 351655
rect 278344 351624 278376 351625
rect 278424 351815 278456 351816
rect 278424 351785 278425 351815
rect 278425 351785 278455 351815
rect 278455 351785 278456 351815
rect 278424 351784 278456 351785
rect 278424 351704 278456 351736
rect 278424 351655 278456 351656
rect 278424 351625 278425 351655
rect 278425 351625 278455 351655
rect 278455 351625 278456 351655
rect 278424 351624 278456 351625
rect 278504 351815 278536 351816
rect 278504 351785 278505 351815
rect 278505 351785 278535 351815
rect 278535 351785 278536 351815
rect 278504 351784 278536 351785
rect 278504 351704 278536 351736
rect 278504 351655 278536 351656
rect 278504 351625 278505 351655
rect 278505 351625 278535 351655
rect 278535 351625 278536 351655
rect 278504 351624 278536 351625
rect 278584 351815 278616 351816
rect 278584 351785 278585 351815
rect 278585 351785 278615 351815
rect 278615 351785 278616 351815
rect 278584 351784 278616 351785
rect 278584 351704 278616 351736
rect 278584 351655 278616 351656
rect 278584 351625 278585 351655
rect 278585 351625 278615 351655
rect 278615 351625 278616 351655
rect 278584 351624 278616 351625
rect 278664 351815 278696 351816
rect 278664 351785 278665 351815
rect 278665 351785 278695 351815
rect 278695 351785 278696 351815
rect 278664 351784 278696 351785
rect 278664 351704 278696 351736
rect 278664 351655 278696 351656
rect 278664 351625 278665 351655
rect 278665 351625 278695 351655
rect 278695 351625 278696 351655
rect 278664 351624 278696 351625
rect 278744 351815 278776 351816
rect 278744 351785 278745 351815
rect 278745 351785 278775 351815
rect 278775 351785 278776 351815
rect 278744 351784 278776 351785
rect 278744 351704 278776 351736
rect 278744 351655 278776 351656
rect 278744 351625 278745 351655
rect 278745 351625 278775 351655
rect 278775 351625 278776 351655
rect 278744 351624 278776 351625
rect 278824 351815 278856 351816
rect 278824 351785 278825 351815
rect 278825 351785 278855 351815
rect 278855 351785 278856 351815
rect 278824 351784 278856 351785
rect 278824 351704 278856 351736
rect 278824 351655 278856 351656
rect 278824 351625 278825 351655
rect 278825 351625 278855 351655
rect 278855 351625 278856 351655
rect 278824 351624 278856 351625
rect 278904 351815 278936 351816
rect 278904 351785 278905 351815
rect 278905 351785 278935 351815
rect 278935 351785 278936 351815
rect 278904 351784 278936 351785
rect 278904 351704 278936 351736
rect 278904 351655 278936 351656
rect 278904 351625 278905 351655
rect 278905 351625 278935 351655
rect 278935 351625 278936 351655
rect 278904 351624 278936 351625
rect 278984 351815 279016 351816
rect 278984 351785 278985 351815
rect 278985 351785 279015 351815
rect 279015 351785 279016 351815
rect 278984 351784 279016 351785
rect 278984 351704 279016 351736
rect 278984 351655 279016 351656
rect 278984 351625 278985 351655
rect 278985 351625 279015 351655
rect 279015 351625 279016 351655
rect 278984 351624 279016 351625
rect 279064 351815 279096 351816
rect 279064 351785 279065 351815
rect 279065 351785 279095 351815
rect 279095 351785 279096 351815
rect 279064 351784 279096 351785
rect 279064 351704 279096 351736
rect 279064 351655 279096 351656
rect 279064 351625 279065 351655
rect 279065 351625 279095 351655
rect 279095 351625 279096 351655
rect 279064 351624 279096 351625
rect 279144 351815 279176 351816
rect 279144 351785 279145 351815
rect 279145 351785 279175 351815
rect 279175 351785 279176 351815
rect 279144 351784 279176 351785
rect 279144 351704 279176 351736
rect 279144 351655 279176 351656
rect 279144 351625 279145 351655
rect 279145 351625 279175 351655
rect 279175 351625 279176 351655
rect 279144 351624 279176 351625
rect 279224 351815 279256 351816
rect 279224 351785 279225 351815
rect 279225 351785 279255 351815
rect 279255 351785 279256 351815
rect 279224 351784 279256 351785
rect 279224 351704 279256 351736
rect 279224 351655 279256 351656
rect 279224 351625 279225 351655
rect 279225 351625 279255 351655
rect 279255 351625 279256 351655
rect 279224 351624 279256 351625
rect 279304 351815 279336 351816
rect 279304 351785 279305 351815
rect 279305 351785 279335 351815
rect 279335 351785 279336 351815
rect 279304 351784 279336 351785
rect 279304 351704 279336 351736
rect 279304 351655 279336 351656
rect 279304 351625 279305 351655
rect 279305 351625 279335 351655
rect 279335 351625 279336 351655
rect 279304 351624 279336 351625
rect 279384 351815 279416 351816
rect 279384 351785 279385 351815
rect 279385 351785 279415 351815
rect 279415 351785 279416 351815
rect 279384 351784 279416 351785
rect 279384 351704 279416 351736
rect 279384 351655 279416 351656
rect 279384 351625 279385 351655
rect 279385 351625 279415 351655
rect 279415 351625 279416 351655
rect 279384 351624 279416 351625
rect 279464 351815 279496 351816
rect 279464 351785 279465 351815
rect 279465 351785 279495 351815
rect 279495 351785 279496 351815
rect 279464 351784 279496 351785
rect 279464 351704 279496 351736
rect 279464 351655 279496 351656
rect 279464 351625 279465 351655
rect 279465 351625 279495 351655
rect 279495 351625 279496 351655
rect 279464 351624 279496 351625
rect 279544 351815 279576 351816
rect 279544 351785 279545 351815
rect 279545 351785 279575 351815
rect 279575 351785 279576 351815
rect 279544 351784 279576 351785
rect 279544 351704 279576 351736
rect 279544 351655 279576 351656
rect 279544 351625 279545 351655
rect 279545 351625 279575 351655
rect 279575 351625 279576 351655
rect 279544 351624 279576 351625
rect 279624 351815 279656 351816
rect 279624 351785 279625 351815
rect 279625 351785 279655 351815
rect 279655 351785 279656 351815
rect 279624 351784 279656 351785
rect 279624 351704 279656 351736
rect 279624 351655 279656 351656
rect 279624 351625 279625 351655
rect 279625 351625 279655 351655
rect 279655 351625 279656 351655
rect 279624 351624 279656 351625
rect 279704 351815 279736 351816
rect 279704 351785 279705 351815
rect 279705 351785 279735 351815
rect 279735 351785 279736 351815
rect 279704 351784 279736 351785
rect 279704 351704 279736 351736
rect 279704 351655 279736 351656
rect 279704 351625 279705 351655
rect 279705 351625 279735 351655
rect 279735 351625 279736 351655
rect 279704 351624 279736 351625
rect 279784 351815 279816 351816
rect 279784 351785 279785 351815
rect 279785 351785 279815 351815
rect 279815 351785 279816 351815
rect 279784 351784 279816 351785
rect 279784 351704 279816 351736
rect 279784 351655 279816 351656
rect 279784 351625 279785 351655
rect 279785 351625 279815 351655
rect 279815 351625 279816 351655
rect 279784 351624 279816 351625
rect 279864 351815 279896 351816
rect 279864 351785 279865 351815
rect 279865 351785 279895 351815
rect 279895 351785 279896 351815
rect 279864 351784 279896 351785
rect 279864 351704 279896 351736
rect 279864 351655 279896 351656
rect 279864 351625 279865 351655
rect 279865 351625 279895 351655
rect 279895 351625 279896 351655
rect 279864 351624 279896 351625
rect 279944 351815 279976 351816
rect 279944 351785 279945 351815
rect 279945 351785 279975 351815
rect 279975 351785 279976 351815
rect 279944 351784 279976 351785
rect 279944 351704 279976 351736
rect 279944 351655 279976 351656
rect 279944 351625 279945 351655
rect 279945 351625 279975 351655
rect 279975 351625 279976 351655
rect 279944 351624 279976 351625
rect 280024 351815 280056 351816
rect 280024 351785 280025 351815
rect 280025 351785 280055 351815
rect 280055 351785 280056 351815
rect 280024 351784 280056 351785
rect 280024 351704 280056 351736
rect 280024 351655 280056 351656
rect 280024 351625 280025 351655
rect 280025 351625 280055 351655
rect 280055 351625 280056 351655
rect 280024 351624 280056 351625
rect 280104 351815 280136 351816
rect 280104 351785 280105 351815
rect 280105 351785 280135 351815
rect 280135 351785 280136 351815
rect 280104 351784 280136 351785
rect 280104 351704 280136 351736
rect 280104 351655 280136 351656
rect 280104 351625 280105 351655
rect 280105 351625 280135 351655
rect 280135 351625 280136 351655
rect 280104 351624 280136 351625
rect 280184 351815 280216 351816
rect 280184 351785 280185 351815
rect 280185 351785 280215 351815
rect 280215 351785 280216 351815
rect 280184 351784 280216 351785
rect 280184 351704 280216 351736
rect 280184 351655 280216 351656
rect 280184 351625 280185 351655
rect 280185 351625 280215 351655
rect 280215 351625 280216 351655
rect 280184 351624 280216 351625
rect 280264 351815 280296 351816
rect 280264 351785 280265 351815
rect 280265 351785 280295 351815
rect 280295 351785 280296 351815
rect 280264 351784 280296 351785
rect 280264 351704 280296 351736
rect 280264 351655 280296 351656
rect 280264 351625 280265 351655
rect 280265 351625 280295 351655
rect 280295 351625 280296 351655
rect 280264 351624 280296 351625
rect 280344 351815 280376 351816
rect 280344 351785 280345 351815
rect 280345 351785 280375 351815
rect 280375 351785 280376 351815
rect 280344 351784 280376 351785
rect 280344 351704 280376 351736
rect 280344 351655 280376 351656
rect 280344 351625 280345 351655
rect 280345 351625 280375 351655
rect 280375 351625 280376 351655
rect 280344 351624 280376 351625
rect 280424 351815 280456 351816
rect 280424 351785 280425 351815
rect 280425 351785 280455 351815
rect 280455 351785 280456 351815
rect 280424 351784 280456 351785
rect 280424 351704 280456 351736
rect 280424 351655 280456 351656
rect 280424 351625 280425 351655
rect 280425 351625 280455 351655
rect 280455 351625 280456 351655
rect 280424 351624 280456 351625
rect 280504 351815 280536 351816
rect 280504 351785 280505 351815
rect 280505 351785 280535 351815
rect 280535 351785 280536 351815
rect 280504 351784 280536 351785
rect 280504 351704 280536 351736
rect 280504 351655 280536 351656
rect 280504 351625 280505 351655
rect 280505 351625 280535 351655
rect 280535 351625 280536 351655
rect 280504 351624 280536 351625
rect 280584 351815 280616 351816
rect 280584 351785 280585 351815
rect 280585 351785 280615 351815
rect 280615 351785 280616 351815
rect 280584 351784 280616 351785
rect 280584 351704 280616 351736
rect 280584 351655 280616 351656
rect 280584 351625 280585 351655
rect 280585 351625 280615 351655
rect 280615 351625 280616 351655
rect 280584 351624 280616 351625
rect 280664 351815 280696 351816
rect 280664 351785 280665 351815
rect 280665 351785 280695 351815
rect 280695 351785 280696 351815
rect 280664 351784 280696 351785
rect 280664 351704 280696 351736
rect 280664 351655 280696 351656
rect 280664 351625 280665 351655
rect 280665 351625 280695 351655
rect 280695 351625 280696 351655
rect 280664 351624 280696 351625
rect 280744 351815 280776 351816
rect 280744 351785 280745 351815
rect 280745 351785 280775 351815
rect 280775 351785 280776 351815
rect 280744 351784 280776 351785
rect 280744 351704 280776 351736
rect 280744 351655 280776 351656
rect 280744 351625 280745 351655
rect 280745 351625 280775 351655
rect 280775 351625 280776 351655
rect 280744 351624 280776 351625
rect 280824 351815 280856 351816
rect 280824 351785 280825 351815
rect 280825 351785 280855 351815
rect 280855 351785 280856 351815
rect 280824 351784 280856 351785
rect 280824 351704 280856 351736
rect 280824 351655 280856 351656
rect 280824 351625 280825 351655
rect 280825 351625 280855 351655
rect 280855 351625 280856 351655
rect 280824 351624 280856 351625
rect 280904 351815 280936 351816
rect 280904 351785 280905 351815
rect 280905 351785 280935 351815
rect 280935 351785 280936 351815
rect 280904 351784 280936 351785
rect 280904 351704 280936 351736
rect 280904 351655 280936 351656
rect 280904 351625 280905 351655
rect 280905 351625 280935 351655
rect 280935 351625 280936 351655
rect 280904 351624 280936 351625
rect 280984 351815 281016 351816
rect 280984 351785 280985 351815
rect 280985 351785 281015 351815
rect 281015 351785 281016 351815
rect 280984 351784 281016 351785
rect 280984 351704 281016 351736
rect 280984 351655 281016 351656
rect 280984 351625 280985 351655
rect 280985 351625 281015 351655
rect 281015 351625 281016 351655
rect 280984 351624 281016 351625
rect 281064 351815 281096 351816
rect 281064 351785 281065 351815
rect 281065 351785 281095 351815
rect 281095 351785 281096 351815
rect 281064 351784 281096 351785
rect 281064 351704 281096 351736
rect 281064 351655 281096 351656
rect 281064 351625 281065 351655
rect 281065 351625 281095 351655
rect 281095 351625 281096 351655
rect 281064 351624 281096 351625
rect 281144 351815 281176 351816
rect 281144 351785 281145 351815
rect 281145 351785 281175 351815
rect 281175 351785 281176 351815
rect 281144 351784 281176 351785
rect 281144 351704 281176 351736
rect 281144 351655 281176 351656
rect 281144 351625 281145 351655
rect 281145 351625 281175 351655
rect 281175 351625 281176 351655
rect 281144 351624 281176 351625
rect 281224 351815 281256 351816
rect 281224 351785 281225 351815
rect 281225 351785 281255 351815
rect 281255 351785 281256 351815
rect 281224 351784 281256 351785
rect 281224 351704 281256 351736
rect 281224 351655 281256 351656
rect 281224 351625 281225 351655
rect 281225 351625 281255 351655
rect 281255 351625 281256 351655
rect 281224 351624 281256 351625
rect 281304 351815 281336 351816
rect 281304 351785 281305 351815
rect 281305 351785 281335 351815
rect 281335 351785 281336 351815
rect 281304 351784 281336 351785
rect 281304 351704 281336 351736
rect 281304 351655 281336 351656
rect 281304 351625 281305 351655
rect 281305 351625 281335 351655
rect 281335 351625 281336 351655
rect 281304 351624 281336 351625
rect 281384 351815 281416 351816
rect 281384 351785 281385 351815
rect 281385 351785 281415 351815
rect 281415 351785 281416 351815
rect 281384 351784 281416 351785
rect 281384 351704 281416 351736
rect 281384 351655 281416 351656
rect 281384 351625 281385 351655
rect 281385 351625 281415 351655
rect 281415 351625 281416 351655
rect 281384 351624 281416 351625
rect 281464 351815 281496 351816
rect 281464 351785 281465 351815
rect 281465 351785 281495 351815
rect 281495 351785 281496 351815
rect 281464 351784 281496 351785
rect 281464 351704 281496 351736
rect 281464 351655 281496 351656
rect 281464 351625 281465 351655
rect 281465 351625 281495 351655
rect 281495 351625 281496 351655
rect 281464 351624 281496 351625
rect 281544 351815 281576 351816
rect 281544 351785 281545 351815
rect 281545 351785 281575 351815
rect 281575 351785 281576 351815
rect 281544 351784 281576 351785
rect 281544 351704 281576 351736
rect 281544 351655 281576 351656
rect 281544 351625 281545 351655
rect 281545 351625 281575 351655
rect 281575 351625 281576 351655
rect 281544 351624 281576 351625
rect 281624 351815 281656 351816
rect 281624 351785 281625 351815
rect 281625 351785 281655 351815
rect 281655 351785 281656 351815
rect 281624 351784 281656 351785
rect 281624 351704 281656 351736
rect 281624 351655 281656 351656
rect 281624 351625 281625 351655
rect 281625 351625 281655 351655
rect 281655 351625 281656 351655
rect 281624 351624 281656 351625
rect 281704 351815 281736 351816
rect 281704 351785 281705 351815
rect 281705 351785 281735 351815
rect 281735 351785 281736 351815
rect 281704 351784 281736 351785
rect 281704 351704 281736 351736
rect 281704 351655 281736 351656
rect 281704 351625 281705 351655
rect 281705 351625 281735 351655
rect 281735 351625 281736 351655
rect 281704 351624 281736 351625
rect 281784 351815 281816 351816
rect 281784 351785 281785 351815
rect 281785 351785 281815 351815
rect 281815 351785 281816 351815
rect 281784 351784 281816 351785
rect 281784 351704 281816 351736
rect 281784 351655 281816 351656
rect 281784 351625 281785 351655
rect 281785 351625 281815 351655
rect 281815 351625 281816 351655
rect 281784 351624 281816 351625
rect 281864 351815 281896 351816
rect 281864 351785 281865 351815
rect 281865 351785 281895 351815
rect 281895 351785 281896 351815
rect 281864 351784 281896 351785
rect 281864 351704 281896 351736
rect 281864 351655 281896 351656
rect 281864 351625 281865 351655
rect 281865 351625 281895 351655
rect 281895 351625 281896 351655
rect 281864 351624 281896 351625
rect 281944 351815 281976 351816
rect 281944 351785 281945 351815
rect 281945 351785 281975 351815
rect 281975 351785 281976 351815
rect 281944 351784 281976 351785
rect 281944 351704 281976 351736
rect 281944 351655 281976 351656
rect 281944 351625 281945 351655
rect 281945 351625 281975 351655
rect 281975 351625 281976 351655
rect 281944 351624 281976 351625
rect 282024 351815 282056 351816
rect 282024 351785 282025 351815
rect 282025 351785 282055 351815
rect 282055 351785 282056 351815
rect 282024 351784 282056 351785
rect 282024 351704 282056 351736
rect 282024 351655 282056 351656
rect 282024 351625 282025 351655
rect 282025 351625 282055 351655
rect 282055 351625 282056 351655
rect 282024 351624 282056 351625
rect 282104 351815 282136 351816
rect 282104 351785 282105 351815
rect 282105 351785 282135 351815
rect 282135 351785 282136 351815
rect 282104 351784 282136 351785
rect 282104 351704 282136 351736
rect 282104 351655 282136 351656
rect 282104 351625 282105 351655
rect 282105 351625 282135 351655
rect 282135 351625 282136 351655
rect 282104 351624 282136 351625
rect 282184 351815 282216 351816
rect 282184 351785 282185 351815
rect 282185 351785 282215 351815
rect 282215 351785 282216 351815
rect 282184 351784 282216 351785
rect 282184 351704 282216 351736
rect 282184 351655 282216 351656
rect 282184 351625 282185 351655
rect 282185 351625 282215 351655
rect 282215 351625 282216 351655
rect 282184 351624 282216 351625
rect 282264 351815 282296 351816
rect 282264 351785 282265 351815
rect 282265 351785 282295 351815
rect 282295 351785 282296 351815
rect 282264 351784 282296 351785
rect 282264 351704 282296 351736
rect 282264 351655 282296 351656
rect 282264 351625 282265 351655
rect 282265 351625 282295 351655
rect 282295 351625 282296 351655
rect 282264 351624 282296 351625
rect 282344 351815 282376 351816
rect 282344 351785 282345 351815
rect 282345 351785 282375 351815
rect 282375 351785 282376 351815
rect 282344 351784 282376 351785
rect 282344 351704 282376 351736
rect 282344 351655 282376 351656
rect 282344 351625 282345 351655
rect 282345 351625 282375 351655
rect 282375 351625 282376 351655
rect 282344 351624 282376 351625
rect 282424 351815 282456 351816
rect 282424 351785 282425 351815
rect 282425 351785 282455 351815
rect 282455 351785 282456 351815
rect 282424 351784 282456 351785
rect 282424 351704 282456 351736
rect 282424 351655 282456 351656
rect 282424 351625 282425 351655
rect 282425 351625 282455 351655
rect 282455 351625 282456 351655
rect 282424 351624 282456 351625
rect 282504 351815 282536 351816
rect 282504 351785 282505 351815
rect 282505 351785 282535 351815
rect 282535 351785 282536 351815
rect 282504 351784 282536 351785
rect 282504 351704 282536 351736
rect 282504 351655 282536 351656
rect 282504 351625 282505 351655
rect 282505 351625 282535 351655
rect 282535 351625 282536 351655
rect 282504 351624 282536 351625
rect 282584 351815 282616 351816
rect 282584 351785 282585 351815
rect 282585 351785 282615 351815
rect 282615 351785 282616 351815
rect 282584 351784 282616 351785
rect 282584 351704 282616 351736
rect 282584 351655 282616 351656
rect 282584 351625 282585 351655
rect 282585 351625 282615 351655
rect 282615 351625 282616 351655
rect 282584 351624 282616 351625
rect 282664 351815 282696 351816
rect 282664 351785 282665 351815
rect 282665 351785 282695 351815
rect 282695 351785 282696 351815
rect 282664 351784 282696 351785
rect 282664 351704 282696 351736
rect 282664 351655 282696 351656
rect 282664 351625 282665 351655
rect 282665 351625 282695 351655
rect 282695 351625 282696 351655
rect 282664 351624 282696 351625
rect 282744 351815 282776 351816
rect 282744 351785 282745 351815
rect 282745 351785 282775 351815
rect 282775 351785 282776 351815
rect 282744 351784 282776 351785
rect 282744 351704 282776 351736
rect 282744 351655 282776 351656
rect 282744 351625 282745 351655
rect 282745 351625 282775 351655
rect 282775 351625 282776 351655
rect 282744 351624 282776 351625
rect 282824 351815 282856 351816
rect 282824 351785 282825 351815
rect 282825 351785 282855 351815
rect 282855 351785 282856 351815
rect 282824 351784 282856 351785
rect 282824 351704 282856 351736
rect 282824 351655 282856 351656
rect 282824 351625 282825 351655
rect 282825 351625 282855 351655
rect 282855 351625 282856 351655
rect 282824 351624 282856 351625
rect 282904 351815 282936 351816
rect 282904 351785 282905 351815
rect 282905 351785 282935 351815
rect 282935 351785 282936 351815
rect 282904 351784 282936 351785
rect 282904 351704 282936 351736
rect 282904 351655 282936 351656
rect 282904 351625 282905 351655
rect 282905 351625 282935 351655
rect 282935 351625 282936 351655
rect 282904 351624 282936 351625
rect 282984 351815 283016 351816
rect 282984 351785 282985 351815
rect 282985 351785 283015 351815
rect 283015 351785 283016 351815
rect 282984 351784 283016 351785
rect 282984 351704 283016 351736
rect 282984 351655 283016 351656
rect 282984 351625 282985 351655
rect 282985 351625 283015 351655
rect 283015 351625 283016 351655
rect 282984 351624 283016 351625
rect 283064 351815 283096 351816
rect 283064 351785 283065 351815
rect 283065 351785 283095 351815
rect 283095 351785 283096 351815
rect 283064 351784 283096 351785
rect 283064 351704 283096 351736
rect 283064 351655 283096 351656
rect 283064 351625 283065 351655
rect 283065 351625 283095 351655
rect 283095 351625 283096 351655
rect 283064 351624 283096 351625
rect 283144 351815 283176 351816
rect 283144 351785 283145 351815
rect 283145 351785 283175 351815
rect 283175 351785 283176 351815
rect 283144 351784 283176 351785
rect 283144 351704 283176 351736
rect 283144 351655 283176 351656
rect 283144 351625 283145 351655
rect 283145 351625 283175 351655
rect 283175 351625 283176 351655
rect 283144 351624 283176 351625
rect 272024 351575 272056 351576
rect 272024 351545 272025 351575
rect 272025 351545 272055 351575
rect 272055 351545 272056 351575
rect 272024 351544 272056 351545
rect 272024 351495 272056 351496
rect 272024 351465 272025 351495
rect 272025 351465 272055 351495
rect 272055 351465 272056 351495
rect 272024 351464 272056 351465
rect 272024 351415 272056 351416
rect 272024 351385 272025 351415
rect 272025 351385 272055 351415
rect 272055 351385 272056 351415
rect 272024 351384 272056 351385
rect 272024 351335 272056 351336
rect 272024 351305 272025 351335
rect 272025 351305 272055 351335
rect 272055 351305 272056 351335
rect 272024 351304 272056 351305
rect 272024 351255 272056 351256
rect 272024 351225 272025 351255
rect 272025 351225 272055 351255
rect 272055 351225 272056 351255
rect 272024 351224 272056 351225
rect 272024 351175 272056 351176
rect 272024 351145 272025 351175
rect 272025 351145 272055 351175
rect 272055 351145 272056 351175
rect 272024 351144 272056 351145
rect 272024 351095 272056 351096
rect 272024 351065 272025 351095
rect 272025 351065 272055 351095
rect 272055 351065 272056 351095
rect 272024 351064 272056 351065
rect 272024 351015 272056 351016
rect 272024 350985 272025 351015
rect 272025 350985 272055 351015
rect 272055 350985 272056 351015
rect 272024 350984 272056 350985
rect 272024 350935 272056 350936
rect 272024 350905 272025 350935
rect 272025 350905 272055 350935
rect 272055 350905 272056 350935
rect 272024 350904 272056 350905
rect 272024 350855 272056 350856
rect 272024 350825 272025 350855
rect 272025 350825 272055 350855
rect 272055 350825 272056 350855
rect 272024 350824 272056 350825
rect 272024 350775 272056 350776
rect 272024 350745 272025 350775
rect 272025 350745 272055 350775
rect 272055 350745 272056 350775
rect 272024 350744 272056 350745
rect 272024 350695 272056 350696
rect 272024 350665 272025 350695
rect 272025 350665 272055 350695
rect 272055 350665 272056 350695
rect 272024 350664 272056 350665
rect 272024 350615 272056 350616
rect 272024 350585 272025 350615
rect 272025 350585 272055 350615
rect 272055 350585 272056 350615
rect 272024 350584 272056 350585
rect 272024 350535 272056 350536
rect 272024 350505 272025 350535
rect 272025 350505 272055 350535
rect 272055 350505 272056 350535
rect 272024 350504 272056 350505
rect 272024 350455 272056 350456
rect 272024 350425 272025 350455
rect 272025 350425 272055 350455
rect 272055 350425 272056 350455
rect 272024 350424 272056 350425
rect 272024 350375 272056 350376
rect 272024 350345 272025 350375
rect 272025 350345 272055 350375
rect 272055 350345 272056 350375
rect 272024 350344 272056 350345
rect 272024 350295 272056 350296
rect 272024 350265 272025 350295
rect 272025 350265 272055 350295
rect 272055 350265 272056 350295
rect 272024 350264 272056 350265
rect 272024 350215 272056 350216
rect 272024 350185 272025 350215
rect 272025 350185 272055 350215
rect 272055 350185 272056 350215
rect 272024 350184 272056 350185
rect 272024 350135 272056 350136
rect 272024 350105 272025 350135
rect 272025 350105 272055 350135
rect 272055 350105 272056 350135
rect 272024 350104 272056 350105
rect 272024 350055 272056 350056
rect 272024 350025 272025 350055
rect 272025 350025 272055 350055
rect 272055 350025 272056 350055
rect 272024 350024 272056 350025
rect 258910 275010 259090 275190
rect 16884 274875 16916 274876
rect 16884 274845 16885 274875
rect 16885 274845 16915 274875
rect 16915 274845 16916 274875
rect 16884 274844 16916 274845
rect 16884 274555 16916 274556
rect 16884 274525 16885 274555
rect 16885 274525 16915 274555
rect 16915 274525 16916 274555
rect 16884 274524 16916 274525
rect 16884 274475 16916 274476
rect 16884 274445 16885 274475
rect 16885 274445 16915 274475
rect 16915 274445 16916 274475
rect 16884 274444 16916 274445
rect 16884 274395 16916 274396
rect 16884 274365 16885 274395
rect 16885 274365 16915 274395
rect 16915 274365 16916 274395
rect 16884 274364 16916 274365
rect 16884 274315 16916 274316
rect 16884 274285 16885 274315
rect 16885 274285 16915 274315
rect 16915 274285 16916 274315
rect 16884 274284 16916 274285
rect 16884 274235 16916 274236
rect 16884 274205 16885 274235
rect 16885 274205 16915 274235
rect 16915 274205 16916 274235
rect 16884 274204 16916 274205
rect 16884 274155 16916 274156
rect 16884 274125 16885 274155
rect 16885 274125 16915 274155
rect 16915 274125 16916 274155
rect 16884 274124 16916 274125
rect 16884 274075 16916 274076
rect 16884 274045 16885 274075
rect 16885 274045 16915 274075
rect 16915 274045 16916 274075
rect 16884 274044 16916 274045
rect 16884 273995 16916 273996
rect 16884 273965 16885 273995
rect 16885 273965 16915 273995
rect 16915 273965 16916 273995
rect 16884 273964 16916 273965
rect 16884 273915 16916 273916
rect 16884 273885 16885 273915
rect 16885 273885 16915 273915
rect 16915 273885 16916 273915
rect 16884 273884 16916 273885
rect 16884 273835 16916 273836
rect 16884 273805 16885 273835
rect 16885 273805 16915 273835
rect 16915 273805 16916 273835
rect 16884 273804 16916 273805
rect 16884 273755 16916 273756
rect 16884 273725 16885 273755
rect 16885 273725 16915 273755
rect 16915 273725 16916 273755
rect 16884 273724 16916 273725
rect 16884 273675 16916 273676
rect 16884 273645 16885 273675
rect 16885 273645 16915 273675
rect 16915 273645 16916 273675
rect 16884 273644 16916 273645
rect 16884 273595 16916 273596
rect 16884 273565 16885 273595
rect 16885 273565 16915 273595
rect 16915 273565 16916 273595
rect 16884 273564 16916 273565
rect 16884 273515 16916 273516
rect 16884 273485 16885 273515
rect 16885 273485 16915 273515
rect 16915 273485 16916 273515
rect 16884 273484 16916 273485
rect 16884 273435 16916 273436
rect 16884 273405 16885 273435
rect 16885 273405 16915 273435
rect 16915 273405 16916 273435
rect 16884 273404 16916 273405
rect 16884 273355 16916 273356
rect 16884 273325 16885 273355
rect 16885 273325 16915 273355
rect 16915 273325 16916 273355
rect 16884 273324 16916 273325
rect 16884 273275 16916 273276
rect 16884 273245 16885 273275
rect 16885 273245 16915 273275
rect 16915 273245 16916 273275
rect 16884 273244 16916 273245
rect 16884 273195 16916 273196
rect 16884 273165 16885 273195
rect 16885 273165 16915 273195
rect 16915 273165 16916 273195
rect 16884 273164 16916 273165
rect 16884 273115 16916 273116
rect 16884 273085 16885 273115
rect 16885 273085 16915 273115
rect 16915 273085 16916 273115
rect 16884 273084 16916 273085
rect 16884 273035 16916 273036
rect 16884 273005 16885 273035
rect 16885 273005 16915 273035
rect 16915 273005 16916 273035
rect 16884 273004 16916 273005
rect 16884 272955 16916 272956
rect 16884 272925 16885 272955
rect 16885 272925 16915 272955
rect 16915 272925 16916 272955
rect 16884 272924 16916 272925
rect 16884 272875 16916 272876
rect 16884 272845 16885 272875
rect 16885 272845 16915 272875
rect 16915 272845 16916 272875
rect 16884 272844 16916 272845
rect 16884 272795 16916 272796
rect 16884 272765 16885 272795
rect 16885 272765 16915 272795
rect 16915 272765 16916 272795
rect 16884 272764 16916 272765
rect 16884 272715 16916 272716
rect 16884 272685 16885 272715
rect 16885 272685 16915 272715
rect 16915 272685 16916 272715
rect 16884 272684 16916 272685
rect 16884 272635 16916 272636
rect 16884 272605 16885 272635
rect 16885 272605 16915 272635
rect 16915 272605 16916 272635
rect 16884 272604 16916 272605
rect 16884 272555 16916 272556
rect 16884 272525 16885 272555
rect 16885 272525 16915 272555
rect 16915 272525 16916 272555
rect 16884 272524 16916 272525
rect 16884 272475 16916 272476
rect 16884 272445 16885 272475
rect 16885 272445 16915 272475
rect 16915 272445 16916 272475
rect 16884 272444 16916 272445
rect 16884 272395 16916 272396
rect 16884 272365 16885 272395
rect 16885 272365 16915 272395
rect 16915 272365 16916 272395
rect 16884 272364 16916 272365
rect 16884 272315 16916 272316
rect 16884 272285 16885 272315
rect 16885 272285 16915 272315
rect 16915 272285 16916 272315
rect 16884 272284 16916 272285
rect 16884 272235 16916 272236
rect 16884 272205 16885 272235
rect 16885 272205 16915 272235
rect 16915 272205 16916 272235
rect 16884 272204 16916 272205
rect 16884 272155 16916 272156
rect 16884 272125 16885 272155
rect 16885 272125 16915 272155
rect 16915 272125 16916 272155
rect 16884 272124 16916 272125
rect 16884 272075 16916 272076
rect 16884 272045 16885 272075
rect 16885 272045 16915 272075
rect 16915 272045 16916 272075
rect 16884 272044 16916 272045
rect 16884 271995 16916 271996
rect 16884 271965 16885 271995
rect 16885 271965 16915 271995
rect 16915 271965 16916 271995
rect 16884 271964 16916 271965
rect 16884 271915 16916 271916
rect 16884 271885 16885 271915
rect 16885 271885 16915 271915
rect 16915 271885 16916 271915
rect 16884 271884 16916 271885
rect 16884 271835 16916 271836
rect 16884 271805 16885 271835
rect 16885 271805 16915 271835
rect 16915 271805 16916 271835
rect 16884 271804 16916 271805
rect 16884 271755 16916 271756
rect 16884 271725 16885 271755
rect 16885 271725 16915 271755
rect 16915 271725 16916 271755
rect 16884 271724 16916 271725
rect 16884 271675 16916 271676
rect 16884 271645 16885 271675
rect 16885 271645 16915 271675
rect 16915 271645 16916 271675
rect 16884 271644 16916 271645
rect 16884 271595 16916 271596
rect 16884 271565 16885 271595
rect 16885 271565 16915 271595
rect 16915 271565 16916 271595
rect 16884 271564 16916 271565
rect 16884 271515 16916 271516
rect 16884 271485 16885 271515
rect 16885 271485 16915 271515
rect 16915 271485 16916 271515
rect 16884 271484 16916 271485
rect 16884 271435 16916 271436
rect 16884 271405 16885 271435
rect 16885 271405 16915 271435
rect 16915 271405 16916 271435
rect 16884 271404 16916 271405
rect 16884 271355 16916 271356
rect 16884 271325 16885 271355
rect 16885 271325 16915 271355
rect 16915 271325 16916 271355
rect 16884 271324 16916 271325
rect 16884 271275 16916 271276
rect 16884 271245 16885 271275
rect 16885 271245 16915 271275
rect 16915 271245 16916 271275
rect 16884 271244 16916 271245
rect 16884 271195 16916 271196
rect 16884 271165 16885 271195
rect 16885 271165 16915 271195
rect 16915 271165 16916 271195
rect 16884 271164 16916 271165
rect 16884 271115 16916 271116
rect 16884 271085 16885 271115
rect 16885 271085 16915 271115
rect 16915 271085 16916 271115
rect 16884 271084 16916 271085
rect 16884 271035 16916 271036
rect 16884 271005 16885 271035
rect 16885 271005 16915 271035
rect 16915 271005 16916 271035
rect 16884 271004 16916 271005
rect 16884 270955 16916 270956
rect 16884 270925 16885 270955
rect 16885 270925 16915 270955
rect 16915 270925 16916 270955
rect 16884 270924 16916 270925
rect 16884 270875 16916 270876
rect 16884 270845 16885 270875
rect 16885 270845 16915 270875
rect 16915 270845 16916 270875
rect 16884 270844 16916 270845
rect 16884 270795 16916 270796
rect 16884 270765 16885 270795
rect 16885 270765 16915 270795
rect 16915 270765 16916 270795
rect 16884 270764 16916 270765
rect 16884 270715 16916 270716
rect 16884 270685 16885 270715
rect 16885 270685 16915 270715
rect 16915 270685 16916 270715
rect 16884 270684 16916 270685
rect 16884 270635 16916 270636
rect 16884 270605 16885 270635
rect 16885 270605 16915 270635
rect 16915 270605 16916 270635
rect 16884 270604 16916 270605
rect 16884 270555 16916 270556
rect 16884 270525 16885 270555
rect 16885 270525 16915 270555
rect 16915 270525 16916 270555
rect 16884 270524 16916 270525
rect 16884 270475 16916 270476
rect 16884 270445 16885 270475
rect 16885 270445 16915 270475
rect 16915 270445 16916 270475
rect 16884 270444 16916 270445
rect 16884 270395 16916 270396
rect 16884 270365 16885 270395
rect 16885 270365 16915 270395
rect 16915 270365 16916 270395
rect 16884 270364 16916 270365
rect 16884 270315 16916 270316
rect 16884 270285 16885 270315
rect 16885 270285 16915 270315
rect 16915 270285 16916 270315
rect 16884 270284 16916 270285
rect 16884 270235 16916 270236
rect 16884 270205 16885 270235
rect 16885 270205 16915 270235
rect 16915 270205 16916 270235
rect 16884 270204 16916 270205
rect 16884 270155 16916 270156
rect 16884 270125 16885 270155
rect 16885 270125 16915 270155
rect 16915 270125 16916 270155
rect 16884 270124 16916 270125
rect 16884 270075 16916 270076
rect 16884 270045 16885 270075
rect 16885 270045 16915 270075
rect 16915 270045 16916 270075
rect 16884 270044 16916 270045
rect 16884 269995 16916 269996
rect 16884 269965 16885 269995
rect 16885 269965 16915 269995
rect 16915 269965 16916 269995
rect 16884 269964 16916 269965
rect 16884 269915 16916 269916
rect 16884 269885 16885 269915
rect 16885 269885 16915 269915
rect 16915 269885 16916 269915
rect 16884 269884 16916 269885
rect 16884 269835 16916 269836
rect 16884 269805 16885 269835
rect 16885 269805 16915 269835
rect 16915 269805 16916 269835
rect 16884 269804 16916 269805
rect 16884 269755 16916 269756
rect 16884 269725 16885 269755
rect 16885 269725 16915 269755
rect 16915 269725 16916 269755
rect 16884 269724 16916 269725
rect 16884 269675 16916 269676
rect 16884 269645 16885 269675
rect 16885 269645 16915 269675
rect 16915 269645 16916 269675
rect 16884 269644 16916 269645
rect 16884 269595 16916 269596
rect 16884 269565 16885 269595
rect 16885 269565 16915 269595
rect 16915 269565 16916 269595
rect 16884 269564 16916 269565
rect 16884 269515 16916 269516
rect 16884 269485 16885 269515
rect 16885 269485 16915 269515
rect 16915 269485 16916 269515
rect 16884 269484 16916 269485
rect 16884 269435 16916 269436
rect 16884 269405 16885 269435
rect 16885 269405 16915 269435
rect 16915 269405 16916 269435
rect 16884 269404 16916 269405
rect 16884 269355 16916 269356
rect 16884 269325 16885 269355
rect 16885 269325 16915 269355
rect 16915 269325 16916 269355
rect 16884 269324 16916 269325
rect 16884 269275 16916 269276
rect 16884 269245 16885 269275
rect 16885 269245 16915 269275
rect 16915 269245 16916 269275
rect 16884 269244 16916 269245
rect 16884 269195 16916 269196
rect 16884 269165 16885 269195
rect 16885 269165 16915 269195
rect 16915 269165 16916 269195
rect 16884 269164 16916 269165
rect 16884 269115 16916 269116
rect 16884 269085 16885 269115
rect 16885 269085 16915 269115
rect 16915 269085 16916 269115
rect 16884 269084 16916 269085
rect 16884 269035 16916 269036
rect 16884 269005 16885 269035
rect 16885 269005 16915 269035
rect 16915 269005 16916 269035
rect 16884 269004 16916 269005
rect 16884 268955 16916 268956
rect 16884 268925 16885 268955
rect 16885 268925 16915 268955
rect 16915 268925 16916 268955
rect 16884 268924 16916 268925
rect 16884 268875 16916 268876
rect 16884 268845 16885 268875
rect 16885 268845 16915 268875
rect 16915 268845 16916 268875
rect 16884 268844 16916 268845
rect 16884 268795 16916 268796
rect 16884 268765 16885 268795
rect 16885 268765 16915 268795
rect 16915 268765 16916 268795
rect 16884 268764 16916 268765
rect 16884 268715 16916 268716
rect 16884 268685 16885 268715
rect 16885 268685 16915 268715
rect 16915 268685 16916 268715
rect 16884 268684 16916 268685
rect 16884 268635 16916 268636
rect 16884 268605 16885 268635
rect 16885 268605 16915 268635
rect 16915 268605 16916 268635
rect 16884 268604 16916 268605
rect 16884 268555 16916 268556
rect 16884 268525 16885 268555
rect 16885 268525 16915 268555
rect 16915 268525 16916 268555
rect 16884 268524 16916 268525
rect 16884 268475 16916 268476
rect 16884 268445 16885 268475
rect 16885 268445 16915 268475
rect 16915 268445 16916 268475
rect 16884 268444 16916 268445
rect 16884 268395 16916 268396
rect 16884 268365 16885 268395
rect 16885 268365 16915 268395
rect 16915 268365 16916 268395
rect 16884 268364 16916 268365
rect 16884 268315 16916 268316
rect 16884 268285 16885 268315
rect 16885 268285 16915 268315
rect 16915 268285 16916 268315
rect 16884 268284 16916 268285
rect 16884 268235 16916 268236
rect 16884 268205 16885 268235
rect 16885 268205 16915 268235
rect 16915 268205 16916 268235
rect 16884 268204 16916 268205
rect 16884 268155 16916 268156
rect 16884 268125 16885 268155
rect 16885 268125 16915 268155
rect 16915 268125 16916 268155
rect 16884 268124 16916 268125
rect 16884 268075 16916 268076
rect 16884 268045 16885 268075
rect 16885 268045 16915 268075
rect 16915 268045 16916 268075
rect 16884 268044 16916 268045
rect 16884 267995 16916 267996
rect 16884 267965 16885 267995
rect 16885 267965 16915 267995
rect 16915 267965 16916 267995
rect 16884 267964 16916 267965
rect 16884 267915 16916 267916
rect 16884 267885 16885 267915
rect 16885 267885 16915 267915
rect 16915 267885 16916 267915
rect 16884 267884 16916 267885
rect 16884 267835 16916 267836
rect 16884 267805 16885 267835
rect 16885 267805 16915 267835
rect 16915 267805 16916 267835
rect 16884 267804 16916 267805
rect 16884 267755 16916 267756
rect 16884 267725 16885 267755
rect 16885 267725 16915 267755
rect 16915 267725 16916 267755
rect 16884 267724 16916 267725
rect 16884 267675 16916 267676
rect 16884 267645 16885 267675
rect 16885 267645 16915 267675
rect 16915 267645 16916 267675
rect 16884 267644 16916 267645
rect 16884 267595 16916 267596
rect 16884 267565 16885 267595
rect 16885 267565 16915 267595
rect 16915 267565 16916 267595
rect 16884 267564 16916 267565
rect 16884 267515 16916 267516
rect 16884 267485 16885 267515
rect 16885 267485 16915 267515
rect 16915 267485 16916 267515
rect 16884 267484 16916 267485
rect 16884 267435 16916 267436
rect 16884 267405 16885 267435
rect 16885 267405 16915 267435
rect 16915 267405 16916 267435
rect 16884 267404 16916 267405
rect 16884 267355 16916 267356
rect 16884 267325 16885 267355
rect 16885 267325 16915 267355
rect 16915 267325 16916 267355
rect 16884 267324 16916 267325
rect 16884 267275 16916 267276
rect 16884 267245 16885 267275
rect 16885 267245 16915 267275
rect 16915 267245 16916 267275
rect 16884 267244 16916 267245
rect 16884 267195 16916 267196
rect 16884 267165 16885 267195
rect 16885 267165 16915 267195
rect 16915 267165 16916 267195
rect 16884 267164 16916 267165
rect 16884 267115 16916 267116
rect 16884 267085 16885 267115
rect 16885 267085 16915 267115
rect 16915 267085 16916 267115
rect 16884 267084 16916 267085
rect 16884 267035 16916 267036
rect 16884 267005 16885 267035
rect 16885 267005 16915 267035
rect 16915 267005 16916 267035
rect 16884 267004 16916 267005
rect 16884 266955 16916 266956
rect 16884 266925 16885 266955
rect 16885 266925 16915 266955
rect 16915 266925 16916 266955
rect 16884 266924 16916 266925
rect 16884 266875 16916 266876
rect 16884 266845 16885 266875
rect 16885 266845 16915 266875
rect 16915 266845 16916 266875
rect 16884 266844 16916 266845
rect 16884 266795 16916 266796
rect 16884 266765 16885 266795
rect 16885 266765 16915 266795
rect 16915 266765 16916 266795
rect 16884 266764 16916 266765
rect 16884 266715 16916 266716
rect 16884 266685 16885 266715
rect 16885 266685 16915 266715
rect 16915 266685 16916 266715
rect 16884 266684 16916 266685
rect 16884 266635 16916 266636
rect 16884 266605 16885 266635
rect 16885 266605 16915 266635
rect 16915 266605 16916 266635
rect 16884 266604 16916 266605
rect 16884 266555 16916 266556
rect 16884 266525 16885 266555
rect 16885 266525 16915 266555
rect 16915 266525 16916 266555
rect 16884 266524 16916 266525
rect 16884 266475 16916 266476
rect 16884 266445 16885 266475
rect 16885 266445 16915 266475
rect 16915 266445 16916 266475
rect 16884 266444 16916 266445
rect 16884 266395 16916 266396
rect 16884 266365 16885 266395
rect 16885 266365 16915 266395
rect 16915 266365 16916 266395
rect 16884 266364 16916 266365
rect 16884 266315 16916 266316
rect 16884 266285 16885 266315
rect 16885 266285 16915 266315
rect 16915 266285 16916 266315
rect 16884 266284 16916 266285
rect 16884 266235 16916 266236
rect 16884 266205 16885 266235
rect 16885 266205 16915 266235
rect 16915 266205 16916 266235
rect 16884 266204 16916 266205
rect 16884 266155 16916 266156
rect 16884 266125 16885 266155
rect 16885 266125 16915 266155
rect 16915 266125 16916 266155
rect 16884 266124 16916 266125
rect 16884 266075 16916 266076
rect 16884 266045 16885 266075
rect 16885 266045 16915 266075
rect 16915 266045 16916 266075
rect 16884 266044 16916 266045
rect 16884 265995 16916 265996
rect 16884 265965 16885 265995
rect 16885 265965 16915 265995
rect 16915 265965 16916 265995
rect 16884 265964 16916 265965
rect 16884 265915 16916 265916
rect 16884 265885 16885 265915
rect 16885 265885 16915 265915
rect 16915 265885 16916 265915
rect 16884 265884 16916 265885
rect 16884 265835 16916 265836
rect 16884 265805 16885 265835
rect 16885 265805 16915 265835
rect 16915 265805 16916 265835
rect 16884 265804 16916 265805
rect 16884 265755 16916 265756
rect 16884 265725 16885 265755
rect 16885 265725 16915 265755
rect 16915 265725 16916 265755
rect 16884 265724 16916 265725
rect 16884 265675 16916 265676
rect 16884 265645 16885 265675
rect 16885 265645 16915 265675
rect 16915 265645 16916 265675
rect 16884 265644 16916 265645
rect 16884 265595 16916 265596
rect 16884 265565 16885 265595
rect 16885 265565 16915 265595
rect 16915 265565 16916 265595
rect 16884 265564 16916 265565
rect 16884 265515 16916 265516
rect 16884 265485 16885 265515
rect 16885 265485 16915 265515
rect 16915 265485 16916 265515
rect 16884 265484 16916 265485
rect 16884 265435 16916 265436
rect 16884 265405 16885 265435
rect 16885 265405 16915 265435
rect 16915 265405 16916 265435
rect 16884 265404 16916 265405
rect 16884 265355 16916 265356
rect 16884 265325 16885 265355
rect 16885 265325 16915 265355
rect 16915 265325 16916 265355
rect 16884 265324 16916 265325
rect 16884 265275 16916 265276
rect 16884 265245 16885 265275
rect 16885 265245 16915 265275
rect 16915 265245 16916 265275
rect 16884 265244 16916 265245
rect 16884 265195 16916 265196
rect 16884 265165 16885 265195
rect 16885 265165 16915 265195
rect 16915 265165 16916 265195
rect 16884 265164 16916 265165
rect 16884 265115 16916 265116
rect 16884 265085 16885 265115
rect 16885 265085 16915 265115
rect 16915 265085 16916 265115
rect 16884 265084 16916 265085
rect 16884 265035 16916 265036
rect 16884 265005 16885 265035
rect 16885 265005 16915 265035
rect 16915 265005 16916 265035
rect 16884 265004 16916 265005
rect 16884 264955 16916 264956
rect 16884 264925 16885 264955
rect 16885 264925 16915 264955
rect 16915 264925 16916 264955
rect 16884 264924 16916 264925
rect 16884 264875 16916 264876
rect 16884 264845 16885 264875
rect 16885 264845 16915 264875
rect 16915 264845 16916 264875
rect 16884 264844 16916 264845
rect 16884 264795 16916 264796
rect 16884 264765 16885 264795
rect 16885 264765 16915 264795
rect 16915 264765 16916 264795
rect 16884 264764 16916 264765
rect 16884 264715 16916 264716
rect 16884 264685 16885 264715
rect 16885 264685 16915 264715
rect 16915 264685 16916 264715
rect 16884 264684 16916 264685
rect 16884 264635 16916 264636
rect 16884 264605 16885 264635
rect 16885 264605 16915 264635
rect 16915 264605 16916 264635
rect 16884 264604 16916 264605
rect 16884 264555 16916 264556
rect 16884 264525 16885 264555
rect 16885 264525 16915 264555
rect 16915 264525 16916 264555
rect 16884 264524 16916 264525
rect 16884 264475 16916 264476
rect 16884 264445 16885 264475
rect 16885 264445 16915 264475
rect 16915 264445 16916 264475
rect 16884 264444 16916 264445
rect 16884 264395 16916 264396
rect 16884 264365 16885 264395
rect 16885 264365 16915 264395
rect 16915 264365 16916 264395
rect 16884 264364 16916 264365
rect 16884 264315 16916 264316
rect 16884 264285 16885 264315
rect 16885 264285 16915 264315
rect 16915 264285 16916 264315
rect 16884 264284 16916 264285
rect 16884 264235 16916 264236
rect 16884 264205 16885 264235
rect 16885 264205 16915 264235
rect 16915 264205 16916 264235
rect 16884 264204 16916 264205
rect 16884 264155 16916 264156
rect 16884 264125 16885 264155
rect 16885 264125 16915 264155
rect 16915 264125 16916 264155
rect 16884 264124 16916 264125
rect 16884 264075 16916 264076
rect 16884 264045 16885 264075
rect 16885 264045 16915 264075
rect 16915 264045 16916 264075
rect 16884 264044 16916 264045
rect 16884 263995 16916 263996
rect 16884 263965 16885 263995
rect 16885 263965 16915 263995
rect 16915 263965 16916 263995
rect 16884 263964 16916 263965
rect 16884 263915 16916 263916
rect 16884 263885 16885 263915
rect 16885 263885 16915 263915
rect 16915 263885 16916 263915
rect 16884 263884 16916 263885
rect 16884 263835 16916 263836
rect 16884 263805 16885 263835
rect 16885 263805 16915 263835
rect 16915 263805 16916 263835
rect 16884 263804 16916 263805
rect 16884 263755 16916 263756
rect 16884 263725 16885 263755
rect 16885 263725 16915 263755
rect 16915 263725 16916 263755
rect 16884 263724 16916 263725
rect 16884 263675 16916 263676
rect 16884 263645 16885 263675
rect 16885 263645 16915 263675
rect 16915 263645 16916 263675
rect 16884 263644 16916 263645
rect 16884 263595 16916 263596
rect 16884 263565 16885 263595
rect 16885 263565 16915 263595
rect 16915 263565 16916 263595
rect 16884 263564 16916 263565
rect 16884 263515 16916 263516
rect 16884 263485 16885 263515
rect 16885 263485 16915 263515
rect 16915 263485 16916 263515
rect 16884 263484 16916 263485
rect 16884 263435 16916 263436
rect 16884 263405 16885 263435
rect 16885 263405 16915 263435
rect 16915 263405 16916 263435
rect 16884 263404 16916 263405
rect 16884 263355 16916 263356
rect 16884 263325 16885 263355
rect 16885 263325 16915 263355
rect 16915 263325 16916 263355
rect 16884 263324 16916 263325
rect 16884 263275 16916 263276
rect 16884 263245 16885 263275
rect 16885 263245 16915 263275
rect 16915 263245 16916 263275
rect 16884 263244 16916 263245
rect 16884 263195 16916 263196
rect 16884 263165 16885 263195
rect 16885 263165 16915 263195
rect 16915 263165 16916 263195
rect 16884 263164 16916 263165
rect 16884 263115 16916 263116
rect 16884 263085 16885 263115
rect 16885 263085 16915 263115
rect 16915 263085 16916 263115
rect 16884 263084 16916 263085
rect 16884 263035 16916 263036
rect 16884 263005 16885 263035
rect 16885 263005 16915 263035
rect 16915 263005 16916 263035
rect 16884 263004 16916 263005
rect 16884 262955 16916 262956
rect 16884 262925 16885 262955
rect 16885 262925 16915 262955
rect 16915 262925 16916 262955
rect 16884 262924 16916 262925
rect 16884 262875 16916 262876
rect 16884 262845 16885 262875
rect 16885 262845 16915 262875
rect 16915 262845 16916 262875
rect 16884 262844 16916 262845
rect 16884 262795 16916 262796
rect 16884 262765 16885 262795
rect 16885 262765 16915 262795
rect 16915 262765 16916 262795
rect 16884 262764 16916 262765
rect 16884 262715 16916 262716
rect 16884 262685 16885 262715
rect 16885 262685 16915 262715
rect 16915 262685 16916 262715
rect 16884 262684 16916 262685
rect 16884 262635 16916 262636
rect 16884 262605 16885 262635
rect 16885 262605 16915 262635
rect 16915 262605 16916 262635
rect 16884 262604 16916 262605
rect 16884 262555 16916 262556
rect 16884 262525 16885 262555
rect 16885 262525 16915 262555
rect 16915 262525 16916 262555
rect 16884 262524 16916 262525
rect 16884 262475 16916 262476
rect 16884 262445 16885 262475
rect 16885 262445 16915 262475
rect 16915 262445 16916 262475
rect 16884 262444 16916 262445
rect 16884 262395 16916 262396
rect 16884 262365 16885 262395
rect 16885 262365 16915 262395
rect 16915 262365 16916 262395
rect 16884 262364 16916 262365
rect 16884 262315 16916 262316
rect 16884 262285 16885 262315
rect 16885 262285 16915 262315
rect 16915 262285 16916 262315
rect 16884 262284 16916 262285
rect 16884 262235 16916 262236
rect 16884 262205 16885 262235
rect 16885 262205 16915 262235
rect 16915 262205 16916 262235
rect 16884 262204 16916 262205
rect 16884 262155 16916 262156
rect 16884 262125 16885 262155
rect 16885 262125 16915 262155
rect 16915 262125 16916 262155
rect 16884 262124 16916 262125
rect 16884 262075 16916 262076
rect 16884 262045 16885 262075
rect 16885 262045 16915 262075
rect 16915 262045 16916 262075
rect 16884 262044 16916 262045
rect 16884 261995 16916 261996
rect 16884 261965 16885 261995
rect 16885 261965 16915 261995
rect 16915 261965 16916 261995
rect 16884 261964 16916 261965
rect 16884 261915 16916 261916
rect 16884 261885 16885 261915
rect 16885 261885 16915 261915
rect 16915 261885 16916 261915
rect 16884 261884 16916 261885
rect 16884 261835 16916 261836
rect 16884 261805 16885 261835
rect 16885 261805 16915 261835
rect 16915 261805 16916 261835
rect 16884 261804 16916 261805
rect 16884 261755 16916 261756
rect 16884 261725 16885 261755
rect 16885 261725 16915 261755
rect 16915 261725 16916 261755
rect 16884 261724 16916 261725
rect 16884 261675 16916 261676
rect 16884 261645 16885 261675
rect 16885 261645 16915 261675
rect 16915 261645 16916 261675
rect 16884 261644 16916 261645
rect 16884 261595 16916 261596
rect 16884 261565 16885 261595
rect 16885 261565 16915 261595
rect 16915 261565 16916 261595
rect 16884 261564 16916 261565
rect 16884 261515 16916 261516
rect 16884 261485 16885 261515
rect 16885 261485 16915 261515
rect 16915 261485 16916 261515
rect 16884 261484 16916 261485
rect 16884 261435 16916 261436
rect 16884 261405 16885 261435
rect 16885 261405 16915 261435
rect 16915 261405 16916 261435
rect 16884 261404 16916 261405
rect 16884 261355 16916 261356
rect 16884 261325 16885 261355
rect 16885 261325 16915 261355
rect 16915 261325 16916 261355
rect 16884 261324 16916 261325
rect 16884 261275 16916 261276
rect 16884 261245 16885 261275
rect 16885 261245 16915 261275
rect 16915 261245 16916 261275
rect 16884 261244 16916 261245
rect 16884 261195 16916 261196
rect 16884 261165 16885 261195
rect 16885 261165 16915 261195
rect 16915 261165 16916 261195
rect 16884 261164 16916 261165
rect 16884 261115 16916 261116
rect 16884 261085 16885 261115
rect 16885 261085 16915 261115
rect 16915 261085 16916 261115
rect 16884 261084 16916 261085
rect 16884 261035 16916 261036
rect 16884 261005 16885 261035
rect 16885 261005 16915 261035
rect 16915 261005 16916 261035
rect 16884 261004 16916 261005
rect 16884 260955 16916 260956
rect 16884 260925 16885 260955
rect 16885 260925 16915 260955
rect 16915 260925 16916 260955
rect 16884 260924 16916 260925
rect 16884 260875 16916 260876
rect 16884 260845 16885 260875
rect 16885 260845 16915 260875
rect 16915 260845 16916 260875
rect 16884 260844 16916 260845
rect 16884 260795 16916 260796
rect 16884 260765 16885 260795
rect 16885 260765 16915 260795
rect 16915 260765 16916 260795
rect 16884 260764 16916 260765
rect 16884 260715 16916 260716
rect 16884 260685 16885 260715
rect 16885 260685 16915 260715
rect 16915 260685 16916 260715
rect 16884 260684 16916 260685
rect 16884 260635 16916 260636
rect 16884 260605 16885 260635
rect 16885 260605 16915 260635
rect 16915 260605 16916 260635
rect 16884 260604 16916 260605
rect 16884 260555 16916 260556
rect 16884 260525 16885 260555
rect 16885 260525 16915 260555
rect 16915 260525 16916 260555
rect 16884 260524 16916 260525
rect 16884 260475 16916 260476
rect 16884 260445 16885 260475
rect 16885 260445 16915 260475
rect 16915 260445 16916 260475
rect 16884 260444 16916 260445
rect 16884 260395 16916 260396
rect 16884 260365 16885 260395
rect 16885 260365 16915 260395
rect 16915 260365 16916 260395
rect 16884 260364 16916 260365
rect 16884 260315 16916 260316
rect 16884 260285 16885 260315
rect 16885 260285 16915 260315
rect 16915 260285 16916 260315
rect 16884 260284 16916 260285
rect 16884 260235 16916 260236
rect 16884 260205 16885 260235
rect 16885 260205 16915 260235
rect 16915 260205 16916 260235
rect 16884 260204 16916 260205
rect 16884 260155 16916 260156
rect 16884 260125 16885 260155
rect 16885 260125 16915 260155
rect 16915 260125 16916 260155
rect 16884 260124 16916 260125
rect 16884 260075 16916 260076
rect 16884 260045 16885 260075
rect 16885 260045 16915 260075
rect 16915 260045 16916 260075
rect 16884 260044 16916 260045
rect 16884 259995 16916 259996
rect 16884 259965 16885 259995
rect 16885 259965 16915 259995
rect 16915 259965 16916 259995
rect 16884 259964 16916 259965
rect 16884 259915 16916 259916
rect 16884 259885 16885 259915
rect 16885 259885 16915 259915
rect 16915 259885 16916 259915
rect 16884 259884 16916 259885
rect 16884 259835 16916 259836
rect 16884 259805 16885 259835
rect 16885 259805 16915 259835
rect 16915 259805 16916 259835
rect 16884 259804 16916 259805
rect 16884 259755 16916 259756
rect 16884 259725 16885 259755
rect 16885 259725 16915 259755
rect 16915 259725 16916 259755
rect 16884 259724 16916 259725
rect 16884 259675 16916 259676
rect 16884 259645 16885 259675
rect 16885 259645 16915 259675
rect 16915 259645 16916 259675
rect 16884 259644 16916 259645
rect 16884 259595 16916 259596
rect 16884 259565 16885 259595
rect 16885 259565 16915 259595
rect 16915 259565 16916 259595
rect 16884 259564 16916 259565
rect 16884 259515 16916 259516
rect 16884 259485 16885 259515
rect 16885 259485 16915 259515
rect 16915 259485 16916 259515
rect 16884 259484 16916 259485
rect 16884 259435 16916 259436
rect 16884 259405 16885 259435
rect 16885 259405 16915 259435
rect 16915 259405 16916 259435
rect 16884 259404 16916 259405
rect 16884 259355 16916 259356
rect 16884 259325 16885 259355
rect 16885 259325 16915 259355
rect 16915 259325 16916 259355
rect 16884 259324 16916 259325
rect 16884 259275 16916 259276
rect 16884 259245 16885 259275
rect 16885 259245 16915 259275
rect 16915 259245 16916 259275
rect 16884 259244 16916 259245
rect 16884 259195 16916 259196
rect 16884 259165 16885 259195
rect 16885 259165 16915 259195
rect 16915 259165 16916 259195
rect 16884 259164 16916 259165
rect 16884 259115 16916 259116
rect 16884 259085 16885 259115
rect 16885 259085 16915 259115
rect 16915 259085 16916 259115
rect 16884 259084 16916 259085
rect 16884 259035 16916 259036
rect 16884 259005 16885 259035
rect 16885 259005 16915 259035
rect 16915 259005 16916 259035
rect 16884 259004 16916 259005
rect 16884 258955 16916 258956
rect 16884 258925 16885 258955
rect 16885 258925 16915 258955
rect 16915 258925 16916 258955
rect 16884 258924 16916 258925
rect 16884 258875 16916 258876
rect 16884 258845 16885 258875
rect 16885 258845 16915 258875
rect 16915 258845 16916 258875
rect 16884 258844 16916 258845
rect 16884 258795 16916 258796
rect 16884 258765 16885 258795
rect 16885 258765 16915 258795
rect 16915 258765 16916 258795
rect 16884 258764 16916 258765
rect 16884 258715 16916 258716
rect 16884 258685 16885 258715
rect 16885 258685 16915 258715
rect 16915 258685 16916 258715
rect 16884 258684 16916 258685
rect 16884 258635 16916 258636
rect 16884 258605 16885 258635
rect 16885 258605 16915 258635
rect 16915 258605 16916 258635
rect 16884 258604 16916 258605
rect 16884 258555 16916 258556
rect 16884 258525 16885 258555
rect 16885 258525 16915 258555
rect 16915 258525 16916 258555
rect 16884 258524 16916 258525
rect 16884 258475 16916 258476
rect 16884 258445 16885 258475
rect 16885 258445 16915 258475
rect 16915 258445 16916 258475
rect 16884 258444 16916 258445
rect 16884 258395 16916 258396
rect 16884 258365 16885 258395
rect 16885 258365 16915 258395
rect 16915 258365 16916 258395
rect 16884 258364 16916 258365
rect 16884 258315 16916 258316
rect 16884 258285 16885 258315
rect 16885 258285 16915 258315
rect 16915 258285 16916 258315
rect 16884 258284 16916 258285
rect 16884 258235 16916 258236
rect 16884 258205 16885 258235
rect 16885 258205 16915 258235
rect 16915 258205 16916 258235
rect 16884 258204 16916 258205
rect 16884 258155 16916 258156
rect 16884 258125 16885 258155
rect 16885 258125 16915 258155
rect 16915 258125 16916 258155
rect 16884 258124 16916 258125
rect 16884 258075 16916 258076
rect 16884 258045 16885 258075
rect 16885 258045 16915 258075
rect 16915 258045 16916 258075
rect 16884 258044 16916 258045
rect 16884 257995 16916 257996
rect 16884 257965 16885 257995
rect 16885 257965 16915 257995
rect 16915 257965 16916 257995
rect 16884 257964 16916 257965
rect 16884 257915 16916 257916
rect 16884 257885 16885 257915
rect 16885 257885 16915 257915
rect 16915 257885 16916 257915
rect 16884 257884 16916 257885
rect 16884 257835 16916 257836
rect 16884 257805 16885 257835
rect 16885 257805 16915 257835
rect 16915 257805 16916 257835
rect 16884 257804 16916 257805
rect 16884 257755 16916 257756
rect 16884 257725 16885 257755
rect 16885 257725 16915 257755
rect 16915 257725 16916 257755
rect 16884 257724 16916 257725
rect 16884 257675 16916 257676
rect 16884 257645 16885 257675
rect 16885 257645 16915 257675
rect 16915 257645 16916 257675
rect 16884 257644 16916 257645
rect 16884 257595 16916 257596
rect 16884 257565 16885 257595
rect 16885 257565 16915 257595
rect 16915 257565 16916 257595
rect 16884 257564 16916 257565
rect 16884 257515 16916 257516
rect 16884 257485 16885 257515
rect 16885 257485 16915 257515
rect 16915 257485 16916 257515
rect 16884 257484 16916 257485
rect 16884 257435 16916 257436
rect 16884 257405 16885 257435
rect 16885 257405 16915 257435
rect 16915 257405 16916 257435
rect 16884 257404 16916 257405
rect 16884 257355 16916 257356
rect 16884 257325 16885 257355
rect 16885 257325 16915 257355
rect 16915 257325 16916 257355
rect 16884 257324 16916 257325
rect 16884 257275 16916 257276
rect 16884 257245 16885 257275
rect 16885 257245 16915 257275
rect 16915 257245 16916 257275
rect 16884 257244 16916 257245
rect 16884 257195 16916 257196
rect 16884 257165 16885 257195
rect 16885 257165 16915 257195
rect 16915 257165 16916 257195
rect 16884 257164 16916 257165
rect 16884 257115 16916 257116
rect 16884 257085 16885 257115
rect 16885 257085 16915 257115
rect 16915 257085 16916 257115
rect 16884 257084 16916 257085
rect 16884 257035 16916 257036
rect 16884 257005 16885 257035
rect 16885 257005 16915 257035
rect 16915 257005 16916 257035
rect 16884 257004 16916 257005
rect 16884 256955 16916 256956
rect 16884 256925 16885 256955
rect 16885 256925 16915 256955
rect 16915 256925 16916 256955
rect 16884 256924 16916 256925
rect 16884 256875 16916 256876
rect 16884 256845 16885 256875
rect 16885 256845 16915 256875
rect 16915 256845 16916 256875
rect 16884 256844 16916 256845
rect 16884 256795 16916 256796
rect 16884 256765 16885 256795
rect 16885 256765 16915 256795
rect 16915 256765 16916 256795
rect 16884 256764 16916 256765
rect 16884 256715 16916 256716
rect 16884 256685 16885 256715
rect 16885 256685 16915 256715
rect 16915 256685 16916 256715
rect 16884 256684 16916 256685
rect 16884 256635 16916 256636
rect 16884 256605 16885 256635
rect 16885 256605 16915 256635
rect 16915 256605 16916 256635
rect 16884 256604 16916 256605
rect 16884 256555 16916 256556
rect 16884 256525 16885 256555
rect 16885 256525 16915 256555
rect 16915 256525 16916 256555
rect 16884 256524 16916 256525
rect 16884 256475 16916 256476
rect 16884 256445 16885 256475
rect 16885 256445 16915 256475
rect 16915 256445 16916 256475
rect 16884 256444 16916 256445
rect 16884 256395 16916 256396
rect 16884 256365 16885 256395
rect 16885 256365 16915 256395
rect 16915 256365 16916 256395
rect 16884 256364 16916 256365
rect 16884 256315 16916 256316
rect 16884 256285 16885 256315
rect 16885 256285 16915 256315
rect 16915 256285 16916 256315
rect 16884 256284 16916 256285
rect 16884 256235 16916 256236
rect 16884 256205 16885 256235
rect 16885 256205 16915 256235
rect 16915 256205 16916 256235
rect 16884 256204 16916 256205
rect 16884 256155 16916 256156
rect 16884 256125 16885 256155
rect 16885 256125 16915 256155
rect 16915 256125 16916 256155
rect 16884 256124 16916 256125
rect 16884 256075 16916 256076
rect 16884 256045 16885 256075
rect 16885 256045 16915 256075
rect 16915 256045 16916 256075
rect 16884 256044 16916 256045
rect 16884 255995 16916 255996
rect 16884 255965 16885 255995
rect 16885 255965 16915 255995
rect 16915 255965 16916 255995
rect 16884 255964 16916 255965
rect 16884 255875 16916 255876
rect 16884 255845 16885 255875
rect 16885 255845 16915 255875
rect 16915 255845 16916 255875
rect 16884 255844 16916 255845
rect 16724 255715 16756 255716
rect 16724 255685 16725 255715
rect 16725 255685 16755 255715
rect 16755 255685 16756 255715
rect 16724 255684 16756 255685
rect 16884 255715 16916 255716
rect 16884 255685 16885 255715
rect 16885 255685 16915 255715
rect 16915 255685 16916 255715
rect 16884 255684 16916 255685
<< metal4 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
rect 271860 351816 283220 351820
rect 271860 351784 271864 351816
rect 271896 351784 272024 351816
rect 272056 351784 272104 351816
rect 272136 351784 272184 351816
rect 272216 351784 272264 351816
rect 272296 351784 272344 351816
rect 272376 351784 272424 351816
rect 272456 351784 272504 351816
rect 272536 351784 272584 351816
rect 272616 351784 272664 351816
rect 272696 351784 272744 351816
rect 272776 351784 272824 351816
rect 272856 351784 272904 351816
rect 272936 351784 272984 351816
rect 273016 351784 273064 351816
rect 273096 351784 273144 351816
rect 273176 351784 273224 351816
rect 273256 351784 273304 351816
rect 273336 351784 273384 351816
rect 273416 351784 273464 351816
rect 273496 351784 273544 351816
rect 273576 351784 273624 351816
rect 273656 351784 273704 351816
rect 273736 351784 273784 351816
rect 273816 351784 273864 351816
rect 273896 351784 273944 351816
rect 273976 351784 274024 351816
rect 274056 351784 274104 351816
rect 274136 351784 274184 351816
rect 274216 351784 274264 351816
rect 274296 351784 274344 351816
rect 274376 351784 274424 351816
rect 274456 351784 274504 351816
rect 274536 351784 274584 351816
rect 274616 351784 274664 351816
rect 274696 351784 274744 351816
rect 274776 351784 274824 351816
rect 274856 351784 274904 351816
rect 274936 351784 274984 351816
rect 275016 351784 275064 351816
rect 275096 351784 275144 351816
rect 275176 351784 275224 351816
rect 275256 351784 275304 351816
rect 275336 351784 275384 351816
rect 275416 351784 275464 351816
rect 275496 351784 275544 351816
rect 275576 351784 275624 351816
rect 275656 351784 275704 351816
rect 275736 351784 275784 351816
rect 275816 351784 275864 351816
rect 275896 351784 275944 351816
rect 275976 351784 276024 351816
rect 276056 351784 276104 351816
rect 276136 351784 276184 351816
rect 276216 351784 276264 351816
rect 276296 351784 276344 351816
rect 276376 351784 276424 351816
rect 276456 351784 276504 351816
rect 276536 351784 276584 351816
rect 276616 351784 276664 351816
rect 276696 351784 276744 351816
rect 276776 351784 276824 351816
rect 276856 351784 276904 351816
rect 276936 351784 276984 351816
rect 277016 351784 277064 351816
rect 277096 351784 277144 351816
rect 277176 351784 277224 351816
rect 277256 351784 277304 351816
rect 277336 351784 277384 351816
rect 277416 351784 277464 351816
rect 277496 351784 277544 351816
rect 277576 351784 277624 351816
rect 277656 351784 277704 351816
rect 277736 351784 277784 351816
rect 277816 351784 277864 351816
rect 277896 351784 277944 351816
rect 277976 351784 278024 351816
rect 278056 351784 278104 351816
rect 278136 351784 278184 351816
rect 278216 351784 278264 351816
rect 278296 351784 278344 351816
rect 278376 351784 278424 351816
rect 278456 351784 278504 351816
rect 278536 351784 278584 351816
rect 278616 351784 278664 351816
rect 278696 351784 278744 351816
rect 278776 351784 278824 351816
rect 278856 351784 278904 351816
rect 278936 351784 278984 351816
rect 279016 351784 279064 351816
rect 279096 351784 279144 351816
rect 279176 351784 279224 351816
rect 279256 351784 279304 351816
rect 279336 351784 279384 351816
rect 279416 351784 279464 351816
rect 279496 351784 279544 351816
rect 279576 351784 279624 351816
rect 279656 351784 279704 351816
rect 279736 351784 279784 351816
rect 279816 351784 279864 351816
rect 279896 351784 279944 351816
rect 279976 351784 280024 351816
rect 280056 351784 280104 351816
rect 280136 351784 280184 351816
rect 280216 351784 280264 351816
rect 280296 351784 280344 351816
rect 280376 351784 280424 351816
rect 280456 351784 280504 351816
rect 280536 351784 280584 351816
rect 280616 351784 280664 351816
rect 280696 351784 280744 351816
rect 280776 351784 280824 351816
rect 280856 351784 280904 351816
rect 280936 351784 280984 351816
rect 281016 351784 281064 351816
rect 281096 351784 281144 351816
rect 281176 351784 281224 351816
rect 281256 351784 281304 351816
rect 281336 351784 281384 351816
rect 281416 351784 281464 351816
rect 281496 351784 281544 351816
rect 281576 351784 281624 351816
rect 281656 351784 281704 351816
rect 281736 351784 281784 351816
rect 281816 351784 281864 351816
rect 281896 351784 281944 351816
rect 281976 351784 282024 351816
rect 282056 351784 282104 351816
rect 282136 351784 282184 351816
rect 282216 351784 282264 351816
rect 282296 351784 282344 351816
rect 282376 351784 282424 351816
rect 282456 351784 282504 351816
rect 282536 351784 282584 351816
rect 282616 351784 282664 351816
rect 282696 351784 282744 351816
rect 282776 351784 282824 351816
rect 282856 351784 282904 351816
rect 282936 351784 282984 351816
rect 283016 351784 283064 351816
rect 283096 351784 283144 351816
rect 283176 351784 283220 351816
rect 271860 351780 283220 351784
rect 271940 351736 283220 351740
rect 271940 351704 272024 351736
rect 272056 351704 272104 351736
rect 272136 351704 272184 351736
rect 272216 351704 272264 351736
rect 272296 351704 272344 351736
rect 272376 351704 272424 351736
rect 272456 351704 272504 351736
rect 272536 351704 272584 351736
rect 272616 351704 272664 351736
rect 272696 351704 272744 351736
rect 272776 351704 272824 351736
rect 272856 351704 272904 351736
rect 272936 351704 272984 351736
rect 273016 351704 273064 351736
rect 273096 351704 273144 351736
rect 273176 351704 273224 351736
rect 273256 351704 273304 351736
rect 273336 351704 273384 351736
rect 273416 351704 273464 351736
rect 273496 351704 273544 351736
rect 273576 351704 273624 351736
rect 273656 351704 273704 351736
rect 273736 351704 273784 351736
rect 273816 351704 273864 351736
rect 273896 351704 273944 351736
rect 273976 351704 274024 351736
rect 274056 351704 274104 351736
rect 274136 351704 274184 351736
rect 274216 351704 274264 351736
rect 274296 351704 274344 351736
rect 274376 351704 274424 351736
rect 274456 351704 274504 351736
rect 274536 351704 274584 351736
rect 274616 351704 274664 351736
rect 274696 351704 274744 351736
rect 274776 351704 274824 351736
rect 274856 351704 274904 351736
rect 274936 351704 274984 351736
rect 275016 351704 275064 351736
rect 275096 351704 275144 351736
rect 275176 351704 275224 351736
rect 275256 351704 275304 351736
rect 275336 351704 275384 351736
rect 275416 351704 275464 351736
rect 275496 351704 275544 351736
rect 275576 351704 275624 351736
rect 275656 351704 275704 351736
rect 275736 351704 275784 351736
rect 275816 351704 275864 351736
rect 275896 351704 275944 351736
rect 275976 351704 276024 351736
rect 276056 351704 276104 351736
rect 276136 351704 276184 351736
rect 276216 351704 276264 351736
rect 276296 351704 276344 351736
rect 276376 351704 276424 351736
rect 276456 351704 276504 351736
rect 276536 351704 276584 351736
rect 276616 351704 276664 351736
rect 276696 351704 276744 351736
rect 276776 351704 276824 351736
rect 276856 351704 276904 351736
rect 276936 351704 276984 351736
rect 277016 351704 277064 351736
rect 277096 351704 277144 351736
rect 277176 351704 277224 351736
rect 277256 351704 277304 351736
rect 277336 351704 277384 351736
rect 277416 351704 277464 351736
rect 277496 351704 277544 351736
rect 277576 351704 277624 351736
rect 277656 351704 277704 351736
rect 277736 351704 277784 351736
rect 277816 351704 277864 351736
rect 277896 351704 277944 351736
rect 277976 351704 278024 351736
rect 278056 351704 278104 351736
rect 278136 351704 278184 351736
rect 278216 351704 278264 351736
rect 278296 351704 278344 351736
rect 278376 351704 278424 351736
rect 278456 351704 278504 351736
rect 278536 351704 278584 351736
rect 278616 351704 278664 351736
rect 278696 351704 278744 351736
rect 278776 351704 278824 351736
rect 278856 351704 278904 351736
rect 278936 351704 278984 351736
rect 279016 351704 279064 351736
rect 279096 351704 279144 351736
rect 279176 351704 279224 351736
rect 279256 351704 279304 351736
rect 279336 351704 279384 351736
rect 279416 351704 279464 351736
rect 279496 351704 279544 351736
rect 279576 351704 279624 351736
rect 279656 351704 279704 351736
rect 279736 351704 279784 351736
rect 279816 351704 279864 351736
rect 279896 351704 279944 351736
rect 279976 351704 280024 351736
rect 280056 351704 280104 351736
rect 280136 351704 280184 351736
rect 280216 351704 280264 351736
rect 280296 351704 280344 351736
rect 280376 351704 280424 351736
rect 280456 351704 280504 351736
rect 280536 351704 280584 351736
rect 280616 351704 280664 351736
rect 280696 351704 280744 351736
rect 280776 351704 280824 351736
rect 280856 351704 280904 351736
rect 280936 351704 280984 351736
rect 281016 351704 281064 351736
rect 281096 351704 281144 351736
rect 281176 351704 281224 351736
rect 281256 351704 281304 351736
rect 281336 351704 281384 351736
rect 281416 351704 281464 351736
rect 281496 351704 281544 351736
rect 281576 351704 281624 351736
rect 281656 351704 281704 351736
rect 281736 351704 281784 351736
rect 281816 351704 281864 351736
rect 281896 351704 281944 351736
rect 281976 351704 282024 351736
rect 282056 351704 282104 351736
rect 282136 351704 282184 351736
rect 282216 351704 282264 351736
rect 282296 351704 282344 351736
rect 282376 351704 282424 351736
rect 282456 351704 282504 351736
rect 282536 351704 282584 351736
rect 282616 351704 282664 351736
rect 282696 351704 282744 351736
rect 282776 351704 282824 351736
rect 282856 351704 282904 351736
rect 282936 351704 282984 351736
rect 283016 351704 283064 351736
rect 283096 351704 283144 351736
rect 283176 351704 283220 351736
rect 271940 351700 283220 351704
rect 271860 351656 283220 351660
rect 271860 351624 271864 351656
rect 271896 351624 272024 351656
rect 272056 351624 272104 351656
rect 272136 351624 272184 351656
rect 272216 351624 272264 351656
rect 272296 351624 272344 351656
rect 272376 351624 272424 351656
rect 272456 351624 272504 351656
rect 272536 351624 272584 351656
rect 272616 351624 272664 351656
rect 272696 351624 272744 351656
rect 272776 351624 272824 351656
rect 272856 351624 272904 351656
rect 272936 351624 272984 351656
rect 273016 351624 273064 351656
rect 273096 351624 273144 351656
rect 273176 351624 273224 351656
rect 273256 351624 273304 351656
rect 273336 351624 273384 351656
rect 273416 351624 273464 351656
rect 273496 351624 273544 351656
rect 273576 351624 273624 351656
rect 273656 351624 273704 351656
rect 273736 351624 273784 351656
rect 273816 351624 273864 351656
rect 273896 351624 273944 351656
rect 273976 351624 274024 351656
rect 274056 351624 274104 351656
rect 274136 351624 274184 351656
rect 274216 351624 274264 351656
rect 274296 351624 274344 351656
rect 274376 351624 274424 351656
rect 274456 351624 274504 351656
rect 274536 351624 274584 351656
rect 274616 351624 274664 351656
rect 274696 351624 274744 351656
rect 274776 351624 274824 351656
rect 274856 351624 274904 351656
rect 274936 351624 274984 351656
rect 275016 351624 275064 351656
rect 275096 351624 275144 351656
rect 275176 351624 275224 351656
rect 275256 351624 275304 351656
rect 275336 351624 275384 351656
rect 275416 351624 275464 351656
rect 275496 351624 275544 351656
rect 275576 351624 275624 351656
rect 275656 351624 275704 351656
rect 275736 351624 275784 351656
rect 275816 351624 275864 351656
rect 275896 351624 275944 351656
rect 275976 351624 276024 351656
rect 276056 351624 276104 351656
rect 276136 351624 276184 351656
rect 276216 351624 276264 351656
rect 276296 351624 276344 351656
rect 276376 351624 276424 351656
rect 276456 351624 276504 351656
rect 276536 351624 276584 351656
rect 276616 351624 276664 351656
rect 276696 351624 276744 351656
rect 276776 351624 276824 351656
rect 276856 351624 276904 351656
rect 276936 351624 276984 351656
rect 277016 351624 277064 351656
rect 277096 351624 277144 351656
rect 277176 351624 277224 351656
rect 277256 351624 277304 351656
rect 277336 351624 277384 351656
rect 277416 351624 277464 351656
rect 277496 351624 277544 351656
rect 277576 351624 277624 351656
rect 277656 351624 277704 351656
rect 277736 351624 277784 351656
rect 277816 351624 277864 351656
rect 277896 351624 277944 351656
rect 277976 351624 278024 351656
rect 278056 351624 278104 351656
rect 278136 351624 278184 351656
rect 278216 351624 278264 351656
rect 278296 351624 278344 351656
rect 278376 351624 278424 351656
rect 278456 351624 278504 351656
rect 278536 351624 278584 351656
rect 278616 351624 278664 351656
rect 278696 351624 278744 351656
rect 278776 351624 278824 351656
rect 278856 351624 278904 351656
rect 278936 351624 278984 351656
rect 279016 351624 279064 351656
rect 279096 351624 279144 351656
rect 279176 351624 279224 351656
rect 279256 351624 279304 351656
rect 279336 351624 279384 351656
rect 279416 351624 279464 351656
rect 279496 351624 279544 351656
rect 279576 351624 279624 351656
rect 279656 351624 279704 351656
rect 279736 351624 279784 351656
rect 279816 351624 279864 351656
rect 279896 351624 279944 351656
rect 279976 351624 280024 351656
rect 280056 351624 280104 351656
rect 280136 351624 280184 351656
rect 280216 351624 280264 351656
rect 280296 351624 280344 351656
rect 280376 351624 280424 351656
rect 280456 351624 280504 351656
rect 280536 351624 280584 351656
rect 280616 351624 280664 351656
rect 280696 351624 280744 351656
rect 280776 351624 280824 351656
rect 280856 351624 280904 351656
rect 280936 351624 280984 351656
rect 281016 351624 281064 351656
rect 281096 351624 281144 351656
rect 281176 351624 281224 351656
rect 281256 351624 281304 351656
rect 281336 351624 281384 351656
rect 281416 351624 281464 351656
rect 281496 351624 281544 351656
rect 281576 351624 281624 351656
rect 281656 351624 281704 351656
rect 281736 351624 281784 351656
rect 281816 351624 281864 351656
rect 281896 351624 281944 351656
rect 281976 351624 282024 351656
rect 282056 351624 282104 351656
rect 282136 351624 282184 351656
rect 282216 351624 282264 351656
rect 282296 351624 282344 351656
rect 282376 351624 282424 351656
rect 282456 351624 282504 351656
rect 282536 351624 282584 351656
rect 282616 351624 282664 351656
rect 282696 351624 282744 351656
rect 282776 351624 282824 351656
rect 282856 351624 282904 351656
rect 282936 351624 282984 351656
rect 283016 351624 283064 351656
rect 283096 351624 283144 351656
rect 283176 351624 283220 351656
rect 271860 351620 283220 351624
rect 271860 351576 272060 351580
rect 271860 351544 271864 351576
rect 271896 351544 272024 351576
rect 272056 351544 272060 351576
rect 271860 351540 272060 351544
rect 271860 351496 272060 351500
rect 271860 351464 271864 351496
rect 271896 351464 272024 351496
rect 272056 351464 272060 351496
rect 271860 351460 272060 351464
rect 271860 351416 272060 351420
rect 271860 351384 271864 351416
rect 271896 351384 272024 351416
rect 272056 351384 272060 351416
rect 271860 351380 272060 351384
rect 271860 351336 272060 351340
rect 271860 351304 271864 351336
rect 271896 351304 272024 351336
rect 272056 351304 272060 351336
rect 271860 351300 272060 351304
rect 271860 351256 272060 351260
rect 271860 351224 271864 351256
rect 271896 351224 272024 351256
rect 272056 351224 272060 351256
rect 271860 351220 272060 351224
rect 271860 351176 272060 351180
rect 271860 351144 271864 351176
rect 271896 351144 272024 351176
rect 272056 351144 272060 351176
rect 271860 351140 272060 351144
rect 271860 351096 272060 351100
rect 271860 351064 271864 351096
rect 271896 351064 272024 351096
rect 272056 351064 272060 351096
rect 271860 351060 272060 351064
rect 271860 351016 272060 351020
rect 271860 350984 271864 351016
rect 271896 350984 272024 351016
rect 272056 350984 272060 351016
rect 271860 350980 272060 350984
rect 271860 350936 272060 350940
rect 271860 350904 271864 350936
rect 271896 350904 272024 350936
rect 272056 350904 272060 350936
rect 271860 350900 272060 350904
rect 271860 350856 272060 350860
rect 271860 350824 271864 350856
rect 271896 350824 272024 350856
rect 272056 350824 272060 350856
rect 271860 350820 272060 350824
rect 271860 350776 272060 350780
rect 271860 350744 271864 350776
rect 271896 350744 272024 350776
rect 272056 350744 272060 350776
rect 271860 350740 272060 350744
rect 271860 350696 272060 350700
rect 271860 350664 271864 350696
rect 271896 350664 272024 350696
rect 272056 350664 272060 350696
rect 271860 350660 272060 350664
rect 271860 350616 272060 350620
rect 271860 350584 271864 350616
rect 271896 350584 272024 350616
rect 272056 350584 272060 350616
rect 271860 350580 272060 350584
rect 271860 350536 272060 350540
rect 271860 350504 271864 350536
rect 271896 350504 272024 350536
rect 272056 350504 272060 350536
rect 271860 350500 272060 350504
rect 271860 350456 272060 350460
rect 271860 350424 271864 350456
rect 271896 350424 272024 350456
rect 272056 350424 272060 350456
rect 271860 350420 272060 350424
rect 271860 350376 272060 350380
rect 271860 350344 271864 350376
rect 271896 350344 272024 350376
rect 272056 350344 272060 350376
rect 271860 350340 272060 350344
rect 271860 350296 272060 350300
rect 271860 350264 271864 350296
rect 271896 350264 272024 350296
rect 272056 350264 272060 350296
rect 271860 350260 272060 350264
rect 271860 350216 272060 350220
rect 271860 350184 271864 350216
rect 271896 350184 272024 350216
rect 272056 350184 272060 350216
rect 271860 350180 272060 350184
rect 271860 350136 272060 350140
rect 271860 350104 271864 350136
rect 271896 350104 272024 350136
rect 272056 350104 272060 350136
rect 271860 350100 272060 350104
rect 271860 350056 272060 350060
rect 271860 350024 271864 350056
rect 271896 350024 272024 350056
rect 272056 350024 272060 350056
rect 271860 350020 272060 350024
rect 1000 317790 16400 317800
rect 1000 317610 1010 317790
rect 1190 317610 16210 317790
rect 16390 317610 16400 317790
rect 1000 317600 16400 317610
rect 16720 275476 17240 275480
rect 16720 275444 16724 275476
rect 16756 275444 16884 275476
rect 16916 275444 16964 275476
rect 16996 275444 17044 275476
rect 17076 275444 17124 275476
rect 17156 275444 17204 275476
rect 17236 275444 17240 275476
rect 16720 275440 17240 275444
rect 16720 275396 17240 275400
rect 16720 275364 16884 275396
rect 16916 275364 16964 275396
rect 16996 275364 17044 275396
rect 17076 275364 17240 275396
rect 16720 275360 17240 275364
rect 28400 275356 28760 275360
rect 28400 275324 28404 275356
rect 28436 275324 28564 275356
rect 28596 275324 28724 275356
rect 28756 275324 28760 275356
rect 28400 275320 28760 275324
rect 16720 275316 17240 275320
rect 16720 275284 16724 275316
rect 16756 275284 16884 275316
rect 16916 275284 16964 275316
rect 16996 275284 17044 275316
rect 17076 275284 17204 275316
rect 17236 275284 17240 275316
rect 16720 275280 17240 275284
rect 28400 275276 28760 275280
rect 28400 275244 28404 275276
rect 28436 275244 28564 275276
rect 28596 275244 28724 275276
rect 28756 275244 28760 275276
rect 28400 275240 28760 275244
rect 1000 275190 259100 275200
rect 1000 275160 258910 275190
rect 1000 275040 1040 275160
rect 1160 275040 258910 275160
rect 1000 275010 258910 275040
rect 259090 275010 259100 275190
rect 1000 275000 259100 275010
rect 16720 274956 16920 274960
rect 16720 274924 16724 274956
rect 16756 274924 16884 274956
rect 16916 274924 16920 274956
rect 16720 274920 16920 274924
rect 16720 274876 16920 274880
rect 16720 274844 16724 274876
rect 16756 274844 16884 274876
rect 16916 274844 16920 274876
rect 16720 274840 16920 274844
rect 17000 274840 17200 274880
rect 17000 274800 17100 274840
rect 16200 274790 17200 274800
rect 16200 274610 16210 274790
rect 16390 274760 17200 274790
rect 16390 274720 17100 274760
rect 16390 274680 17200 274720
rect 16390 274640 17100 274680
rect 16390 274610 17200 274640
rect 16200 274600 17200 274610
rect 17000 274560 17100 274600
rect 16720 274556 16920 274560
rect 16720 274524 16724 274556
rect 16756 274524 16884 274556
rect 16916 274524 16920 274556
rect 16720 274520 16920 274524
rect 17000 274520 17200 274560
rect 16720 274476 16920 274480
rect 16720 274444 16724 274476
rect 16756 274444 16884 274476
rect 16916 274444 16920 274476
rect 16720 274440 16920 274444
rect 16720 274396 16920 274400
rect 16720 274364 16724 274396
rect 16756 274364 16884 274396
rect 16916 274364 16920 274396
rect 16720 274360 16920 274364
rect 16720 274316 16920 274320
rect 16720 274284 16724 274316
rect 16756 274284 16884 274316
rect 16916 274284 16920 274316
rect 16720 274280 16920 274284
rect 16720 274236 16920 274240
rect 16720 274204 16724 274236
rect 16756 274204 16884 274236
rect 16916 274204 16920 274236
rect 16720 274200 16920 274204
rect 16720 274156 16920 274160
rect 16720 274124 16724 274156
rect 16756 274124 16884 274156
rect 16916 274124 16920 274156
rect 16720 274120 16920 274124
rect 16720 274076 16920 274080
rect 16720 274044 16724 274076
rect 16756 274044 16884 274076
rect 16916 274044 16920 274076
rect 16720 274040 16920 274044
rect 16720 273996 16920 274000
rect 16720 273964 16724 273996
rect 16756 273964 16884 273996
rect 16916 273964 16920 273996
rect 16720 273960 16920 273964
rect 16720 273916 16920 273920
rect 16720 273884 16724 273916
rect 16756 273884 16884 273916
rect 16916 273884 16920 273916
rect 16720 273880 16920 273884
rect 16720 273836 16920 273840
rect 16720 273804 16724 273836
rect 16756 273804 16884 273836
rect 16916 273804 16920 273836
rect 16720 273800 16920 273804
rect 16720 273756 16920 273760
rect 16720 273724 16724 273756
rect 16756 273724 16884 273756
rect 16916 273724 16920 273756
rect 16720 273720 16920 273724
rect 16720 273676 16920 273680
rect 16720 273644 16724 273676
rect 16756 273644 16884 273676
rect 16916 273644 16920 273676
rect 16720 273640 16920 273644
rect 16720 273596 16920 273600
rect 16720 273564 16724 273596
rect 16756 273564 16884 273596
rect 16916 273564 16920 273596
rect 16720 273560 16920 273564
rect 16720 273516 16920 273520
rect 16720 273484 16724 273516
rect 16756 273484 16884 273516
rect 16916 273484 16920 273516
rect 16720 273480 16920 273484
rect 16720 273436 16920 273440
rect 16720 273404 16724 273436
rect 16756 273404 16884 273436
rect 16916 273404 16920 273436
rect 16720 273400 16920 273404
rect 16720 273356 16920 273360
rect 16720 273324 16724 273356
rect 16756 273324 16884 273356
rect 16916 273324 16920 273356
rect 16720 273320 16920 273324
rect 16720 273276 16920 273280
rect 16720 273244 16724 273276
rect 16756 273244 16884 273276
rect 16916 273244 16920 273276
rect 16720 273240 16920 273244
rect 16720 273196 16920 273200
rect 16720 273164 16724 273196
rect 16756 273164 16884 273196
rect 16916 273164 16920 273196
rect 16720 273160 16920 273164
rect 16720 273116 16920 273120
rect 16720 273084 16724 273116
rect 16756 273084 16884 273116
rect 16916 273084 16920 273116
rect 16720 273080 16920 273084
rect 16720 273036 16920 273040
rect 16720 273004 16724 273036
rect 16756 273004 16884 273036
rect 16916 273004 16920 273036
rect 16720 273000 16920 273004
rect 16720 272956 16920 272960
rect 16720 272924 16724 272956
rect 16756 272924 16884 272956
rect 16916 272924 16920 272956
rect 16720 272920 16920 272924
rect 16720 272876 16920 272880
rect 16720 272844 16724 272876
rect 16756 272844 16884 272876
rect 16916 272844 16920 272876
rect 16720 272840 16920 272844
rect 16720 272796 16920 272800
rect 16720 272764 16724 272796
rect 16756 272764 16884 272796
rect 16916 272764 16920 272796
rect 16720 272760 16920 272764
rect 16720 272716 16920 272720
rect 16720 272684 16724 272716
rect 16756 272684 16884 272716
rect 16916 272684 16920 272716
rect 16720 272680 16920 272684
rect 16720 272636 16920 272640
rect 16720 272604 16724 272636
rect 16756 272604 16884 272636
rect 16916 272604 16920 272636
rect 16720 272600 16920 272604
rect 16720 272556 16920 272560
rect 16720 272524 16724 272556
rect 16756 272524 16884 272556
rect 16916 272524 16920 272556
rect 16720 272520 16920 272524
rect 16720 272476 16920 272480
rect 16720 272444 16724 272476
rect 16756 272444 16884 272476
rect 16916 272444 16920 272476
rect 16720 272440 16920 272444
rect 16720 272396 16920 272400
rect 16720 272364 16724 272396
rect 16756 272364 16884 272396
rect 16916 272364 16920 272396
rect 16720 272360 16920 272364
rect 16720 272316 16920 272320
rect 16720 272284 16724 272316
rect 16756 272284 16884 272316
rect 16916 272284 16920 272316
rect 16720 272280 16920 272284
rect 16720 272236 16920 272240
rect 16720 272204 16724 272236
rect 16756 272204 16884 272236
rect 16916 272204 16920 272236
rect 16720 272200 16920 272204
rect 16720 272156 16920 272160
rect 16720 272124 16724 272156
rect 16756 272124 16884 272156
rect 16916 272124 16920 272156
rect 16720 272120 16920 272124
rect 16720 272076 16920 272080
rect 16720 272044 16724 272076
rect 16756 272044 16884 272076
rect 16916 272044 16920 272076
rect 16720 272040 16920 272044
rect 16720 271996 16920 272000
rect 16720 271964 16724 271996
rect 16756 271964 16884 271996
rect 16916 271964 16920 271996
rect 16720 271960 16920 271964
rect 16720 271916 16920 271920
rect 16720 271884 16724 271916
rect 16756 271884 16884 271916
rect 16916 271884 16920 271916
rect 16720 271880 16920 271884
rect 16720 271836 16920 271840
rect 16720 271804 16724 271836
rect 16756 271804 16884 271836
rect 16916 271804 16920 271836
rect 16720 271800 16920 271804
rect 16720 271756 16920 271760
rect 16720 271724 16724 271756
rect 16756 271724 16884 271756
rect 16916 271724 16920 271756
rect 16720 271720 16920 271724
rect 16720 271676 16920 271680
rect 16720 271644 16724 271676
rect 16756 271644 16884 271676
rect 16916 271644 16920 271676
rect 16720 271640 16920 271644
rect 16720 271596 16920 271600
rect 16720 271564 16724 271596
rect 16756 271564 16884 271596
rect 16916 271564 16920 271596
rect 16720 271560 16920 271564
rect 16720 271516 16920 271520
rect 16720 271484 16724 271516
rect 16756 271484 16884 271516
rect 16916 271484 16920 271516
rect 16720 271480 16920 271484
rect 16720 271436 16920 271440
rect 16720 271404 16724 271436
rect 16756 271404 16884 271436
rect 16916 271404 16920 271436
rect 16720 271400 16920 271404
rect 16720 271356 16920 271360
rect 16720 271324 16724 271356
rect 16756 271324 16884 271356
rect 16916 271324 16920 271356
rect 16720 271320 16920 271324
rect 16720 271276 16920 271280
rect 16720 271244 16724 271276
rect 16756 271244 16884 271276
rect 16916 271244 16920 271276
rect 16720 271240 16920 271244
rect 16720 271196 16920 271200
rect 16720 271164 16724 271196
rect 16756 271164 16884 271196
rect 16916 271164 16920 271196
rect 16720 271160 16920 271164
rect 16720 271116 16920 271120
rect 16720 271084 16724 271116
rect 16756 271084 16884 271116
rect 16916 271084 16920 271116
rect 16720 271080 16920 271084
rect 16720 271036 16920 271040
rect 16720 271004 16724 271036
rect 16756 271004 16884 271036
rect 16916 271004 16920 271036
rect 16720 271000 16920 271004
rect 16720 270956 16920 270960
rect 16720 270924 16724 270956
rect 16756 270924 16884 270956
rect 16916 270924 16920 270956
rect 16720 270920 16920 270924
rect 16720 270876 16920 270880
rect 16720 270844 16724 270876
rect 16756 270844 16884 270876
rect 16916 270844 16920 270876
rect 16720 270840 16920 270844
rect 16720 270796 16920 270800
rect 16720 270764 16724 270796
rect 16756 270764 16884 270796
rect 16916 270764 16920 270796
rect 16720 270760 16920 270764
rect 16720 270716 16920 270720
rect 16720 270684 16724 270716
rect 16756 270684 16884 270716
rect 16916 270684 16920 270716
rect 16720 270680 16920 270684
rect 16720 270636 16920 270640
rect 16720 270604 16724 270636
rect 16756 270604 16884 270636
rect 16916 270604 16920 270636
rect 16720 270600 16920 270604
rect 16720 270556 16920 270560
rect 16720 270524 16724 270556
rect 16756 270524 16884 270556
rect 16916 270524 16920 270556
rect 16720 270520 16920 270524
rect 16720 270476 16920 270480
rect 16720 270444 16724 270476
rect 16756 270444 16884 270476
rect 16916 270444 16920 270476
rect 16720 270440 16920 270444
rect 16720 270396 16920 270400
rect 16720 270364 16724 270396
rect 16756 270364 16884 270396
rect 16916 270364 16920 270396
rect 16720 270360 16920 270364
rect 16720 270316 16920 270320
rect 16720 270284 16724 270316
rect 16756 270284 16884 270316
rect 16916 270284 16920 270316
rect 16720 270280 16920 270284
rect 16720 270236 16920 270240
rect 16720 270204 16724 270236
rect 16756 270204 16884 270236
rect 16916 270204 16920 270236
rect 16720 270200 16920 270204
rect 16720 270156 16920 270160
rect 16720 270124 16724 270156
rect 16756 270124 16884 270156
rect 16916 270124 16920 270156
rect 16720 270120 16920 270124
rect 16720 270076 16920 270080
rect 16720 270044 16724 270076
rect 16756 270044 16884 270076
rect 16916 270044 16920 270076
rect 16720 270040 16920 270044
rect 16720 269996 16920 270000
rect 16720 269964 16724 269996
rect 16756 269964 16884 269996
rect 16916 269964 16920 269996
rect 16720 269960 16920 269964
rect 16720 269916 16920 269920
rect 16720 269884 16724 269916
rect 16756 269884 16884 269916
rect 16916 269884 16920 269916
rect 16720 269880 16920 269884
rect 16720 269836 16920 269840
rect 16720 269804 16724 269836
rect 16756 269804 16884 269836
rect 16916 269804 16920 269836
rect 16720 269800 16920 269804
rect 16720 269756 16920 269760
rect 16720 269724 16724 269756
rect 16756 269724 16884 269756
rect 16916 269724 16920 269756
rect 16720 269720 16920 269724
rect 16720 269676 16920 269680
rect 16720 269644 16724 269676
rect 16756 269644 16884 269676
rect 16916 269644 16920 269676
rect 16720 269640 16920 269644
rect 16720 269596 16920 269600
rect 16720 269564 16724 269596
rect 16756 269564 16884 269596
rect 16916 269564 16920 269596
rect 16720 269560 16920 269564
rect 16720 269516 16920 269520
rect 16720 269484 16724 269516
rect 16756 269484 16884 269516
rect 16916 269484 16920 269516
rect 16720 269480 16920 269484
rect 16720 269436 16920 269440
rect 16720 269404 16724 269436
rect 16756 269404 16884 269436
rect 16916 269404 16920 269436
rect 16720 269400 16920 269404
rect 16720 269356 16920 269360
rect 16720 269324 16724 269356
rect 16756 269324 16884 269356
rect 16916 269324 16920 269356
rect 16720 269320 16920 269324
rect 16720 269276 16920 269280
rect 16720 269244 16724 269276
rect 16756 269244 16884 269276
rect 16916 269244 16920 269276
rect 16720 269240 16920 269244
rect 16720 269196 16920 269200
rect 16720 269164 16724 269196
rect 16756 269164 16884 269196
rect 16916 269164 16920 269196
rect 16720 269160 16920 269164
rect 16720 269116 16920 269120
rect 16720 269084 16724 269116
rect 16756 269084 16884 269116
rect 16916 269084 16920 269116
rect 16720 269080 16920 269084
rect 16720 269036 16920 269040
rect 16720 269004 16724 269036
rect 16756 269004 16884 269036
rect 16916 269004 16920 269036
rect 16720 269000 16920 269004
rect 16720 268956 16920 268960
rect 16720 268924 16724 268956
rect 16756 268924 16884 268956
rect 16916 268924 16920 268956
rect 16720 268920 16920 268924
rect 16720 268876 16920 268880
rect 16720 268844 16724 268876
rect 16756 268844 16884 268876
rect 16916 268844 16920 268876
rect 16720 268840 16920 268844
rect 16720 268796 16920 268800
rect 16720 268764 16724 268796
rect 16756 268764 16884 268796
rect 16916 268764 16920 268796
rect 16720 268760 16920 268764
rect 16720 268716 16920 268720
rect 16720 268684 16724 268716
rect 16756 268684 16884 268716
rect 16916 268684 16920 268716
rect 16720 268680 16920 268684
rect 16720 268636 16920 268640
rect 16720 268604 16724 268636
rect 16756 268604 16884 268636
rect 16916 268604 16920 268636
rect 16720 268600 16920 268604
rect 16720 268556 16920 268560
rect 16720 268524 16724 268556
rect 16756 268524 16884 268556
rect 16916 268524 16920 268556
rect 16720 268520 16920 268524
rect 16720 268476 16920 268480
rect 16720 268444 16724 268476
rect 16756 268444 16884 268476
rect 16916 268444 16920 268476
rect 16720 268440 16920 268444
rect 16720 268396 16920 268400
rect 16720 268364 16724 268396
rect 16756 268364 16884 268396
rect 16916 268364 16920 268396
rect 16720 268360 16920 268364
rect 16720 268316 16920 268320
rect 16720 268284 16724 268316
rect 16756 268284 16884 268316
rect 16916 268284 16920 268316
rect 16720 268280 16920 268284
rect 16720 268236 16920 268240
rect 16720 268204 16724 268236
rect 16756 268204 16884 268236
rect 16916 268204 16920 268236
rect 16720 268200 16920 268204
rect 16720 268156 16920 268160
rect 16720 268124 16724 268156
rect 16756 268124 16884 268156
rect 16916 268124 16920 268156
rect 16720 268120 16920 268124
rect 16720 268076 16920 268080
rect 16720 268044 16724 268076
rect 16756 268044 16884 268076
rect 16916 268044 16920 268076
rect 16720 268040 16920 268044
rect 16720 267996 16920 268000
rect 16720 267964 16724 267996
rect 16756 267964 16884 267996
rect 16916 267964 16920 267996
rect 16720 267960 16920 267964
rect 16720 267916 16920 267920
rect 16720 267884 16724 267916
rect 16756 267884 16884 267916
rect 16916 267884 16920 267916
rect 16720 267880 16920 267884
rect 16720 267836 16920 267840
rect 16720 267804 16724 267836
rect 16756 267804 16884 267836
rect 16916 267804 16920 267836
rect 16720 267800 16920 267804
rect 16720 267756 16920 267760
rect 16720 267724 16724 267756
rect 16756 267724 16884 267756
rect 16916 267724 16920 267756
rect 16720 267720 16920 267724
rect 16720 267676 16920 267680
rect 16720 267644 16724 267676
rect 16756 267644 16884 267676
rect 16916 267644 16920 267676
rect 16720 267640 16920 267644
rect 16720 267596 16920 267600
rect 16720 267564 16724 267596
rect 16756 267564 16884 267596
rect 16916 267564 16920 267596
rect 16720 267560 16920 267564
rect 16720 267516 16920 267520
rect 16720 267484 16724 267516
rect 16756 267484 16884 267516
rect 16916 267484 16920 267516
rect 16720 267480 16920 267484
rect 16720 267436 16920 267440
rect 16720 267404 16724 267436
rect 16756 267404 16884 267436
rect 16916 267404 16920 267436
rect 16720 267400 16920 267404
rect 16720 267356 16920 267360
rect 16720 267324 16724 267356
rect 16756 267324 16884 267356
rect 16916 267324 16920 267356
rect 16720 267320 16920 267324
rect 16720 267276 16920 267280
rect 16720 267244 16724 267276
rect 16756 267244 16884 267276
rect 16916 267244 16920 267276
rect 16720 267240 16920 267244
rect 16720 267196 16920 267200
rect 16720 267164 16724 267196
rect 16756 267164 16884 267196
rect 16916 267164 16920 267196
rect 16720 267160 16920 267164
rect 16720 267116 16920 267120
rect 16720 267084 16724 267116
rect 16756 267084 16884 267116
rect 16916 267084 16920 267116
rect 16720 267080 16920 267084
rect 16720 267036 16920 267040
rect 16720 267004 16724 267036
rect 16756 267004 16884 267036
rect 16916 267004 16920 267036
rect 16720 267000 16920 267004
rect 16720 266956 16920 266960
rect 16720 266924 16724 266956
rect 16756 266924 16884 266956
rect 16916 266924 16920 266956
rect 16720 266920 16920 266924
rect 16720 266876 16920 266880
rect 16720 266844 16724 266876
rect 16756 266844 16884 266876
rect 16916 266844 16920 266876
rect 16720 266840 16920 266844
rect 16720 266796 16920 266800
rect 16720 266764 16724 266796
rect 16756 266764 16884 266796
rect 16916 266764 16920 266796
rect 16720 266760 16920 266764
rect 16720 266716 16920 266720
rect 16720 266684 16724 266716
rect 16756 266684 16884 266716
rect 16916 266684 16920 266716
rect 16720 266680 16920 266684
rect 16720 266636 16920 266640
rect 16720 266604 16724 266636
rect 16756 266604 16884 266636
rect 16916 266604 16920 266636
rect 16720 266600 16920 266604
rect 16720 266556 16920 266560
rect 16720 266524 16724 266556
rect 16756 266524 16884 266556
rect 16916 266524 16920 266556
rect 16720 266520 16920 266524
rect 16720 266476 16920 266480
rect 16720 266444 16724 266476
rect 16756 266444 16884 266476
rect 16916 266444 16920 266476
rect 16720 266440 16920 266444
rect 16720 266396 16920 266400
rect 16720 266364 16724 266396
rect 16756 266364 16884 266396
rect 16916 266364 16920 266396
rect 16720 266360 16920 266364
rect 16720 266316 16920 266320
rect 16720 266284 16724 266316
rect 16756 266284 16884 266316
rect 16916 266284 16920 266316
rect 16720 266280 16920 266284
rect 16720 266236 16920 266240
rect 16720 266204 16724 266236
rect 16756 266204 16884 266236
rect 16916 266204 16920 266236
rect 16720 266200 16920 266204
rect 16720 266156 16920 266160
rect 16720 266124 16724 266156
rect 16756 266124 16884 266156
rect 16916 266124 16920 266156
rect 16720 266120 16920 266124
rect 16720 266076 16920 266080
rect 16720 266044 16724 266076
rect 16756 266044 16884 266076
rect 16916 266044 16920 266076
rect 16720 266040 16920 266044
rect 16720 265996 16920 266000
rect 16720 265964 16724 265996
rect 16756 265964 16884 265996
rect 16916 265964 16920 265996
rect 16720 265960 16920 265964
rect 16720 265916 16920 265920
rect 16720 265884 16724 265916
rect 16756 265884 16884 265916
rect 16916 265884 16920 265916
rect 16720 265880 16920 265884
rect 16720 265836 16920 265840
rect 16720 265804 16724 265836
rect 16756 265804 16884 265836
rect 16916 265804 16920 265836
rect 16720 265800 16920 265804
rect 16720 265756 16920 265760
rect 16720 265724 16724 265756
rect 16756 265724 16884 265756
rect 16916 265724 16920 265756
rect 16720 265720 16920 265724
rect 16720 265676 16920 265680
rect 16720 265644 16724 265676
rect 16756 265644 16884 265676
rect 16916 265644 16920 265676
rect 16720 265640 16920 265644
rect 16720 265596 16920 265600
rect 16720 265564 16724 265596
rect 16756 265564 16884 265596
rect 16916 265564 16920 265596
rect 16720 265560 16920 265564
rect 16720 265516 16920 265520
rect 16720 265484 16724 265516
rect 16756 265484 16884 265516
rect 16916 265484 16920 265516
rect 16720 265480 16920 265484
rect 16720 265436 16920 265440
rect 16720 265404 16724 265436
rect 16756 265404 16884 265436
rect 16916 265404 16920 265436
rect 16720 265400 16920 265404
rect 16720 265356 16920 265360
rect 16720 265324 16724 265356
rect 16756 265324 16884 265356
rect 16916 265324 16920 265356
rect 16720 265320 16920 265324
rect 16720 265276 16920 265280
rect 16720 265244 16724 265276
rect 16756 265244 16884 265276
rect 16916 265244 16920 265276
rect 16720 265240 16920 265244
rect 16720 265196 16920 265200
rect 16720 265164 16724 265196
rect 16756 265164 16884 265196
rect 16916 265164 16920 265196
rect 16720 265160 16920 265164
rect 16720 265116 16920 265120
rect 16720 265084 16724 265116
rect 16756 265084 16884 265116
rect 16916 265084 16920 265116
rect 16720 265080 16920 265084
rect 16720 265036 16920 265040
rect 16720 265004 16724 265036
rect 16756 265004 16884 265036
rect 16916 265004 16920 265036
rect 16720 265000 16920 265004
rect 16720 264956 16920 264960
rect 16720 264924 16724 264956
rect 16756 264924 16884 264956
rect 16916 264924 16920 264956
rect 16720 264920 16920 264924
rect 16720 264876 16920 264880
rect 16720 264844 16724 264876
rect 16756 264844 16884 264876
rect 16916 264844 16920 264876
rect 16720 264840 16920 264844
rect 16720 264796 16920 264800
rect 16720 264764 16724 264796
rect 16756 264764 16884 264796
rect 16916 264764 16920 264796
rect 16720 264760 16920 264764
rect 16720 264716 16920 264720
rect 16720 264684 16724 264716
rect 16756 264684 16884 264716
rect 16916 264684 16920 264716
rect 16720 264680 16920 264684
rect 16720 264636 16920 264640
rect 16720 264604 16724 264636
rect 16756 264604 16884 264636
rect 16916 264604 16920 264636
rect 16720 264600 16920 264604
rect 16720 264556 16920 264560
rect 16720 264524 16724 264556
rect 16756 264524 16884 264556
rect 16916 264524 16920 264556
rect 16720 264520 16920 264524
rect 16720 264476 16920 264480
rect 16720 264444 16724 264476
rect 16756 264444 16884 264476
rect 16916 264444 16920 264476
rect 16720 264440 16920 264444
rect 16720 264396 16920 264400
rect 16720 264364 16724 264396
rect 16756 264364 16884 264396
rect 16916 264364 16920 264396
rect 16720 264360 16920 264364
rect 16720 264316 16920 264320
rect 16720 264284 16724 264316
rect 16756 264284 16884 264316
rect 16916 264284 16920 264316
rect 16720 264280 16920 264284
rect 16720 264236 16920 264240
rect 16720 264204 16724 264236
rect 16756 264204 16884 264236
rect 16916 264204 16920 264236
rect 16720 264200 16920 264204
rect 16720 264156 16920 264160
rect 16720 264124 16724 264156
rect 16756 264124 16884 264156
rect 16916 264124 16920 264156
rect 16720 264120 16920 264124
rect 16720 264076 16920 264080
rect 16720 264044 16724 264076
rect 16756 264044 16884 264076
rect 16916 264044 16920 264076
rect 16720 264040 16920 264044
rect 16720 263996 16920 264000
rect 16720 263964 16724 263996
rect 16756 263964 16884 263996
rect 16916 263964 16920 263996
rect 16720 263960 16920 263964
rect 16720 263916 16920 263920
rect 16720 263884 16724 263916
rect 16756 263884 16884 263916
rect 16916 263884 16920 263916
rect 16720 263880 16920 263884
rect 16720 263836 16920 263840
rect 16720 263804 16724 263836
rect 16756 263804 16884 263836
rect 16916 263804 16920 263836
rect 16720 263800 16920 263804
rect 16720 263756 16920 263760
rect 16720 263724 16724 263756
rect 16756 263724 16884 263756
rect 16916 263724 16920 263756
rect 16720 263720 16920 263724
rect 16720 263676 16920 263680
rect 16720 263644 16724 263676
rect 16756 263644 16884 263676
rect 16916 263644 16920 263676
rect 16720 263640 16920 263644
rect 16720 263596 16920 263600
rect 16720 263564 16724 263596
rect 16756 263564 16884 263596
rect 16916 263564 16920 263596
rect 16720 263560 16920 263564
rect 16720 263516 16920 263520
rect 16720 263484 16724 263516
rect 16756 263484 16884 263516
rect 16916 263484 16920 263516
rect 16720 263480 16920 263484
rect 16720 263436 16920 263440
rect 16720 263404 16724 263436
rect 16756 263404 16884 263436
rect 16916 263404 16920 263436
rect 16720 263400 16920 263404
rect 16720 263356 16920 263360
rect 16720 263324 16724 263356
rect 16756 263324 16884 263356
rect 16916 263324 16920 263356
rect 16720 263320 16920 263324
rect 16720 263276 16920 263280
rect 16720 263244 16724 263276
rect 16756 263244 16884 263276
rect 16916 263244 16920 263276
rect 16720 263240 16920 263244
rect 16720 263196 16920 263200
rect 16720 263164 16724 263196
rect 16756 263164 16884 263196
rect 16916 263164 16920 263196
rect 16720 263160 16920 263164
rect 16720 263116 16920 263120
rect 16720 263084 16724 263116
rect 16756 263084 16884 263116
rect 16916 263084 16920 263116
rect 16720 263080 16920 263084
rect 16720 263036 16920 263040
rect 16720 263004 16724 263036
rect 16756 263004 16884 263036
rect 16916 263004 16920 263036
rect 16720 263000 16920 263004
rect 16720 262956 16920 262960
rect 16720 262924 16724 262956
rect 16756 262924 16884 262956
rect 16916 262924 16920 262956
rect 16720 262920 16920 262924
rect 16720 262876 16920 262880
rect 16720 262844 16724 262876
rect 16756 262844 16884 262876
rect 16916 262844 16920 262876
rect 16720 262840 16920 262844
rect 16720 262796 16920 262800
rect 16720 262764 16724 262796
rect 16756 262764 16884 262796
rect 16916 262764 16920 262796
rect 16720 262760 16920 262764
rect 16720 262716 16920 262720
rect 16720 262684 16724 262716
rect 16756 262684 16884 262716
rect 16916 262684 16920 262716
rect 16720 262680 16920 262684
rect 16720 262636 16920 262640
rect 16720 262604 16724 262636
rect 16756 262604 16884 262636
rect 16916 262604 16920 262636
rect 16720 262600 16920 262604
rect 16720 262556 16920 262560
rect 16720 262524 16724 262556
rect 16756 262524 16884 262556
rect 16916 262524 16920 262556
rect 16720 262520 16920 262524
rect 16720 262476 16920 262480
rect 16720 262444 16724 262476
rect 16756 262444 16884 262476
rect 16916 262444 16920 262476
rect 16720 262440 16920 262444
rect 16720 262396 16920 262400
rect 16720 262364 16724 262396
rect 16756 262364 16884 262396
rect 16916 262364 16920 262396
rect 16720 262360 16920 262364
rect 16720 262316 16920 262320
rect 16720 262284 16724 262316
rect 16756 262284 16884 262316
rect 16916 262284 16920 262316
rect 16720 262280 16920 262284
rect 16720 262236 16920 262240
rect 16720 262204 16724 262236
rect 16756 262204 16884 262236
rect 16916 262204 16920 262236
rect 16720 262200 16920 262204
rect 16720 262156 16920 262160
rect 16720 262124 16724 262156
rect 16756 262124 16884 262156
rect 16916 262124 16920 262156
rect 16720 262120 16920 262124
rect 16720 262076 16920 262080
rect 16720 262044 16724 262076
rect 16756 262044 16884 262076
rect 16916 262044 16920 262076
rect 16720 262040 16920 262044
rect 16720 261996 16920 262000
rect 16720 261964 16724 261996
rect 16756 261964 16884 261996
rect 16916 261964 16920 261996
rect 16720 261960 16920 261964
rect 16720 261916 16920 261920
rect 16720 261884 16724 261916
rect 16756 261884 16884 261916
rect 16916 261884 16920 261916
rect 16720 261880 16920 261884
rect 16720 261836 16920 261840
rect 16720 261804 16724 261836
rect 16756 261804 16884 261836
rect 16916 261804 16920 261836
rect 16720 261800 16920 261804
rect 16720 261756 16920 261760
rect 16720 261724 16724 261756
rect 16756 261724 16884 261756
rect 16916 261724 16920 261756
rect 16720 261720 16920 261724
rect 16720 261676 16920 261680
rect 16720 261644 16724 261676
rect 16756 261644 16884 261676
rect 16916 261644 16920 261676
rect 16720 261640 16920 261644
rect 16720 261596 16920 261600
rect 16720 261564 16724 261596
rect 16756 261564 16884 261596
rect 16916 261564 16920 261596
rect 16720 261560 16920 261564
rect 16720 261516 16920 261520
rect 16720 261484 16724 261516
rect 16756 261484 16884 261516
rect 16916 261484 16920 261516
rect 16720 261480 16920 261484
rect 16720 261436 16920 261440
rect 16720 261404 16724 261436
rect 16756 261404 16884 261436
rect 16916 261404 16920 261436
rect 16720 261400 16920 261404
rect 16720 261356 16920 261360
rect 16720 261324 16724 261356
rect 16756 261324 16884 261356
rect 16916 261324 16920 261356
rect 16720 261320 16920 261324
rect 16720 261276 16920 261280
rect 16720 261244 16724 261276
rect 16756 261244 16884 261276
rect 16916 261244 16920 261276
rect 16720 261240 16920 261244
rect 16720 261196 16920 261200
rect 16720 261164 16724 261196
rect 16756 261164 16884 261196
rect 16916 261164 16920 261196
rect 16720 261160 16920 261164
rect 16720 261116 16920 261120
rect 16720 261084 16724 261116
rect 16756 261084 16884 261116
rect 16916 261084 16920 261116
rect 16720 261080 16920 261084
rect 16720 261036 16920 261040
rect 16720 261004 16724 261036
rect 16756 261004 16884 261036
rect 16916 261004 16920 261036
rect 16720 261000 16920 261004
rect 16720 260956 16920 260960
rect 16720 260924 16724 260956
rect 16756 260924 16884 260956
rect 16916 260924 16920 260956
rect 16720 260920 16920 260924
rect 16720 260876 16920 260880
rect 16720 260844 16724 260876
rect 16756 260844 16884 260876
rect 16916 260844 16920 260876
rect 16720 260840 16920 260844
rect 16720 260796 16920 260800
rect 16720 260764 16724 260796
rect 16756 260764 16884 260796
rect 16916 260764 16920 260796
rect 16720 260760 16920 260764
rect 16720 260716 16920 260720
rect 16720 260684 16724 260716
rect 16756 260684 16884 260716
rect 16916 260684 16920 260716
rect 16720 260680 16920 260684
rect 16720 260636 16920 260640
rect 16720 260604 16724 260636
rect 16756 260604 16884 260636
rect 16916 260604 16920 260636
rect 16720 260600 16920 260604
rect 16720 260556 16920 260560
rect 16720 260524 16724 260556
rect 16756 260524 16884 260556
rect 16916 260524 16920 260556
rect 16720 260520 16920 260524
rect 16720 260476 16920 260480
rect 16720 260444 16724 260476
rect 16756 260444 16884 260476
rect 16916 260444 16920 260476
rect 16720 260440 16920 260444
rect 16720 260396 16920 260400
rect 16720 260364 16724 260396
rect 16756 260364 16884 260396
rect 16916 260364 16920 260396
rect 16720 260360 16920 260364
rect 16720 260316 16920 260320
rect 16720 260284 16724 260316
rect 16756 260284 16884 260316
rect 16916 260284 16920 260316
rect 16720 260280 16920 260284
rect 16720 260236 16920 260240
rect 16720 260204 16724 260236
rect 16756 260204 16884 260236
rect 16916 260204 16920 260236
rect 16720 260200 16920 260204
rect 16720 260156 16920 260160
rect 16720 260124 16724 260156
rect 16756 260124 16884 260156
rect 16916 260124 16920 260156
rect 16720 260120 16920 260124
rect 16720 260076 16920 260080
rect 16720 260044 16724 260076
rect 16756 260044 16884 260076
rect 16916 260044 16920 260076
rect 16720 260040 16920 260044
rect 16720 259996 16920 260000
rect 16720 259964 16724 259996
rect 16756 259964 16884 259996
rect 16916 259964 16920 259996
rect 16720 259960 16920 259964
rect 16720 259916 16920 259920
rect 16720 259884 16724 259916
rect 16756 259884 16884 259916
rect 16916 259884 16920 259916
rect 16720 259880 16920 259884
rect 16720 259836 16920 259840
rect 16720 259804 16724 259836
rect 16756 259804 16884 259836
rect 16916 259804 16920 259836
rect 16720 259800 16920 259804
rect 16720 259756 16920 259760
rect 16720 259724 16724 259756
rect 16756 259724 16884 259756
rect 16916 259724 16920 259756
rect 16720 259720 16920 259724
rect 16720 259676 16920 259680
rect 16720 259644 16724 259676
rect 16756 259644 16884 259676
rect 16916 259644 16920 259676
rect 16720 259640 16920 259644
rect 16720 259596 16920 259600
rect 16720 259564 16724 259596
rect 16756 259564 16884 259596
rect 16916 259564 16920 259596
rect 16720 259560 16920 259564
rect 16720 259516 16920 259520
rect 16720 259484 16724 259516
rect 16756 259484 16884 259516
rect 16916 259484 16920 259516
rect 16720 259480 16920 259484
rect 16720 259436 16920 259440
rect 16720 259404 16724 259436
rect 16756 259404 16884 259436
rect 16916 259404 16920 259436
rect 16720 259400 16920 259404
rect 16720 259356 16920 259360
rect 16720 259324 16724 259356
rect 16756 259324 16884 259356
rect 16916 259324 16920 259356
rect 16720 259320 16920 259324
rect 16720 259276 16920 259280
rect 16720 259244 16724 259276
rect 16756 259244 16884 259276
rect 16916 259244 16920 259276
rect 16720 259240 16920 259244
rect 16720 259196 16920 259200
rect 16720 259164 16724 259196
rect 16756 259164 16884 259196
rect 16916 259164 16920 259196
rect 16720 259160 16920 259164
rect 16720 259116 16920 259120
rect 16720 259084 16724 259116
rect 16756 259084 16884 259116
rect 16916 259084 16920 259116
rect 16720 259080 16920 259084
rect 16720 259036 16920 259040
rect 16720 259004 16724 259036
rect 16756 259004 16884 259036
rect 16916 259004 16920 259036
rect 16720 259000 16920 259004
rect 16720 258956 16920 258960
rect 16720 258924 16724 258956
rect 16756 258924 16884 258956
rect 16916 258924 16920 258956
rect 16720 258920 16920 258924
rect 16720 258876 16920 258880
rect 16720 258844 16724 258876
rect 16756 258844 16884 258876
rect 16916 258844 16920 258876
rect 16720 258840 16920 258844
rect 16720 258796 16920 258800
rect 16720 258764 16724 258796
rect 16756 258764 16884 258796
rect 16916 258764 16920 258796
rect 16720 258760 16920 258764
rect 16720 258716 16920 258720
rect 16720 258684 16724 258716
rect 16756 258684 16884 258716
rect 16916 258684 16920 258716
rect 16720 258680 16920 258684
rect 16720 258636 16920 258640
rect 16720 258604 16724 258636
rect 16756 258604 16884 258636
rect 16916 258604 16920 258636
rect 16720 258600 16920 258604
rect 16720 258556 16920 258560
rect 16720 258524 16724 258556
rect 16756 258524 16884 258556
rect 16916 258524 16920 258556
rect 16720 258520 16920 258524
rect 16720 258476 16920 258480
rect 16720 258444 16724 258476
rect 16756 258444 16884 258476
rect 16916 258444 16920 258476
rect 16720 258440 16920 258444
rect 16720 258396 16920 258400
rect 16720 258364 16724 258396
rect 16756 258364 16884 258396
rect 16916 258364 16920 258396
rect 16720 258360 16920 258364
rect 16720 258316 16920 258320
rect 16720 258284 16724 258316
rect 16756 258284 16884 258316
rect 16916 258284 16920 258316
rect 16720 258280 16920 258284
rect 16720 258236 16920 258240
rect 16720 258204 16724 258236
rect 16756 258204 16884 258236
rect 16916 258204 16920 258236
rect 16720 258200 16920 258204
rect 16720 258156 16920 258160
rect 16720 258124 16724 258156
rect 16756 258124 16884 258156
rect 16916 258124 16920 258156
rect 16720 258120 16920 258124
rect 16720 258076 16920 258080
rect 16720 258044 16724 258076
rect 16756 258044 16884 258076
rect 16916 258044 16920 258076
rect 16720 258040 16920 258044
rect 16720 257996 16920 258000
rect 16720 257964 16724 257996
rect 16756 257964 16884 257996
rect 16916 257964 16920 257996
rect 16720 257960 16920 257964
rect 16720 257916 16920 257920
rect 16720 257884 16724 257916
rect 16756 257884 16884 257916
rect 16916 257884 16920 257916
rect 16720 257880 16920 257884
rect 16720 257836 16920 257840
rect 16720 257804 16724 257836
rect 16756 257804 16884 257836
rect 16916 257804 16920 257836
rect 16720 257800 16920 257804
rect 16720 257756 16920 257760
rect 16720 257724 16724 257756
rect 16756 257724 16884 257756
rect 16916 257724 16920 257756
rect 16720 257720 16920 257724
rect 16720 257676 16920 257680
rect 16720 257644 16724 257676
rect 16756 257644 16884 257676
rect 16916 257644 16920 257676
rect 16720 257640 16920 257644
rect 16720 257596 16920 257600
rect 16720 257564 16724 257596
rect 16756 257564 16884 257596
rect 16916 257564 16920 257596
rect 16720 257560 16920 257564
rect 16720 257516 16920 257520
rect 16720 257484 16724 257516
rect 16756 257484 16884 257516
rect 16916 257484 16920 257516
rect 16720 257480 16920 257484
rect 16720 257436 16920 257440
rect 16720 257404 16724 257436
rect 16756 257404 16884 257436
rect 16916 257404 16920 257436
rect 16720 257400 16920 257404
rect 16720 257356 16920 257360
rect 16720 257324 16724 257356
rect 16756 257324 16884 257356
rect 16916 257324 16920 257356
rect 16720 257320 16920 257324
rect 16720 257276 16920 257280
rect 16720 257244 16724 257276
rect 16756 257244 16884 257276
rect 16916 257244 16920 257276
rect 16720 257240 16920 257244
rect 16720 257196 16920 257200
rect 16720 257164 16724 257196
rect 16756 257164 16884 257196
rect 16916 257164 16920 257196
rect 16720 257160 16920 257164
rect 16720 257116 16920 257120
rect 16720 257084 16724 257116
rect 16756 257084 16884 257116
rect 16916 257084 16920 257116
rect 16720 257080 16920 257084
rect 16720 257036 16920 257040
rect 16720 257004 16724 257036
rect 16756 257004 16884 257036
rect 16916 257004 16920 257036
rect 16720 257000 16920 257004
rect 16720 256956 16920 256960
rect 16720 256924 16724 256956
rect 16756 256924 16884 256956
rect 16916 256924 16920 256956
rect 16720 256920 16920 256924
rect 16720 256876 16920 256880
rect 16720 256844 16724 256876
rect 16756 256844 16884 256876
rect 16916 256844 16920 256876
rect 16720 256840 16920 256844
rect 16720 256796 16920 256800
rect 16720 256764 16724 256796
rect 16756 256764 16884 256796
rect 16916 256764 16920 256796
rect 16720 256760 16920 256764
rect 16720 256716 16920 256720
rect 16720 256684 16724 256716
rect 16756 256684 16884 256716
rect 16916 256684 16920 256716
rect 16720 256680 16920 256684
rect 16720 256636 16920 256640
rect 16720 256604 16724 256636
rect 16756 256604 16884 256636
rect 16916 256604 16920 256636
rect 16720 256600 16920 256604
rect 16720 256556 16920 256560
rect 16720 256524 16724 256556
rect 16756 256524 16884 256556
rect 16916 256524 16920 256556
rect 16720 256520 16920 256524
rect 16720 256476 16920 256480
rect 16720 256444 16724 256476
rect 16756 256444 16884 256476
rect 16916 256444 16920 256476
rect 16720 256440 16920 256444
rect 16720 256396 16920 256400
rect 16720 256364 16724 256396
rect 16756 256364 16884 256396
rect 16916 256364 16920 256396
rect 16720 256360 16920 256364
rect 16720 256316 16920 256320
rect 16720 256284 16724 256316
rect 16756 256284 16884 256316
rect 16916 256284 16920 256316
rect 16720 256280 16920 256284
rect 16720 256236 16920 256240
rect 16720 256204 16724 256236
rect 16756 256204 16884 256236
rect 16916 256204 16920 256236
rect 16720 256200 16920 256204
rect 16720 256156 16920 256160
rect 16720 256124 16724 256156
rect 16756 256124 16884 256156
rect 16916 256124 16920 256156
rect 16720 256120 16920 256124
rect 16720 256076 16920 256080
rect 16720 256044 16724 256076
rect 16756 256044 16884 256076
rect 16916 256044 16920 256076
rect 16720 256040 16920 256044
rect 16720 255996 16920 256000
rect 16720 255964 16724 255996
rect 16756 255964 16884 255996
rect 16916 255964 16920 255996
rect 16720 255960 16920 255964
rect 400 255876 16920 255880
rect 400 255844 404 255876
rect 436 255844 484 255876
rect 516 255844 564 255876
rect 596 255844 644 255876
rect 676 255844 724 255876
rect 756 255844 804 255876
rect 836 255844 884 255876
rect 916 255844 964 255876
rect 996 255844 1044 255876
rect 1076 255844 1124 255876
rect 1156 255844 1204 255876
rect 1236 255844 1284 255876
rect 1316 255844 1364 255876
rect 1396 255844 1444 255876
rect 1476 255844 1524 255876
rect 1556 255844 1604 255876
rect 1636 255844 1684 255876
rect 1716 255844 1764 255876
rect 1796 255844 1844 255876
rect 1876 255844 1924 255876
rect 1956 255844 2004 255876
rect 2036 255844 2084 255876
rect 2116 255844 2164 255876
rect 2196 255844 2244 255876
rect 2276 255844 2324 255876
rect 2356 255844 2404 255876
rect 2436 255844 2484 255876
rect 2516 255844 2564 255876
rect 2596 255844 2644 255876
rect 2676 255844 2724 255876
rect 2756 255844 3044 255876
rect 3076 255844 3124 255876
rect 3156 255844 3204 255876
rect 3236 255844 3284 255876
rect 3316 255844 3364 255876
rect 3396 255844 3444 255876
rect 3476 255844 3524 255876
rect 3556 255844 3604 255876
rect 3636 255844 3684 255876
rect 3716 255844 3764 255876
rect 3796 255844 3844 255876
rect 3876 255844 3924 255876
rect 3956 255844 4004 255876
rect 4036 255844 4084 255876
rect 4116 255844 4164 255876
rect 4196 255844 4244 255876
rect 4276 255844 4324 255876
rect 4356 255844 4404 255876
rect 4436 255844 4484 255876
rect 4516 255844 4564 255876
rect 4596 255844 4644 255876
rect 4676 255844 4724 255876
rect 4756 255844 4804 255876
rect 4836 255844 4884 255876
rect 4916 255844 4964 255876
rect 4996 255844 5044 255876
rect 5076 255844 5124 255876
rect 5156 255844 5204 255876
rect 5236 255844 5284 255876
rect 5316 255844 5364 255876
rect 5396 255844 5444 255876
rect 5476 255844 5524 255876
rect 5556 255844 5604 255876
rect 5636 255844 5684 255876
rect 5716 255844 5764 255876
rect 5796 255844 5844 255876
rect 5876 255844 5924 255876
rect 5956 255844 6004 255876
rect 6036 255844 6084 255876
rect 6116 255844 6164 255876
rect 6196 255844 6244 255876
rect 6276 255844 6324 255876
rect 6356 255844 6404 255876
rect 6436 255844 6484 255876
rect 6516 255844 6564 255876
rect 6596 255844 6644 255876
rect 6676 255844 6724 255876
rect 6756 255844 6804 255876
rect 6836 255844 6884 255876
rect 6916 255844 6964 255876
rect 6996 255844 7044 255876
rect 7076 255844 7124 255876
rect 7156 255844 7204 255876
rect 7236 255844 7284 255876
rect 7316 255844 7364 255876
rect 7396 255844 7444 255876
rect 7476 255844 7524 255876
rect 7556 255844 7604 255876
rect 7636 255844 7684 255876
rect 7716 255844 7764 255876
rect 7796 255844 7844 255876
rect 7876 255844 7924 255876
rect 7956 255844 8004 255876
rect 8036 255844 8084 255876
rect 8116 255844 8164 255876
rect 8196 255844 8244 255876
rect 8276 255844 8324 255876
rect 8356 255844 8404 255876
rect 8436 255844 8484 255876
rect 8516 255844 8564 255876
rect 8596 255844 8644 255876
rect 8676 255844 8724 255876
rect 8756 255844 8804 255876
rect 8836 255844 8884 255876
rect 8916 255844 8964 255876
rect 8996 255844 9044 255876
rect 9076 255844 9124 255876
rect 9156 255844 9204 255876
rect 9236 255844 9284 255876
rect 9316 255844 9364 255876
rect 9396 255844 9444 255876
rect 9476 255844 9524 255876
rect 9556 255844 9604 255876
rect 9636 255844 9684 255876
rect 9716 255844 9764 255876
rect 9796 255844 9844 255876
rect 9876 255844 9924 255876
rect 9956 255844 10004 255876
rect 10036 255844 10084 255876
rect 10116 255844 10164 255876
rect 10196 255844 10244 255876
rect 10276 255844 10324 255876
rect 10356 255844 10404 255876
rect 10436 255844 10484 255876
rect 10516 255844 10564 255876
rect 10596 255844 10644 255876
rect 10676 255844 10724 255876
rect 10756 255844 10804 255876
rect 10836 255844 10884 255876
rect 10916 255844 10964 255876
rect 10996 255844 11044 255876
rect 11076 255844 11124 255876
rect 11156 255844 11204 255876
rect 11236 255844 11284 255876
rect 11316 255844 11364 255876
rect 11396 255844 11444 255876
rect 11476 255844 11524 255876
rect 11556 255844 11604 255876
rect 11636 255844 11684 255876
rect 11716 255844 11764 255876
rect 11796 255844 11844 255876
rect 11876 255844 11924 255876
rect 11956 255844 12004 255876
rect 12036 255844 12084 255876
rect 12116 255844 12164 255876
rect 12196 255844 12244 255876
rect 12276 255844 12324 255876
rect 12356 255844 12404 255876
rect 12436 255844 12484 255876
rect 12516 255844 12564 255876
rect 12596 255844 12644 255876
rect 12676 255844 12724 255876
rect 12756 255844 12804 255876
rect 12836 255844 12884 255876
rect 12916 255844 12964 255876
rect 12996 255844 13044 255876
rect 13076 255844 13124 255876
rect 13156 255844 13204 255876
rect 13236 255844 13284 255876
rect 13316 255844 13364 255876
rect 13396 255844 13444 255876
rect 13476 255844 13524 255876
rect 13556 255844 13604 255876
rect 13636 255844 13684 255876
rect 13716 255844 13764 255876
rect 13796 255844 13844 255876
rect 13876 255844 13924 255876
rect 13956 255844 14004 255876
rect 14036 255844 14084 255876
rect 14116 255844 14164 255876
rect 14196 255844 14244 255876
rect 14276 255844 14324 255876
rect 14356 255844 14404 255876
rect 14436 255844 14484 255876
rect 14516 255844 14564 255876
rect 14596 255844 14644 255876
rect 14676 255844 14724 255876
rect 14756 255844 14804 255876
rect 14836 255844 14884 255876
rect 14916 255844 14964 255876
rect 14996 255844 15044 255876
rect 15076 255844 15124 255876
rect 15156 255844 15204 255876
rect 15236 255844 15284 255876
rect 15316 255844 15364 255876
rect 15396 255844 15444 255876
rect 15476 255844 15524 255876
rect 15556 255844 15604 255876
rect 15636 255844 15684 255876
rect 15716 255844 15764 255876
rect 15796 255844 15844 255876
rect 15876 255844 15924 255876
rect 15956 255844 16004 255876
rect 16036 255844 16084 255876
rect 16116 255844 16164 255876
rect 16196 255844 16244 255876
rect 16276 255844 16324 255876
rect 16356 255844 16404 255876
rect 16436 255844 16484 255876
rect 16516 255844 16564 255876
rect 16596 255844 16644 255876
rect 16676 255844 16724 255876
rect 16756 255844 16884 255876
rect 16916 255844 16920 255876
rect 400 255840 16920 255844
rect 400 255796 16840 255800
rect 400 255764 404 255796
rect 436 255764 484 255796
rect 516 255764 564 255796
rect 596 255764 644 255796
rect 676 255764 724 255796
rect 756 255764 804 255796
rect 836 255764 884 255796
rect 916 255764 964 255796
rect 996 255764 1044 255796
rect 1076 255764 1124 255796
rect 1156 255764 1204 255796
rect 1236 255764 1284 255796
rect 1316 255764 1364 255796
rect 1396 255764 1444 255796
rect 1476 255764 1524 255796
rect 1556 255764 1604 255796
rect 1636 255764 1684 255796
rect 1716 255764 1764 255796
rect 1796 255764 1844 255796
rect 1876 255764 1924 255796
rect 1956 255764 2004 255796
rect 2036 255764 2084 255796
rect 2116 255764 2164 255796
rect 2196 255764 2244 255796
rect 2276 255764 2324 255796
rect 2356 255764 2404 255796
rect 2436 255764 2484 255796
rect 2516 255764 2564 255796
rect 2596 255764 2644 255796
rect 2676 255764 2724 255796
rect 2756 255764 3044 255796
rect 3076 255764 3124 255796
rect 3156 255764 3204 255796
rect 3236 255764 3284 255796
rect 3316 255764 3364 255796
rect 3396 255764 3444 255796
rect 3476 255764 3524 255796
rect 3556 255764 3604 255796
rect 3636 255764 3684 255796
rect 3716 255764 3764 255796
rect 3796 255764 3844 255796
rect 3876 255764 3924 255796
rect 3956 255764 4004 255796
rect 4036 255764 4084 255796
rect 4116 255764 4164 255796
rect 4196 255764 4244 255796
rect 4276 255764 4324 255796
rect 4356 255764 4404 255796
rect 4436 255764 4484 255796
rect 4516 255764 4564 255796
rect 4596 255764 4644 255796
rect 4676 255764 4724 255796
rect 4756 255764 4804 255796
rect 4836 255764 4884 255796
rect 4916 255764 4964 255796
rect 4996 255764 5044 255796
rect 5076 255764 5124 255796
rect 5156 255764 5204 255796
rect 5236 255764 5284 255796
rect 5316 255764 5364 255796
rect 5396 255764 5444 255796
rect 5476 255764 5524 255796
rect 5556 255764 5604 255796
rect 5636 255764 5684 255796
rect 5716 255764 5764 255796
rect 5796 255764 5844 255796
rect 5876 255764 5924 255796
rect 5956 255764 6004 255796
rect 6036 255764 6084 255796
rect 6116 255764 6164 255796
rect 6196 255764 6244 255796
rect 6276 255764 6324 255796
rect 6356 255764 6404 255796
rect 6436 255764 6484 255796
rect 6516 255764 6564 255796
rect 6596 255764 6644 255796
rect 6676 255764 6724 255796
rect 6756 255764 6804 255796
rect 6836 255764 6884 255796
rect 6916 255764 6964 255796
rect 6996 255764 7044 255796
rect 7076 255764 7124 255796
rect 7156 255764 7204 255796
rect 7236 255764 7284 255796
rect 7316 255764 7364 255796
rect 7396 255764 7444 255796
rect 7476 255764 7524 255796
rect 7556 255764 7604 255796
rect 7636 255764 7684 255796
rect 7716 255764 7764 255796
rect 7796 255764 7844 255796
rect 7876 255764 7924 255796
rect 7956 255764 8004 255796
rect 8036 255764 8084 255796
rect 8116 255764 8164 255796
rect 8196 255764 8244 255796
rect 8276 255764 8324 255796
rect 8356 255764 8404 255796
rect 8436 255764 8484 255796
rect 8516 255764 8564 255796
rect 8596 255764 8644 255796
rect 8676 255764 8724 255796
rect 8756 255764 8804 255796
rect 8836 255764 8884 255796
rect 8916 255764 8964 255796
rect 8996 255764 9044 255796
rect 9076 255764 9124 255796
rect 9156 255764 9204 255796
rect 9236 255764 9284 255796
rect 9316 255764 9364 255796
rect 9396 255764 9444 255796
rect 9476 255764 9524 255796
rect 9556 255764 9604 255796
rect 9636 255764 9684 255796
rect 9716 255764 9764 255796
rect 9796 255764 9844 255796
rect 9876 255764 9924 255796
rect 9956 255764 10004 255796
rect 10036 255764 10084 255796
rect 10116 255764 10164 255796
rect 10196 255764 10244 255796
rect 10276 255764 10324 255796
rect 10356 255764 10404 255796
rect 10436 255764 10484 255796
rect 10516 255764 10564 255796
rect 10596 255764 10644 255796
rect 10676 255764 10724 255796
rect 10756 255764 10804 255796
rect 10836 255764 10884 255796
rect 10916 255764 10964 255796
rect 10996 255764 11044 255796
rect 11076 255764 11124 255796
rect 11156 255764 11204 255796
rect 11236 255764 11284 255796
rect 11316 255764 11364 255796
rect 11396 255764 11444 255796
rect 11476 255764 11524 255796
rect 11556 255764 11604 255796
rect 11636 255764 11684 255796
rect 11716 255764 11764 255796
rect 11796 255764 11844 255796
rect 11876 255764 11924 255796
rect 11956 255764 12004 255796
rect 12036 255764 12084 255796
rect 12116 255764 12164 255796
rect 12196 255764 12244 255796
rect 12276 255764 12324 255796
rect 12356 255764 12404 255796
rect 12436 255764 12484 255796
rect 12516 255764 12564 255796
rect 12596 255764 12644 255796
rect 12676 255764 12724 255796
rect 12756 255764 12804 255796
rect 12836 255764 12884 255796
rect 12916 255764 12964 255796
rect 12996 255764 13044 255796
rect 13076 255764 13124 255796
rect 13156 255764 13204 255796
rect 13236 255764 13284 255796
rect 13316 255764 13364 255796
rect 13396 255764 13444 255796
rect 13476 255764 13524 255796
rect 13556 255764 13604 255796
rect 13636 255764 13684 255796
rect 13716 255764 13764 255796
rect 13796 255764 13844 255796
rect 13876 255764 13924 255796
rect 13956 255764 14004 255796
rect 14036 255764 14084 255796
rect 14116 255764 14164 255796
rect 14196 255764 14244 255796
rect 14276 255764 14324 255796
rect 14356 255764 14404 255796
rect 14436 255764 14484 255796
rect 14516 255764 14564 255796
rect 14596 255764 14644 255796
rect 14676 255764 14724 255796
rect 14756 255764 14804 255796
rect 14836 255764 14884 255796
rect 14916 255764 14964 255796
rect 14996 255764 15044 255796
rect 15076 255764 15124 255796
rect 15156 255764 15204 255796
rect 15236 255764 15284 255796
rect 15316 255764 15364 255796
rect 15396 255764 15444 255796
rect 15476 255764 15524 255796
rect 15556 255764 15604 255796
rect 15636 255764 15684 255796
rect 15716 255764 15764 255796
rect 15796 255764 15844 255796
rect 15876 255764 15924 255796
rect 15956 255764 16004 255796
rect 16036 255764 16084 255796
rect 16116 255764 16164 255796
rect 16196 255764 16244 255796
rect 16276 255764 16324 255796
rect 16356 255764 16404 255796
rect 16436 255764 16484 255796
rect 16516 255764 16564 255796
rect 16596 255764 16644 255796
rect 16676 255764 16724 255796
rect 16756 255764 16840 255796
rect 400 255760 16840 255764
rect 400 255716 16920 255720
rect 400 255684 404 255716
rect 436 255684 484 255716
rect 516 255684 564 255716
rect 596 255684 644 255716
rect 676 255684 724 255716
rect 756 255684 804 255716
rect 836 255684 884 255716
rect 916 255684 964 255716
rect 996 255684 1044 255716
rect 1076 255684 1124 255716
rect 1156 255684 1204 255716
rect 1236 255684 1284 255716
rect 1316 255684 1364 255716
rect 1396 255684 1444 255716
rect 1476 255684 1524 255716
rect 1556 255684 1604 255716
rect 1636 255684 1684 255716
rect 1716 255684 1764 255716
rect 1796 255684 1844 255716
rect 1876 255684 1924 255716
rect 1956 255684 2004 255716
rect 2036 255684 2084 255716
rect 2116 255684 2164 255716
rect 2196 255684 2244 255716
rect 2276 255684 2324 255716
rect 2356 255684 2404 255716
rect 2436 255684 2484 255716
rect 2516 255684 2564 255716
rect 2596 255684 2644 255716
rect 2676 255684 2724 255716
rect 2756 255684 3044 255716
rect 3076 255684 3124 255716
rect 3156 255684 3204 255716
rect 3236 255684 3284 255716
rect 3316 255684 3364 255716
rect 3396 255684 3444 255716
rect 3476 255684 3524 255716
rect 3556 255684 3604 255716
rect 3636 255684 3684 255716
rect 3716 255684 3764 255716
rect 3796 255684 3844 255716
rect 3876 255684 3924 255716
rect 3956 255684 4004 255716
rect 4036 255684 4084 255716
rect 4116 255684 4164 255716
rect 4196 255684 4244 255716
rect 4276 255684 4324 255716
rect 4356 255684 4404 255716
rect 4436 255684 4484 255716
rect 4516 255684 4564 255716
rect 4596 255684 4644 255716
rect 4676 255684 4724 255716
rect 4756 255684 4804 255716
rect 4836 255684 4884 255716
rect 4916 255684 4964 255716
rect 4996 255684 5044 255716
rect 5076 255684 5124 255716
rect 5156 255684 5204 255716
rect 5236 255684 5284 255716
rect 5316 255684 5364 255716
rect 5396 255684 5444 255716
rect 5476 255684 5524 255716
rect 5556 255684 5604 255716
rect 5636 255684 5684 255716
rect 5716 255684 5764 255716
rect 5796 255684 5844 255716
rect 5876 255684 5924 255716
rect 5956 255684 6004 255716
rect 6036 255684 6084 255716
rect 6116 255684 6164 255716
rect 6196 255684 6244 255716
rect 6276 255684 6324 255716
rect 6356 255684 6404 255716
rect 6436 255684 6484 255716
rect 6516 255684 6564 255716
rect 6596 255684 6644 255716
rect 6676 255684 6724 255716
rect 6756 255684 6804 255716
rect 6836 255684 6884 255716
rect 6916 255684 6964 255716
rect 6996 255684 7044 255716
rect 7076 255684 7124 255716
rect 7156 255684 7204 255716
rect 7236 255684 7284 255716
rect 7316 255684 7364 255716
rect 7396 255684 7444 255716
rect 7476 255684 7524 255716
rect 7556 255684 7604 255716
rect 7636 255684 7684 255716
rect 7716 255684 7764 255716
rect 7796 255684 7844 255716
rect 7876 255684 7924 255716
rect 7956 255684 8004 255716
rect 8036 255684 8084 255716
rect 8116 255684 8164 255716
rect 8196 255684 8244 255716
rect 8276 255684 8324 255716
rect 8356 255684 8404 255716
rect 8436 255684 8484 255716
rect 8516 255684 8564 255716
rect 8596 255684 8644 255716
rect 8676 255684 8724 255716
rect 8756 255684 8804 255716
rect 8836 255684 8884 255716
rect 8916 255684 8964 255716
rect 8996 255684 9044 255716
rect 9076 255684 9124 255716
rect 9156 255684 9204 255716
rect 9236 255684 9284 255716
rect 9316 255684 9364 255716
rect 9396 255684 9444 255716
rect 9476 255684 9524 255716
rect 9556 255684 9604 255716
rect 9636 255684 9684 255716
rect 9716 255684 9764 255716
rect 9796 255684 9844 255716
rect 9876 255684 9924 255716
rect 9956 255684 10004 255716
rect 10036 255684 10084 255716
rect 10116 255684 10164 255716
rect 10196 255684 10244 255716
rect 10276 255684 10324 255716
rect 10356 255684 10404 255716
rect 10436 255684 10484 255716
rect 10516 255684 10564 255716
rect 10596 255684 10644 255716
rect 10676 255684 10724 255716
rect 10756 255684 10804 255716
rect 10836 255684 10884 255716
rect 10916 255684 10964 255716
rect 10996 255684 11044 255716
rect 11076 255684 11124 255716
rect 11156 255684 11204 255716
rect 11236 255684 11284 255716
rect 11316 255684 11364 255716
rect 11396 255684 11444 255716
rect 11476 255684 11524 255716
rect 11556 255684 11604 255716
rect 11636 255684 11684 255716
rect 11716 255684 11764 255716
rect 11796 255684 11844 255716
rect 11876 255684 11924 255716
rect 11956 255684 12004 255716
rect 12036 255684 12084 255716
rect 12116 255684 12164 255716
rect 12196 255684 12244 255716
rect 12276 255684 12324 255716
rect 12356 255684 12404 255716
rect 12436 255684 12484 255716
rect 12516 255684 12564 255716
rect 12596 255684 12644 255716
rect 12676 255684 12724 255716
rect 12756 255684 12804 255716
rect 12836 255684 12884 255716
rect 12916 255684 12964 255716
rect 12996 255684 13044 255716
rect 13076 255684 13124 255716
rect 13156 255684 13204 255716
rect 13236 255684 13284 255716
rect 13316 255684 13364 255716
rect 13396 255684 13444 255716
rect 13476 255684 13524 255716
rect 13556 255684 13604 255716
rect 13636 255684 13684 255716
rect 13716 255684 13764 255716
rect 13796 255684 13844 255716
rect 13876 255684 13924 255716
rect 13956 255684 14004 255716
rect 14036 255684 14084 255716
rect 14116 255684 14164 255716
rect 14196 255684 14244 255716
rect 14276 255684 14324 255716
rect 14356 255684 14404 255716
rect 14436 255684 14484 255716
rect 14516 255684 14564 255716
rect 14596 255684 14644 255716
rect 14676 255684 14724 255716
rect 14756 255684 14804 255716
rect 14836 255684 14884 255716
rect 14916 255684 14964 255716
rect 14996 255684 15044 255716
rect 15076 255684 15124 255716
rect 15156 255684 15204 255716
rect 15236 255684 15284 255716
rect 15316 255684 15364 255716
rect 15396 255684 15444 255716
rect 15476 255684 15524 255716
rect 15556 255684 15604 255716
rect 15636 255684 15684 255716
rect 15716 255684 15764 255716
rect 15796 255684 15844 255716
rect 15876 255684 15924 255716
rect 15956 255684 16004 255716
rect 16036 255684 16084 255716
rect 16116 255684 16164 255716
rect 16196 255684 16244 255716
rect 16276 255684 16324 255716
rect 16356 255684 16404 255716
rect 16436 255684 16484 255716
rect 16516 255684 16564 255716
rect 16596 255684 16644 255716
rect 16676 255684 16724 255716
rect 16756 255684 16884 255716
rect 16916 255684 16920 255716
rect 400 255680 16920 255684
<< metal5 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
<< comment >>
rect -50 352000 292050 352050
rect -50 0 0 352000
rect 292000 0 292050 352000
rect -50 -50 292050 0
use sbcs5v0  sbcs5v0_0 ../lib/sbcs5v0/mag
timestamp 1640892658
transform 1 0 262020 0 1 344380
box -1520 -5880 10040 5640
use sbcs1v8  sbcs1v8_1 ../lib/sbcs1v8/mag
timestamp 1640892658
transform 1 0 18720 0 1 269280
box -1520 -5880 10040 5640
use sbcs1v8  sbcs1v8_0
timestamp 1640892658
transform 1 0 4320 0 1 269280
box -1520 -5880 10040 5640
use vref1v8  vref1v8_0 ../lib/vref1v8/mag
timestamp 1641007606
transform -1 0 28040 0 -1 276480
box -720 -3720 11000 1080
<< labels >>
flabel metal3 s 291760 134615 292400 134671 0 FreeSans 560 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -400 190932 240 190988 0 FreeSans 560 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -400 169321 240 169377 0 FreeSans 560 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -400 147710 240 147766 0 FreeSans 560 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -400 126199 240 126255 0 FreeSans 560 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -400 62388 240 62444 0 FreeSans 560 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -400 40777 240 40833 0 FreeSans 560 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -400 19166 240 19222 0 FreeSans 560 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -400 8455 240 8511 0 FreeSans 560 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 291760 156826 292400 156882 0 FreeSans 560 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 291760 179437 292400 179493 0 FreeSans 560 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 291760 202648 292400 202704 0 FreeSans 560 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 291760 224859 292400 224915 0 FreeSans 560 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 291760 247070 292400 247126 0 FreeSans 560 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 291760 291781 292400 291837 0 FreeSans 560 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -400 255765 240 255821 0 FreeSans 560 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -400 234154 240 234210 0 FreeSans 560 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -400 212543 240 212599 0 FreeSans 560 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 291760 135206 292400 135262 0 FreeSans 560 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -400 190341 240 190397 0 FreeSans 560 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -400 168730 240 168786 0 FreeSans 560 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -400 147119 240 147175 0 FreeSans 560 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -400 125608 240 125664 0 FreeSans 560 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -400 61797 240 61853 0 FreeSans 560 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -400 40186 240 40242 0 FreeSans 560 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -400 18575 240 18631 0 FreeSans 560 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -400 7864 240 7920 0 FreeSans 560 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 291760 157417 292400 157473 0 FreeSans 560 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 291760 180028 292400 180084 0 FreeSans 560 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 291760 203239 292400 203295 0 FreeSans 560 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 291760 225450 292400 225506 0 FreeSans 560 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 291760 247661 292400 247717 0 FreeSans 560 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 291760 292372 292400 292428 0 FreeSans 560 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -400 255174 240 255230 0 FreeSans 560 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -400 233563 240 233619 0 FreeSans 560 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -400 211952 240 212008 0 FreeSans 560 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 291150 338992 292400 341492 0 FreeSans 560 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 340121 850 342621 0 FreeSans 560 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 283297 351150 285797 352400 0 FreeSans 960 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 232697 351150 235197 352400 0 FreeSans 960 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 206697 351150 209197 352400 0 FreeSans 960 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 60097 351150 62597 352400 0 FreeSans 960 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 34097 351150 36597 352400 0 FreeSans 960 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 8097 351150 10597 352400 0 FreeSans 960 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 163397 351150 164497 352400 0 FreeSans 960 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 112547 351150 113647 352400 0 FreeSans 960 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 86697 351150 87797 352400 0 FreeSans 960 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 162147 351150 163247 352400 0 FreeSans 960 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 111297 351150 112397 352400 0 FreeSans 960 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 85447 351150 86547 352400 0 FreeSans 960 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 291760 1363 292400 1419 0 FreeSans 560 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 291760 204421 292400 204477 0 FreeSans 560 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 291760 226632 292400 226688 0 FreeSans 560 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 291760 248843 292400 248899 0 FreeSans 560 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 291760 293554 292400 293610 0 FreeSans 560 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -400 253992 240 254048 0 FreeSans 560 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -400 232381 240 232437 0 FreeSans 560 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -400 210770 240 210826 0 FreeSans 560 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -400 189159 240 189215 0 FreeSans 560 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -400 167548 240 167604 0 FreeSans 560 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -400 145937 240 145993 0 FreeSans 560 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 291760 3727 292400 3783 0 FreeSans 560 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -400 124426 240 124482 0 FreeSans 560 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -400 60615 240 60671 0 FreeSans 560 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -400 39004 240 39060 0 FreeSans 560 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -400 17393 240 17449 0 FreeSans 560 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -400 6682 240 6738 0 FreeSans 560 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -400 4318 240 4374 0 FreeSans 560 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -400 1954 240 2010 0 FreeSans 560 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 291760 6091 292400 6147 0 FreeSans 560 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 291760 8455 292400 8511 0 FreeSans 560 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 291760 10819 292400 10875 0 FreeSans 560 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 291760 24048 292400 24104 0 FreeSans 560 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 291760 46377 292400 46433 0 FreeSans 560 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 291760 136388 292400 136444 0 FreeSans 560 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 291760 158599 292400 158655 0 FreeSans 560 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 291760 181210 292400 181266 0 FreeSans 560 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 291760 772 292400 828 0 FreeSans 560 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 291760 203830 292400 203886 0 FreeSans 560 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 291760 226041 292400 226097 0 FreeSans 560 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 291760 248252 292400 248308 0 FreeSans 560 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 291760 292963 292400 293019 0 FreeSans 560 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -400 254583 240 254639 0 FreeSans 560 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -400 232972 240 233028 0 FreeSans 560 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -400 211361 240 211417 0 FreeSans 560 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -400 189750 240 189806 0 FreeSans 560 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -400 168139 240 168195 0 FreeSans 560 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -400 146528 240 146584 0 FreeSans 560 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 291760 3136 292400 3192 0 FreeSans 560 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -400 125017 240 125073 0 FreeSans 560 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -400 61206 240 61262 0 FreeSans 560 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -400 39595 240 39651 0 FreeSans 560 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -400 17984 240 18040 0 FreeSans 560 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -400 7273 240 7329 0 FreeSans 560 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -400 4909 240 4965 0 FreeSans 560 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -400 2545 240 2601 0 FreeSans 560 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 291760 5500 292400 5556 0 FreeSans 560 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 291760 7864 292400 7920 0 FreeSans 560 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 291760 10228 292400 10284 0 FreeSans 560 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 291760 23457 292400 23513 0 FreeSans 560 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 291760 45786 292400 45842 0 FreeSans 560 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 291760 135797 292400 135853 0 FreeSans 560 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 291760 158008 292400 158064 0 FreeSans 560 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 291760 180619 292400 180675 0 FreeSans 560 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 291760 2545 292400 2601 0 FreeSans 560 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 291760 205603 292400 205659 0 FreeSans 560 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 291760 227814 292400 227870 0 FreeSans 560 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 291760 250025 292400 250081 0 FreeSans 560 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 291760 294736 292400 294792 0 FreeSans 560 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -400 252810 240 252866 0 FreeSans 560 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -400 231199 240 231255 0 FreeSans 560 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -400 209588 240 209644 0 FreeSans 560 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -400 187977 240 188033 0 FreeSans 560 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -400 166366 240 166422 0 FreeSans 560 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -400 144755 240 144811 0 FreeSans 560 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 291760 4909 292400 4965 0 FreeSans 560 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -400 123244 240 123300 0 FreeSans 560 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -400 59433 240 59489 0 FreeSans 560 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -400 37822 240 37878 0 FreeSans 560 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -400 16211 240 16267 0 FreeSans 560 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -400 5500 240 5556 0 FreeSans 560 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -400 3136 240 3192 0 FreeSans 560 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -400 772 240 828 0 FreeSans 560 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 291760 7273 292400 7329 0 FreeSans 560 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 291760 9637 292400 9693 0 FreeSans 560 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 291760 12001 292400 12057 0 FreeSans 560 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 291760 25230 292400 25286 0 FreeSans 560 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 291760 47559 292400 47615 0 FreeSans 560 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 291760 137570 292400 137626 0 FreeSans 560 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 291760 159781 292400 159837 0 FreeSans 560 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 291760 182392 292400 182448 0 FreeSans 560 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 291760 1954 292400 2010 0 FreeSans 560 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 291760 205012 292400 205068 0 FreeSans 560 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 291760 227223 292400 227279 0 FreeSans 560 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 291760 249434 292400 249490 0 FreeSans 560 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 291760 294145 292400 294201 0 FreeSans 560 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -400 253401 240 253457 0 FreeSans 560 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -400 231790 240 231846 0 FreeSans 560 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -400 210179 240 210235 0 FreeSans 560 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -400 188568 240 188624 0 FreeSans 560 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -400 166957 240 167013 0 FreeSans 560 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -400 145346 240 145402 0 FreeSans 560 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 291760 4318 292400 4374 0 FreeSans 560 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -400 123835 240 123891 0 FreeSans 560 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -400 60024 240 60080 0 FreeSans 560 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -400 38413 240 38469 0 FreeSans 560 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -400 16802 240 16858 0 FreeSans 560 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -400 6091 240 6147 0 FreeSans 560 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -400 3727 240 3783 0 FreeSans 560 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -400 1363 240 1419 0 FreeSans 560 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 291760 6682 292400 6738 0 FreeSans 560 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 291760 9046 292400 9102 0 FreeSans 560 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 291760 11410 292400 11466 0 FreeSans 560 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 291760 24639 292400 24695 0 FreeSans 560 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 291760 46968 292400 47024 0 FreeSans 560 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 291760 136979 292400 137035 0 FreeSans 560 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 291760 159190 292400 159246 0 FreeSans 560 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 291760 181801 292400 181857 0 FreeSans 560 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 62908 -400 62964 240 0 FreeSans 560 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 240208 -400 240264 240 0 FreeSans 560 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 241981 -400 242037 240 0 FreeSans 560 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 243754 -400 243810 240 0 FreeSans 560 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 245527 -400 245583 240 0 FreeSans 560 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 247300 -400 247356 240 0 FreeSans 560 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 249073 -400 249129 240 0 FreeSans 560 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 250846 -400 250902 240 0 FreeSans 560 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 252619 -400 252675 240 0 FreeSans 560 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 254392 -400 254448 240 0 FreeSans 560 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 256165 -400 256221 240 0 FreeSans 560 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 80638 -400 80694 240 0 FreeSans 560 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 257938 -400 257994 240 0 FreeSans 560 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 259711 -400 259767 240 0 FreeSans 560 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 261484 -400 261540 240 0 FreeSans 560 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 263257 -400 263313 240 0 FreeSans 560 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 265030 -400 265086 240 0 FreeSans 560 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 266803 -400 266859 240 0 FreeSans 560 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 268576 -400 268632 240 0 FreeSans 560 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 270349 -400 270405 240 0 FreeSans 560 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 272122 -400 272178 240 0 FreeSans 560 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 273895 -400 273951 240 0 FreeSans 560 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 82411 -400 82467 240 0 FreeSans 560 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 275668 -400 275724 240 0 FreeSans 560 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 277441 -400 277497 240 0 FreeSans 560 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 279214 -400 279270 240 0 FreeSans 560 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 280987 -400 281043 240 0 FreeSans 560 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 282760 -400 282816 240 0 FreeSans 560 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 284533 -400 284589 240 0 FreeSans 560 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 286306 -400 286362 240 0 FreeSans 560 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 288079 -400 288135 240 0 FreeSans 560 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 84184 -400 84240 240 0 FreeSans 560 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 85957 -400 86013 240 0 FreeSans 560 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 87730 -400 87786 240 0 FreeSans 560 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 89503 -400 89559 240 0 FreeSans 560 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 91276 -400 91332 240 0 FreeSans 560 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 93049 -400 93105 240 0 FreeSans 560 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 94822 -400 94878 240 0 FreeSans 560 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 96595 -400 96651 240 0 FreeSans 560 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 64681 -400 64737 240 0 FreeSans 560 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 98368 -400 98424 240 0 FreeSans 560 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 100141 -400 100197 240 0 FreeSans 560 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 101914 -400 101970 240 0 FreeSans 560 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 103687 -400 103743 240 0 FreeSans 560 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 105460 -400 105516 240 0 FreeSans 560 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 107233 -400 107289 240 0 FreeSans 560 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 109006 -400 109062 240 0 FreeSans 560 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 110779 -400 110835 240 0 FreeSans 560 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 112552 -400 112608 240 0 FreeSans 560 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 114325 -400 114381 240 0 FreeSans 560 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 66454 -400 66510 240 0 FreeSans 560 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 116098 -400 116154 240 0 FreeSans 560 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 117871 -400 117927 240 0 FreeSans 560 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 119644 -400 119700 240 0 FreeSans 560 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 121417 -400 121473 240 0 FreeSans 560 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 123190 -400 123246 240 0 FreeSans 560 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 124963 -400 125019 240 0 FreeSans 560 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 126736 -400 126792 240 0 FreeSans 560 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 128509 -400 128565 240 0 FreeSans 560 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 130282 -400 130338 240 0 FreeSans 560 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 132055 -400 132111 240 0 FreeSans 560 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 68227 -400 68283 240 0 FreeSans 560 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 133828 -400 133884 240 0 FreeSans 560 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 135601 -400 135657 240 0 FreeSans 560 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 137374 -400 137430 240 0 FreeSans 560 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 139147 -400 139203 240 0 FreeSans 560 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 140920 -400 140976 240 0 FreeSans 560 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 142693 -400 142749 240 0 FreeSans 560 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 144466 -400 144522 240 0 FreeSans 560 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 146239 -400 146295 240 0 FreeSans 560 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 148012 -400 148068 240 0 FreeSans 560 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 149785 -400 149841 240 0 FreeSans 560 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 70000 -400 70056 240 0 FreeSans 560 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 151558 -400 151614 240 0 FreeSans 560 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 153331 -400 153387 240 0 FreeSans 560 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 155104 -400 155160 240 0 FreeSans 560 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 156877 -400 156933 240 0 FreeSans 560 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 158650 -400 158706 240 0 FreeSans 560 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 160423 -400 160479 240 0 FreeSans 560 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 162196 -400 162252 240 0 FreeSans 560 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 163969 -400 164025 240 0 FreeSans 560 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 165742 -400 165798 240 0 FreeSans 560 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 167515 -400 167571 240 0 FreeSans 560 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 71773 -400 71829 240 0 FreeSans 560 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 169288 -400 169344 240 0 FreeSans 560 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 171061 -400 171117 240 0 FreeSans 560 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 172834 -400 172890 240 0 FreeSans 560 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 174607 -400 174663 240 0 FreeSans 560 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 176380 -400 176436 240 0 FreeSans 560 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 178153 -400 178209 240 0 FreeSans 560 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 179926 -400 179982 240 0 FreeSans 560 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 181699 -400 181755 240 0 FreeSans 560 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 183472 -400 183528 240 0 FreeSans 560 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 185245 -400 185301 240 0 FreeSans 560 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 73546 -400 73602 240 0 FreeSans 560 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 187018 -400 187074 240 0 FreeSans 560 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 188791 -400 188847 240 0 FreeSans 560 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 190564 -400 190620 240 0 FreeSans 560 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 192337 -400 192393 240 0 FreeSans 560 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 194110 -400 194166 240 0 FreeSans 560 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 195883 -400 195939 240 0 FreeSans 560 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 197656 -400 197712 240 0 FreeSans 560 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 199429 -400 199485 240 0 FreeSans 560 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 201202 -400 201258 240 0 FreeSans 560 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 202975 -400 203031 240 0 FreeSans 560 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 75319 -400 75375 240 0 FreeSans 560 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 204748 -400 204804 240 0 FreeSans 560 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 206521 -400 206577 240 0 FreeSans 560 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 208294 -400 208350 240 0 FreeSans 560 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 210067 -400 210123 240 0 FreeSans 560 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 211840 -400 211896 240 0 FreeSans 560 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 213613 -400 213669 240 0 FreeSans 560 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 215386 -400 215442 240 0 FreeSans 560 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 217159 -400 217215 240 0 FreeSans 560 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 218932 -400 218988 240 0 FreeSans 560 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 220705 -400 220761 240 0 FreeSans 560 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 77092 -400 77148 240 0 FreeSans 560 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 222478 -400 222534 240 0 FreeSans 560 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 224251 -400 224307 240 0 FreeSans 560 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 226024 -400 226080 240 0 FreeSans 560 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 227797 -400 227853 240 0 FreeSans 560 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 229570 -400 229626 240 0 FreeSans 560 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 231343 -400 231399 240 0 FreeSans 560 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 233116 -400 233172 240 0 FreeSans 560 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 234889 -400 234945 240 0 FreeSans 560 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 236662 -400 236718 240 0 FreeSans 560 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 238435 -400 238491 240 0 FreeSans 560 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 78865 -400 78921 240 0 FreeSans 560 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 63499 -400 63555 240 0 FreeSans 560 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 240799 -400 240855 240 0 FreeSans 560 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 242572 -400 242628 240 0 FreeSans 560 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 244345 -400 244401 240 0 FreeSans 560 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 246118 -400 246174 240 0 FreeSans 560 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 247891 -400 247947 240 0 FreeSans 560 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 249664 -400 249720 240 0 FreeSans 560 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 251437 -400 251493 240 0 FreeSans 560 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 253210 -400 253266 240 0 FreeSans 560 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 254983 -400 255039 240 0 FreeSans 560 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 256756 -400 256812 240 0 FreeSans 560 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 81229 -400 81285 240 0 FreeSans 560 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 258529 -400 258585 240 0 FreeSans 560 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 260302 -400 260358 240 0 FreeSans 560 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 262075 -400 262131 240 0 FreeSans 560 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 263848 -400 263904 240 0 FreeSans 560 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 265621 -400 265677 240 0 FreeSans 560 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 267394 -400 267450 240 0 FreeSans 560 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 269167 -400 269223 240 0 FreeSans 560 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 270940 -400 270996 240 0 FreeSans 560 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 272713 -400 272769 240 0 FreeSans 560 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 274486 -400 274542 240 0 FreeSans 560 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 83002 -400 83058 240 0 FreeSans 560 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 276259 -400 276315 240 0 FreeSans 560 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 278032 -400 278088 240 0 FreeSans 560 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 279805 -400 279861 240 0 FreeSans 560 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 281578 -400 281634 240 0 FreeSans 560 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 283351 -400 283407 240 0 FreeSans 560 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 285124 -400 285180 240 0 FreeSans 560 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 286897 -400 286953 240 0 FreeSans 560 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 288670 -400 288726 240 0 FreeSans 560 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 84775 -400 84831 240 0 FreeSans 560 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 86548 -400 86604 240 0 FreeSans 560 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 88321 -400 88377 240 0 FreeSans 560 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 90094 -400 90150 240 0 FreeSans 560 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 91867 -400 91923 240 0 FreeSans 560 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 93640 -400 93696 240 0 FreeSans 560 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 95413 -400 95469 240 0 FreeSans 560 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 97186 -400 97242 240 0 FreeSans 560 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 65272 -400 65328 240 0 FreeSans 560 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 98959 -400 99015 240 0 FreeSans 560 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 100732 -400 100788 240 0 FreeSans 560 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 102505 -400 102561 240 0 FreeSans 560 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 104278 -400 104334 240 0 FreeSans 560 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 106051 -400 106107 240 0 FreeSans 560 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 107824 -400 107880 240 0 FreeSans 560 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 109597 -400 109653 240 0 FreeSans 560 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 111370 -400 111426 240 0 FreeSans 560 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 113143 -400 113199 240 0 FreeSans 560 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 114916 -400 114972 240 0 FreeSans 560 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 67045 -400 67101 240 0 FreeSans 560 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 116689 -400 116745 240 0 FreeSans 560 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 118462 -400 118518 240 0 FreeSans 560 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 120235 -400 120291 240 0 FreeSans 560 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 122008 -400 122064 240 0 FreeSans 560 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 123781 -400 123837 240 0 FreeSans 560 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 125554 -400 125610 240 0 FreeSans 560 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 127327 -400 127383 240 0 FreeSans 560 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 129100 -400 129156 240 0 FreeSans 560 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 130873 -400 130929 240 0 FreeSans 560 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 132646 -400 132702 240 0 FreeSans 560 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 68818 -400 68874 240 0 FreeSans 560 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 134419 -400 134475 240 0 FreeSans 560 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 136192 -400 136248 240 0 FreeSans 560 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 137965 -400 138021 240 0 FreeSans 560 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 139738 -400 139794 240 0 FreeSans 560 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 141511 -400 141567 240 0 FreeSans 560 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 143284 -400 143340 240 0 FreeSans 560 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 145057 -400 145113 240 0 FreeSans 560 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 146830 -400 146886 240 0 FreeSans 560 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 148603 -400 148659 240 0 FreeSans 560 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 150376 -400 150432 240 0 FreeSans 560 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 70591 -400 70647 240 0 FreeSans 560 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 152149 -400 152205 240 0 FreeSans 560 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 153922 -400 153978 240 0 FreeSans 560 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 155695 -400 155751 240 0 FreeSans 560 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 157468 -400 157524 240 0 FreeSans 560 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 159241 -400 159297 240 0 FreeSans 560 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 161014 -400 161070 240 0 FreeSans 560 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 162787 -400 162843 240 0 FreeSans 560 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 164560 -400 164616 240 0 FreeSans 560 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 166333 -400 166389 240 0 FreeSans 560 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 168106 -400 168162 240 0 FreeSans 560 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 72364 -400 72420 240 0 FreeSans 560 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 169879 -400 169935 240 0 FreeSans 560 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 171652 -400 171708 240 0 FreeSans 560 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 173425 -400 173481 240 0 FreeSans 560 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 175198 -400 175254 240 0 FreeSans 560 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 176971 -400 177027 240 0 FreeSans 560 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 178744 -400 178800 240 0 FreeSans 560 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 180517 -400 180573 240 0 FreeSans 560 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 182290 -400 182346 240 0 FreeSans 560 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 184063 -400 184119 240 0 FreeSans 560 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 185836 -400 185892 240 0 FreeSans 560 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 74137 -400 74193 240 0 FreeSans 560 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 187609 -400 187665 240 0 FreeSans 560 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 189382 -400 189438 240 0 FreeSans 560 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 191155 -400 191211 240 0 FreeSans 560 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 192928 -400 192984 240 0 FreeSans 560 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 194701 -400 194757 240 0 FreeSans 560 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 196474 -400 196530 240 0 FreeSans 560 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 198247 -400 198303 240 0 FreeSans 560 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 200020 -400 200076 240 0 FreeSans 560 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 201793 -400 201849 240 0 FreeSans 560 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 203566 -400 203622 240 0 FreeSans 560 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 75910 -400 75966 240 0 FreeSans 560 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 205339 -400 205395 240 0 FreeSans 560 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 207112 -400 207168 240 0 FreeSans 560 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 208885 -400 208941 240 0 FreeSans 560 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 210658 -400 210714 240 0 FreeSans 560 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 212431 -400 212487 240 0 FreeSans 560 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 214204 -400 214260 240 0 FreeSans 560 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 215977 -400 216033 240 0 FreeSans 560 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 217750 -400 217806 240 0 FreeSans 560 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 219523 -400 219579 240 0 FreeSans 560 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 221296 -400 221352 240 0 FreeSans 560 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 77683 -400 77739 240 0 FreeSans 560 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 223069 -400 223125 240 0 FreeSans 560 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 224842 -400 224898 240 0 FreeSans 560 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 226615 -400 226671 240 0 FreeSans 560 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 228388 -400 228444 240 0 FreeSans 560 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 230161 -400 230217 240 0 FreeSans 560 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 231934 -400 231990 240 0 FreeSans 560 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 233707 -400 233763 240 0 FreeSans 560 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 235480 -400 235536 240 0 FreeSans 560 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 237253 -400 237309 240 0 FreeSans 560 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 239026 -400 239082 240 0 FreeSans 560 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 79456 -400 79512 240 0 FreeSans 560 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 64090 -400 64146 240 0 FreeSans 560 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 241390 -400 241446 240 0 FreeSans 560 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 243163 -400 243219 240 0 FreeSans 560 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 244936 -400 244992 240 0 FreeSans 560 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 246709 -400 246765 240 0 FreeSans 560 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 248482 -400 248538 240 0 FreeSans 560 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 250255 -400 250311 240 0 FreeSans 560 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 252028 -400 252084 240 0 FreeSans 560 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 253801 -400 253857 240 0 FreeSans 560 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 255574 -400 255630 240 0 FreeSans 560 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 257347 -400 257403 240 0 FreeSans 560 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 81820 -400 81876 240 0 FreeSans 560 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 259120 -400 259176 240 0 FreeSans 560 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 260893 -400 260949 240 0 FreeSans 560 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 262666 -400 262722 240 0 FreeSans 560 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 264439 -400 264495 240 0 FreeSans 560 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 266212 -400 266268 240 0 FreeSans 560 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 267985 -400 268041 240 0 FreeSans 560 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 269758 -400 269814 240 0 FreeSans 560 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 271531 -400 271587 240 0 FreeSans 560 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 273304 -400 273360 240 0 FreeSans 560 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 275077 -400 275133 240 0 FreeSans 560 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 83593 -400 83649 240 0 FreeSans 560 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 276850 -400 276906 240 0 FreeSans 560 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 278623 -400 278679 240 0 FreeSans 560 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 280396 -400 280452 240 0 FreeSans 560 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 282169 -400 282225 240 0 FreeSans 560 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 283942 -400 283998 240 0 FreeSans 560 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 285715 -400 285771 240 0 FreeSans 560 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 287488 -400 287544 240 0 FreeSans 560 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 289261 -400 289317 240 0 FreeSans 560 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 85366 -400 85422 240 0 FreeSans 560 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 87139 -400 87195 240 0 FreeSans 560 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 88912 -400 88968 240 0 FreeSans 560 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 90685 -400 90741 240 0 FreeSans 560 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 92458 -400 92514 240 0 FreeSans 560 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 94231 -400 94287 240 0 FreeSans 560 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 96004 -400 96060 240 0 FreeSans 560 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 97777 -400 97833 240 0 FreeSans 560 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 65863 -400 65919 240 0 FreeSans 560 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 99550 -400 99606 240 0 FreeSans 560 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 101323 -400 101379 240 0 FreeSans 560 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 103096 -400 103152 240 0 FreeSans 560 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 104869 -400 104925 240 0 FreeSans 560 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 106642 -400 106698 240 0 FreeSans 560 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 108415 -400 108471 240 0 FreeSans 560 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 110188 -400 110244 240 0 FreeSans 560 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 111961 -400 112017 240 0 FreeSans 560 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 113734 -400 113790 240 0 FreeSans 560 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 115507 -400 115563 240 0 FreeSans 560 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 67636 -400 67692 240 0 FreeSans 560 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 117280 -400 117336 240 0 FreeSans 560 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 119053 -400 119109 240 0 FreeSans 560 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 120826 -400 120882 240 0 FreeSans 560 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 122599 -400 122655 240 0 FreeSans 560 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 124372 -400 124428 240 0 FreeSans 560 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 126145 -400 126201 240 0 FreeSans 560 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 127918 -400 127974 240 0 FreeSans 560 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 129691 -400 129747 240 0 FreeSans 560 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 131464 -400 131520 240 0 FreeSans 560 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 133237 -400 133293 240 0 FreeSans 560 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 69409 -400 69465 240 0 FreeSans 560 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 135010 -400 135066 240 0 FreeSans 560 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 136783 -400 136839 240 0 FreeSans 560 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 138556 -400 138612 240 0 FreeSans 560 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 140329 -400 140385 240 0 FreeSans 560 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 142102 -400 142158 240 0 FreeSans 560 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 143875 -400 143931 240 0 FreeSans 560 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 145648 -400 145704 240 0 FreeSans 560 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 147421 -400 147477 240 0 FreeSans 560 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 149194 -400 149250 240 0 FreeSans 560 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 150967 -400 151023 240 0 FreeSans 560 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 71182 -400 71238 240 0 FreeSans 560 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 152740 -400 152796 240 0 FreeSans 560 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 154513 -400 154569 240 0 FreeSans 560 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 156286 -400 156342 240 0 FreeSans 560 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 158059 -400 158115 240 0 FreeSans 560 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 159832 -400 159888 240 0 FreeSans 560 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 161605 -400 161661 240 0 FreeSans 560 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 163378 -400 163434 240 0 FreeSans 560 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 165151 -400 165207 240 0 FreeSans 560 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 166924 -400 166980 240 0 FreeSans 560 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 168697 -400 168753 240 0 FreeSans 560 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 72955 -400 73011 240 0 FreeSans 560 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 170470 -400 170526 240 0 FreeSans 560 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 172243 -400 172299 240 0 FreeSans 560 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 174016 -400 174072 240 0 FreeSans 560 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 175789 -400 175845 240 0 FreeSans 560 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 177562 -400 177618 240 0 FreeSans 560 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 179335 -400 179391 240 0 FreeSans 560 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 181108 -400 181164 240 0 FreeSans 560 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 182881 -400 182937 240 0 FreeSans 560 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 184654 -400 184710 240 0 FreeSans 560 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 186427 -400 186483 240 0 FreeSans 560 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 74728 -400 74784 240 0 FreeSans 560 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 188200 -400 188256 240 0 FreeSans 560 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 189973 -400 190029 240 0 FreeSans 560 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 191746 -400 191802 240 0 FreeSans 560 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 193519 -400 193575 240 0 FreeSans 560 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 195292 -400 195348 240 0 FreeSans 560 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 197065 -400 197121 240 0 FreeSans 560 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 198838 -400 198894 240 0 FreeSans 560 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 200611 -400 200667 240 0 FreeSans 560 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 202384 -400 202440 240 0 FreeSans 560 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 204157 -400 204213 240 0 FreeSans 560 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 76501 -400 76557 240 0 FreeSans 560 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 205930 -400 205986 240 0 FreeSans 560 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 207703 -400 207759 240 0 FreeSans 560 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 209476 -400 209532 240 0 FreeSans 560 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 211249 -400 211305 240 0 FreeSans 560 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 213022 -400 213078 240 0 FreeSans 560 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 214795 -400 214851 240 0 FreeSans 560 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 216568 -400 216624 240 0 FreeSans 560 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 218341 -400 218397 240 0 FreeSans 560 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 220114 -400 220170 240 0 FreeSans 560 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 221887 -400 221943 240 0 FreeSans 560 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 78274 -400 78330 240 0 FreeSans 560 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 223660 -400 223716 240 0 FreeSans 560 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 225433 -400 225489 240 0 FreeSans 560 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 227206 -400 227262 240 0 FreeSans 560 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 228979 -400 229035 240 0 FreeSans 560 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 230752 -400 230808 240 0 FreeSans 560 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 232525 -400 232581 240 0 FreeSans 560 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 234298 -400 234354 240 0 FreeSans 560 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 236071 -400 236127 240 0 FreeSans 560 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 237844 -400 237900 240 0 FreeSans 560 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 239617 -400 239673 240 0 FreeSans 560 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 80047 -400 80103 240 0 FreeSans 560 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 289852 -400 289908 240 0 FreeSans 560 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 290443 -400 290499 240 0 FreeSans 560 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 291034 -400 291090 240 0 FreeSans 560 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 291625 -400 291681 240 0 FreeSans 560 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 291170 319892 292400 322292 0 FreeSans 560 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 291170 314892 292400 317292 0 FreeSans 560 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 321921 830 324321 0 FreeSans 560 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 316921 830 319321 0 FreeSans 560 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 291170 270281 292400 272681 0 FreeSans 560 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 291170 275281 292400 277681 0 FreeSans 560 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 291170 117615 292400 120015 0 FreeSans 560 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 291170 112615 292400 115015 0 FreeSans 560 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 102444 830 104844 0 FreeSans 560 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 107444 830 109844 0 FreeSans 560 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 260297 351170 262697 352400 0 FreeSans 960 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 255297 351170 257697 352400 0 FreeSans 960 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 291170 73415 292400 75815 0 FreeSans 560 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 291170 68415 292400 70815 0 FreeSans 560 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 279721 830 282121 0 FreeSans 560 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 274721 830 277121 0 FreeSans 560 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 291170 95715 292400 98115 0 FreeSans 560 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 291170 90715 292400 93115 0 FreeSans 560 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 86444 830 88844 0 FreeSans 560 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 81444 830 83844 0 FreeSans 560 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 262 -400 318 240 0 FreeSans 560 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 853 -400 909 240 0 FreeSans 560 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 1444 -400 1500 240 0 FreeSans 560 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 3808 -400 3864 240 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 23902 -400 23958 240 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 25675 -400 25731 240 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 27448 -400 27504 240 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 29221 -400 29277 240 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 30994 -400 31050 240 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 32767 -400 32823 240 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 34540 -400 34596 240 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 36313 -400 36369 240 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 38086 -400 38142 240 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 39859 -400 39915 240 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 6172 -400 6228 240 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 41632 -400 41688 240 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 43405 -400 43461 240 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 45178 -400 45234 240 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 46951 -400 47007 240 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 48724 -400 48780 240 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 50497 -400 50553 240 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 52270 -400 52326 240 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 54043 -400 54099 240 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 55816 -400 55872 240 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 57589 -400 57645 240 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 8536 -400 8592 240 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 59362 -400 59418 240 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 61135 -400 61191 240 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 10900 -400 10956 240 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 13264 -400 13320 240 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 15037 -400 15093 240 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 16810 -400 16866 240 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 18583 -400 18639 240 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 20356 -400 20412 240 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 22129 -400 22185 240 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 2035 -400 2091 240 0 FreeSans 560 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 4399 -400 4455 240 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 24493 -400 24549 240 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 26266 -400 26322 240 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 28039 -400 28095 240 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 29812 -400 29868 240 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 31585 -400 31641 240 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 33358 -400 33414 240 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 35131 -400 35187 240 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 36904 -400 36960 240 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 38677 -400 38733 240 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 40450 -400 40506 240 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 6763 -400 6819 240 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 42223 -400 42279 240 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 43996 -400 44052 240 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 45769 -400 45825 240 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 47542 -400 47598 240 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 49315 -400 49371 240 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 51088 -400 51144 240 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 52861 -400 52917 240 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 54634 -400 54690 240 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 56407 -400 56463 240 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 58180 -400 58236 240 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 9127 -400 9183 240 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 59953 -400 60009 240 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 61726 -400 61782 240 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 11491 -400 11547 240 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 13855 -400 13911 240 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 15628 -400 15684 240 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 17401 -400 17457 240 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 19174 -400 19230 240 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 20947 -400 21003 240 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 22720 -400 22776 240 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 4990 -400 5046 240 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 25084 -400 25140 240 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 26857 -400 26913 240 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 28630 -400 28686 240 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 30403 -400 30459 240 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 32176 -400 32232 240 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 33949 -400 34005 240 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 35722 -400 35778 240 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 37495 -400 37551 240 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 39268 -400 39324 240 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 41041 -400 41097 240 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 7354 -400 7410 240 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 42814 -400 42870 240 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 44587 -400 44643 240 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 46360 -400 46416 240 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 48133 -400 48189 240 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 49906 -400 49962 240 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 51679 -400 51735 240 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 53452 -400 53508 240 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 55225 -400 55281 240 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 56998 -400 57054 240 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 58771 -400 58827 240 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 9718 -400 9774 240 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 60544 -400 60600 240 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 62317 -400 62373 240 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 12082 -400 12138 240 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 14446 -400 14502 240 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 16219 -400 16275 240 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 17992 -400 18048 240 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 19765 -400 19821 240 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 21538 -400 21594 240 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 23311 -400 23367 240 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 5581 -400 5637 240 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 7945 -400 8001 240 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 10309 -400 10365 240 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 12673 -400 12729 240 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 2626 -400 2682 240 0 FreeSans 560 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 3217 -400 3273 240 0 FreeSans 560 90 0 0 wbs_we_i
port 677 nsew signal input
rlabel metal3 28640 274920 28680 274960 1 ii
rlabel metal3 28640 275360 28680 275400 1 ii
rlabel metal3 28480 275360 28520 275400 1 vi
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
