magic
tech sky130A
timestamp 1640820182
<< nwell >>
rect -680 4800 4720 5480
rect -680 2880 4720 3560
rect -680 960 4720 1640
<< mvnmos >>
rect -480 3840 -280 3940
rect 0 3840 200 3940
rect 320 3840 520 3940
rect 640 3840 840 3940
rect 960 3840 1160 3940
rect 1440 3840 1640 3940
rect 1760 3840 1960 3940
rect 2080 3840 2280 3940
rect 2400 3840 2600 3940
rect 2880 3840 3080 3940
rect 3200 3840 3400 3940
rect 3520 3840 3720 3940
rect 3840 3840 4040 3940
rect 4320 3840 4520 3940
rect -480 1920 -280 2020
rect 0 1920 200 2020
rect 320 1920 520 2020
rect 640 1920 840 2020
rect 960 1920 1160 2020
rect 1440 1920 1640 2020
rect 1760 1920 1960 2020
rect 2080 1920 2280 2020
rect 2400 1920 2600 2020
rect 2880 1920 3080 2020
rect 3200 1920 3400 2020
rect 3520 1920 3720 2020
rect 3840 1920 4040 2020
rect 4320 1920 4520 2020
rect -480 0 -280 100
rect 0 0 200 100
rect 320 0 520 100
rect 640 0 840 100
rect 960 0 1160 100
rect 1440 0 1640 100
rect 1760 0 1960 100
rect 2080 0 2280 100
rect 2400 0 2600 100
rect 2880 0 3080 100
rect 3200 0 3400 100
rect 3520 0 3720 100
rect 3840 0 4040 100
rect 4320 0 4520 100
<< mvpmos >>
rect -480 5200 -280 5300
rect -480 4980 -280 5080
rect 0 5200 200 5300
rect 320 5200 520 5300
rect 640 5200 840 5300
rect 960 5200 1160 5300
rect 0 4980 200 5080
rect 320 4980 520 5080
rect 640 4980 840 5080
rect 960 4980 1160 5080
rect 1440 5200 1640 5300
rect 1760 5200 1960 5300
rect 2080 5200 2280 5300
rect 2400 5200 2600 5300
rect 1440 4980 1640 5080
rect 1760 4980 1960 5080
rect 2080 4980 2280 5080
rect 2400 4980 2600 5080
rect 2880 5200 3080 5300
rect 3200 5200 3400 5300
rect 3520 5200 3720 5300
rect 3840 5200 4040 5300
rect 2880 4980 3080 5080
rect 3200 4980 3400 5080
rect 3520 4980 3720 5080
rect 3840 4980 4040 5080
rect 4320 5200 4520 5300
rect 4320 4980 4520 5080
rect -480 3280 -280 3380
rect -480 3060 -280 3160
rect 0 3280 200 3380
rect 320 3280 520 3380
rect 640 3280 840 3380
rect 960 3280 1160 3380
rect 0 3060 200 3160
rect 320 3060 520 3160
rect 640 3060 840 3160
rect 960 3060 1160 3160
rect 1440 3280 1640 3380
rect 1760 3280 1960 3380
rect 2080 3280 2280 3380
rect 2400 3280 2600 3380
rect 1440 3060 1640 3160
rect 1760 3060 1960 3160
rect 2080 3060 2280 3160
rect 2400 3060 2600 3160
rect 2880 3280 3080 3380
rect 3200 3280 3400 3380
rect 3520 3280 3720 3380
rect 3840 3280 4040 3380
rect 2880 3060 3080 3160
rect 3200 3060 3400 3160
rect 3520 3060 3720 3160
rect 3840 3060 4040 3160
rect 4320 3280 4520 3380
rect 4320 3060 4520 3160
rect -480 1360 -280 1460
rect -480 1140 -280 1240
rect 0 1360 200 1460
rect 320 1360 520 1460
rect 640 1360 840 1460
rect 960 1360 1160 1460
rect 0 1140 200 1240
rect 320 1140 520 1240
rect 640 1140 840 1240
rect 960 1140 1160 1240
rect 1440 1360 1640 1460
rect 1760 1360 1960 1460
rect 2080 1360 2280 1460
rect 2400 1360 2600 1460
rect 1440 1140 1640 1240
rect 1760 1140 1960 1240
rect 2080 1140 2280 1240
rect 2400 1140 2600 1240
rect 2880 1360 3080 1460
rect 3200 1360 3400 1460
rect 3520 1360 3720 1460
rect 3840 1360 4040 1460
rect 2880 1140 3080 1240
rect 3200 1140 3400 1240
rect 3520 1140 3720 1240
rect 3840 1140 4040 1240
rect 4320 1360 4520 1460
rect 4320 1140 4520 1240
<< mvndiff >>
rect -560 3930 -480 3940
rect -560 3850 -555 3930
rect -525 3850 -480 3930
rect -560 3840 -480 3850
rect -280 3930 -200 3940
rect -280 3850 -235 3930
rect -205 3850 -200 3930
rect -280 3840 -200 3850
rect -80 3930 0 3940
rect -80 3850 -75 3930
rect -45 3850 0 3930
rect -80 3840 0 3850
rect 200 3930 320 3940
rect 200 3850 245 3930
rect 275 3850 320 3930
rect 200 3840 320 3850
rect 520 3930 640 3940
rect 520 3850 565 3930
rect 595 3850 640 3930
rect 520 3840 640 3850
rect 840 3930 960 3940
rect 840 3850 885 3930
rect 915 3850 960 3930
rect 840 3840 960 3850
rect 1160 3930 1240 3940
rect 1160 3850 1205 3930
rect 1235 3850 1240 3930
rect 1160 3840 1240 3850
rect 1360 3930 1440 3940
rect 1360 3850 1365 3930
rect 1395 3850 1440 3930
rect 1360 3840 1440 3850
rect 1640 3930 1760 3940
rect 1640 3850 1685 3930
rect 1715 3850 1760 3930
rect 1640 3840 1760 3850
rect 1960 3930 2080 3940
rect 1960 3850 2005 3930
rect 2035 3850 2080 3930
rect 1960 3840 2080 3850
rect 2280 3930 2400 3940
rect 2280 3850 2325 3930
rect 2355 3850 2400 3930
rect 2280 3840 2400 3850
rect 2600 3930 2680 3940
rect 2600 3850 2645 3930
rect 2675 3850 2680 3930
rect 2600 3840 2680 3850
rect 2800 3930 2880 3940
rect 2800 3850 2805 3930
rect 2835 3850 2880 3930
rect 2800 3840 2880 3850
rect 3080 3930 3200 3940
rect 3080 3850 3125 3930
rect 3155 3850 3200 3930
rect 3080 3840 3200 3850
rect 3400 3930 3520 3940
rect 3400 3850 3445 3930
rect 3475 3850 3520 3930
rect 3400 3840 3520 3850
rect 3720 3930 3840 3940
rect 3720 3850 3765 3930
rect 3795 3850 3840 3930
rect 3720 3840 3840 3850
rect 4040 3930 4120 3940
rect 4040 3850 4085 3930
rect 4115 3850 4120 3930
rect 4040 3840 4120 3850
rect 4240 3930 4320 3940
rect 4240 3850 4245 3930
rect 4275 3850 4320 3930
rect 4240 3840 4320 3850
rect 4520 3930 4600 3940
rect 4520 3850 4565 3930
rect 4595 3850 4600 3930
rect 4520 3840 4600 3850
rect -560 2010 -480 2020
rect -560 1930 -555 2010
rect -525 1930 -480 2010
rect -560 1920 -480 1930
rect -280 2010 -200 2020
rect -280 1930 -235 2010
rect -205 1930 -200 2010
rect -280 1920 -200 1930
rect -80 2010 0 2020
rect -80 1930 -75 2010
rect -45 1930 0 2010
rect -80 1920 0 1930
rect 200 2010 320 2020
rect 200 1930 245 2010
rect 275 1930 320 2010
rect 200 1920 320 1930
rect 520 2010 640 2020
rect 520 1930 565 2010
rect 595 1930 640 2010
rect 520 1920 640 1930
rect 840 2010 960 2020
rect 840 1930 885 2010
rect 915 1930 960 2010
rect 840 1920 960 1930
rect 1160 2010 1240 2020
rect 1160 1930 1205 2010
rect 1235 1930 1240 2010
rect 1160 1920 1240 1930
rect 1360 2010 1440 2020
rect 1360 1930 1365 2010
rect 1395 1930 1440 2010
rect 1360 1920 1440 1930
rect 1640 2010 1760 2020
rect 1640 1930 1685 2010
rect 1715 1930 1760 2010
rect 1640 1920 1760 1930
rect 1960 2010 2080 2020
rect 1960 1930 2005 2010
rect 2035 1930 2080 2010
rect 1960 1920 2080 1930
rect 2280 2010 2400 2020
rect 2280 1930 2325 2010
rect 2355 1930 2400 2010
rect 2280 1920 2400 1930
rect 2600 2010 2680 2020
rect 2600 1930 2645 2010
rect 2675 1930 2680 2010
rect 2600 1920 2680 1930
rect 2800 2010 2880 2020
rect 2800 1930 2805 2010
rect 2835 1930 2880 2010
rect 2800 1920 2880 1930
rect 3080 2010 3200 2020
rect 3080 1930 3125 2010
rect 3155 1930 3200 2010
rect 3080 1920 3200 1930
rect 3400 2010 3520 2020
rect 3400 1930 3445 2010
rect 3475 1930 3520 2010
rect 3400 1920 3520 1930
rect 3720 2010 3840 2020
rect 3720 1930 3765 2010
rect 3795 1930 3840 2010
rect 3720 1920 3840 1930
rect 4040 2010 4120 2020
rect 4040 1930 4085 2010
rect 4115 1930 4120 2010
rect 4040 1920 4120 1930
rect 4240 2010 4320 2020
rect 4240 1930 4245 2010
rect 4275 1930 4320 2010
rect 4240 1920 4320 1930
rect 4520 2010 4600 2020
rect 4520 1930 4565 2010
rect 4595 1930 4600 2010
rect 4520 1920 4600 1930
rect -560 90 -480 100
rect -560 10 -555 90
rect -525 10 -480 90
rect -560 0 -480 10
rect -280 90 -200 100
rect -280 10 -235 90
rect -205 10 -200 90
rect -280 0 -200 10
rect -80 90 0 100
rect -80 10 -75 90
rect -45 10 0 90
rect -80 0 0 10
rect 200 90 320 100
rect 200 10 245 90
rect 275 10 320 90
rect 200 0 320 10
rect 520 90 640 100
rect 520 10 565 90
rect 595 10 640 90
rect 520 0 640 10
rect 840 90 960 100
rect 840 10 885 90
rect 915 10 960 90
rect 840 0 960 10
rect 1160 90 1240 100
rect 1160 10 1205 90
rect 1235 10 1240 90
rect 1160 0 1240 10
rect 1360 90 1440 100
rect 1360 10 1365 90
rect 1395 10 1440 90
rect 1360 0 1440 10
rect 1640 90 1760 100
rect 1640 10 1685 90
rect 1715 10 1760 90
rect 1640 0 1760 10
rect 1960 90 2080 100
rect 1960 10 2005 90
rect 2035 10 2080 90
rect 1960 0 2080 10
rect 2280 90 2400 100
rect 2280 10 2325 90
rect 2355 10 2400 90
rect 2280 0 2400 10
rect 2600 90 2680 100
rect 2600 10 2645 90
rect 2675 10 2680 90
rect 2600 0 2680 10
rect 2800 90 2880 100
rect 2800 10 2805 90
rect 2835 10 2880 90
rect 2800 0 2880 10
rect 3080 90 3200 100
rect 3080 10 3125 90
rect 3155 10 3200 90
rect 3080 0 3200 10
rect 3400 90 3520 100
rect 3400 10 3445 90
rect 3475 10 3520 90
rect 3400 0 3520 10
rect 3720 90 3840 100
rect 3720 10 3765 90
rect 3795 10 3840 90
rect 3720 0 3840 10
rect 4040 90 4120 100
rect 4040 10 4085 90
rect 4115 10 4120 90
rect 4040 0 4120 10
rect 4240 90 4320 100
rect 4240 10 4245 90
rect 4275 10 4320 90
rect 4240 0 4320 10
rect 4520 90 4600 100
rect 4520 10 4565 90
rect 4595 10 4600 90
rect 4520 0 4600 10
<< mvpdiff >>
rect -560 5290 -480 5300
rect -560 5210 -555 5290
rect -525 5210 -480 5290
rect -560 5200 -480 5210
rect -280 5290 -200 5300
rect -280 5210 -235 5290
rect -205 5210 -200 5290
rect -280 5200 -200 5210
rect -560 5070 -480 5080
rect -560 4990 -555 5070
rect -525 4990 -480 5070
rect -560 4980 -480 4990
rect -280 5070 -200 5080
rect -280 4990 -235 5070
rect -205 4990 -200 5070
rect -280 4980 -200 4990
rect -80 5290 0 5300
rect -80 5210 -75 5290
rect -45 5210 0 5290
rect -80 5200 0 5210
rect 200 5290 320 5300
rect 200 5210 245 5290
rect 275 5210 320 5290
rect 200 5200 320 5210
rect 520 5290 640 5300
rect 520 5210 565 5290
rect 595 5210 640 5290
rect 520 5200 640 5210
rect 840 5290 960 5300
rect 840 5210 885 5290
rect 915 5210 960 5290
rect 840 5200 960 5210
rect 1160 5290 1240 5300
rect 1160 5210 1205 5290
rect 1235 5210 1240 5290
rect 1160 5200 1240 5210
rect -80 5070 0 5080
rect -80 4990 -75 5070
rect -45 4990 0 5070
rect -80 4980 0 4990
rect 200 5070 320 5080
rect 200 4990 245 5070
rect 275 4990 320 5070
rect 200 4980 320 4990
rect 520 5070 640 5080
rect 520 4990 565 5070
rect 595 4990 640 5070
rect 520 4980 640 4990
rect 840 5070 960 5080
rect 840 4990 885 5070
rect 915 4990 960 5070
rect 840 4980 960 4990
rect 1160 5070 1240 5080
rect 1160 4990 1205 5070
rect 1235 4990 1240 5070
rect 1160 4980 1240 4990
rect 1360 5290 1440 5300
rect 1360 5210 1365 5290
rect 1395 5210 1440 5290
rect 1360 5200 1440 5210
rect 1640 5290 1760 5300
rect 1640 5210 1685 5290
rect 1715 5210 1760 5290
rect 1640 5200 1760 5210
rect 1960 5290 2080 5300
rect 1960 5210 2005 5290
rect 2035 5210 2080 5290
rect 1960 5200 2080 5210
rect 2280 5290 2400 5300
rect 2280 5210 2325 5290
rect 2355 5210 2400 5290
rect 2280 5200 2400 5210
rect 2600 5290 2680 5300
rect 2600 5210 2645 5290
rect 2675 5210 2680 5290
rect 2600 5200 2680 5210
rect 1360 5070 1440 5080
rect 1360 4990 1365 5070
rect 1395 4990 1440 5070
rect 1360 4980 1440 4990
rect 1640 5070 1760 5080
rect 1640 4990 1685 5070
rect 1715 4990 1760 5070
rect 1640 4980 1760 4990
rect 1960 5070 2080 5080
rect 1960 4990 2005 5070
rect 2035 4990 2080 5070
rect 1960 4980 2080 4990
rect 2280 5070 2400 5080
rect 2280 4990 2325 5070
rect 2355 4990 2400 5070
rect 2280 4980 2400 4990
rect 2600 5070 2680 5080
rect 2600 4990 2645 5070
rect 2675 4990 2680 5070
rect 2600 4980 2680 4990
rect 2800 5290 2880 5300
rect 2800 5210 2805 5290
rect 2835 5210 2880 5290
rect 2800 5200 2880 5210
rect 3080 5290 3200 5300
rect 3080 5210 3125 5290
rect 3155 5210 3200 5290
rect 3080 5200 3200 5210
rect 3400 5290 3520 5300
rect 3400 5210 3445 5290
rect 3475 5210 3520 5290
rect 3400 5200 3520 5210
rect 3720 5290 3840 5300
rect 3720 5210 3765 5290
rect 3795 5210 3840 5290
rect 3720 5200 3840 5210
rect 4040 5290 4120 5300
rect 4040 5210 4085 5290
rect 4115 5210 4120 5290
rect 4040 5200 4120 5210
rect 2800 5070 2880 5080
rect 2800 4990 2805 5070
rect 2835 4990 2880 5070
rect 2800 4980 2880 4990
rect 3080 5070 3200 5080
rect 3080 4990 3125 5070
rect 3155 4990 3200 5070
rect 3080 4980 3200 4990
rect 3400 5070 3520 5080
rect 3400 4990 3445 5070
rect 3475 4990 3520 5070
rect 3400 4980 3520 4990
rect 3720 5070 3840 5080
rect 3720 4990 3765 5070
rect 3795 4990 3840 5070
rect 3720 4980 3840 4990
rect 4040 5070 4120 5080
rect 4040 4990 4085 5070
rect 4115 4990 4120 5070
rect 4040 4980 4120 4990
rect 4240 5290 4320 5300
rect 4240 5210 4245 5290
rect 4275 5210 4320 5290
rect 4240 5200 4320 5210
rect 4520 5290 4600 5300
rect 4520 5210 4565 5290
rect 4595 5210 4600 5290
rect 4520 5200 4600 5210
rect 4240 5070 4320 5080
rect 4240 4990 4245 5070
rect 4275 4990 4320 5070
rect 4240 4980 4320 4990
rect 4520 5070 4600 5080
rect 4520 4990 4565 5070
rect 4595 4990 4600 5070
rect 4520 4980 4600 4990
rect -560 3370 -480 3380
rect -560 3290 -555 3370
rect -525 3290 -480 3370
rect -560 3280 -480 3290
rect -280 3370 -200 3380
rect -280 3290 -235 3370
rect -205 3290 -200 3370
rect -280 3280 -200 3290
rect -560 3150 -480 3160
rect -560 3070 -555 3150
rect -525 3070 -480 3150
rect -560 3060 -480 3070
rect -280 3150 -200 3160
rect -280 3070 -235 3150
rect -205 3070 -200 3150
rect -280 3060 -200 3070
rect -80 3370 0 3380
rect -80 3290 -75 3370
rect -45 3290 0 3370
rect -80 3280 0 3290
rect 200 3370 320 3380
rect 200 3290 245 3370
rect 275 3290 320 3370
rect 200 3280 320 3290
rect 520 3370 640 3380
rect 520 3290 565 3370
rect 595 3290 640 3370
rect 520 3280 640 3290
rect 840 3370 960 3380
rect 840 3290 885 3370
rect 915 3290 960 3370
rect 840 3280 960 3290
rect 1160 3370 1240 3380
rect 1160 3290 1205 3370
rect 1235 3290 1240 3370
rect 1160 3280 1240 3290
rect -80 3150 0 3160
rect -80 3070 -75 3150
rect -45 3070 0 3150
rect -80 3060 0 3070
rect 200 3150 320 3160
rect 200 3070 245 3150
rect 275 3070 320 3150
rect 200 3060 320 3070
rect 520 3150 640 3160
rect 520 3070 565 3150
rect 595 3070 640 3150
rect 520 3060 640 3070
rect 840 3150 960 3160
rect 840 3070 885 3150
rect 915 3070 960 3150
rect 840 3060 960 3070
rect 1160 3150 1240 3160
rect 1160 3070 1205 3150
rect 1235 3070 1240 3150
rect 1160 3060 1240 3070
rect 1360 3370 1440 3380
rect 1360 3290 1365 3370
rect 1395 3290 1440 3370
rect 1360 3280 1440 3290
rect 1640 3370 1760 3380
rect 1640 3290 1685 3370
rect 1715 3290 1760 3370
rect 1640 3280 1760 3290
rect 1960 3370 2080 3380
rect 1960 3290 2005 3370
rect 2035 3290 2080 3370
rect 1960 3280 2080 3290
rect 2280 3370 2400 3380
rect 2280 3290 2325 3370
rect 2355 3290 2400 3370
rect 2280 3280 2400 3290
rect 2600 3370 2680 3380
rect 2600 3290 2645 3370
rect 2675 3290 2680 3370
rect 2600 3280 2680 3290
rect 1360 3150 1440 3160
rect 1360 3070 1365 3150
rect 1395 3070 1440 3150
rect 1360 3060 1440 3070
rect 1640 3150 1760 3160
rect 1640 3070 1685 3150
rect 1715 3070 1760 3150
rect 1640 3060 1760 3070
rect 1960 3150 2080 3160
rect 1960 3070 2005 3150
rect 2035 3070 2080 3150
rect 1960 3060 2080 3070
rect 2280 3150 2400 3160
rect 2280 3070 2325 3150
rect 2355 3070 2400 3150
rect 2280 3060 2400 3070
rect 2600 3150 2680 3160
rect 2600 3070 2645 3150
rect 2675 3070 2680 3150
rect 2600 3060 2680 3070
rect 2800 3370 2880 3380
rect 2800 3290 2805 3370
rect 2835 3290 2880 3370
rect 2800 3280 2880 3290
rect 3080 3370 3200 3380
rect 3080 3290 3125 3370
rect 3155 3290 3200 3370
rect 3080 3280 3200 3290
rect 3400 3370 3520 3380
rect 3400 3290 3445 3370
rect 3475 3290 3520 3370
rect 3400 3280 3520 3290
rect 3720 3370 3840 3380
rect 3720 3290 3765 3370
rect 3795 3290 3840 3370
rect 3720 3280 3840 3290
rect 4040 3370 4120 3380
rect 4040 3290 4085 3370
rect 4115 3290 4120 3370
rect 4040 3280 4120 3290
rect 2800 3150 2880 3160
rect 2800 3070 2805 3150
rect 2835 3070 2880 3150
rect 2800 3060 2880 3070
rect 3080 3150 3200 3160
rect 3080 3070 3125 3150
rect 3155 3070 3200 3150
rect 3080 3060 3200 3070
rect 3400 3150 3520 3160
rect 3400 3070 3445 3150
rect 3475 3070 3520 3150
rect 3400 3060 3520 3070
rect 3720 3150 3840 3160
rect 3720 3070 3765 3150
rect 3795 3070 3840 3150
rect 3720 3060 3840 3070
rect 4040 3150 4120 3160
rect 4040 3070 4085 3150
rect 4115 3070 4120 3150
rect 4040 3060 4120 3070
rect 4240 3370 4320 3380
rect 4240 3290 4245 3370
rect 4275 3290 4320 3370
rect 4240 3280 4320 3290
rect 4520 3370 4600 3380
rect 4520 3290 4565 3370
rect 4595 3290 4600 3370
rect 4520 3280 4600 3290
rect 4240 3150 4320 3160
rect 4240 3070 4245 3150
rect 4275 3070 4320 3150
rect 4240 3060 4320 3070
rect 4520 3150 4600 3160
rect 4520 3070 4565 3150
rect 4595 3070 4600 3150
rect 4520 3060 4600 3070
rect -560 1450 -480 1460
rect -560 1370 -555 1450
rect -525 1370 -480 1450
rect -560 1360 -480 1370
rect -280 1450 -200 1460
rect -280 1370 -235 1450
rect -205 1370 -200 1450
rect -280 1360 -200 1370
rect -560 1230 -480 1240
rect -560 1150 -555 1230
rect -525 1150 -480 1230
rect -560 1140 -480 1150
rect -280 1230 -200 1240
rect -280 1150 -235 1230
rect -205 1150 -200 1230
rect -280 1140 -200 1150
rect -80 1450 0 1460
rect -80 1370 -75 1450
rect -45 1370 0 1450
rect -80 1360 0 1370
rect 200 1450 320 1460
rect 200 1370 245 1450
rect 275 1370 320 1450
rect 200 1360 320 1370
rect 520 1450 640 1460
rect 520 1370 565 1450
rect 595 1370 640 1450
rect 520 1360 640 1370
rect 840 1450 960 1460
rect 840 1370 885 1450
rect 915 1370 960 1450
rect 840 1360 960 1370
rect 1160 1450 1240 1460
rect 1160 1370 1205 1450
rect 1235 1370 1240 1450
rect 1160 1360 1240 1370
rect -80 1230 0 1240
rect -80 1150 -75 1230
rect -45 1150 0 1230
rect -80 1140 0 1150
rect 200 1230 320 1240
rect 200 1150 245 1230
rect 275 1150 320 1230
rect 200 1140 320 1150
rect 520 1230 640 1240
rect 520 1150 565 1230
rect 595 1150 640 1230
rect 520 1140 640 1150
rect 840 1230 960 1240
rect 840 1150 885 1230
rect 915 1150 960 1230
rect 840 1140 960 1150
rect 1160 1230 1240 1240
rect 1160 1150 1205 1230
rect 1235 1150 1240 1230
rect 1160 1140 1240 1150
rect 1360 1450 1440 1460
rect 1360 1370 1365 1450
rect 1395 1370 1440 1450
rect 1360 1360 1440 1370
rect 1640 1450 1760 1460
rect 1640 1370 1685 1450
rect 1715 1370 1760 1450
rect 1640 1360 1760 1370
rect 1960 1450 2080 1460
rect 1960 1370 2005 1450
rect 2035 1370 2080 1450
rect 1960 1360 2080 1370
rect 2280 1450 2400 1460
rect 2280 1370 2325 1450
rect 2355 1370 2400 1450
rect 2280 1360 2400 1370
rect 2600 1450 2680 1460
rect 2600 1370 2645 1450
rect 2675 1370 2680 1450
rect 2600 1360 2680 1370
rect 1360 1230 1440 1240
rect 1360 1150 1365 1230
rect 1395 1150 1440 1230
rect 1360 1140 1440 1150
rect 1640 1230 1760 1240
rect 1640 1150 1685 1230
rect 1715 1150 1760 1230
rect 1640 1140 1760 1150
rect 1960 1230 2080 1240
rect 1960 1150 2005 1230
rect 2035 1150 2080 1230
rect 1960 1140 2080 1150
rect 2280 1230 2400 1240
rect 2280 1150 2325 1230
rect 2355 1150 2400 1230
rect 2280 1140 2400 1150
rect 2600 1230 2680 1240
rect 2600 1150 2645 1230
rect 2675 1150 2680 1230
rect 2600 1140 2680 1150
rect 2800 1450 2880 1460
rect 2800 1370 2805 1450
rect 2835 1370 2880 1450
rect 2800 1360 2880 1370
rect 3080 1450 3200 1460
rect 3080 1370 3125 1450
rect 3155 1370 3200 1450
rect 3080 1360 3200 1370
rect 3400 1450 3520 1460
rect 3400 1370 3445 1450
rect 3475 1370 3520 1450
rect 3400 1360 3520 1370
rect 3720 1450 3840 1460
rect 3720 1370 3765 1450
rect 3795 1370 3840 1450
rect 3720 1360 3840 1370
rect 4040 1450 4120 1460
rect 4040 1370 4085 1450
rect 4115 1370 4120 1450
rect 4040 1360 4120 1370
rect 2800 1230 2880 1240
rect 2800 1150 2805 1230
rect 2835 1150 2880 1230
rect 2800 1140 2880 1150
rect 3080 1230 3200 1240
rect 3080 1150 3125 1230
rect 3155 1150 3200 1230
rect 3080 1140 3200 1150
rect 3400 1230 3520 1240
rect 3400 1150 3445 1230
rect 3475 1150 3520 1230
rect 3400 1140 3520 1150
rect 3720 1230 3840 1240
rect 3720 1150 3765 1230
rect 3795 1150 3840 1230
rect 3720 1140 3840 1150
rect 4040 1230 4120 1240
rect 4040 1150 4085 1230
rect 4115 1150 4120 1230
rect 4040 1140 4120 1150
rect 4240 1450 4320 1460
rect 4240 1370 4245 1450
rect 4275 1370 4320 1450
rect 4240 1360 4320 1370
rect 4520 1450 4600 1460
rect 4520 1370 4565 1450
rect 4595 1370 4600 1450
rect 4520 1360 4600 1370
rect 4240 1230 4320 1240
rect 4240 1150 4245 1230
rect 4275 1150 4320 1230
rect 4240 1140 4320 1150
rect 4520 1230 4600 1240
rect 4520 1150 4565 1230
rect 4595 1150 4600 1230
rect 4520 1140 4600 1150
<< mvndiffc >>
rect -555 3850 -525 3930
rect -235 3850 -205 3930
rect -75 3850 -45 3930
rect 245 3850 275 3930
rect 565 3850 595 3930
rect 885 3850 915 3930
rect 1205 3850 1235 3930
rect 1365 3850 1395 3930
rect 1685 3850 1715 3930
rect 2005 3850 2035 3930
rect 2325 3850 2355 3930
rect 2645 3850 2675 3930
rect 2805 3850 2835 3930
rect 3125 3850 3155 3930
rect 3445 3850 3475 3930
rect 3765 3850 3795 3930
rect 4085 3850 4115 3930
rect 4245 3850 4275 3930
rect 4565 3850 4595 3930
rect -555 1930 -525 2010
rect -235 1930 -205 2010
rect -75 1930 -45 2010
rect 245 1930 275 2010
rect 565 1930 595 2010
rect 885 1930 915 2010
rect 1205 1930 1235 2010
rect 1365 1930 1395 2010
rect 1685 1930 1715 2010
rect 2005 1930 2035 2010
rect 2325 1930 2355 2010
rect 2645 1930 2675 2010
rect 2805 1930 2835 2010
rect 3125 1930 3155 2010
rect 3445 1930 3475 2010
rect 3765 1930 3795 2010
rect 4085 1930 4115 2010
rect 4245 1930 4275 2010
rect 4565 1930 4595 2010
rect -555 10 -525 90
rect -235 10 -205 90
rect -75 10 -45 90
rect 245 10 275 90
rect 565 10 595 90
rect 885 10 915 90
rect 1205 10 1235 90
rect 1365 10 1395 90
rect 1685 10 1715 90
rect 2005 10 2035 90
rect 2325 10 2355 90
rect 2645 10 2675 90
rect 2805 10 2835 90
rect 3125 10 3155 90
rect 3445 10 3475 90
rect 3765 10 3795 90
rect 4085 10 4115 90
rect 4245 10 4275 90
rect 4565 10 4595 90
<< mvpdiffc >>
rect -555 5210 -525 5290
rect -235 5210 -205 5290
rect -555 4990 -525 5070
rect -235 4990 -205 5070
rect -75 5210 -45 5290
rect 245 5210 275 5290
rect 565 5210 595 5290
rect 885 5210 915 5290
rect 1205 5210 1235 5290
rect -75 4990 -45 5070
rect 245 4990 275 5070
rect 565 4990 595 5070
rect 885 4990 915 5070
rect 1205 4990 1235 5070
rect 1365 5210 1395 5290
rect 1685 5210 1715 5290
rect 2005 5210 2035 5290
rect 2325 5210 2355 5290
rect 2645 5210 2675 5290
rect 1365 4990 1395 5070
rect 1685 4990 1715 5070
rect 2005 4990 2035 5070
rect 2325 4990 2355 5070
rect 2645 4990 2675 5070
rect 2805 5210 2835 5290
rect 3125 5210 3155 5290
rect 3445 5210 3475 5290
rect 3765 5210 3795 5290
rect 4085 5210 4115 5290
rect 2805 4990 2835 5070
rect 3125 4990 3155 5070
rect 3445 4990 3475 5070
rect 3765 4990 3795 5070
rect 4085 4990 4115 5070
rect 4245 5210 4275 5290
rect 4565 5210 4595 5290
rect 4245 4990 4275 5070
rect 4565 4990 4595 5070
rect -555 3290 -525 3370
rect -235 3290 -205 3370
rect -555 3070 -525 3150
rect -235 3070 -205 3150
rect -75 3290 -45 3370
rect 245 3290 275 3370
rect 565 3290 595 3370
rect 885 3290 915 3370
rect 1205 3290 1235 3370
rect -75 3070 -45 3150
rect 245 3070 275 3150
rect 565 3070 595 3150
rect 885 3070 915 3150
rect 1205 3070 1235 3150
rect 1365 3290 1395 3370
rect 1685 3290 1715 3370
rect 2005 3290 2035 3370
rect 2325 3290 2355 3370
rect 2645 3290 2675 3370
rect 1365 3070 1395 3150
rect 1685 3070 1715 3150
rect 2005 3070 2035 3150
rect 2325 3070 2355 3150
rect 2645 3070 2675 3150
rect 2805 3290 2835 3370
rect 3125 3290 3155 3370
rect 3445 3290 3475 3370
rect 3765 3290 3795 3370
rect 4085 3290 4115 3370
rect 2805 3070 2835 3150
rect 3125 3070 3155 3150
rect 3445 3070 3475 3150
rect 3765 3070 3795 3150
rect 4085 3070 4115 3150
rect 4245 3290 4275 3370
rect 4565 3290 4595 3370
rect 4245 3070 4275 3150
rect 4565 3070 4595 3150
rect -555 1370 -525 1450
rect -235 1370 -205 1450
rect -555 1150 -525 1230
rect -235 1150 -205 1230
rect -75 1370 -45 1450
rect 245 1370 275 1450
rect 565 1370 595 1450
rect 885 1370 915 1450
rect 1205 1370 1235 1450
rect -75 1150 -45 1230
rect 245 1150 275 1230
rect 565 1150 595 1230
rect 885 1150 915 1230
rect 1205 1150 1235 1230
rect 1365 1370 1395 1450
rect 1685 1370 1715 1450
rect 2005 1370 2035 1450
rect 2325 1370 2355 1450
rect 2645 1370 2675 1450
rect 1365 1150 1395 1230
rect 1685 1150 1715 1230
rect 2005 1150 2035 1230
rect 2325 1150 2355 1230
rect 2645 1150 2675 1230
rect 2805 1370 2835 1450
rect 3125 1370 3155 1450
rect 3445 1370 3475 1450
rect 3765 1370 3795 1450
rect 4085 1370 4115 1450
rect 2805 1150 2835 1230
rect 3125 1150 3155 1230
rect 3445 1150 3475 1230
rect 3765 1150 3795 1230
rect 4085 1150 4115 1230
rect 4245 1370 4275 1450
rect 4565 1370 4595 1450
rect 4245 1150 4275 1230
rect 4565 1150 4595 1230
<< mvpsubdiff >>
rect -800 5560 -680 5600
rect 4760 5560 4840 5600
rect -800 4680 -680 4720
rect 4760 4680 4840 4720
rect -800 4040 -560 4080
rect -200 4040 -80 4080
rect 1240 4040 1360 4080
rect 2680 4040 2800 4080
rect 4120 4040 4240 4080
rect 4600 4040 4840 4080
rect -800 3720 -560 3760
rect -200 3720 -80 3760
rect 1240 3720 1360 3760
rect 2680 3720 2800 3760
rect 4120 3720 4240 3760
rect 4600 3720 4840 3760
rect -800 3680 -760 3720
rect 4800 3680 4840 3720
rect -800 3640 -680 3680
rect 4760 3640 4840 3680
rect -800 2760 -680 2800
rect 4760 2760 4840 2800
rect -800 2120 -560 2160
rect -200 2120 -80 2160
rect 1240 2120 1360 2160
rect 2680 2120 2800 2160
rect 4120 2120 4240 2160
rect 4600 2120 4840 2160
rect -800 1800 -560 1840
rect -200 1800 -80 1840
rect 1240 1800 1360 1840
rect 2680 1800 2800 1840
rect 4120 1800 4240 1840
rect 4600 1800 4840 1840
rect -800 1760 -760 1800
rect 4800 1760 4840 1800
rect -800 1720 -680 1760
rect 4760 1720 4840 1760
rect -800 840 -680 880
rect 4760 840 4840 880
rect -800 200 -560 240
rect -200 200 -80 240
rect 1240 200 1360 240
rect 2680 200 2800 240
rect 4120 200 4240 240
rect 4600 200 4840 240
rect -800 -120 -560 -80
rect -200 -120 -80 -80
rect 1240 -120 1360 -80
rect 2680 -120 2800 -80
rect 4120 -120 4240 -80
rect 4600 -120 4840 -80
<< mvnsubdiff >>
rect -640 5400 -560 5440
rect -200 5400 -80 5440
rect 1240 5400 1360 5440
rect 2680 5400 2800 5440
rect 4120 5400 4240 5440
rect 4600 5400 4680 5440
rect -640 4840 -560 4880
rect -200 4840 -80 4880
rect 1240 4840 1360 4880
rect 2680 4840 2800 4880
rect 4120 4840 4240 4880
rect 4600 4840 4680 4880
rect -640 3480 -560 3520
rect -200 3480 -80 3520
rect 1240 3480 1360 3520
rect 2680 3480 2800 3520
rect 4120 3480 4240 3520
rect 4600 3480 4680 3520
rect -640 2920 -560 2960
rect -200 2920 -80 2960
rect 1240 2920 1360 2960
rect 2680 2920 2800 2960
rect 4120 2920 4240 2960
rect 4600 2920 4680 2960
rect -640 1560 -560 1600
rect -200 1560 -80 1600
rect 1240 1560 1360 1600
rect 2680 1560 2800 1600
rect 4120 1560 4240 1600
rect 4600 1560 4680 1600
rect -640 1000 -560 1040
rect -200 1000 -80 1040
rect 1240 1000 1360 1040
rect 2680 1000 2800 1040
rect 4120 1000 4240 1040
rect 4600 1000 4680 1040
<< mvpsubdiffcont >>
rect -680 5560 4760 5600
rect -800 4720 -760 5560
rect 4800 4720 4840 5560
rect -680 4680 4760 4720
rect -800 4080 -760 4680
rect 4800 4080 4840 4680
rect -560 4040 -200 4080
rect -80 4040 1240 4080
rect 1360 4040 2680 4080
rect 2800 4040 4120 4080
rect 4240 4040 4600 4080
rect -800 3760 -760 4040
rect -640 3760 -600 4040
rect -160 3760 -120 4040
rect 1280 3760 1320 4040
rect 2720 3760 2760 4040
rect 4160 3760 4200 4040
rect 4640 3760 4680 4040
rect 4800 3760 4840 4040
rect -560 3720 -200 3760
rect -80 3720 1240 3760
rect 1360 3720 2680 3760
rect 2800 3720 4120 3760
rect 4240 3720 4600 3760
rect -680 3640 4760 3680
rect -800 2800 -760 3640
rect 4800 2800 4840 3640
rect -680 2760 4760 2800
rect -800 2160 -760 2760
rect 4800 2160 4840 2760
rect -560 2120 -200 2160
rect -80 2120 1240 2160
rect 1360 2120 2680 2160
rect 2800 2120 4120 2160
rect 4240 2120 4600 2160
rect -800 1840 -760 2120
rect -640 1840 -600 2120
rect -160 1840 -120 2120
rect 1280 1840 1320 2120
rect 2720 1840 2760 2120
rect 4160 1840 4200 2120
rect 4640 1840 4680 2120
rect 4800 1840 4840 2120
rect -560 1800 -200 1840
rect -80 1800 1240 1840
rect 1360 1800 2680 1840
rect 2800 1800 4120 1840
rect 4240 1800 4600 1840
rect -680 1720 4760 1760
rect -800 880 -760 1720
rect 4800 880 4840 1720
rect -680 840 4760 880
rect -800 240 -760 840
rect 4800 240 4840 840
rect -560 200 -200 240
rect -80 200 1240 240
rect 1360 200 2680 240
rect 2800 200 4120 240
rect 4240 200 4600 240
rect -800 -80 -760 200
rect -640 -80 -600 200
rect -160 -80 -120 200
rect 1280 -80 1320 200
rect 2720 -80 2760 200
rect 4160 -80 4200 200
rect 4640 -80 4680 200
rect 4800 -80 4840 200
rect -560 -120 -200 -80
rect -80 -120 1240 -80
rect 1360 -120 2680 -80
rect 2800 -120 4120 -80
rect 4240 -120 4600 -80
<< mvnsubdiffcont >>
rect -560 5400 -200 5440
rect -80 5400 1240 5440
rect 1360 5400 2680 5440
rect 2800 5400 4120 5440
rect 4240 5400 4600 5440
rect -640 4880 -600 5400
rect -160 4880 -120 5400
rect 1280 4880 1320 5400
rect 2720 4880 2760 5400
rect 4160 4880 4200 5400
rect 4640 4880 4680 5400
rect -560 4840 -200 4880
rect -80 4840 1240 4880
rect 1360 4840 2680 4880
rect 2800 4840 4120 4880
rect 4240 4840 4600 4880
rect -560 3480 -200 3520
rect -80 3480 1240 3520
rect 1360 3480 2680 3520
rect 2800 3480 4120 3520
rect 4240 3480 4600 3520
rect -640 2960 -600 3480
rect -160 2960 -120 3480
rect 1280 2960 1320 3480
rect 2720 2960 2760 3480
rect 4160 2960 4200 3480
rect 4640 2960 4680 3480
rect -560 2920 -200 2960
rect -80 2920 1240 2960
rect 1360 2920 2680 2960
rect 2800 2920 4120 2960
rect 4240 2920 4600 2960
rect -560 1560 -200 1600
rect -80 1560 1240 1600
rect 1360 1560 2680 1600
rect 2800 1560 4120 1600
rect 4240 1560 4600 1600
rect -640 1040 -600 1560
rect -160 1040 -120 1560
rect 1280 1040 1320 1560
rect 2720 1040 2760 1560
rect 4160 1040 4200 1560
rect 4640 1040 4680 1560
rect -560 1000 -200 1040
rect -80 1000 1240 1040
rect 1360 1000 2680 1040
rect 2800 1000 4120 1040
rect 4240 1000 4600 1040
<< poly >>
rect -480 5355 -280 5360
rect -480 5325 -470 5355
rect -290 5325 -280 5355
rect -480 5300 -280 5325
rect -480 5180 -280 5200
rect -480 5080 -280 5100
rect -480 4955 -280 4980
rect -480 4925 -470 4955
rect -290 4925 -280 4955
rect -480 4920 -280 4925
rect 0 5355 200 5360
rect 0 5325 10 5355
rect 190 5325 200 5355
rect 0 5300 200 5325
rect 320 5355 520 5360
rect 320 5325 330 5355
rect 510 5325 520 5355
rect 320 5300 520 5325
rect 640 5355 840 5360
rect 640 5325 650 5355
rect 830 5325 840 5355
rect 640 5300 840 5325
rect 960 5355 1160 5360
rect 960 5325 970 5355
rect 1150 5325 1160 5355
rect 960 5300 1160 5325
rect 0 5180 200 5200
rect 320 5180 520 5200
rect 640 5180 840 5200
rect 960 5180 1160 5200
rect 0 5080 200 5100
rect 320 5080 520 5100
rect 640 5080 840 5100
rect 960 5080 1160 5100
rect 0 4955 200 4980
rect 0 4925 10 4955
rect 190 4925 200 4955
rect 0 4920 200 4925
rect 320 4955 520 4980
rect 320 4925 330 4955
rect 510 4925 520 4955
rect 320 4920 520 4925
rect 640 4955 840 4980
rect 640 4925 650 4955
rect 830 4925 840 4955
rect 640 4920 840 4925
rect 960 4955 1160 4980
rect 960 4925 970 4955
rect 1150 4925 1160 4955
rect 960 4920 1160 4925
rect 1440 5355 1640 5360
rect 1440 5325 1450 5355
rect 1630 5325 1640 5355
rect 1440 5300 1640 5325
rect 1760 5355 1960 5360
rect 1760 5325 1770 5355
rect 1950 5325 1960 5355
rect 1760 5300 1960 5325
rect 2080 5355 2280 5360
rect 2080 5325 2090 5355
rect 2270 5325 2280 5355
rect 2080 5300 2280 5325
rect 2400 5355 2600 5360
rect 2400 5325 2410 5355
rect 2590 5325 2600 5355
rect 2400 5300 2600 5325
rect 1440 5180 1640 5200
rect 1760 5180 1960 5200
rect 2080 5180 2280 5200
rect 2400 5180 2600 5200
rect 1440 5080 1640 5100
rect 1760 5080 1960 5100
rect 2080 5080 2280 5100
rect 2400 5080 2600 5100
rect 1440 4955 1640 4980
rect 1440 4925 1450 4955
rect 1630 4925 1640 4955
rect 1440 4920 1640 4925
rect 1760 4955 1960 4980
rect 1760 4925 1770 4955
rect 1950 4925 1960 4955
rect 1760 4920 1960 4925
rect 2080 4955 2280 4980
rect 2080 4925 2090 4955
rect 2270 4925 2280 4955
rect 2080 4920 2280 4925
rect 2400 4955 2600 4980
rect 2400 4925 2410 4955
rect 2590 4925 2600 4955
rect 2400 4920 2600 4925
rect 2880 5355 3080 5360
rect 2880 5325 2890 5355
rect 3070 5325 3080 5355
rect 2880 5300 3080 5325
rect 3200 5355 3400 5360
rect 3200 5325 3210 5355
rect 3390 5325 3400 5355
rect 3200 5300 3400 5325
rect 3520 5355 3720 5360
rect 3520 5325 3530 5355
rect 3710 5325 3720 5355
rect 3520 5300 3720 5325
rect 3840 5355 4040 5360
rect 3840 5325 3850 5355
rect 4030 5325 4040 5355
rect 3840 5300 4040 5325
rect 2880 5180 3080 5200
rect 3200 5180 3400 5200
rect 3520 5180 3720 5200
rect 3840 5180 4040 5200
rect 2880 5080 3080 5100
rect 3200 5080 3400 5100
rect 3520 5080 3720 5100
rect 3840 5080 4040 5100
rect 2880 4955 3080 4980
rect 2880 4925 2890 4955
rect 3070 4925 3080 4955
rect 2880 4920 3080 4925
rect 3200 4955 3400 4980
rect 3200 4925 3210 4955
rect 3390 4925 3400 4955
rect 3200 4920 3400 4925
rect 3520 4955 3720 4980
rect 3520 4925 3530 4955
rect 3710 4925 3720 4955
rect 3520 4920 3720 4925
rect 3840 4955 4040 4980
rect 3840 4925 3850 4955
rect 4030 4925 4040 4955
rect 3840 4920 4040 4925
rect 4320 5355 4520 5360
rect 4320 5325 4330 5355
rect 4510 5325 4520 5355
rect 4320 5300 4520 5325
rect 4320 5180 4520 5200
rect 4320 5080 4520 5100
rect 4320 4955 4520 4980
rect 4320 4925 4330 4955
rect 4510 4925 4520 4955
rect 4320 4920 4520 4925
rect -480 3995 -280 4000
rect -480 3965 -470 3995
rect -290 3965 -280 3995
rect -480 3940 -280 3965
rect -480 3820 -280 3840
rect 0 3995 200 4000
rect 0 3965 10 3995
rect 190 3965 200 3995
rect 0 3940 200 3965
rect 320 3995 520 4000
rect 320 3965 330 3995
rect 510 3965 520 3995
rect 320 3940 520 3965
rect 640 3995 840 4000
rect 640 3965 650 3995
rect 830 3965 840 3995
rect 640 3940 840 3965
rect 960 3995 1160 4000
rect 960 3965 970 3995
rect 1150 3965 1160 3995
rect 960 3940 1160 3965
rect 0 3820 200 3840
rect 320 3820 520 3840
rect 640 3820 840 3840
rect 960 3820 1160 3840
rect 1440 3995 1640 4000
rect 1440 3965 1450 3995
rect 1630 3965 1640 3995
rect 1440 3940 1640 3965
rect 1760 3995 1960 4000
rect 1760 3965 1770 3995
rect 1950 3965 1960 3995
rect 1760 3940 1960 3965
rect 2080 3995 2280 4000
rect 2080 3965 2090 3995
rect 2270 3965 2280 3995
rect 2080 3940 2280 3965
rect 2400 3995 2600 4000
rect 2400 3965 2410 3995
rect 2590 3965 2600 3995
rect 2400 3940 2600 3965
rect 1440 3820 1640 3840
rect 1760 3820 1960 3840
rect 2080 3820 2280 3840
rect 2400 3820 2600 3840
rect 2880 3995 3080 4000
rect 2880 3965 2890 3995
rect 3070 3965 3080 3995
rect 2880 3940 3080 3965
rect 3200 3995 3400 4000
rect 3200 3965 3210 3995
rect 3390 3965 3400 3995
rect 3200 3940 3400 3965
rect 3520 3995 3720 4000
rect 3520 3965 3530 3995
rect 3710 3965 3720 3995
rect 3520 3940 3720 3965
rect 3840 3995 4040 4000
rect 3840 3965 3850 3995
rect 4030 3965 4040 3995
rect 3840 3940 4040 3965
rect 2880 3820 3080 3840
rect 3200 3820 3400 3840
rect 3520 3820 3720 3840
rect 3840 3820 4040 3840
rect 4320 3995 4520 4000
rect 4320 3965 4330 3995
rect 4510 3965 4520 3995
rect 4320 3940 4520 3965
rect 4320 3820 4520 3840
rect -480 3435 -280 3440
rect -480 3405 -470 3435
rect -290 3405 -280 3435
rect -480 3380 -280 3405
rect -480 3260 -280 3280
rect -480 3160 -280 3180
rect -480 3035 -280 3060
rect -480 3005 -470 3035
rect -290 3005 -280 3035
rect -480 3000 -280 3005
rect 0 3435 200 3440
rect 0 3405 10 3435
rect 190 3405 200 3435
rect 0 3380 200 3405
rect 320 3435 520 3440
rect 320 3405 330 3435
rect 510 3405 520 3435
rect 320 3380 520 3405
rect 640 3435 840 3440
rect 640 3405 650 3435
rect 830 3405 840 3435
rect 640 3380 840 3405
rect 960 3435 1160 3440
rect 960 3405 970 3435
rect 1150 3405 1160 3435
rect 960 3380 1160 3405
rect 0 3260 200 3280
rect 320 3260 520 3280
rect 640 3260 840 3280
rect 960 3260 1160 3280
rect 0 3160 200 3180
rect 320 3160 520 3180
rect 640 3160 840 3180
rect 960 3160 1160 3180
rect 0 3035 200 3060
rect 0 3005 10 3035
rect 190 3005 200 3035
rect 0 3000 200 3005
rect 320 3035 520 3060
rect 320 3005 330 3035
rect 510 3005 520 3035
rect 320 3000 520 3005
rect 640 3035 840 3060
rect 640 3005 650 3035
rect 830 3005 840 3035
rect 640 3000 840 3005
rect 960 3035 1160 3060
rect 960 3005 970 3035
rect 1150 3005 1160 3035
rect 960 3000 1160 3005
rect 1440 3435 1640 3440
rect 1440 3405 1450 3435
rect 1630 3405 1640 3435
rect 1440 3380 1640 3405
rect 1760 3435 1960 3440
rect 1760 3405 1770 3435
rect 1950 3405 1960 3435
rect 1760 3380 1960 3405
rect 2080 3435 2280 3440
rect 2080 3405 2090 3435
rect 2270 3405 2280 3435
rect 2080 3380 2280 3405
rect 2400 3435 2600 3440
rect 2400 3405 2410 3435
rect 2590 3405 2600 3435
rect 2400 3380 2600 3405
rect 1440 3260 1640 3280
rect 1760 3260 1960 3280
rect 2080 3260 2280 3280
rect 2400 3260 2600 3280
rect 1440 3160 1640 3180
rect 1760 3160 1960 3180
rect 2080 3160 2280 3180
rect 2400 3160 2600 3180
rect 1440 3035 1640 3060
rect 1440 3005 1450 3035
rect 1630 3005 1640 3035
rect 1440 3000 1640 3005
rect 1760 3035 1960 3060
rect 1760 3005 1770 3035
rect 1950 3005 1960 3035
rect 1760 3000 1960 3005
rect 2080 3035 2280 3060
rect 2080 3005 2090 3035
rect 2270 3005 2280 3035
rect 2080 3000 2280 3005
rect 2400 3035 2600 3060
rect 2400 3005 2410 3035
rect 2590 3005 2600 3035
rect 2400 3000 2600 3005
rect 2880 3435 3080 3440
rect 2880 3405 2890 3435
rect 3070 3405 3080 3435
rect 2880 3380 3080 3405
rect 3200 3435 3400 3440
rect 3200 3405 3210 3435
rect 3390 3405 3400 3435
rect 3200 3380 3400 3405
rect 3520 3435 3720 3440
rect 3520 3405 3530 3435
rect 3710 3405 3720 3435
rect 3520 3380 3720 3405
rect 3840 3435 4040 3440
rect 3840 3405 3850 3435
rect 4030 3405 4040 3435
rect 3840 3380 4040 3405
rect 2880 3260 3080 3280
rect 3200 3260 3400 3280
rect 3520 3260 3720 3280
rect 3840 3260 4040 3280
rect 2880 3160 3080 3180
rect 3200 3160 3400 3180
rect 3520 3160 3720 3180
rect 3840 3160 4040 3180
rect 2880 3035 3080 3060
rect 2880 3005 2890 3035
rect 3070 3005 3080 3035
rect 2880 3000 3080 3005
rect 3200 3035 3400 3060
rect 3200 3005 3210 3035
rect 3390 3005 3400 3035
rect 3200 3000 3400 3005
rect 3520 3035 3720 3060
rect 3520 3005 3530 3035
rect 3710 3005 3720 3035
rect 3520 3000 3720 3005
rect 3840 3035 4040 3060
rect 3840 3005 3850 3035
rect 4030 3005 4040 3035
rect 3840 3000 4040 3005
rect 4320 3435 4520 3440
rect 4320 3405 4330 3435
rect 4510 3405 4520 3435
rect 4320 3380 4520 3405
rect 4320 3260 4520 3280
rect 4320 3160 4520 3180
rect 4320 3035 4520 3060
rect 4320 3005 4330 3035
rect 4510 3005 4520 3035
rect 4320 3000 4520 3005
rect -480 2075 -280 2080
rect -480 2045 -470 2075
rect -290 2045 -280 2075
rect -480 2020 -280 2045
rect -480 1900 -280 1920
rect 0 2075 200 2080
rect 0 2045 10 2075
rect 190 2045 200 2075
rect 0 2020 200 2045
rect 320 2075 520 2080
rect 320 2045 330 2075
rect 510 2045 520 2075
rect 320 2020 520 2045
rect 640 2075 840 2080
rect 640 2045 650 2075
rect 830 2045 840 2075
rect 640 2020 840 2045
rect 960 2075 1160 2080
rect 960 2045 970 2075
rect 1150 2045 1160 2075
rect 960 2020 1160 2045
rect 0 1900 200 1920
rect 320 1900 520 1920
rect 640 1900 840 1920
rect 960 1900 1160 1920
rect 1440 2075 1640 2080
rect 1440 2045 1450 2075
rect 1630 2045 1640 2075
rect 1440 2020 1640 2045
rect 1760 2075 1960 2080
rect 1760 2045 1770 2075
rect 1950 2045 1960 2075
rect 1760 2020 1960 2045
rect 2080 2075 2280 2080
rect 2080 2045 2090 2075
rect 2270 2045 2280 2075
rect 2080 2020 2280 2045
rect 2400 2075 2600 2080
rect 2400 2045 2410 2075
rect 2590 2045 2600 2075
rect 2400 2020 2600 2045
rect 1440 1900 1640 1920
rect 1760 1900 1960 1920
rect 2080 1900 2280 1920
rect 2400 1900 2600 1920
rect 2880 2075 3080 2080
rect 2880 2045 2890 2075
rect 3070 2045 3080 2075
rect 2880 2020 3080 2045
rect 3200 2075 3400 2080
rect 3200 2045 3210 2075
rect 3390 2045 3400 2075
rect 3200 2020 3400 2045
rect 3520 2075 3720 2080
rect 3520 2045 3530 2075
rect 3710 2045 3720 2075
rect 3520 2020 3720 2045
rect 3840 2075 4040 2080
rect 3840 2045 3850 2075
rect 4030 2045 4040 2075
rect 3840 2020 4040 2045
rect 2880 1900 3080 1920
rect 3200 1900 3400 1920
rect 3520 1900 3720 1920
rect 3840 1900 4040 1920
rect 4320 2075 4520 2080
rect 4320 2045 4330 2075
rect 4510 2045 4520 2075
rect 4320 2020 4520 2045
rect 4320 1900 4520 1920
rect -480 1515 -280 1520
rect -480 1485 -470 1515
rect -290 1485 -280 1515
rect -480 1460 -280 1485
rect -480 1340 -280 1360
rect -480 1240 -280 1260
rect -480 1115 -280 1140
rect -480 1085 -470 1115
rect -290 1085 -280 1115
rect -480 1080 -280 1085
rect 0 1515 200 1520
rect 0 1485 10 1515
rect 190 1485 200 1515
rect 0 1460 200 1485
rect 320 1515 520 1520
rect 320 1485 330 1515
rect 510 1485 520 1515
rect 320 1460 520 1485
rect 640 1515 840 1520
rect 640 1485 650 1515
rect 830 1485 840 1515
rect 640 1460 840 1485
rect 960 1515 1160 1520
rect 960 1485 970 1515
rect 1150 1485 1160 1515
rect 960 1460 1160 1485
rect 0 1340 200 1360
rect 320 1340 520 1360
rect 640 1340 840 1360
rect 960 1340 1160 1360
rect 0 1240 200 1260
rect 320 1240 520 1260
rect 640 1240 840 1260
rect 960 1240 1160 1260
rect 0 1115 200 1140
rect 0 1085 10 1115
rect 190 1085 200 1115
rect 0 1080 200 1085
rect 320 1115 520 1140
rect 320 1085 330 1115
rect 510 1085 520 1115
rect 320 1080 520 1085
rect 640 1115 840 1140
rect 640 1085 650 1115
rect 830 1085 840 1115
rect 640 1080 840 1085
rect 960 1115 1160 1140
rect 960 1085 970 1115
rect 1150 1085 1160 1115
rect 960 1080 1160 1085
rect 1440 1515 1640 1520
rect 1440 1485 1450 1515
rect 1630 1485 1640 1515
rect 1440 1460 1640 1485
rect 1760 1515 1960 1520
rect 1760 1485 1770 1515
rect 1950 1485 1960 1515
rect 1760 1460 1960 1485
rect 2080 1515 2280 1520
rect 2080 1485 2090 1515
rect 2270 1485 2280 1515
rect 2080 1460 2280 1485
rect 2400 1515 2600 1520
rect 2400 1485 2410 1515
rect 2590 1485 2600 1515
rect 2400 1460 2600 1485
rect 1440 1340 1640 1360
rect 1760 1340 1960 1360
rect 2080 1340 2280 1360
rect 2400 1340 2600 1360
rect 1440 1240 1640 1260
rect 1760 1240 1960 1260
rect 2080 1240 2280 1260
rect 2400 1240 2600 1260
rect 1440 1115 1640 1140
rect 1440 1085 1450 1115
rect 1630 1085 1640 1115
rect 1440 1080 1640 1085
rect 1760 1115 1960 1140
rect 1760 1085 1770 1115
rect 1950 1085 1960 1115
rect 1760 1080 1960 1085
rect 2080 1115 2280 1140
rect 2080 1085 2090 1115
rect 2270 1085 2280 1115
rect 2080 1080 2280 1085
rect 2400 1115 2600 1140
rect 2400 1085 2410 1115
rect 2590 1085 2600 1115
rect 2400 1080 2600 1085
rect 2880 1515 3080 1520
rect 2880 1485 2890 1515
rect 3070 1485 3080 1515
rect 2880 1460 3080 1485
rect 3200 1515 3400 1520
rect 3200 1485 3210 1515
rect 3390 1485 3400 1515
rect 3200 1460 3400 1485
rect 3520 1515 3720 1520
rect 3520 1485 3530 1515
rect 3710 1485 3720 1515
rect 3520 1460 3720 1485
rect 3840 1515 4040 1520
rect 3840 1485 3850 1515
rect 4030 1485 4040 1515
rect 3840 1460 4040 1485
rect 2880 1340 3080 1360
rect 3200 1340 3400 1360
rect 3520 1340 3720 1360
rect 3840 1340 4040 1360
rect 2880 1240 3080 1260
rect 3200 1240 3400 1260
rect 3520 1240 3720 1260
rect 3840 1240 4040 1260
rect 2880 1115 3080 1140
rect 2880 1085 2890 1115
rect 3070 1085 3080 1115
rect 2880 1080 3080 1085
rect 3200 1115 3400 1140
rect 3200 1085 3210 1115
rect 3390 1085 3400 1115
rect 3200 1080 3400 1085
rect 3520 1115 3720 1140
rect 3520 1085 3530 1115
rect 3710 1085 3720 1115
rect 3520 1080 3720 1085
rect 3840 1115 4040 1140
rect 3840 1085 3850 1115
rect 4030 1085 4040 1115
rect 3840 1080 4040 1085
rect 4320 1515 4520 1520
rect 4320 1485 4330 1515
rect 4510 1485 4520 1515
rect 4320 1460 4520 1485
rect 4320 1340 4520 1360
rect 4320 1240 4520 1260
rect 4320 1115 4520 1140
rect 4320 1085 4330 1115
rect 4510 1085 4520 1115
rect 4320 1080 4520 1085
rect -480 155 -280 160
rect -480 125 -470 155
rect -290 125 -280 155
rect -480 100 -280 125
rect -480 -20 -280 0
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 100 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 100 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 100 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 100 1160 125
rect 0 -20 200 0
rect 320 -20 520 0
rect 640 -20 840 0
rect 960 -20 1160 0
rect 1440 155 1640 160
rect 1440 125 1450 155
rect 1630 125 1640 155
rect 1440 100 1640 125
rect 1760 155 1960 160
rect 1760 125 1770 155
rect 1950 125 1960 155
rect 1760 100 1960 125
rect 2080 155 2280 160
rect 2080 125 2090 155
rect 2270 125 2280 155
rect 2080 100 2280 125
rect 2400 155 2600 160
rect 2400 125 2410 155
rect 2590 125 2600 155
rect 2400 100 2600 125
rect 1440 -20 1640 0
rect 1760 -20 1960 0
rect 2080 -20 2280 0
rect 2400 -20 2600 0
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 100 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 100 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 100 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 100 4040 125
rect 2880 -20 3080 0
rect 3200 -20 3400 0
rect 3520 -20 3720 0
rect 3840 -20 4040 0
rect 4320 155 4520 160
rect 4320 125 4330 155
rect 4510 125 4520 155
rect 4320 100 4520 125
rect 4320 -20 4520 0
<< polycont >>
rect -470 5325 -290 5355
rect -470 4925 -290 4955
rect 10 5325 190 5355
rect 330 5325 510 5355
rect 650 5325 830 5355
rect 970 5325 1150 5355
rect 10 4925 190 4955
rect 330 4925 510 4955
rect 650 4925 830 4955
rect 970 4925 1150 4955
rect 1450 5325 1630 5355
rect 1770 5325 1950 5355
rect 2090 5325 2270 5355
rect 2410 5325 2590 5355
rect 1450 4925 1630 4955
rect 1770 4925 1950 4955
rect 2090 4925 2270 4955
rect 2410 4925 2590 4955
rect 2890 5325 3070 5355
rect 3210 5325 3390 5355
rect 3530 5325 3710 5355
rect 3850 5325 4030 5355
rect 2890 4925 3070 4955
rect 3210 4925 3390 4955
rect 3530 4925 3710 4955
rect 3850 4925 4030 4955
rect 4330 5325 4510 5355
rect 4330 4925 4510 4955
rect -470 3965 -290 3995
rect 10 3965 190 3995
rect 330 3965 510 3995
rect 650 3965 830 3995
rect 970 3965 1150 3995
rect 1450 3965 1630 3995
rect 1770 3965 1950 3995
rect 2090 3965 2270 3995
rect 2410 3965 2590 3995
rect 2890 3965 3070 3995
rect 3210 3965 3390 3995
rect 3530 3965 3710 3995
rect 3850 3965 4030 3995
rect 4330 3965 4510 3995
rect -470 3405 -290 3435
rect -470 3005 -290 3035
rect 10 3405 190 3435
rect 330 3405 510 3435
rect 650 3405 830 3435
rect 970 3405 1150 3435
rect 10 3005 190 3035
rect 330 3005 510 3035
rect 650 3005 830 3035
rect 970 3005 1150 3035
rect 1450 3405 1630 3435
rect 1770 3405 1950 3435
rect 2090 3405 2270 3435
rect 2410 3405 2590 3435
rect 1450 3005 1630 3035
rect 1770 3005 1950 3035
rect 2090 3005 2270 3035
rect 2410 3005 2590 3035
rect 2890 3405 3070 3435
rect 3210 3405 3390 3435
rect 3530 3405 3710 3435
rect 3850 3405 4030 3435
rect 2890 3005 3070 3035
rect 3210 3005 3390 3035
rect 3530 3005 3710 3035
rect 3850 3005 4030 3035
rect 4330 3405 4510 3435
rect 4330 3005 4510 3035
rect -470 2045 -290 2075
rect 10 2045 190 2075
rect 330 2045 510 2075
rect 650 2045 830 2075
rect 970 2045 1150 2075
rect 1450 2045 1630 2075
rect 1770 2045 1950 2075
rect 2090 2045 2270 2075
rect 2410 2045 2590 2075
rect 2890 2045 3070 2075
rect 3210 2045 3390 2075
rect 3530 2045 3710 2075
rect 3850 2045 4030 2075
rect 4330 2045 4510 2075
rect -470 1485 -290 1515
rect -470 1085 -290 1115
rect 10 1485 190 1515
rect 330 1485 510 1515
rect 650 1485 830 1515
rect 970 1485 1150 1515
rect 10 1085 190 1115
rect 330 1085 510 1115
rect 650 1085 830 1115
rect 970 1085 1150 1115
rect 1450 1485 1630 1515
rect 1770 1485 1950 1515
rect 2090 1485 2270 1515
rect 2410 1485 2590 1515
rect 1450 1085 1630 1115
rect 1770 1085 1950 1115
rect 2090 1085 2270 1115
rect 2410 1085 2590 1115
rect 2890 1485 3070 1515
rect 3210 1485 3390 1515
rect 3530 1485 3710 1515
rect 3850 1485 4030 1515
rect 2890 1085 3070 1115
rect 3210 1085 3390 1115
rect 3530 1085 3710 1115
rect 3850 1085 4030 1115
rect 4330 1485 4510 1515
rect 4330 1085 4510 1115
rect -470 125 -290 155
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect 1450 125 1630 155
rect 1770 125 1950 155
rect 2090 125 2270 155
rect 2410 125 2590 155
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3850 125 4030 155
rect 4330 125 4510 155
<< locali >>
rect -800 5560 -680 5600
rect 4760 5560 4840 5600
rect -640 5400 -560 5440
rect -200 5400 -80 5440
rect 1240 5400 1360 5440
rect 2680 5400 2800 5440
rect 4120 5400 4240 5440
rect 4600 5400 4680 5440
rect -560 5290 -520 5400
rect -480 5355 -280 5360
rect -480 5325 -470 5355
rect -290 5325 -280 5355
rect -480 5320 -280 5325
rect -560 5210 -555 5290
rect -525 5210 -520 5290
rect -560 5070 -520 5210
rect -560 4990 -555 5070
rect -525 4990 -520 5070
rect -560 4880 -520 4990
rect -240 5290 -200 5400
rect -240 5210 -235 5290
rect -205 5210 -200 5290
rect -240 5070 -200 5210
rect -240 4990 -235 5070
rect -205 4990 -200 5070
rect -480 4955 -280 4960
rect -480 4925 -470 4955
rect -290 4925 -280 4955
rect -480 4920 -280 4925
rect -240 4880 -200 4990
rect 0 5355 200 5360
rect 0 5325 10 5355
rect 190 5325 200 5355
rect 0 5320 200 5325
rect 320 5355 520 5360
rect 320 5325 330 5355
rect 510 5325 520 5355
rect 320 5320 520 5325
rect 640 5355 840 5360
rect 640 5325 650 5355
rect 830 5325 840 5355
rect 640 5320 840 5325
rect 960 5355 1160 5360
rect 960 5325 970 5355
rect 1150 5325 1160 5355
rect 960 5320 1160 5325
rect -80 5290 -40 5300
rect -80 5210 -75 5290
rect -45 5210 -40 5290
rect -80 5200 -40 5210
rect 240 5290 280 5300
rect 240 5210 245 5290
rect 275 5210 280 5290
rect 240 5200 280 5210
rect 560 5290 600 5300
rect 560 5210 565 5290
rect 595 5210 600 5290
rect 560 5200 600 5210
rect 880 5290 920 5300
rect 880 5210 885 5290
rect 915 5210 920 5290
rect 880 5200 920 5210
rect 1200 5290 1240 5300
rect 1200 5210 1205 5290
rect 1235 5210 1240 5290
rect 1200 5200 1240 5210
rect -80 5070 -40 5080
rect -80 4990 -75 5070
rect -45 4990 -40 5070
rect -80 4980 -40 4990
rect 240 5070 280 5080
rect 240 4990 245 5070
rect 275 4990 280 5070
rect 240 4980 280 4990
rect 560 5070 600 5080
rect 560 4990 565 5070
rect 595 4990 600 5070
rect 560 4980 600 4990
rect 880 5070 920 5080
rect 880 4990 885 5070
rect 915 4990 920 5070
rect 880 4980 920 4990
rect 1200 5070 1240 5080
rect 1200 4990 1205 5070
rect 1235 4990 1240 5070
rect 1200 4980 1240 4990
rect 0 4955 200 4960
rect 0 4925 10 4955
rect 190 4925 200 4955
rect 0 4920 200 4925
rect 320 4955 520 4960
rect 320 4925 330 4955
rect 510 4925 520 4955
rect 320 4920 520 4925
rect 640 4955 840 4960
rect 640 4925 650 4955
rect 830 4925 840 4955
rect 640 4920 840 4925
rect 960 4955 1160 4960
rect 960 4925 970 4955
rect 1150 4925 1160 4955
rect 960 4920 1160 4925
rect 1440 5355 1640 5360
rect 1440 5325 1450 5355
rect 1630 5325 1640 5355
rect 1440 5320 1640 5325
rect 1760 5355 1960 5360
rect 1760 5325 1770 5355
rect 1950 5325 1960 5355
rect 1760 5320 1960 5325
rect 2080 5355 2280 5360
rect 2080 5325 2090 5355
rect 2270 5325 2280 5355
rect 2080 5320 2280 5325
rect 2400 5355 2600 5360
rect 2400 5325 2410 5355
rect 2590 5325 2600 5355
rect 2400 5320 2600 5325
rect 1360 5290 1400 5300
rect 1360 5210 1365 5290
rect 1395 5210 1400 5290
rect 1360 5200 1400 5210
rect 1680 5290 1720 5300
rect 1680 5210 1685 5290
rect 1715 5210 1720 5290
rect 1680 5200 1720 5210
rect 2000 5290 2040 5300
rect 2000 5210 2005 5290
rect 2035 5210 2040 5290
rect 2000 5200 2040 5210
rect 2320 5290 2360 5300
rect 2320 5210 2325 5290
rect 2355 5210 2360 5290
rect 2320 5200 2360 5210
rect 2640 5290 2680 5300
rect 2640 5210 2645 5290
rect 2675 5210 2680 5290
rect 2640 5200 2680 5210
rect 1360 5070 1400 5080
rect 1360 4990 1365 5070
rect 1395 4990 1400 5070
rect 1360 4980 1400 4990
rect 1680 5070 1720 5080
rect 1680 4990 1685 5070
rect 1715 4990 1720 5070
rect 1680 4980 1720 4990
rect 2000 5070 2040 5080
rect 2000 4990 2005 5070
rect 2035 4990 2040 5070
rect 2000 4980 2040 4990
rect 2320 5070 2360 5080
rect 2320 4990 2325 5070
rect 2355 4990 2360 5070
rect 2320 4980 2360 4990
rect 2640 5070 2680 5080
rect 2640 4990 2645 5070
rect 2675 4990 2680 5070
rect 2640 4980 2680 4990
rect 1440 4955 1640 4960
rect 1440 4925 1450 4955
rect 1630 4925 1640 4955
rect 1440 4920 1640 4925
rect 1760 4955 1960 4960
rect 1760 4925 1770 4955
rect 1950 4925 1960 4955
rect 1760 4920 1960 4925
rect 2080 4955 2280 4960
rect 2080 4925 2090 4955
rect 2270 4925 2280 4955
rect 2080 4920 2280 4925
rect 2400 4955 2600 4960
rect 2400 4925 2410 4955
rect 2590 4925 2600 4955
rect 2400 4920 2600 4925
rect 2880 5355 3080 5360
rect 2880 5325 2890 5355
rect 3070 5325 3080 5355
rect 2880 5320 3080 5325
rect 3200 5355 3400 5360
rect 3200 5325 3210 5355
rect 3390 5325 3400 5355
rect 3200 5320 3400 5325
rect 3520 5355 3720 5360
rect 3520 5325 3530 5355
rect 3710 5325 3720 5355
rect 3520 5320 3720 5325
rect 3840 5355 4040 5360
rect 3840 5325 3850 5355
rect 4030 5325 4040 5355
rect 3840 5320 4040 5325
rect 2800 5290 2840 5300
rect 2800 5210 2805 5290
rect 2835 5210 2840 5290
rect 2800 5200 2840 5210
rect 3120 5290 3160 5300
rect 3120 5210 3125 5290
rect 3155 5210 3160 5290
rect 3120 5200 3160 5210
rect 3440 5290 3480 5300
rect 3440 5210 3445 5290
rect 3475 5210 3480 5290
rect 3440 5200 3480 5210
rect 3760 5290 3800 5300
rect 3760 5210 3765 5290
rect 3795 5210 3800 5290
rect 3760 5200 3800 5210
rect 4080 5290 4120 5300
rect 4080 5210 4085 5290
rect 4115 5210 4120 5290
rect 4080 5200 4120 5210
rect 2800 5070 2840 5080
rect 2800 4990 2805 5070
rect 2835 4990 2840 5070
rect 2800 4980 2840 4990
rect 3120 5070 3160 5080
rect 3120 4990 3125 5070
rect 3155 4990 3160 5070
rect 3120 4980 3160 4990
rect 3440 5070 3480 5080
rect 3440 4990 3445 5070
rect 3475 4990 3480 5070
rect 3440 4980 3480 4990
rect 3760 5070 3800 5080
rect 3760 4990 3765 5070
rect 3795 4990 3800 5070
rect 3760 4980 3800 4990
rect 4080 5070 4120 5080
rect 4080 4990 4085 5070
rect 4115 4990 4120 5070
rect 4080 4980 4120 4990
rect 2880 4955 3080 4960
rect 2880 4925 2890 4955
rect 3070 4925 3080 4955
rect 2880 4920 3080 4925
rect 3200 4955 3400 4960
rect 3200 4925 3210 4955
rect 3390 4925 3400 4955
rect 3200 4920 3400 4925
rect 3520 4955 3720 4960
rect 3520 4925 3530 4955
rect 3710 4925 3720 4955
rect 3520 4920 3720 4925
rect 3840 4955 4040 4960
rect 3840 4925 3850 4955
rect 4030 4925 4040 4955
rect 3840 4920 4040 4925
rect 4240 5290 4280 5400
rect 4320 5355 4520 5360
rect 4320 5325 4330 5355
rect 4510 5325 4520 5355
rect 4320 5320 4520 5325
rect 4240 5210 4245 5290
rect 4275 5210 4280 5290
rect 4240 5070 4280 5210
rect 4240 4990 4245 5070
rect 4275 4990 4280 5070
rect 4240 4880 4280 4990
rect 4560 5290 4600 5400
rect 4560 5210 4565 5290
rect 4595 5210 4600 5290
rect 4560 5070 4600 5210
rect 4560 4990 4565 5070
rect 4595 4990 4600 5070
rect 4320 4955 4520 4960
rect 4320 4925 4330 4955
rect 4510 4925 4520 4955
rect 4320 4920 4520 4925
rect 4560 4880 4600 4990
rect -640 4840 -560 4880
rect -200 4840 -80 4880
rect 1240 4840 1360 4880
rect 2680 4840 2800 4880
rect 4120 4840 4240 4880
rect 4600 4840 4680 4880
rect -800 4680 -680 4720
rect 4760 4680 4840 4720
rect -800 4040 -560 4080
rect -200 4040 -80 4080
rect 1240 4040 1360 4080
rect 2680 4040 2800 4080
rect 4120 4040 4240 4080
rect 4600 4040 4840 4080
rect -560 3930 -520 4040
rect -480 3995 -280 4000
rect -480 3965 -470 3995
rect -290 3965 -280 3995
rect -480 3960 -280 3965
rect -560 3850 -555 3930
rect -525 3850 -520 3930
rect -560 3760 -520 3850
rect -240 3930 -200 4040
rect -240 3850 -235 3930
rect -205 3850 -200 3930
rect -240 3760 -200 3850
rect 0 3995 200 4000
rect 0 3965 10 3995
rect 190 3965 200 3995
rect 0 3960 200 3965
rect 320 3995 520 4000
rect 320 3965 330 3995
rect 510 3965 520 3995
rect 320 3960 520 3965
rect 640 3995 840 4000
rect 640 3965 650 3995
rect 830 3965 840 3995
rect 640 3960 840 3965
rect 960 3995 1160 4000
rect 960 3965 970 3995
rect 1150 3965 1160 3995
rect 960 3960 1160 3965
rect -80 3930 -40 3940
rect -80 3850 -75 3930
rect -45 3850 -40 3930
rect -80 3840 -40 3850
rect 240 3930 280 3940
rect 240 3850 245 3930
rect 275 3850 280 3930
rect 240 3840 280 3850
rect 560 3930 600 3940
rect 560 3850 565 3930
rect 595 3850 600 3930
rect 560 3840 600 3850
rect 880 3930 920 3940
rect 880 3850 885 3930
rect 915 3850 920 3930
rect 880 3840 920 3850
rect 1200 3930 1240 3940
rect 1200 3850 1205 3930
rect 1235 3850 1240 3930
rect 1200 3840 1240 3850
rect 1440 3995 1640 4000
rect 1440 3965 1450 3995
rect 1630 3965 1640 3995
rect 1440 3960 1640 3965
rect 1760 3995 1960 4000
rect 1760 3965 1770 3995
rect 1950 3965 1960 3995
rect 1760 3960 1960 3965
rect 2080 3995 2280 4000
rect 2080 3965 2090 3995
rect 2270 3965 2280 3995
rect 2080 3960 2280 3965
rect 2400 3995 2600 4000
rect 2400 3965 2410 3995
rect 2590 3965 2600 3995
rect 2400 3960 2600 3965
rect 1360 3930 1400 3940
rect 1360 3850 1365 3930
rect 1395 3850 1400 3930
rect 1360 3840 1400 3850
rect 1680 3930 1720 3940
rect 1680 3850 1685 3930
rect 1715 3850 1720 3930
rect 1680 3840 1720 3850
rect 2000 3930 2040 3940
rect 2000 3850 2005 3930
rect 2035 3850 2040 3930
rect 2000 3840 2040 3850
rect 2320 3930 2360 3940
rect 2320 3850 2325 3930
rect 2355 3850 2360 3930
rect 2320 3840 2360 3850
rect 2640 3930 2680 3940
rect 2640 3850 2645 3930
rect 2675 3850 2680 3930
rect 2640 3840 2680 3850
rect 2880 3995 3080 4000
rect 2880 3965 2890 3995
rect 3070 3965 3080 3995
rect 2880 3960 3080 3965
rect 3200 3995 3400 4000
rect 3200 3965 3210 3995
rect 3390 3965 3400 3995
rect 3200 3960 3400 3965
rect 3520 3995 3720 4000
rect 3520 3965 3530 3995
rect 3710 3965 3720 3995
rect 3520 3960 3720 3965
rect 3840 3995 4040 4000
rect 3840 3965 3850 3995
rect 4030 3965 4040 3995
rect 3840 3960 4040 3965
rect 2800 3930 2840 3940
rect 2800 3850 2805 3930
rect 2835 3850 2840 3930
rect 2800 3840 2840 3850
rect 3120 3930 3160 3940
rect 3120 3850 3125 3930
rect 3155 3850 3160 3930
rect 3120 3840 3160 3850
rect 3440 3930 3480 3940
rect 3440 3850 3445 3930
rect 3475 3850 3480 3930
rect 3440 3840 3480 3850
rect 3760 3930 3800 3940
rect 3760 3850 3765 3930
rect 3795 3850 3800 3930
rect 3760 3840 3800 3850
rect 4080 3930 4120 3940
rect 4080 3850 4085 3930
rect 4115 3850 4120 3930
rect 4080 3840 4120 3850
rect 4240 3930 4280 4040
rect 4320 3995 4520 4000
rect 4320 3965 4330 3995
rect 4510 3965 4520 3995
rect 4320 3960 4520 3965
rect 4240 3850 4245 3930
rect 4275 3850 4280 3930
rect 4240 3760 4280 3850
rect 4560 3930 4600 4040
rect 4560 3850 4565 3930
rect 4595 3850 4600 3930
rect 4560 3760 4600 3850
rect -800 3720 -560 3760
rect -200 3720 -80 3760
rect 1240 3720 1360 3760
rect 2680 3720 2800 3760
rect 4120 3720 4240 3760
rect 4600 3720 4840 3760
rect -800 3680 -760 3720
rect 4800 3680 4840 3720
rect -800 3640 -680 3680
rect 4760 3640 4840 3680
rect -640 3480 -560 3520
rect -200 3480 -80 3520
rect 1240 3480 1360 3520
rect 2680 3480 2800 3520
rect 4120 3480 4240 3520
rect 4600 3480 4680 3520
rect -560 3370 -520 3480
rect -480 3435 -280 3440
rect -480 3405 -470 3435
rect -290 3405 -280 3435
rect -480 3400 -280 3405
rect -560 3290 -555 3370
rect -525 3290 -520 3370
rect -560 3150 -520 3290
rect -560 3070 -555 3150
rect -525 3070 -520 3150
rect -560 2960 -520 3070
rect -240 3370 -200 3480
rect -240 3290 -235 3370
rect -205 3290 -200 3370
rect -240 3150 -200 3290
rect -240 3070 -235 3150
rect -205 3070 -200 3150
rect -480 3035 -280 3040
rect -480 3005 -470 3035
rect -290 3005 -280 3035
rect -480 3000 -280 3005
rect -240 2960 -200 3070
rect 0 3435 200 3440
rect 0 3405 10 3435
rect 190 3405 200 3435
rect 0 3400 200 3405
rect 320 3435 520 3440
rect 320 3405 330 3435
rect 510 3405 520 3435
rect 320 3400 520 3405
rect 640 3435 840 3440
rect 640 3405 650 3435
rect 830 3405 840 3435
rect 640 3400 840 3405
rect 960 3435 1160 3440
rect 960 3405 970 3435
rect 1150 3405 1160 3435
rect 960 3400 1160 3405
rect -80 3370 -40 3380
rect -80 3290 -75 3370
rect -45 3290 -40 3370
rect -80 3280 -40 3290
rect 240 3370 280 3380
rect 240 3290 245 3370
rect 275 3290 280 3370
rect 240 3280 280 3290
rect 560 3370 600 3380
rect 560 3290 565 3370
rect 595 3290 600 3370
rect 560 3280 600 3290
rect 880 3370 920 3380
rect 880 3290 885 3370
rect 915 3290 920 3370
rect 880 3280 920 3290
rect 1200 3370 1240 3380
rect 1200 3290 1205 3370
rect 1235 3290 1240 3370
rect 1200 3280 1240 3290
rect -80 3150 -40 3160
rect -80 3070 -75 3150
rect -45 3070 -40 3150
rect -80 3060 -40 3070
rect 240 3150 280 3160
rect 240 3070 245 3150
rect 275 3070 280 3150
rect 240 3060 280 3070
rect 560 3150 600 3160
rect 560 3070 565 3150
rect 595 3070 600 3150
rect 560 3060 600 3070
rect 880 3150 920 3160
rect 880 3070 885 3150
rect 915 3070 920 3150
rect 880 3060 920 3070
rect 1200 3150 1240 3160
rect 1200 3070 1205 3150
rect 1235 3070 1240 3150
rect 1200 3060 1240 3070
rect 0 3035 200 3040
rect 0 3005 10 3035
rect 190 3005 200 3035
rect 0 3000 200 3005
rect 320 3035 520 3040
rect 320 3005 330 3035
rect 510 3005 520 3035
rect 320 3000 520 3005
rect 640 3035 840 3040
rect 640 3005 650 3035
rect 830 3005 840 3035
rect 640 3000 840 3005
rect 960 3035 1160 3040
rect 960 3005 970 3035
rect 1150 3005 1160 3035
rect 960 3000 1160 3005
rect 1440 3435 1640 3440
rect 1440 3405 1450 3435
rect 1630 3405 1640 3435
rect 1440 3400 1640 3405
rect 1760 3435 1960 3440
rect 1760 3405 1770 3435
rect 1950 3405 1960 3435
rect 1760 3400 1960 3405
rect 2080 3435 2280 3440
rect 2080 3405 2090 3435
rect 2270 3405 2280 3435
rect 2080 3400 2280 3405
rect 2400 3435 2600 3440
rect 2400 3405 2410 3435
rect 2590 3405 2600 3435
rect 2400 3400 2600 3405
rect 1360 3370 1400 3380
rect 1360 3290 1365 3370
rect 1395 3290 1400 3370
rect 1360 3280 1400 3290
rect 1680 3370 1720 3380
rect 1680 3290 1685 3370
rect 1715 3290 1720 3370
rect 1680 3280 1720 3290
rect 2000 3370 2040 3380
rect 2000 3290 2005 3370
rect 2035 3290 2040 3370
rect 2000 3280 2040 3290
rect 2320 3370 2360 3380
rect 2320 3290 2325 3370
rect 2355 3290 2360 3370
rect 2320 3280 2360 3290
rect 2640 3370 2680 3380
rect 2640 3290 2645 3370
rect 2675 3290 2680 3370
rect 2640 3280 2680 3290
rect 1360 3150 1400 3160
rect 1360 3070 1365 3150
rect 1395 3070 1400 3150
rect 1360 3060 1400 3070
rect 1680 3150 1720 3160
rect 1680 3070 1685 3150
rect 1715 3070 1720 3150
rect 1680 3060 1720 3070
rect 2000 3150 2040 3160
rect 2000 3070 2005 3150
rect 2035 3070 2040 3150
rect 2000 3060 2040 3070
rect 2320 3150 2360 3160
rect 2320 3070 2325 3150
rect 2355 3070 2360 3150
rect 2320 3060 2360 3070
rect 2640 3150 2680 3160
rect 2640 3070 2645 3150
rect 2675 3070 2680 3150
rect 2640 3060 2680 3070
rect 1440 3035 1640 3040
rect 1440 3005 1450 3035
rect 1630 3005 1640 3035
rect 1440 3000 1640 3005
rect 1760 3035 1960 3040
rect 1760 3005 1770 3035
rect 1950 3005 1960 3035
rect 1760 3000 1960 3005
rect 2080 3035 2280 3040
rect 2080 3005 2090 3035
rect 2270 3005 2280 3035
rect 2080 3000 2280 3005
rect 2400 3035 2600 3040
rect 2400 3005 2410 3035
rect 2590 3005 2600 3035
rect 2400 3000 2600 3005
rect 2880 3435 3080 3440
rect 2880 3405 2890 3435
rect 3070 3405 3080 3435
rect 2880 3400 3080 3405
rect 3200 3435 3400 3440
rect 3200 3405 3210 3435
rect 3390 3405 3400 3435
rect 3200 3400 3400 3405
rect 3520 3435 3720 3440
rect 3520 3405 3530 3435
rect 3710 3405 3720 3435
rect 3520 3400 3720 3405
rect 3840 3435 4040 3440
rect 3840 3405 3850 3435
rect 4030 3405 4040 3435
rect 3840 3400 4040 3405
rect 2800 3370 2840 3380
rect 2800 3290 2805 3370
rect 2835 3290 2840 3370
rect 2800 3280 2840 3290
rect 3120 3370 3160 3380
rect 3120 3290 3125 3370
rect 3155 3290 3160 3370
rect 3120 3280 3160 3290
rect 3440 3370 3480 3380
rect 3440 3290 3445 3370
rect 3475 3290 3480 3370
rect 3440 3280 3480 3290
rect 3760 3370 3800 3380
rect 3760 3290 3765 3370
rect 3795 3290 3800 3370
rect 3760 3280 3800 3290
rect 4080 3370 4120 3380
rect 4080 3290 4085 3370
rect 4115 3290 4120 3370
rect 4080 3280 4120 3290
rect 2800 3150 2840 3160
rect 2800 3070 2805 3150
rect 2835 3070 2840 3150
rect 2800 3060 2840 3070
rect 3120 3150 3160 3160
rect 3120 3070 3125 3150
rect 3155 3070 3160 3150
rect 3120 3060 3160 3070
rect 3440 3150 3480 3160
rect 3440 3070 3445 3150
rect 3475 3070 3480 3150
rect 3440 3060 3480 3070
rect 3760 3150 3800 3160
rect 3760 3070 3765 3150
rect 3795 3070 3800 3150
rect 3760 3060 3800 3070
rect 4080 3150 4120 3160
rect 4080 3070 4085 3150
rect 4115 3070 4120 3150
rect 4080 3060 4120 3070
rect 2880 3035 3080 3040
rect 2880 3005 2890 3035
rect 3070 3005 3080 3035
rect 2880 3000 3080 3005
rect 3200 3035 3400 3040
rect 3200 3005 3210 3035
rect 3390 3005 3400 3035
rect 3200 3000 3400 3005
rect 3520 3035 3720 3040
rect 3520 3005 3530 3035
rect 3710 3005 3720 3035
rect 3520 3000 3720 3005
rect 3840 3035 4040 3040
rect 3840 3005 3850 3035
rect 4030 3005 4040 3035
rect 3840 3000 4040 3005
rect 4240 3370 4280 3480
rect 4320 3435 4520 3440
rect 4320 3405 4330 3435
rect 4510 3405 4520 3435
rect 4320 3400 4520 3405
rect 4240 3290 4245 3370
rect 4275 3290 4280 3370
rect 4240 3150 4280 3290
rect 4240 3070 4245 3150
rect 4275 3070 4280 3150
rect 4240 2960 4280 3070
rect 4560 3370 4600 3480
rect 4560 3290 4565 3370
rect 4595 3290 4600 3370
rect 4560 3150 4600 3290
rect 4560 3070 4565 3150
rect 4595 3070 4600 3150
rect 4320 3035 4520 3040
rect 4320 3005 4330 3035
rect 4510 3005 4520 3035
rect 4320 3000 4520 3005
rect 4560 2960 4600 3070
rect -640 2920 -560 2960
rect -200 2920 -80 2960
rect 1240 2920 1360 2960
rect 2680 2920 2800 2960
rect 4120 2920 4240 2960
rect 4600 2920 4680 2960
rect -800 2760 -680 2800
rect 4760 2760 4840 2800
rect -800 2120 -560 2160
rect -200 2120 -80 2160
rect 1240 2120 1360 2160
rect 2680 2120 2800 2160
rect 4120 2120 4240 2160
rect 4600 2120 4840 2160
rect -560 2010 -520 2120
rect -480 2075 -280 2080
rect -480 2045 -470 2075
rect -290 2045 -280 2075
rect -480 2040 -280 2045
rect -560 1930 -555 2010
rect -525 1930 -520 2010
rect -560 1840 -520 1930
rect -240 2010 -200 2120
rect -240 1930 -235 2010
rect -205 1930 -200 2010
rect -240 1840 -200 1930
rect 0 2075 200 2080
rect 0 2045 10 2075
rect 190 2045 200 2075
rect 0 2040 200 2045
rect 320 2075 520 2080
rect 320 2045 330 2075
rect 510 2045 520 2075
rect 320 2040 520 2045
rect 640 2075 840 2080
rect 640 2045 650 2075
rect 830 2045 840 2075
rect 640 2040 840 2045
rect 960 2075 1160 2080
rect 960 2045 970 2075
rect 1150 2045 1160 2075
rect 960 2040 1160 2045
rect -80 2010 -40 2020
rect -80 1930 -75 2010
rect -45 1930 -40 2010
rect -80 1920 -40 1930
rect 240 2010 280 2020
rect 240 1930 245 2010
rect 275 1930 280 2010
rect 240 1920 280 1930
rect 560 2010 600 2020
rect 560 1930 565 2010
rect 595 1930 600 2010
rect 560 1920 600 1930
rect 880 2010 920 2020
rect 880 1930 885 2010
rect 915 1930 920 2010
rect 880 1920 920 1930
rect 1200 2010 1240 2020
rect 1200 1930 1205 2010
rect 1235 1930 1240 2010
rect 1200 1920 1240 1930
rect 1440 2075 1640 2080
rect 1440 2045 1450 2075
rect 1630 2045 1640 2075
rect 1440 2040 1640 2045
rect 1760 2075 1960 2080
rect 1760 2045 1770 2075
rect 1950 2045 1960 2075
rect 1760 2040 1960 2045
rect 2080 2075 2280 2080
rect 2080 2045 2090 2075
rect 2270 2045 2280 2075
rect 2080 2040 2280 2045
rect 2400 2075 2600 2080
rect 2400 2045 2410 2075
rect 2590 2045 2600 2075
rect 2400 2040 2600 2045
rect 1360 2010 1400 2020
rect 1360 1930 1365 2010
rect 1395 1930 1400 2010
rect 1360 1920 1400 1930
rect 1680 2010 1720 2020
rect 1680 1930 1685 2010
rect 1715 1930 1720 2010
rect 1680 1920 1720 1930
rect 2000 2010 2040 2020
rect 2000 1930 2005 2010
rect 2035 1930 2040 2010
rect 2000 1920 2040 1930
rect 2320 2010 2360 2020
rect 2320 1930 2325 2010
rect 2355 1930 2360 2010
rect 2320 1920 2360 1930
rect 2640 2010 2680 2020
rect 2640 1930 2645 2010
rect 2675 1930 2680 2010
rect 2640 1920 2680 1930
rect 2880 2075 3080 2080
rect 2880 2045 2890 2075
rect 3070 2045 3080 2075
rect 2880 2040 3080 2045
rect 3200 2075 3400 2080
rect 3200 2045 3210 2075
rect 3390 2045 3400 2075
rect 3200 2040 3400 2045
rect 3520 2075 3720 2080
rect 3520 2045 3530 2075
rect 3710 2045 3720 2075
rect 3520 2040 3720 2045
rect 3840 2075 4040 2080
rect 3840 2045 3850 2075
rect 4030 2045 4040 2075
rect 3840 2040 4040 2045
rect 2800 2010 2840 2020
rect 2800 1930 2805 2010
rect 2835 1930 2840 2010
rect 2800 1920 2840 1930
rect 3120 2010 3160 2020
rect 3120 1930 3125 2010
rect 3155 1930 3160 2010
rect 3120 1920 3160 1930
rect 3440 2010 3480 2020
rect 3440 1930 3445 2010
rect 3475 1930 3480 2010
rect 3440 1920 3480 1930
rect 3760 2010 3800 2020
rect 3760 1930 3765 2010
rect 3795 1930 3800 2010
rect 3760 1920 3800 1930
rect 4080 2010 4120 2020
rect 4080 1930 4085 2010
rect 4115 1930 4120 2010
rect 4080 1920 4120 1930
rect 4240 2010 4280 2120
rect 4320 2075 4520 2080
rect 4320 2045 4330 2075
rect 4510 2045 4520 2075
rect 4320 2040 4520 2045
rect 4240 1930 4245 2010
rect 4275 1930 4280 2010
rect 4240 1840 4280 1930
rect 4560 2010 4600 2120
rect 4560 1930 4565 2010
rect 4595 1930 4600 2010
rect 4560 1840 4600 1930
rect -800 1800 -560 1840
rect -200 1800 -80 1840
rect 1240 1800 1360 1840
rect 2680 1800 2800 1840
rect 4120 1800 4240 1840
rect 4600 1800 4840 1840
rect -800 1760 -760 1800
rect 4800 1760 4840 1800
rect -800 1720 -680 1760
rect 4760 1720 4840 1760
rect -640 1560 -560 1600
rect -200 1560 -80 1600
rect 1240 1560 1360 1600
rect 2680 1560 2800 1600
rect 4120 1560 4240 1600
rect 4600 1560 4680 1600
rect -560 1450 -520 1560
rect -480 1515 -280 1520
rect -480 1485 -470 1515
rect -290 1485 -280 1515
rect -480 1480 -280 1485
rect -560 1370 -555 1450
rect -525 1370 -520 1450
rect -560 1230 -520 1370
rect -560 1150 -555 1230
rect -525 1150 -520 1230
rect -560 1040 -520 1150
rect -240 1450 -200 1560
rect -240 1370 -235 1450
rect -205 1370 -200 1450
rect -240 1230 -200 1370
rect -240 1150 -235 1230
rect -205 1150 -200 1230
rect -480 1115 -280 1120
rect -480 1085 -470 1115
rect -290 1085 -280 1115
rect -480 1080 -280 1085
rect -240 1040 -200 1150
rect 0 1515 200 1520
rect 0 1485 10 1515
rect 190 1485 200 1515
rect 0 1480 200 1485
rect 320 1515 520 1520
rect 320 1485 330 1515
rect 510 1485 520 1515
rect 320 1480 520 1485
rect 640 1515 840 1520
rect 640 1485 650 1515
rect 830 1485 840 1515
rect 640 1480 840 1485
rect 960 1515 1160 1520
rect 960 1485 970 1515
rect 1150 1485 1160 1515
rect 960 1480 1160 1485
rect -80 1450 -40 1460
rect -80 1370 -75 1450
rect -45 1370 -40 1450
rect -80 1360 -40 1370
rect 240 1450 280 1460
rect 240 1370 245 1450
rect 275 1370 280 1450
rect 240 1360 280 1370
rect 560 1450 600 1460
rect 560 1370 565 1450
rect 595 1370 600 1450
rect 560 1360 600 1370
rect 880 1450 920 1460
rect 880 1370 885 1450
rect 915 1370 920 1450
rect 880 1360 920 1370
rect 1200 1450 1240 1460
rect 1200 1370 1205 1450
rect 1235 1370 1240 1450
rect 1200 1360 1240 1370
rect -80 1230 -40 1240
rect -80 1150 -75 1230
rect -45 1150 -40 1230
rect -80 1140 -40 1150
rect 240 1230 280 1240
rect 240 1150 245 1230
rect 275 1150 280 1230
rect 240 1140 280 1150
rect 560 1230 600 1240
rect 560 1150 565 1230
rect 595 1150 600 1230
rect 560 1140 600 1150
rect 880 1230 920 1240
rect 880 1150 885 1230
rect 915 1150 920 1230
rect 880 1140 920 1150
rect 1200 1230 1240 1240
rect 1200 1150 1205 1230
rect 1235 1150 1240 1230
rect 1200 1140 1240 1150
rect 0 1115 200 1120
rect 0 1085 10 1115
rect 190 1085 200 1115
rect 0 1080 200 1085
rect 320 1115 520 1120
rect 320 1085 330 1115
rect 510 1085 520 1115
rect 320 1080 520 1085
rect 640 1115 840 1120
rect 640 1085 650 1115
rect 830 1085 840 1115
rect 640 1080 840 1085
rect 960 1115 1160 1120
rect 960 1085 970 1115
rect 1150 1085 1160 1115
rect 960 1080 1160 1085
rect 1440 1515 1640 1520
rect 1440 1485 1450 1515
rect 1630 1485 1640 1515
rect 1440 1480 1640 1485
rect 1760 1515 1960 1520
rect 1760 1485 1770 1515
rect 1950 1485 1960 1515
rect 1760 1480 1960 1485
rect 2080 1515 2280 1520
rect 2080 1485 2090 1515
rect 2270 1485 2280 1515
rect 2080 1480 2280 1485
rect 2400 1515 2600 1520
rect 2400 1485 2410 1515
rect 2590 1485 2600 1515
rect 2400 1480 2600 1485
rect 1360 1450 1400 1460
rect 1360 1370 1365 1450
rect 1395 1370 1400 1450
rect 1360 1360 1400 1370
rect 1680 1450 1720 1460
rect 1680 1370 1685 1450
rect 1715 1370 1720 1450
rect 1680 1360 1720 1370
rect 2000 1450 2040 1460
rect 2000 1370 2005 1450
rect 2035 1370 2040 1450
rect 2000 1360 2040 1370
rect 2320 1450 2360 1460
rect 2320 1370 2325 1450
rect 2355 1370 2360 1450
rect 2320 1360 2360 1370
rect 2640 1450 2680 1460
rect 2640 1370 2645 1450
rect 2675 1370 2680 1450
rect 2640 1360 2680 1370
rect 1360 1230 1400 1240
rect 1360 1150 1365 1230
rect 1395 1150 1400 1230
rect 1360 1140 1400 1150
rect 1680 1230 1720 1240
rect 1680 1150 1685 1230
rect 1715 1150 1720 1230
rect 1680 1140 1720 1150
rect 2000 1230 2040 1240
rect 2000 1150 2005 1230
rect 2035 1150 2040 1230
rect 2000 1140 2040 1150
rect 2320 1230 2360 1240
rect 2320 1150 2325 1230
rect 2355 1150 2360 1230
rect 2320 1140 2360 1150
rect 2640 1230 2680 1240
rect 2640 1150 2645 1230
rect 2675 1150 2680 1230
rect 2640 1140 2680 1150
rect 1440 1115 1640 1120
rect 1440 1085 1450 1115
rect 1630 1085 1640 1115
rect 1440 1080 1640 1085
rect 1760 1115 1960 1120
rect 1760 1085 1770 1115
rect 1950 1085 1960 1115
rect 1760 1080 1960 1085
rect 2080 1115 2280 1120
rect 2080 1085 2090 1115
rect 2270 1085 2280 1115
rect 2080 1080 2280 1085
rect 2400 1115 2600 1120
rect 2400 1085 2410 1115
rect 2590 1085 2600 1115
rect 2400 1080 2600 1085
rect 2880 1515 3080 1520
rect 2880 1485 2890 1515
rect 3070 1485 3080 1515
rect 2880 1480 3080 1485
rect 3200 1515 3400 1520
rect 3200 1485 3210 1515
rect 3390 1485 3400 1515
rect 3200 1480 3400 1485
rect 3520 1515 3720 1520
rect 3520 1485 3530 1515
rect 3710 1485 3720 1515
rect 3520 1480 3720 1485
rect 3840 1515 4040 1520
rect 3840 1485 3850 1515
rect 4030 1485 4040 1515
rect 3840 1480 4040 1485
rect 2800 1450 2840 1460
rect 2800 1370 2805 1450
rect 2835 1370 2840 1450
rect 2800 1360 2840 1370
rect 3120 1450 3160 1460
rect 3120 1370 3125 1450
rect 3155 1370 3160 1450
rect 3120 1360 3160 1370
rect 3440 1450 3480 1460
rect 3440 1370 3445 1450
rect 3475 1370 3480 1450
rect 3440 1360 3480 1370
rect 3760 1450 3800 1460
rect 3760 1370 3765 1450
rect 3795 1370 3800 1450
rect 3760 1360 3800 1370
rect 4080 1450 4120 1460
rect 4080 1370 4085 1450
rect 4115 1370 4120 1450
rect 4080 1360 4120 1370
rect 2800 1230 2840 1240
rect 2800 1150 2805 1230
rect 2835 1150 2840 1230
rect 2800 1140 2840 1150
rect 3120 1230 3160 1240
rect 3120 1150 3125 1230
rect 3155 1150 3160 1230
rect 3120 1140 3160 1150
rect 3440 1230 3480 1240
rect 3440 1150 3445 1230
rect 3475 1150 3480 1230
rect 3440 1140 3480 1150
rect 3760 1230 3800 1240
rect 3760 1150 3765 1230
rect 3795 1150 3800 1230
rect 3760 1140 3800 1150
rect 4080 1230 4120 1240
rect 4080 1150 4085 1230
rect 4115 1150 4120 1230
rect 4080 1140 4120 1150
rect 2880 1115 3080 1120
rect 2880 1085 2890 1115
rect 3070 1085 3080 1115
rect 2880 1080 3080 1085
rect 3200 1115 3400 1120
rect 3200 1085 3210 1115
rect 3390 1085 3400 1115
rect 3200 1080 3400 1085
rect 3520 1115 3720 1120
rect 3520 1085 3530 1115
rect 3710 1085 3720 1115
rect 3520 1080 3720 1085
rect 3840 1115 4040 1120
rect 3840 1085 3850 1115
rect 4030 1085 4040 1115
rect 3840 1080 4040 1085
rect 4240 1450 4280 1560
rect 4320 1515 4520 1520
rect 4320 1485 4330 1515
rect 4510 1485 4520 1515
rect 4320 1480 4520 1485
rect 4240 1370 4245 1450
rect 4275 1370 4280 1450
rect 4240 1230 4280 1370
rect 4240 1150 4245 1230
rect 4275 1150 4280 1230
rect 4240 1040 4280 1150
rect 4560 1450 4600 1560
rect 4560 1370 4565 1450
rect 4595 1370 4600 1450
rect 4560 1230 4600 1370
rect 4560 1150 4565 1230
rect 4595 1150 4600 1230
rect 4320 1115 4520 1120
rect 4320 1085 4330 1115
rect 4510 1085 4520 1115
rect 4320 1080 4520 1085
rect 4560 1040 4600 1150
rect -640 1000 -560 1040
rect -200 1000 -80 1040
rect 1240 1000 1360 1040
rect 2680 1000 2800 1040
rect 4120 1000 4240 1040
rect 4600 1000 4680 1040
rect -800 840 -680 880
rect 4760 840 4840 880
rect -800 200 -560 240
rect -200 200 -80 240
rect 1240 200 1360 240
rect 2680 200 2800 240
rect 4120 200 4240 240
rect 4600 200 4840 240
rect -560 90 -520 200
rect -480 155 -280 160
rect -480 125 -470 155
rect -290 125 -280 155
rect -480 120 -280 125
rect -560 10 -555 90
rect -525 10 -520 90
rect -560 -80 -520 10
rect -240 90 -200 200
rect -240 10 -235 90
rect -205 10 -200 90
rect -240 -80 -200 10
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 120 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 120 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 120 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 120 1160 125
rect -80 90 -40 100
rect -80 10 -75 90
rect -45 10 -40 90
rect -80 0 -40 10
rect 240 90 280 100
rect 240 10 245 90
rect 275 10 280 90
rect 240 0 280 10
rect 560 90 600 100
rect 560 10 565 90
rect 595 10 600 90
rect 560 0 600 10
rect 880 90 920 100
rect 880 10 885 90
rect 915 10 920 90
rect 880 0 920 10
rect 1200 90 1240 100
rect 1200 10 1205 90
rect 1235 10 1240 90
rect 1200 0 1240 10
rect 1440 155 1640 160
rect 1440 125 1450 155
rect 1630 125 1640 155
rect 1440 120 1640 125
rect 1760 155 1960 160
rect 1760 125 1770 155
rect 1950 125 1960 155
rect 1760 120 1960 125
rect 2080 155 2280 160
rect 2080 125 2090 155
rect 2270 125 2280 155
rect 2080 120 2280 125
rect 2400 155 2600 160
rect 2400 125 2410 155
rect 2590 125 2600 155
rect 2400 120 2600 125
rect 1360 90 1400 100
rect 1360 10 1365 90
rect 1395 10 1400 90
rect 1360 0 1400 10
rect 1680 90 1720 100
rect 1680 10 1685 90
rect 1715 10 1720 90
rect 1680 0 1720 10
rect 2000 90 2040 100
rect 2000 10 2005 90
rect 2035 10 2040 90
rect 2000 0 2040 10
rect 2320 90 2360 100
rect 2320 10 2325 90
rect 2355 10 2360 90
rect 2320 0 2360 10
rect 2640 90 2680 100
rect 2640 10 2645 90
rect 2675 10 2680 90
rect 2640 0 2680 10
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 120 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 120 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 120 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 120 4040 125
rect 2800 90 2840 100
rect 2800 10 2805 90
rect 2835 10 2840 90
rect 2800 0 2840 10
rect 3120 90 3160 100
rect 3120 10 3125 90
rect 3155 10 3160 90
rect 3120 0 3160 10
rect 3440 90 3480 100
rect 3440 10 3445 90
rect 3475 10 3480 90
rect 3440 0 3480 10
rect 3760 90 3800 100
rect 3760 10 3765 90
rect 3795 10 3800 90
rect 3760 0 3800 10
rect 4080 90 4120 100
rect 4080 10 4085 90
rect 4115 10 4120 90
rect 4080 0 4120 10
rect 4240 90 4280 200
rect 4320 155 4520 160
rect 4320 125 4330 155
rect 4510 125 4520 155
rect 4320 120 4520 125
rect 4240 10 4245 90
rect 4275 10 4280 90
rect 4240 -80 4280 10
rect 4560 90 4600 200
rect 4560 10 4565 90
rect 4595 10 4600 90
rect 4560 -80 4600 10
rect -800 -120 -560 -80
rect -200 -120 -80 -80
rect 1240 -120 1360 -80
rect 2680 -120 2800 -80
rect 4120 -120 4240 -80
rect 4600 -120 4840 -80
<< viali >>
rect -470 5325 -290 5355
rect -555 5210 -525 5290
rect -555 4990 -525 5070
rect -235 5210 -205 5290
rect -235 4990 -205 5070
rect -470 4925 -290 4955
rect 10 5325 190 5355
rect 330 5325 510 5355
rect 650 5325 830 5355
rect 970 5325 1150 5355
rect -75 5210 -45 5290
rect 245 5210 275 5290
rect 565 5210 595 5290
rect 885 5210 915 5290
rect 1205 5210 1235 5290
rect -75 4990 -45 5070
rect 245 4990 275 5070
rect 565 4990 595 5070
rect 885 4990 915 5070
rect 1205 4990 1235 5070
rect 10 4925 190 4955
rect 330 4925 510 4955
rect 650 4925 830 4955
rect 970 4925 1150 4955
rect 1450 5325 1630 5355
rect 1770 5325 1950 5355
rect 2090 5325 2270 5355
rect 2410 5325 2590 5355
rect 1365 5210 1395 5290
rect 1685 5210 1715 5290
rect 2005 5210 2035 5290
rect 2325 5210 2355 5290
rect 2645 5210 2675 5290
rect 1365 4990 1395 5070
rect 1685 4990 1715 5070
rect 2005 4990 2035 5070
rect 2325 4990 2355 5070
rect 2645 4990 2675 5070
rect 1450 4925 1630 4955
rect 1770 4925 1950 4955
rect 2090 4925 2270 4955
rect 2410 4925 2590 4955
rect 2890 5325 3070 5355
rect 3210 5325 3390 5355
rect 3530 5325 3710 5355
rect 3850 5325 4030 5355
rect 2805 5210 2835 5290
rect 3125 5210 3155 5290
rect 3445 5210 3475 5290
rect 3765 5210 3795 5290
rect 4085 5210 4115 5290
rect 2805 4990 2835 5070
rect 3125 4990 3155 5070
rect 3445 4990 3475 5070
rect 3765 4990 3795 5070
rect 4085 4990 4115 5070
rect 2890 4925 3070 4955
rect 3210 4925 3390 4955
rect 3530 4925 3710 4955
rect 3850 4925 4030 4955
rect 4330 5325 4510 5355
rect 4245 5210 4275 5290
rect 4245 4990 4275 5070
rect 4565 5210 4595 5290
rect 4565 4990 4595 5070
rect 4330 4925 4510 4955
rect -470 3965 -290 3995
rect -555 3850 -525 3930
rect -235 3850 -205 3930
rect 10 3965 190 3995
rect 330 3965 510 3995
rect 650 3965 830 3995
rect 970 3965 1150 3995
rect -75 3850 -45 3930
rect 245 3850 275 3930
rect 565 3850 595 3930
rect 885 3850 915 3930
rect 1205 3850 1235 3930
rect 1450 3965 1630 3995
rect 1770 3965 1950 3995
rect 2090 3965 2270 3995
rect 2410 3965 2590 3995
rect 1365 3850 1395 3930
rect 1685 3850 1715 3930
rect 2005 3850 2035 3930
rect 2325 3850 2355 3930
rect 2645 3850 2675 3930
rect 2890 3965 3070 3995
rect 3210 3965 3390 3995
rect 3530 3965 3710 3995
rect 3850 3965 4030 3995
rect 2805 3850 2835 3930
rect 3125 3850 3155 3930
rect 3445 3850 3475 3930
rect 3765 3850 3795 3930
rect 4085 3850 4115 3930
rect 4330 3965 4510 3995
rect 4245 3850 4275 3930
rect 4565 3850 4595 3930
rect -470 3405 -290 3435
rect -555 3290 -525 3370
rect -555 3070 -525 3150
rect -235 3290 -205 3370
rect -235 3070 -205 3150
rect -470 3005 -290 3035
rect 10 3405 190 3435
rect 330 3405 510 3435
rect 650 3405 830 3435
rect 970 3405 1150 3435
rect -75 3290 -45 3370
rect 245 3290 275 3370
rect 565 3290 595 3370
rect 885 3290 915 3370
rect 1205 3290 1235 3370
rect -75 3070 -45 3150
rect 245 3070 275 3150
rect 565 3070 595 3150
rect 885 3070 915 3150
rect 1205 3070 1235 3150
rect 10 3005 190 3035
rect 330 3005 510 3035
rect 650 3005 830 3035
rect 970 3005 1150 3035
rect 1450 3405 1630 3435
rect 1770 3405 1950 3435
rect 2090 3405 2270 3435
rect 2410 3405 2590 3435
rect 1365 3290 1395 3370
rect 1685 3290 1715 3370
rect 2005 3290 2035 3370
rect 2325 3290 2355 3370
rect 2645 3290 2675 3370
rect 1365 3070 1395 3150
rect 1685 3070 1715 3150
rect 2005 3070 2035 3150
rect 2325 3070 2355 3150
rect 2645 3070 2675 3150
rect 1450 3005 1630 3035
rect 1770 3005 1950 3035
rect 2090 3005 2270 3035
rect 2410 3005 2590 3035
rect 2890 3405 3070 3435
rect 3210 3405 3390 3435
rect 3530 3405 3710 3435
rect 3850 3405 4030 3435
rect 2805 3290 2835 3370
rect 3125 3290 3155 3370
rect 3445 3290 3475 3370
rect 3765 3290 3795 3370
rect 4085 3290 4115 3370
rect 2805 3070 2835 3150
rect 3125 3070 3155 3150
rect 3445 3070 3475 3150
rect 3765 3070 3795 3150
rect 4085 3070 4115 3150
rect 2890 3005 3070 3035
rect 3210 3005 3390 3035
rect 3530 3005 3710 3035
rect 3850 3005 4030 3035
rect 4330 3405 4510 3435
rect 4245 3290 4275 3370
rect 4245 3070 4275 3150
rect 4565 3290 4595 3370
rect 4565 3070 4595 3150
rect 4330 3005 4510 3035
rect -470 2045 -290 2075
rect -555 1930 -525 2010
rect -235 1930 -205 2010
rect 10 2045 190 2075
rect 330 2045 510 2075
rect 650 2045 830 2075
rect 970 2045 1150 2075
rect -75 1930 -45 2010
rect 245 1930 275 2010
rect 565 1930 595 2010
rect 885 1930 915 2010
rect 1205 1930 1235 2010
rect 1450 2045 1630 2075
rect 1770 2045 1950 2075
rect 2090 2045 2270 2075
rect 2410 2045 2590 2075
rect 1365 1930 1395 2010
rect 1685 1930 1715 2010
rect 2005 1930 2035 2010
rect 2325 1930 2355 2010
rect 2645 1930 2675 2010
rect 2890 2045 3070 2075
rect 3210 2045 3390 2075
rect 3530 2045 3710 2075
rect 3850 2045 4030 2075
rect 2805 1930 2835 2010
rect 3125 1930 3155 2010
rect 3445 1930 3475 2010
rect 3765 1930 3795 2010
rect 4085 1930 4115 2010
rect 4330 2045 4510 2075
rect 4245 1930 4275 2010
rect 4565 1930 4595 2010
rect -470 1485 -290 1515
rect -555 1370 -525 1450
rect -555 1150 -525 1230
rect -235 1370 -205 1450
rect -235 1150 -205 1230
rect -470 1085 -290 1115
rect 10 1485 190 1515
rect 330 1485 510 1515
rect 650 1485 830 1515
rect 970 1485 1150 1515
rect -75 1370 -45 1450
rect 245 1370 275 1450
rect 565 1370 595 1450
rect 885 1370 915 1450
rect 1205 1370 1235 1450
rect -75 1150 -45 1230
rect 245 1150 275 1230
rect 565 1150 595 1230
rect 885 1150 915 1230
rect 1205 1150 1235 1230
rect 10 1085 190 1115
rect 330 1085 510 1115
rect 650 1085 830 1115
rect 970 1085 1150 1115
rect 1450 1485 1630 1515
rect 1770 1485 1950 1515
rect 2090 1485 2270 1515
rect 2410 1485 2590 1515
rect 1365 1370 1395 1450
rect 1685 1370 1715 1450
rect 2005 1370 2035 1450
rect 2325 1370 2355 1450
rect 2645 1370 2675 1450
rect 1365 1150 1395 1230
rect 1685 1150 1715 1230
rect 2005 1150 2035 1230
rect 2325 1150 2355 1230
rect 2645 1150 2675 1230
rect 1450 1085 1630 1115
rect 1770 1085 1950 1115
rect 2090 1085 2270 1115
rect 2410 1085 2590 1115
rect 2890 1485 3070 1515
rect 3210 1485 3390 1515
rect 3530 1485 3710 1515
rect 3850 1485 4030 1515
rect 2805 1370 2835 1450
rect 3125 1370 3155 1450
rect 3445 1370 3475 1450
rect 3765 1370 3795 1450
rect 4085 1370 4115 1450
rect 2805 1150 2835 1230
rect 3125 1150 3155 1230
rect 3445 1150 3475 1230
rect 3765 1150 3795 1230
rect 4085 1150 4115 1230
rect 2890 1085 3070 1115
rect 3210 1085 3390 1115
rect 3530 1085 3710 1115
rect 3850 1085 4030 1115
rect 4330 1485 4510 1515
rect 4245 1370 4275 1450
rect 4245 1150 4275 1230
rect 4565 1370 4595 1450
rect 4565 1150 4595 1230
rect 4330 1085 4510 1115
rect -470 125 -290 155
rect -555 10 -525 90
rect -235 10 -205 90
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect -75 10 -45 90
rect 245 10 275 90
rect 565 10 595 90
rect 885 10 915 90
rect 1205 10 1235 90
rect 1450 125 1630 155
rect 1770 125 1950 155
rect 2090 125 2270 155
rect 2410 125 2590 155
rect 1365 10 1395 90
rect 1685 10 1715 90
rect 2005 10 2035 90
rect 2325 10 2355 90
rect 2645 10 2675 90
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3850 125 4030 155
rect 2805 10 2835 90
rect 3125 10 3155 90
rect 3445 10 3475 90
rect 3765 10 3795 90
rect 4085 10 4115 90
rect 4330 125 4510 155
rect 4245 10 4275 90
rect 4565 10 4595 90
<< metal1 >>
rect -800 5595 -760 5600
rect -800 5565 -795 5595
rect -765 5565 -760 5595
rect -800 5560 -760 5565
rect -480 5355 -280 5360
rect -480 5325 -470 5355
rect -290 5325 -280 5355
rect -480 5320 -280 5325
rect 0 5355 200 5360
rect 0 5325 10 5355
rect 190 5325 200 5355
rect 0 5320 200 5325
rect 320 5355 520 5360
rect 320 5325 330 5355
rect 510 5325 520 5355
rect 320 5320 520 5325
rect 640 5355 840 5360
rect 640 5325 650 5355
rect 830 5325 840 5355
rect 640 5320 840 5325
rect 960 5355 1160 5360
rect 960 5325 970 5355
rect 1150 5325 1160 5355
rect 960 5320 1160 5325
rect 1440 5355 1640 5360
rect 1440 5325 1450 5355
rect 1630 5325 1640 5355
rect 1440 5320 1640 5325
rect 1760 5355 1960 5360
rect 1760 5325 1770 5355
rect 1950 5325 1960 5355
rect 1760 5320 1960 5325
rect 2080 5355 2280 5360
rect 2080 5325 2090 5355
rect 2270 5325 2280 5355
rect 2080 5320 2280 5325
rect 2400 5355 2600 5360
rect 2400 5325 2410 5355
rect 2590 5325 2600 5355
rect 2400 5320 2600 5325
rect 2880 5355 3080 5360
rect 2880 5325 2890 5355
rect 3070 5325 3080 5355
rect 2880 5320 3080 5325
rect 3200 5355 3400 5360
rect 3200 5325 3210 5355
rect 3390 5325 3400 5355
rect 3200 5320 3400 5325
rect 3520 5355 3720 5360
rect 3520 5325 3530 5355
rect 3710 5325 3720 5355
rect 3520 5320 3720 5325
rect 3840 5355 4040 5360
rect 3840 5325 3850 5355
rect 4030 5325 4040 5355
rect 3840 5320 4040 5325
rect 4320 5355 4520 5360
rect 4320 5325 4330 5355
rect 4510 5325 4520 5355
rect 4320 5320 4520 5325
rect -560 5290 -520 5300
rect -560 5210 -555 5290
rect -525 5210 -520 5290
rect -560 5195 -520 5210
rect -560 5165 -555 5195
rect -525 5165 -520 5195
rect -560 5115 -520 5165
rect -560 5085 -555 5115
rect -525 5085 -520 5115
rect -560 5070 -520 5085
rect -560 4990 -555 5070
rect -525 4990 -520 5070
rect -560 4980 -520 4990
rect -240 5290 -200 5300
rect -240 5210 -235 5290
rect -205 5210 -200 5290
rect -240 5195 -200 5210
rect -240 5165 -235 5195
rect -205 5165 -200 5195
rect -240 5115 -200 5165
rect -240 5085 -235 5115
rect -205 5085 -200 5115
rect -240 5070 -200 5085
rect -240 4990 -235 5070
rect -205 4990 -200 5070
rect -240 4980 -200 4990
rect -80 5290 -40 5300
rect -80 5210 -75 5290
rect -45 5210 -40 5290
rect -80 5070 -40 5210
rect 240 5290 280 5300
rect 240 5210 245 5290
rect 275 5210 280 5290
rect 240 5200 280 5210
rect 560 5290 600 5300
rect 560 5210 565 5290
rect 595 5210 600 5290
rect 560 5195 600 5210
rect 880 5290 920 5300
rect 880 5210 885 5290
rect 915 5210 920 5290
rect 880 5200 920 5210
rect 1200 5290 1240 5300
rect 1200 5210 1205 5290
rect 1235 5210 1240 5290
rect 560 5165 565 5195
rect 595 5165 600 5195
rect 560 5160 600 5165
rect -80 4990 -75 5070
rect -45 4990 -40 5070
rect -80 4980 -40 4990
rect 240 5070 280 5080
rect 240 4990 245 5070
rect 275 4990 280 5070
rect 240 4980 280 4990
rect 560 5070 600 5080
rect 560 4990 565 5070
rect 595 4990 600 5070
rect -480 4955 -280 4960
rect -480 4925 -470 4955
rect -290 4925 -280 4955
rect -480 4920 -280 4925
rect 0 4955 200 4960
rect 0 4925 10 4955
rect 190 4925 200 4955
rect 0 4920 200 4925
rect 320 4955 520 4960
rect 320 4925 330 4955
rect 510 4925 520 4955
rect 320 4920 520 4925
rect 80 4795 120 4800
rect 80 4765 85 4795
rect 115 4765 120 4795
rect -400 4155 -360 4160
rect -400 4125 -395 4155
rect -365 4125 -360 4155
rect -800 4075 -760 4080
rect -800 4045 -795 4075
rect -765 4045 -760 4075
rect -800 3915 -760 4045
rect -400 4000 -360 4125
rect -80 4155 -40 4160
rect -80 4125 -75 4155
rect -45 4125 -40 4155
rect -480 3995 -280 4000
rect -480 3965 -470 3995
rect -290 3965 -280 3995
rect -480 3960 -280 3965
rect -800 3885 -795 3915
rect -765 3885 -760 3915
rect -800 3835 -760 3885
rect -800 3805 -795 3835
rect -765 3805 -760 3835
rect -800 3755 -760 3805
rect -560 3930 -520 3940
rect -560 3850 -555 3930
rect -525 3850 -520 3930
rect -560 3835 -520 3850
rect -560 3805 -555 3835
rect -525 3805 -520 3835
rect -560 3800 -520 3805
rect -240 3930 -200 3940
rect -240 3850 -235 3930
rect -205 3850 -200 3930
rect -240 3835 -200 3850
rect -240 3805 -235 3835
rect -205 3805 -200 3835
rect -240 3800 -200 3805
rect -160 3915 -120 4000
rect -160 3885 -155 3915
rect -125 3885 -120 3915
rect -160 3835 -120 3885
rect -80 3930 -40 4125
rect 80 4000 120 4765
rect 400 4795 440 4800
rect 400 4765 405 4795
rect 435 4765 440 4795
rect 240 4555 280 4560
rect 240 4525 245 4555
rect 275 4525 280 4555
rect 0 3995 200 4000
rect 0 3965 10 3995
rect 190 3965 200 3995
rect 0 3960 200 3965
rect -80 3850 -75 3930
rect -45 3850 -40 3930
rect -80 3840 -40 3850
rect 240 3930 280 4525
rect 400 4000 440 4765
rect 560 4315 600 4990
rect 880 5070 920 5080
rect 880 4990 885 5070
rect 915 4990 920 5070
rect 880 4980 920 4990
rect 1200 5070 1240 5210
rect 1200 4990 1205 5070
rect 1235 4990 1240 5070
rect 1200 4980 1240 4990
rect 1360 5290 1400 5300
rect 1360 5210 1365 5290
rect 1395 5210 1400 5290
rect 1360 5195 1400 5210
rect 1360 5165 1365 5195
rect 1395 5165 1400 5195
rect 1360 5115 1400 5165
rect 1360 5085 1365 5115
rect 1395 5085 1400 5115
rect 1360 5070 1400 5085
rect 1360 4990 1365 5070
rect 1395 4990 1400 5070
rect 1360 4980 1400 4990
rect 1680 5290 1720 5300
rect 1680 5210 1685 5290
rect 1715 5210 1720 5290
rect 1680 5195 1720 5210
rect 1680 5165 1685 5195
rect 1715 5165 1720 5195
rect 1680 5115 1720 5165
rect 1680 5085 1685 5115
rect 1715 5085 1720 5115
rect 1680 5070 1720 5085
rect 1680 4990 1685 5070
rect 1715 4990 1720 5070
rect 1680 4980 1720 4990
rect 2000 5290 2040 5300
rect 2000 5210 2005 5290
rect 2035 5210 2040 5290
rect 2000 5195 2040 5210
rect 2000 5165 2005 5195
rect 2035 5165 2040 5195
rect 2000 5115 2040 5165
rect 2000 5085 2005 5115
rect 2035 5085 2040 5115
rect 2000 5070 2040 5085
rect 2000 4990 2005 5070
rect 2035 4990 2040 5070
rect 2000 4980 2040 4990
rect 2320 5290 2360 5300
rect 2320 5210 2325 5290
rect 2355 5210 2360 5290
rect 2320 5195 2360 5210
rect 2320 5165 2325 5195
rect 2355 5165 2360 5195
rect 2320 5115 2360 5165
rect 2320 5085 2325 5115
rect 2355 5085 2360 5115
rect 2320 5070 2360 5085
rect 2320 4990 2325 5070
rect 2355 4990 2360 5070
rect 2320 4980 2360 4990
rect 2640 5290 2680 5300
rect 2640 5210 2645 5290
rect 2675 5210 2680 5290
rect 2640 5195 2680 5210
rect 2640 5165 2645 5195
rect 2675 5165 2680 5195
rect 2640 5115 2680 5165
rect 2640 5085 2645 5115
rect 2675 5085 2680 5115
rect 2640 5070 2680 5085
rect 2640 4990 2645 5070
rect 2675 4990 2680 5070
rect 2640 4980 2680 4990
rect 2800 5290 2840 5300
rect 2800 5210 2805 5290
rect 2835 5210 2840 5290
rect 2800 5195 2840 5210
rect 2800 5165 2805 5195
rect 2835 5165 2840 5195
rect 2800 5115 2840 5165
rect 2800 5085 2805 5115
rect 2835 5085 2840 5115
rect 2800 5070 2840 5085
rect 2800 4990 2805 5070
rect 2835 4990 2840 5070
rect 2800 4980 2840 4990
rect 3120 5290 3160 5300
rect 3120 5210 3125 5290
rect 3155 5210 3160 5290
rect 3120 5195 3160 5210
rect 3120 5165 3125 5195
rect 3155 5165 3160 5195
rect 3120 5115 3160 5165
rect 3120 5085 3125 5115
rect 3155 5085 3160 5115
rect 3120 5070 3160 5085
rect 3120 4990 3125 5070
rect 3155 4990 3160 5070
rect 3120 4980 3160 4990
rect 3440 5290 3480 5300
rect 3440 5210 3445 5290
rect 3475 5210 3480 5290
rect 3440 5195 3480 5210
rect 3440 5165 3445 5195
rect 3475 5165 3480 5195
rect 3440 5115 3480 5165
rect 3440 5085 3445 5115
rect 3475 5085 3480 5115
rect 3440 5070 3480 5085
rect 3440 4990 3445 5070
rect 3475 4990 3480 5070
rect 3440 4980 3480 4990
rect 3760 5290 3800 5300
rect 3760 5210 3765 5290
rect 3795 5210 3800 5290
rect 3760 5195 3800 5210
rect 3760 5165 3765 5195
rect 3795 5165 3800 5195
rect 3760 5115 3800 5165
rect 3760 5085 3765 5115
rect 3795 5085 3800 5115
rect 3760 5070 3800 5085
rect 3760 4990 3765 5070
rect 3795 4990 3800 5070
rect 3760 4980 3800 4990
rect 4080 5290 4120 5300
rect 4080 5210 4085 5290
rect 4115 5210 4120 5290
rect 4080 5195 4120 5210
rect 4080 5165 4085 5195
rect 4115 5165 4120 5195
rect 4080 5115 4120 5165
rect 4080 5085 4085 5115
rect 4115 5085 4120 5115
rect 4080 5070 4120 5085
rect 4080 4990 4085 5070
rect 4115 4990 4120 5070
rect 4080 4980 4120 4990
rect 4240 5290 4280 5300
rect 4240 5210 4245 5290
rect 4275 5210 4280 5290
rect 4240 5195 4280 5210
rect 4240 5165 4245 5195
rect 4275 5165 4280 5195
rect 4240 5115 4280 5165
rect 4240 5085 4245 5115
rect 4275 5085 4280 5115
rect 4240 5070 4280 5085
rect 4240 4990 4245 5070
rect 4275 4990 4280 5070
rect 4240 4980 4280 4990
rect 4560 5290 4600 5300
rect 4560 5210 4565 5290
rect 4595 5210 4600 5290
rect 4560 5195 4600 5210
rect 4560 5165 4565 5195
rect 4595 5165 4600 5195
rect 4560 5115 4600 5165
rect 4560 5085 4565 5115
rect 4595 5085 4600 5115
rect 4560 5070 4600 5085
rect 4560 4990 4565 5070
rect 4595 4990 4600 5070
rect 4560 4980 4600 4990
rect 640 4955 840 4960
rect 640 4925 650 4955
rect 830 4925 840 4955
rect 640 4920 840 4925
rect 960 4955 1160 4960
rect 960 4925 970 4955
rect 1150 4925 1160 4955
rect 960 4920 1160 4925
rect 1440 4955 1640 4960
rect 1440 4925 1450 4955
rect 1630 4925 1640 4955
rect 1440 4920 1640 4925
rect 1760 4955 1960 4960
rect 1760 4925 1770 4955
rect 1950 4925 1960 4955
rect 1760 4920 1960 4925
rect 2080 4955 2280 4960
rect 2080 4925 2090 4955
rect 2270 4925 2280 4955
rect 2080 4920 2280 4925
rect 2400 4955 2600 4960
rect 2400 4925 2410 4955
rect 2590 4925 2600 4955
rect 2400 4920 2600 4925
rect 2880 4955 3080 4960
rect 2880 4925 2890 4955
rect 3070 4925 3080 4955
rect 2880 4920 3080 4925
rect 3200 4955 3400 4960
rect 3200 4925 3210 4955
rect 3390 4925 3400 4955
rect 3200 4920 3400 4925
rect 3520 4955 3720 4960
rect 3520 4925 3530 4955
rect 3710 4925 3720 4955
rect 3520 4920 3720 4925
rect 3840 4955 4040 4960
rect 3840 4925 3850 4955
rect 4030 4925 4040 4955
rect 3840 4920 4040 4925
rect 4320 4955 4520 4960
rect 4320 4925 4330 4955
rect 4510 4925 4520 4955
rect 4320 4920 4520 4925
rect 560 4285 565 4315
rect 595 4285 600 4315
rect 560 4280 600 4285
rect 720 4795 760 4800
rect 720 4765 725 4795
rect 755 4765 760 4795
rect 560 4155 600 4160
rect 560 4125 565 4155
rect 595 4125 600 4155
rect 320 3995 520 4000
rect 320 3965 330 3995
rect 510 3965 520 3995
rect 320 3960 520 3965
rect 560 3960 600 4125
rect 720 4000 760 4765
rect 1040 4795 1080 4800
rect 1040 4765 1045 4795
rect 1075 4765 1080 4795
rect 880 4555 920 4560
rect 880 4525 885 4555
rect 915 4525 920 4555
rect 640 3995 840 4000
rect 640 3965 650 3995
rect 830 3965 840 3995
rect 640 3960 840 3965
rect 240 3850 245 3930
rect 275 3850 280 3930
rect 240 3840 280 3850
rect 560 3930 600 3940
rect 560 3850 565 3930
rect 595 3850 600 3930
rect 560 3840 600 3850
rect 880 3930 920 4525
rect 1040 4000 1080 4765
rect 1520 4795 1560 4800
rect 1520 4765 1525 4795
rect 1555 4765 1560 4795
rect 1200 4155 1240 4160
rect 1200 4125 1205 4155
rect 1235 4125 1240 4155
rect 960 3995 1160 4000
rect 960 3965 970 3995
rect 1150 3965 1160 3995
rect 960 3960 1160 3965
rect 880 3850 885 3930
rect 915 3850 920 3930
rect 880 3840 920 3850
rect 1200 3930 1240 4125
rect 1360 4155 1400 4160
rect 1360 4125 1365 4155
rect 1395 4125 1400 4155
rect 1200 3850 1205 3930
rect 1235 3850 1240 3930
rect 1200 3840 1240 3850
rect 1280 3915 1320 4000
rect 1280 3885 1285 3915
rect 1315 3885 1320 3915
rect -160 3805 -155 3835
rect -125 3805 -120 3835
rect -800 3725 -795 3755
rect -765 3725 -760 3755
rect -800 3720 -760 3725
rect -160 3755 -120 3805
rect -160 3725 -155 3755
rect -125 3725 -120 3755
rect -160 3720 -120 3725
rect 1280 3835 1320 3885
rect 1280 3805 1285 3835
rect 1315 3805 1320 3835
rect 1280 3755 1320 3805
rect 1360 3930 1400 4125
rect 1520 4000 1560 4765
rect 1840 4795 1880 4800
rect 1840 4765 1845 4795
rect 1875 4765 1880 4795
rect 1680 4555 1720 4560
rect 1680 4525 1685 4555
rect 1715 4525 1720 4555
rect 1440 3995 1640 4000
rect 1440 3965 1450 3995
rect 1630 3965 1640 3995
rect 1440 3960 1640 3965
rect 1360 3850 1365 3930
rect 1395 3850 1400 3930
rect 1360 3800 1400 3850
rect 1680 3930 1720 4525
rect 1840 4000 1880 4765
rect 2160 4795 2200 4800
rect 2160 4765 2165 4795
rect 2195 4765 2200 4795
rect 2000 4155 2040 4160
rect 2000 4125 2005 4155
rect 2035 4125 2040 4155
rect 1760 3995 1960 4000
rect 1760 3965 1770 3995
rect 1950 3965 1960 3995
rect 1760 3960 1960 3965
rect 1680 3850 1685 3930
rect 1715 3850 1720 3930
rect 1680 3840 1720 3850
rect 2000 3930 2040 4125
rect 2160 4000 2200 4765
rect 2480 4795 2520 4800
rect 2480 4765 2485 4795
rect 2515 4765 2520 4795
rect 2320 4555 2360 4560
rect 2320 4525 2325 4555
rect 2355 4525 2360 4555
rect 2080 3995 2280 4000
rect 2080 3965 2090 3995
rect 2270 3965 2280 3995
rect 2080 3960 2280 3965
rect 2000 3850 2005 3930
rect 2035 3850 2040 3930
rect 2000 3840 2040 3850
rect 2320 3930 2360 4525
rect 2480 4000 2520 4765
rect 4080 4795 4120 4800
rect 4080 4765 4085 4795
rect 4115 4765 4120 4795
rect 2640 4155 2680 4160
rect 2640 4125 2645 4155
rect 2675 4125 2680 4155
rect 2400 3995 2600 4000
rect 2400 3965 2410 3995
rect 2590 3965 2600 3995
rect 2400 3960 2600 3965
rect 2320 3850 2325 3930
rect 2355 3850 2360 3930
rect 2320 3840 2360 3850
rect 2640 3930 2680 4125
rect 2960 4155 3000 4160
rect 2960 4125 2965 4155
rect 2995 4125 3000 4155
rect 2960 4000 3000 4125
rect 3280 4155 3320 4160
rect 3280 4125 3285 4155
rect 3315 4125 3320 4155
rect 3280 4000 3320 4125
rect 3600 4155 3640 4160
rect 3600 4125 3605 4155
rect 3635 4125 3640 4155
rect 3600 4000 3640 4125
rect 3920 4155 3960 4160
rect 3920 4125 3925 4155
rect 3955 4125 3960 4155
rect 3920 4000 3960 4125
rect 2640 3850 2645 3930
rect 2675 3850 2680 3930
rect 2640 3840 2680 3850
rect 2720 3915 2760 4000
rect 2880 3995 3080 4000
rect 2880 3965 2890 3995
rect 3070 3965 3080 3995
rect 2880 3960 3080 3965
rect 3200 3995 3400 4000
rect 3200 3965 3210 3995
rect 3390 3965 3400 3995
rect 3200 3960 3400 3965
rect 2720 3885 2725 3915
rect 2755 3885 2760 3915
rect 2720 3835 2760 3885
rect 2720 3805 2725 3835
rect 2755 3805 2760 3835
rect 1280 3725 1285 3755
rect 1315 3725 1320 3755
rect 1280 3720 1320 3725
rect 2720 3755 2760 3805
rect 2800 3930 2840 3940
rect 2800 3850 2805 3930
rect 2835 3850 2840 3930
rect 2800 3835 2840 3850
rect 3120 3930 3160 3940
rect 3120 3850 3125 3930
rect 3155 3850 3160 3930
rect 3120 3840 3160 3850
rect 3440 3930 3480 4000
rect 3520 3995 3720 4000
rect 3520 3965 3530 3995
rect 3710 3965 3720 3995
rect 3520 3960 3720 3965
rect 3840 3995 4040 4000
rect 3840 3965 3850 3995
rect 4030 3965 4040 3995
rect 3840 3960 4040 3965
rect 3440 3850 3445 3930
rect 3475 3850 3480 3930
rect 3440 3840 3480 3850
rect 3760 3930 3800 3940
rect 3760 3850 3765 3930
rect 3795 3850 3800 3930
rect 3760 3840 3800 3850
rect 4080 3930 4120 4765
rect 4400 4155 4440 4160
rect 4400 4125 4405 4155
rect 4435 4125 4440 4155
rect 4400 4000 4440 4125
rect 4080 3850 4085 3930
rect 4115 3850 4120 3930
rect 4080 3840 4120 3850
rect 4160 3915 4200 4000
rect 4320 3995 4520 4000
rect 4320 3965 4330 3995
rect 4510 3965 4520 3995
rect 4320 3960 4520 3965
rect 4160 3885 4165 3915
rect 4195 3885 4200 3915
rect 2800 3805 2805 3835
rect 2835 3805 2840 3835
rect 2800 3800 2840 3805
rect 4160 3835 4200 3885
rect 4160 3805 4165 3835
rect 4195 3805 4200 3835
rect 2720 3725 2725 3755
rect 2755 3725 2760 3755
rect 2720 3720 2760 3725
rect 4160 3755 4200 3805
rect 4240 3930 4280 3940
rect 4240 3850 4245 3930
rect 4275 3850 4280 3930
rect 4240 3835 4280 3850
rect 4240 3805 4245 3835
rect 4275 3805 4280 3835
rect 4240 3800 4280 3805
rect 4560 3930 4600 3940
rect 4560 3850 4565 3930
rect 4595 3850 4600 3930
rect 4560 3835 4600 3850
rect 4560 3805 4565 3835
rect 4595 3805 4600 3835
rect 4560 3800 4600 3805
rect 4640 3915 4680 4000
rect 4640 3885 4645 3915
rect 4675 3885 4680 3915
rect 4640 3835 4680 3885
rect 4640 3805 4645 3835
rect 4675 3805 4680 3835
rect 4160 3725 4165 3755
rect 4195 3725 4200 3755
rect 4160 3720 4200 3725
rect 4640 3755 4680 3805
rect 4640 3725 4645 3755
rect 4675 3725 4680 3755
rect 4640 3720 4680 3725
rect -800 3675 -760 3680
rect -800 3645 -795 3675
rect -765 3645 -760 3675
rect -800 3640 -760 3645
rect -480 3435 -280 3440
rect -480 3405 -470 3435
rect -290 3405 -280 3435
rect -480 3400 -280 3405
rect 0 3435 200 3440
rect 0 3405 10 3435
rect 190 3405 200 3435
rect 0 3400 200 3405
rect 320 3435 520 3440
rect 320 3405 330 3435
rect 510 3405 520 3435
rect 320 3400 520 3405
rect 640 3435 840 3440
rect 640 3405 650 3435
rect 830 3405 840 3435
rect 640 3400 840 3405
rect 960 3435 1160 3440
rect 960 3405 970 3435
rect 1150 3405 1160 3435
rect 960 3400 1160 3405
rect 1440 3435 1640 3440
rect 1440 3405 1450 3435
rect 1630 3405 1640 3435
rect 1440 3400 1640 3405
rect 1760 3435 1960 3440
rect 1760 3405 1770 3435
rect 1950 3405 1960 3435
rect 1760 3400 1960 3405
rect 2080 3435 2280 3440
rect 2080 3405 2090 3435
rect 2270 3405 2280 3435
rect 2080 3400 2280 3405
rect 2400 3435 2600 3440
rect 2400 3405 2410 3435
rect 2590 3405 2600 3435
rect 2400 3400 2600 3405
rect 2880 3435 3080 3440
rect 2880 3405 2890 3435
rect 3070 3405 3080 3435
rect 2880 3400 3080 3405
rect 3200 3435 3400 3440
rect 3200 3405 3210 3435
rect 3390 3405 3400 3435
rect 3200 3400 3400 3405
rect 3520 3435 3720 3440
rect 3520 3405 3530 3435
rect 3710 3405 3720 3435
rect 3520 3400 3720 3405
rect 3840 3435 4040 3440
rect 3840 3405 3850 3435
rect 4030 3405 4040 3435
rect 3840 3400 4040 3405
rect 4080 3435 4120 3440
rect 4080 3405 4085 3435
rect 4115 3405 4120 3435
rect -560 3370 -520 3380
rect -560 3290 -555 3370
rect -525 3290 -520 3370
rect -560 3275 -520 3290
rect -560 3245 -555 3275
rect -525 3245 -520 3275
rect -560 3195 -520 3245
rect -560 3165 -555 3195
rect -525 3165 -520 3195
rect -560 3150 -520 3165
rect -560 3070 -555 3150
rect -525 3070 -520 3150
rect -560 3060 -520 3070
rect -240 3370 -200 3380
rect -240 3290 -235 3370
rect -205 3290 -200 3370
rect -240 3275 -200 3290
rect -240 3245 -235 3275
rect -205 3245 -200 3275
rect -240 3195 -200 3245
rect -240 3165 -235 3195
rect -205 3165 -200 3195
rect -240 3150 -200 3165
rect -240 3070 -235 3150
rect -205 3070 -200 3150
rect -240 3060 -200 3070
rect -80 3370 -40 3380
rect -80 3290 -75 3370
rect -45 3290 -40 3370
rect -80 3150 -40 3290
rect 240 3370 280 3380
rect 240 3290 245 3370
rect 275 3290 280 3370
rect 240 3280 280 3290
rect 560 3370 600 3380
rect 560 3290 565 3370
rect 595 3290 600 3370
rect 560 3275 600 3290
rect 880 3370 920 3380
rect 880 3290 885 3370
rect 915 3290 920 3370
rect 880 3280 920 3290
rect 1200 3370 1240 3380
rect 1200 3290 1205 3370
rect 1235 3290 1240 3370
rect 560 3245 565 3275
rect 595 3245 600 3275
rect 560 3240 600 3245
rect -80 3070 -75 3150
rect -45 3070 -40 3150
rect -80 3060 -40 3070
rect 240 3150 280 3160
rect 240 3070 245 3150
rect 275 3070 280 3150
rect 240 3060 280 3070
rect 560 3150 600 3160
rect 560 3070 565 3150
rect 595 3070 600 3150
rect -480 3035 -280 3040
rect -480 3005 -470 3035
rect -290 3005 -280 3035
rect -480 3000 -280 3005
rect 0 3035 200 3040
rect 0 3005 10 3035
rect 190 3005 200 3035
rect 0 3000 200 3005
rect 320 3035 520 3040
rect 320 3005 330 3035
rect 510 3005 520 3035
rect 320 3000 520 3005
rect 560 2635 600 3070
rect 880 3150 920 3160
rect 880 3070 885 3150
rect 915 3070 920 3150
rect 880 3060 920 3070
rect 1200 3150 1240 3290
rect 1200 3070 1205 3150
rect 1235 3070 1240 3150
rect 1200 3060 1240 3070
rect 1360 3370 1400 3380
rect 1360 3290 1365 3370
rect 1395 3290 1400 3370
rect 1360 3150 1400 3290
rect 1680 3370 1720 3380
rect 1680 3290 1685 3370
rect 1715 3290 1720 3370
rect 1680 3280 1720 3290
rect 2000 3370 2040 3380
rect 2000 3290 2005 3370
rect 2035 3290 2040 3370
rect 2000 3275 2040 3290
rect 2320 3370 2360 3380
rect 2320 3290 2325 3370
rect 2355 3290 2360 3370
rect 2320 3280 2360 3290
rect 2640 3370 2680 3380
rect 2640 3290 2645 3370
rect 2675 3290 2680 3370
rect 2000 3245 2005 3275
rect 2035 3245 2040 3275
rect 2000 3240 2040 3245
rect 1360 3070 1365 3150
rect 1395 3070 1400 3150
rect 1360 3060 1400 3070
rect 1680 3150 1720 3160
rect 1680 3070 1685 3150
rect 1715 3070 1720 3150
rect 1680 3060 1720 3070
rect 2000 3150 2040 3160
rect 2000 3070 2005 3150
rect 2035 3070 2040 3150
rect 640 3035 840 3040
rect 640 3005 650 3035
rect 830 3005 840 3035
rect 640 3000 840 3005
rect 960 3035 1160 3040
rect 960 3005 970 3035
rect 1150 3005 1160 3035
rect 960 3000 1160 3005
rect 1440 3035 1640 3040
rect 1440 3005 1450 3035
rect 1630 3005 1640 3035
rect 1440 3000 1640 3005
rect 1760 3035 1960 3040
rect 1760 3005 1770 3035
rect 1950 3005 1960 3035
rect 1760 3000 1960 3005
rect 2000 2875 2040 3070
rect 2320 3150 2360 3160
rect 2320 3070 2325 3150
rect 2355 3070 2360 3150
rect 2320 3060 2360 3070
rect 2640 3150 2680 3290
rect 2640 3070 2645 3150
rect 2675 3070 2680 3150
rect 2640 3060 2680 3070
rect 2800 3370 2840 3380
rect 2800 3290 2805 3370
rect 2835 3290 2840 3370
rect 2800 3275 2840 3290
rect 3120 3370 3160 3380
rect 3120 3290 3125 3370
rect 3155 3290 3160 3370
rect 3120 3280 3160 3290
rect 3440 3370 3480 3380
rect 3440 3290 3445 3370
rect 3475 3290 3480 3370
rect 3440 3280 3480 3290
rect 3760 3370 3800 3380
rect 3760 3290 3765 3370
rect 3795 3290 3800 3370
rect 3760 3280 3800 3290
rect 4080 3370 4120 3405
rect 4320 3435 4520 3440
rect 4320 3405 4330 3435
rect 4510 3405 4520 3435
rect 4320 3400 4520 3405
rect 4080 3290 4085 3370
rect 4115 3290 4120 3370
rect 2800 3245 2805 3275
rect 2835 3245 2840 3275
rect 2800 3195 2840 3245
rect 2800 3165 2805 3195
rect 2835 3165 2840 3195
rect 2800 3150 2840 3165
rect 2800 3070 2805 3150
rect 2835 3070 2840 3150
rect 2800 3060 2840 3070
rect 3120 3150 3160 3160
rect 3120 3070 3125 3150
rect 3155 3070 3160 3150
rect 3120 3060 3160 3070
rect 3440 3150 3480 3160
rect 3440 3070 3445 3150
rect 3475 3070 3480 3150
rect 3440 3060 3480 3070
rect 3760 3150 3800 3160
rect 3760 3070 3765 3150
rect 3795 3070 3800 3150
rect 3760 3060 3800 3070
rect 4080 3150 4120 3290
rect 4080 3070 4085 3150
rect 4115 3070 4120 3150
rect 2080 3035 2280 3040
rect 2080 3005 2090 3035
rect 2270 3005 2280 3035
rect 2080 3000 2280 3005
rect 2400 3035 2600 3040
rect 2400 3005 2410 3035
rect 2590 3005 2600 3035
rect 2400 3000 2600 3005
rect 2880 3035 3080 3040
rect 2880 3005 2890 3035
rect 3070 3005 3080 3035
rect 2880 3000 3080 3005
rect 3200 3035 3400 3040
rect 3200 3005 3210 3035
rect 3390 3005 3400 3035
rect 3200 3000 3400 3005
rect 3440 3035 3480 3040
rect 3440 3005 3445 3035
rect 3475 3005 3480 3035
rect 2000 2845 2005 2875
rect 2035 2845 2040 2875
rect 2000 2840 2040 2845
rect 2640 2875 2680 2880
rect 2640 2845 2645 2875
rect 2675 2845 2680 2875
rect 560 2605 565 2635
rect 595 2605 600 2635
rect 560 2600 600 2605
rect 1200 2635 1240 2640
rect 1200 2605 1205 2635
rect 1235 2605 1240 2635
rect -160 2475 -120 2480
rect -160 2445 -155 2475
rect -125 2445 -120 2475
rect -160 2315 -120 2445
rect -160 2285 -155 2315
rect -125 2285 -120 2315
rect -400 2235 -360 2240
rect -400 2205 -395 2235
rect -365 2205 -360 2235
rect -400 2080 -360 2205
rect -160 2155 -120 2285
rect -160 2125 -155 2155
rect -125 2125 -120 2155
rect -480 2075 -280 2080
rect -480 2045 -470 2075
rect -290 2045 -280 2075
rect -480 2040 -280 2045
rect -560 2010 -520 2020
rect -560 1930 -555 2010
rect -525 1930 -520 2010
rect -560 1915 -520 1930
rect -560 1885 -555 1915
rect -525 1885 -520 1915
rect -560 1880 -520 1885
rect -240 2010 -200 2020
rect -240 1930 -235 2010
rect -205 1930 -200 2010
rect -240 1915 -200 1930
rect -240 1885 -235 1915
rect -205 1885 -200 1915
rect -240 1880 -200 1885
rect -160 1995 -120 2125
rect 80 2395 120 2400
rect 80 2365 85 2395
rect 115 2365 120 2395
rect 80 2080 120 2365
rect 400 2395 440 2400
rect 400 2365 405 2395
rect 435 2365 440 2395
rect 400 2080 440 2365
rect 720 2395 760 2400
rect 720 2365 725 2395
rect 755 2365 760 2395
rect 720 2080 760 2365
rect 1040 2395 1080 2400
rect 1040 2365 1045 2395
rect 1075 2365 1080 2395
rect 1040 2080 1080 2365
rect 0 2075 200 2080
rect 0 2045 10 2075
rect 190 2045 200 2075
rect 0 2040 200 2045
rect 320 2075 520 2080
rect 320 2045 330 2075
rect 510 2045 520 2075
rect 320 2040 520 2045
rect 640 2075 840 2080
rect 640 2045 650 2075
rect 830 2045 840 2075
rect 640 2040 840 2045
rect 960 2075 1160 2080
rect 960 2045 970 2075
rect 1150 2045 1160 2075
rect 960 2040 1160 2045
rect -160 1965 -155 1995
rect -125 1965 -120 1995
rect -160 1915 -120 1965
rect -160 1885 -155 1915
rect -125 1885 -120 1915
rect -160 1835 -120 1885
rect -80 2010 -40 2020
rect -80 1930 -75 2010
rect -45 1930 -40 2010
rect -80 1915 -40 1930
rect 240 2010 280 2020
rect 240 1930 245 2010
rect 275 1930 280 2010
rect 240 1920 280 1930
rect 560 2010 600 2020
rect 560 1930 565 2010
rect 595 1930 600 2010
rect 560 1920 600 1930
rect 880 2010 920 2020
rect 880 1930 885 2010
rect 915 1930 920 2010
rect 880 1920 920 1930
rect 1200 2010 1240 2605
rect 1200 1930 1205 2010
rect 1235 1930 1240 2010
rect 1200 1920 1240 1930
rect 1280 2475 1320 2480
rect 1280 2445 1285 2475
rect 1315 2445 1320 2475
rect 1280 2315 1320 2445
rect 1280 2285 1285 2315
rect 1315 2285 1320 2315
rect 1280 2155 1320 2285
rect 1280 2125 1285 2155
rect 1315 2125 1320 2155
rect 1280 1995 1320 2125
rect 1520 2235 1560 2240
rect 1520 2205 1525 2235
rect 1555 2205 1560 2235
rect 1520 2080 1560 2205
rect 1840 2235 1880 2240
rect 1840 2205 1845 2235
rect 1875 2205 1880 2235
rect 1840 2080 1880 2205
rect 2160 2235 2200 2240
rect 2160 2205 2165 2235
rect 2195 2205 2200 2235
rect 2160 2080 2200 2205
rect 2480 2235 2520 2240
rect 2480 2205 2485 2235
rect 2515 2205 2520 2235
rect 2480 2080 2520 2205
rect 1440 2075 1640 2080
rect 1440 2045 1450 2075
rect 1630 2045 1640 2075
rect 1440 2040 1640 2045
rect 1760 2075 1960 2080
rect 1760 2045 1770 2075
rect 1950 2045 1960 2075
rect 1760 2040 1960 2045
rect 2080 2075 2280 2080
rect 2080 2045 2090 2075
rect 2270 2045 2280 2075
rect 2080 2040 2280 2045
rect 2400 2075 2600 2080
rect 2400 2045 2410 2075
rect 2590 2045 2600 2075
rect 2400 2040 2600 2045
rect 1280 1965 1285 1995
rect 1315 1965 1320 1995
rect -80 1885 -75 1915
rect -45 1885 -40 1915
rect -80 1880 -40 1885
rect 1280 1915 1320 1965
rect 1280 1885 1285 1915
rect 1315 1885 1320 1915
rect -160 1805 -155 1835
rect -125 1805 -120 1835
rect -160 1800 -120 1805
rect 1280 1835 1320 1885
rect 1360 2010 1400 2020
rect 1360 1930 1365 2010
rect 1395 1930 1400 2010
rect 1360 1915 1400 1930
rect 1680 2010 1720 2020
rect 1680 1930 1685 2010
rect 1715 1930 1720 2010
rect 1680 1920 1720 1930
rect 2000 2010 2040 2020
rect 2000 1930 2005 2010
rect 2035 1930 2040 2010
rect 2000 1920 2040 1930
rect 2320 2010 2360 2020
rect 2320 1930 2325 2010
rect 2355 1930 2360 2010
rect 2320 1920 2360 1930
rect 2640 2010 2680 2845
rect 2640 1930 2645 2010
rect 2675 1930 2680 2010
rect 2640 1920 2680 1930
rect 2720 2475 2760 2480
rect 2720 2445 2725 2475
rect 2755 2445 2760 2475
rect 2720 2315 2760 2445
rect 2720 2285 2725 2315
rect 2755 2285 2760 2315
rect 2720 2155 2760 2285
rect 2720 2125 2725 2155
rect 2755 2125 2760 2155
rect 2720 1995 2760 2125
rect 2960 2235 3000 2240
rect 2960 2205 2965 2235
rect 2995 2205 3000 2235
rect 2960 2080 3000 2205
rect 3280 2235 3320 2240
rect 3280 2205 3285 2235
rect 3315 2205 3320 2235
rect 3280 2080 3320 2205
rect 2880 2075 3080 2080
rect 2880 2045 2890 2075
rect 3070 2045 3080 2075
rect 2880 2040 3080 2045
rect 3200 2075 3400 2080
rect 3200 2045 3210 2075
rect 3390 2045 3400 2075
rect 3200 2040 3400 2045
rect 2720 1965 2725 1995
rect 2755 1965 2760 1995
rect 1360 1885 1365 1915
rect 1395 1885 1400 1915
rect 1360 1880 1400 1885
rect 2720 1915 2760 1965
rect 2720 1885 2725 1915
rect 2755 1885 2760 1915
rect 1280 1805 1285 1835
rect 1315 1805 1320 1835
rect 1280 1800 1320 1805
rect 2720 1835 2760 1885
rect 2800 2010 2840 2020
rect 2800 1930 2805 2010
rect 2835 1930 2840 2010
rect 2800 1915 2840 1930
rect 3120 2010 3160 2020
rect 3120 1930 3125 2010
rect 3155 1930 3160 2010
rect 3120 1920 3160 1930
rect 3440 2010 3480 3005
rect 3520 3035 3720 3040
rect 3520 3005 3530 3035
rect 3710 3005 3720 3035
rect 3520 3000 3720 3005
rect 3840 3035 4040 3040
rect 3840 3005 3850 3035
rect 4030 3005 4040 3035
rect 3840 3000 4040 3005
rect 4080 3035 4120 3070
rect 4240 3370 4280 3380
rect 4240 3290 4245 3370
rect 4275 3290 4280 3370
rect 4240 3275 4280 3290
rect 4240 3245 4245 3275
rect 4275 3245 4280 3275
rect 4240 3195 4280 3245
rect 4240 3165 4245 3195
rect 4275 3165 4280 3195
rect 4240 3150 4280 3165
rect 4240 3070 4245 3150
rect 4275 3070 4280 3150
rect 4240 3060 4280 3070
rect 4560 3370 4600 3380
rect 4560 3290 4565 3370
rect 4595 3290 4600 3370
rect 4560 3275 4600 3290
rect 4560 3245 4565 3275
rect 4595 3245 4600 3275
rect 4560 3195 4600 3245
rect 4560 3165 4565 3195
rect 4595 3165 4600 3195
rect 4560 3150 4600 3165
rect 4560 3070 4565 3150
rect 4595 3070 4600 3150
rect 4560 3060 4600 3070
rect 4080 3005 4085 3035
rect 4115 3005 4120 3035
rect 4080 3000 4120 3005
rect 4320 3035 4520 3040
rect 4320 3005 4330 3035
rect 4510 3005 4520 3035
rect 4320 3000 4520 3005
rect 4160 2475 4200 2480
rect 4160 2445 4165 2475
rect 4195 2445 4200 2475
rect 4160 2315 4200 2445
rect 4160 2285 4165 2315
rect 4195 2285 4200 2315
rect 3600 2235 3640 2240
rect 3600 2205 3605 2235
rect 3635 2205 3640 2235
rect 3600 2080 3640 2205
rect 3920 2235 3960 2240
rect 3920 2205 3925 2235
rect 3955 2205 3960 2235
rect 3920 2080 3960 2205
rect 4160 2155 4200 2285
rect 4640 2475 4680 2480
rect 4640 2445 4645 2475
rect 4675 2445 4680 2475
rect 4640 2315 4680 2445
rect 4640 2285 4645 2315
rect 4675 2285 4680 2315
rect 4160 2125 4165 2155
rect 4195 2125 4200 2155
rect 3520 2075 3720 2080
rect 3520 2045 3530 2075
rect 3710 2045 3720 2075
rect 3520 2040 3720 2045
rect 3840 2075 4040 2080
rect 3840 2045 3850 2075
rect 4030 2045 4040 2075
rect 3840 2040 4040 2045
rect 3440 1930 3445 2010
rect 3475 1930 3480 2010
rect 3440 1920 3480 1930
rect 3760 2010 3800 2020
rect 3760 1930 3765 2010
rect 3795 1930 3800 2010
rect 3760 1920 3800 1930
rect 4080 2010 4120 2020
rect 4080 1930 4085 2010
rect 4115 1930 4120 2010
rect 2800 1885 2805 1915
rect 2835 1885 2840 1915
rect 2800 1880 2840 1885
rect 4080 1915 4120 1930
rect 4080 1885 4085 1915
rect 4115 1885 4120 1915
rect 4080 1880 4120 1885
rect 4160 1995 4200 2125
rect 4400 2235 4440 2240
rect 4400 2205 4405 2235
rect 4435 2205 4440 2235
rect 4400 2080 4440 2205
rect 4640 2155 4680 2285
rect 4640 2125 4645 2155
rect 4675 2125 4680 2155
rect 4320 2075 4520 2080
rect 4320 2045 4330 2075
rect 4510 2045 4520 2075
rect 4320 2040 4520 2045
rect 4160 1965 4165 1995
rect 4195 1965 4200 1995
rect 4160 1915 4200 1965
rect 4160 1885 4165 1915
rect 4195 1885 4200 1915
rect 2720 1805 2725 1835
rect 2755 1805 2760 1835
rect 2720 1800 2760 1805
rect 4160 1835 4200 1885
rect 4240 2010 4280 2020
rect 4240 1930 4245 2010
rect 4275 1930 4280 2010
rect 4240 1915 4280 1930
rect 4240 1885 4245 1915
rect 4275 1885 4280 1915
rect 4240 1880 4280 1885
rect 4560 2010 4600 2020
rect 4560 1930 4565 2010
rect 4595 1930 4600 2010
rect 4560 1915 4600 1930
rect 4560 1885 4565 1915
rect 4595 1885 4600 1915
rect 4560 1880 4600 1885
rect 4640 1995 4680 2125
rect 4640 1965 4645 1995
rect 4675 1965 4680 1995
rect 4640 1915 4680 1965
rect 4640 1885 4645 1915
rect 4675 1885 4680 1915
rect 4160 1805 4165 1835
rect 4195 1805 4200 1835
rect 4160 1800 4200 1805
rect 4640 1835 4680 1885
rect 4640 1805 4645 1835
rect 4675 1805 4680 1835
rect 4640 1800 4680 1805
rect -480 1515 -280 1520
rect -480 1485 -470 1515
rect -290 1485 -280 1515
rect -480 1480 -280 1485
rect 0 1515 200 1520
rect 0 1485 10 1515
rect 190 1485 200 1515
rect 0 1480 200 1485
rect 320 1515 520 1520
rect 320 1485 330 1515
rect 510 1485 520 1515
rect 320 1480 520 1485
rect 640 1515 840 1520
rect 640 1485 650 1515
rect 830 1485 840 1515
rect 640 1480 840 1485
rect 960 1515 1160 1520
rect 960 1485 970 1515
rect 1150 1485 1160 1515
rect 960 1480 1160 1485
rect 1440 1515 1640 1520
rect 1440 1485 1450 1515
rect 1630 1485 1640 1515
rect 1440 1480 1640 1485
rect 1760 1515 1960 1520
rect 1760 1485 1770 1515
rect 1950 1485 1960 1515
rect 1760 1480 1960 1485
rect 2080 1515 2280 1520
rect 2080 1485 2090 1515
rect 2270 1485 2280 1515
rect 2080 1480 2280 1485
rect 2400 1515 2600 1520
rect 2400 1485 2410 1515
rect 2590 1485 2600 1515
rect 2400 1480 2600 1485
rect 2880 1515 3080 1520
rect 2880 1485 2890 1515
rect 3070 1485 3080 1515
rect 2880 1480 3080 1485
rect 3200 1515 3400 1520
rect 3200 1485 3210 1515
rect 3390 1485 3400 1515
rect 3200 1480 3400 1485
rect 3520 1515 3720 1520
rect 3520 1485 3530 1515
rect 3710 1485 3720 1515
rect 3520 1480 3720 1485
rect 3840 1515 4040 1520
rect 3840 1485 3850 1515
rect 4030 1485 4040 1515
rect 3840 1480 4040 1485
rect 4320 1515 4520 1520
rect 4320 1485 4330 1515
rect 4510 1485 4520 1515
rect 4320 1480 4520 1485
rect -560 1450 -520 1460
rect -560 1370 -555 1450
rect -525 1370 -520 1450
rect -560 1355 -520 1370
rect -560 1325 -555 1355
rect -525 1325 -520 1355
rect -560 1275 -520 1325
rect -560 1245 -555 1275
rect -525 1245 -520 1275
rect -560 1230 -520 1245
rect -560 1150 -555 1230
rect -525 1150 -520 1230
rect -560 1140 -520 1150
rect -240 1450 -200 1460
rect -240 1370 -235 1450
rect -205 1370 -200 1450
rect -240 1355 -200 1370
rect -240 1325 -235 1355
rect -205 1325 -200 1355
rect -240 1275 -200 1325
rect -240 1245 -235 1275
rect -205 1245 -200 1275
rect -240 1230 -200 1245
rect -240 1150 -235 1230
rect -205 1150 -200 1230
rect -240 1140 -200 1150
rect -80 1450 -40 1460
rect -80 1370 -75 1450
rect -45 1370 -40 1450
rect -80 1230 -40 1370
rect 240 1450 280 1460
rect 240 1370 245 1450
rect 275 1370 280 1450
rect 240 1355 280 1370
rect 240 1325 245 1355
rect 275 1325 280 1355
rect 240 1320 280 1325
rect 560 1450 600 1460
rect 560 1370 565 1450
rect 595 1370 600 1450
rect -80 1150 -75 1230
rect -45 1150 -40 1230
rect -80 1140 -40 1150
rect 240 1230 280 1240
rect 240 1150 245 1230
rect 275 1150 280 1230
rect -480 1115 -280 1120
rect -480 1085 -470 1115
rect -290 1085 -280 1115
rect -480 1080 -280 1085
rect 0 1115 200 1120
rect 0 1085 10 1115
rect 190 1085 200 1115
rect 0 1080 200 1085
rect -160 875 -120 880
rect -160 845 -155 875
rect -125 845 -120 875
rect -160 715 -120 845
rect -160 685 -155 715
rect -125 685 -120 715
rect -160 555 -120 685
rect -160 525 -155 555
rect -125 525 -120 555
rect -160 395 -120 525
rect -160 365 -155 395
rect -125 365 -120 395
rect -400 315 -360 320
rect -400 285 -395 315
rect -365 285 -360 315
rect -400 160 -360 285
rect -160 235 -120 365
rect -160 205 -155 235
rect -125 205 -120 235
rect -480 155 -280 160
rect -480 125 -470 155
rect -290 125 -280 155
rect -480 120 -280 125
rect -560 90 -520 100
rect -560 10 -555 90
rect -525 10 -520 90
rect -560 -5 -520 10
rect -560 -35 -555 -5
rect -525 -35 -520 -5
rect -560 -40 -520 -35
rect -240 90 -200 100
rect -240 10 -235 90
rect -205 10 -200 90
rect -240 -5 -200 10
rect -240 -35 -235 -5
rect -205 -35 -200 -5
rect -240 -40 -200 -35
rect -160 75 -120 205
rect 80 795 120 800
rect 80 765 85 795
rect 115 765 120 795
rect 80 160 120 765
rect 240 795 280 1150
rect 560 1230 600 1370
rect 880 1450 920 1460
rect 880 1370 885 1450
rect 915 1370 920 1450
rect 880 1355 920 1370
rect 880 1325 885 1355
rect 915 1325 920 1355
rect 880 1320 920 1325
rect 1200 1450 1240 1460
rect 1200 1370 1205 1450
rect 1235 1370 1240 1450
rect 560 1150 565 1230
rect 595 1150 600 1230
rect 560 1140 600 1150
rect 880 1230 920 1240
rect 880 1150 885 1230
rect 915 1150 920 1230
rect 320 1115 520 1120
rect 320 1085 330 1115
rect 510 1085 520 1115
rect 320 1080 520 1085
rect 640 1115 840 1120
rect 640 1085 650 1115
rect 830 1085 840 1115
rect 640 1080 840 1085
rect 240 765 245 795
rect 275 765 280 795
rect 240 760 280 765
rect 400 795 440 800
rect 400 765 405 795
rect 435 765 440 795
rect 400 160 440 765
rect 720 795 760 800
rect 720 765 725 795
rect 755 765 760 795
rect 560 475 600 480
rect 560 445 565 475
rect 595 445 600 475
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 120 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 120 520 125
rect -160 45 -155 75
rect -125 45 -120 75
rect -160 -5 -120 45
rect -160 -35 -155 -5
rect -125 -35 -120 -5
rect -160 -85 -120 -35
rect -80 90 -40 100
rect -80 10 -75 90
rect -45 10 -40 90
rect -80 -5 -40 10
rect 240 90 280 100
rect 240 10 245 90
rect 275 10 280 90
rect 240 0 280 10
rect 560 90 600 445
rect 720 160 760 765
rect 880 795 920 1150
rect 1200 1230 1240 1370
rect 1200 1150 1205 1230
rect 1235 1150 1240 1230
rect 1200 1140 1240 1150
rect 1360 1450 1400 1460
rect 1360 1370 1365 1450
rect 1395 1370 1400 1450
rect 1360 1230 1400 1370
rect 1680 1450 1720 1460
rect 1680 1370 1685 1450
rect 1715 1370 1720 1450
rect 1680 1360 1720 1370
rect 2000 1450 2040 1460
rect 2000 1370 2005 1450
rect 2035 1370 2040 1450
rect 2000 1355 2040 1370
rect 2320 1450 2360 1460
rect 2320 1370 2325 1450
rect 2355 1370 2360 1450
rect 2320 1360 2360 1370
rect 2640 1450 2680 1460
rect 2640 1370 2645 1450
rect 2675 1370 2680 1450
rect 2000 1325 2005 1355
rect 2035 1325 2040 1355
rect 2000 1320 2040 1325
rect 1360 1150 1365 1230
rect 1395 1150 1400 1230
rect 1360 1140 1400 1150
rect 1680 1230 1720 1240
rect 1680 1150 1685 1230
rect 1715 1150 1720 1230
rect 1680 1140 1720 1150
rect 2000 1230 2040 1240
rect 2000 1150 2005 1230
rect 2035 1150 2040 1230
rect 960 1115 1160 1120
rect 960 1085 970 1115
rect 1150 1085 1160 1115
rect 960 1080 1160 1085
rect 1440 1115 1640 1120
rect 1440 1085 1450 1115
rect 1630 1085 1640 1115
rect 1440 1080 1640 1085
rect 1760 1115 1960 1120
rect 1760 1085 1770 1115
rect 1950 1085 1960 1115
rect 1760 1080 1960 1085
rect 1280 875 1320 880
rect 1280 845 1285 875
rect 1315 845 1320 875
rect 880 765 885 795
rect 915 765 920 795
rect 880 760 920 765
rect 1040 795 1080 800
rect 1040 765 1045 795
rect 1075 765 1080 795
rect 1040 160 1080 765
rect 1200 795 1240 800
rect 1200 765 1205 795
rect 1235 765 1240 795
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 120 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 120 1160 125
rect 560 10 565 90
rect 595 10 600 90
rect 560 0 600 10
rect 880 90 920 100
rect 880 10 885 90
rect 915 10 920 90
rect 880 0 920 10
rect 1200 90 1240 765
rect 1200 10 1205 90
rect 1235 10 1240 90
rect 1200 0 1240 10
rect 1280 715 1320 845
rect 1280 685 1285 715
rect 1315 685 1320 715
rect 1280 555 1320 685
rect 1280 525 1285 555
rect 1315 525 1320 555
rect 1280 395 1320 525
rect 1280 365 1285 395
rect 1315 365 1320 395
rect 1280 235 1320 365
rect 1280 205 1285 235
rect 1315 205 1320 235
rect 1280 75 1320 205
rect 1520 795 1560 800
rect 1520 765 1525 795
rect 1555 765 1560 795
rect 1520 160 1560 765
rect 1840 795 1880 800
rect 1840 765 1845 795
rect 1875 765 1880 795
rect 1840 160 1880 765
rect 2000 635 2040 1150
rect 2320 1230 2360 1240
rect 2320 1150 2325 1230
rect 2355 1150 2360 1230
rect 2320 1140 2360 1150
rect 2640 1230 2680 1370
rect 2640 1150 2645 1230
rect 2675 1150 2680 1230
rect 2640 1140 2680 1150
rect 2800 1450 2840 1460
rect 2800 1370 2805 1450
rect 2835 1370 2840 1450
rect 2800 1230 2840 1370
rect 3120 1450 3160 1460
rect 3120 1370 3125 1450
rect 3155 1370 3160 1450
rect 3120 1360 3160 1370
rect 3440 1450 3480 1460
rect 3440 1370 3445 1450
rect 3475 1370 3480 1450
rect 3440 1355 3480 1370
rect 3760 1450 3800 1460
rect 3760 1370 3765 1450
rect 3795 1370 3800 1450
rect 3760 1360 3800 1370
rect 4080 1450 4120 1460
rect 4080 1370 4085 1450
rect 4115 1370 4120 1450
rect 3440 1325 3445 1355
rect 3475 1325 3480 1355
rect 3440 1320 3480 1325
rect 2800 1150 2805 1230
rect 2835 1150 2840 1230
rect 2800 1140 2840 1150
rect 3120 1230 3160 1240
rect 3120 1150 3125 1230
rect 3155 1150 3160 1230
rect 3120 1140 3160 1150
rect 3440 1230 3480 1240
rect 3440 1150 3445 1230
rect 3475 1150 3480 1230
rect 2080 1115 2280 1120
rect 2080 1085 2090 1115
rect 2270 1085 2280 1115
rect 2080 1080 2280 1085
rect 2400 1115 2600 1120
rect 2400 1085 2410 1115
rect 2590 1085 2600 1115
rect 2400 1080 2600 1085
rect 2880 1115 3080 1120
rect 2880 1085 2890 1115
rect 3070 1085 3080 1115
rect 2880 1080 3080 1085
rect 3200 1115 3400 1120
rect 3200 1085 3210 1115
rect 3390 1085 3400 1115
rect 3200 1080 3400 1085
rect 2720 875 2760 880
rect 2720 845 2725 875
rect 2755 845 2760 875
rect 2720 715 2760 845
rect 2720 685 2725 715
rect 2755 685 2760 715
rect 2000 605 2005 635
rect 2035 605 2040 635
rect 2000 600 2040 605
rect 2160 635 2200 640
rect 2160 605 2165 635
rect 2195 605 2200 635
rect 2000 475 2040 480
rect 2000 445 2005 475
rect 2035 445 2040 475
rect 1440 155 1640 160
rect 1440 125 1450 155
rect 1630 125 1640 155
rect 1440 120 1640 125
rect 1760 155 1960 160
rect 1760 125 1770 155
rect 1950 125 1960 155
rect 1760 120 1960 125
rect 1280 45 1285 75
rect 1315 45 1320 75
rect -80 -35 -75 -5
rect -45 -35 -40 -5
rect -80 -40 -40 -35
rect 1280 -5 1320 45
rect 1280 -35 1285 -5
rect 1315 -35 1320 -5
rect -160 -115 -155 -85
rect -125 -115 -120 -85
rect -160 -120 -120 -115
rect 1280 -85 1320 -35
rect 1360 90 1400 100
rect 1360 10 1365 90
rect 1395 10 1400 90
rect 1360 -5 1400 10
rect 1680 90 1720 100
rect 1680 10 1685 90
rect 1715 10 1720 90
rect 1680 0 1720 10
rect 2000 90 2040 445
rect 2160 160 2200 605
rect 2480 635 2520 640
rect 2480 605 2485 635
rect 2515 605 2520 635
rect 2480 160 2520 605
rect 2640 635 2680 640
rect 2640 605 2645 635
rect 2675 605 2680 635
rect 2080 155 2280 160
rect 2080 125 2090 155
rect 2270 125 2280 155
rect 2080 120 2280 125
rect 2400 155 2600 160
rect 2400 125 2410 155
rect 2590 125 2600 155
rect 2400 120 2600 125
rect 2000 10 2005 90
rect 2035 10 2040 90
rect 2000 0 2040 10
rect 2320 90 2360 100
rect 2320 10 2325 90
rect 2355 10 2360 90
rect 2320 0 2360 10
rect 2640 90 2680 605
rect 2640 10 2645 90
rect 2675 10 2680 90
rect 2640 0 2680 10
rect 2720 555 2760 685
rect 2720 525 2725 555
rect 2755 525 2760 555
rect 2720 395 2760 525
rect 2720 365 2725 395
rect 2755 365 2760 395
rect 2720 235 2760 365
rect 2720 205 2725 235
rect 2755 205 2760 235
rect 2720 75 2760 205
rect 2960 315 3000 320
rect 2960 285 2965 315
rect 2995 285 3000 315
rect 2960 160 3000 285
rect 3280 315 3320 320
rect 3280 285 3285 315
rect 3315 285 3320 315
rect 3280 160 3320 285
rect 3440 315 3480 1150
rect 3760 1230 3800 1240
rect 3760 1150 3765 1230
rect 3795 1150 3800 1230
rect 3760 1140 3800 1150
rect 4080 1230 4120 1370
rect 4080 1150 4085 1230
rect 4115 1150 4120 1230
rect 4080 1140 4120 1150
rect 4240 1450 4280 1460
rect 4240 1370 4245 1450
rect 4275 1370 4280 1450
rect 4240 1355 4280 1370
rect 4240 1325 4245 1355
rect 4275 1325 4280 1355
rect 4240 1275 4280 1325
rect 4240 1245 4245 1275
rect 4275 1245 4280 1275
rect 4240 1230 4280 1245
rect 4240 1150 4245 1230
rect 4275 1150 4280 1230
rect 4240 1140 4280 1150
rect 4560 1450 4600 1460
rect 4560 1370 4565 1450
rect 4595 1370 4600 1450
rect 4560 1355 4600 1370
rect 4560 1325 4565 1355
rect 4595 1325 4600 1355
rect 4560 1275 4600 1325
rect 4560 1245 4565 1275
rect 4595 1245 4600 1275
rect 4560 1230 4600 1245
rect 4560 1150 4565 1230
rect 4595 1150 4600 1230
rect 4560 1140 4600 1150
rect 3520 1115 3720 1120
rect 3520 1085 3530 1115
rect 3710 1085 3720 1115
rect 3520 1080 3720 1085
rect 3840 1115 4040 1120
rect 3840 1085 3850 1115
rect 4030 1085 4040 1115
rect 3840 1080 4040 1085
rect 4320 1115 4520 1120
rect 4320 1085 4330 1115
rect 4510 1085 4520 1115
rect 4320 1080 4520 1085
rect 4160 875 4200 880
rect 4160 845 4165 875
rect 4195 845 4200 875
rect 4160 715 4200 845
rect 4160 685 4165 715
rect 4195 685 4200 715
rect 4160 555 4200 685
rect 4160 525 4165 555
rect 4195 525 4200 555
rect 4160 395 4200 525
rect 4160 365 4165 395
rect 4195 365 4200 395
rect 3440 285 3445 315
rect 3475 285 3480 315
rect 3440 280 3480 285
rect 3600 315 3640 320
rect 3600 285 3605 315
rect 3635 285 3640 315
rect 3600 160 3640 285
rect 3920 315 3960 320
rect 3920 285 3925 315
rect 3955 285 3960 315
rect 3920 160 3960 285
rect 4080 315 4120 320
rect 4080 285 4085 315
rect 4115 285 4120 315
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 120 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 120 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 120 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 120 4040 125
rect 2720 45 2725 75
rect 2755 45 2760 75
rect 1360 -35 1365 -5
rect 1395 -35 1400 -5
rect 1360 -40 1400 -35
rect 2720 -5 2760 45
rect 2720 -35 2725 -5
rect 2755 -35 2760 -5
rect 1280 -115 1285 -85
rect 1315 -115 1320 -85
rect 1280 -120 1320 -115
rect 2720 -85 2760 -35
rect 2800 90 2840 100
rect 2800 10 2805 90
rect 2835 10 2840 90
rect 2800 -5 2840 10
rect 3120 90 3160 100
rect 3120 10 3125 90
rect 3155 10 3160 90
rect 3120 0 3160 10
rect 3440 90 3480 100
rect 3440 10 3445 90
rect 3475 10 3480 90
rect 3440 0 3480 10
rect 3760 90 3800 100
rect 3760 10 3765 90
rect 3795 10 3800 90
rect 3760 0 3800 10
rect 4080 90 4120 285
rect 4080 10 4085 90
rect 4115 10 4120 90
rect 4080 0 4120 10
rect 4160 235 4200 365
rect 4640 875 4680 880
rect 4640 845 4645 875
rect 4675 845 4680 875
rect 4640 715 4680 845
rect 4640 685 4645 715
rect 4675 685 4680 715
rect 4640 555 4680 685
rect 4640 525 4645 555
rect 4675 525 4680 555
rect 4640 395 4680 525
rect 4640 365 4645 395
rect 4675 365 4680 395
rect 4160 205 4165 235
rect 4195 205 4200 235
rect 4160 75 4200 205
rect 4400 315 4440 320
rect 4400 285 4405 315
rect 4435 285 4440 315
rect 4400 160 4440 285
rect 4640 235 4680 365
rect 4640 205 4645 235
rect 4675 205 4680 235
rect 4320 155 4520 160
rect 4320 125 4330 155
rect 4510 125 4520 155
rect 4320 120 4520 125
rect 4160 45 4165 75
rect 4195 45 4200 75
rect 2800 -35 2805 -5
rect 2835 -35 2840 -5
rect 2800 -40 2840 -35
rect 4160 -5 4200 45
rect 4160 -35 4165 -5
rect 4195 -35 4200 -5
rect 2720 -115 2725 -85
rect 2755 -115 2760 -85
rect 2720 -120 2760 -115
rect 4160 -85 4200 -35
rect 4240 90 4280 100
rect 4240 10 4245 90
rect 4275 10 4280 90
rect 4240 -5 4280 10
rect 4240 -35 4245 -5
rect 4275 -35 4280 -5
rect 4240 -40 4280 -35
rect 4560 90 4600 100
rect 4560 10 4565 90
rect 4595 10 4600 90
rect 4560 -5 4600 10
rect 4560 -35 4565 -5
rect 4595 -35 4600 -5
rect 4560 -40 4600 -35
rect 4640 75 4680 205
rect 4640 45 4645 75
rect 4675 45 4680 75
rect 4640 -5 4680 45
rect 4640 -35 4645 -5
rect 4675 -35 4680 -5
rect 4160 -115 4165 -85
rect 4195 -115 4200 -85
rect 4160 -120 4200 -115
rect 4640 -85 4680 -35
rect 4640 -115 4645 -85
rect 4675 -115 4680 -85
rect 4640 -120 4680 -115
<< via1 >>
rect -795 5565 -765 5595
rect -470 5325 -290 5355
rect 10 5325 190 5355
rect 330 5325 510 5355
rect 650 5325 830 5355
rect 970 5325 1150 5355
rect 1450 5325 1630 5355
rect 1770 5325 1950 5355
rect 2090 5325 2270 5355
rect 2410 5325 2590 5355
rect 2890 5325 3070 5355
rect 3210 5325 3390 5355
rect 3530 5325 3710 5355
rect 3850 5325 4030 5355
rect 4330 5325 4510 5355
rect -555 5165 -525 5195
rect -555 5085 -525 5115
rect -235 5165 -205 5195
rect -235 5085 -205 5115
rect 565 5245 595 5275
rect 565 5165 595 5195
rect -470 4925 -290 4955
rect 10 4925 190 4955
rect 330 4925 510 4955
rect 85 4765 115 4795
rect -395 4125 -365 4155
rect -795 4045 -765 4075
rect -75 4125 -45 4155
rect -795 3885 -765 3915
rect -795 3805 -765 3835
rect -555 3885 -525 3915
rect -555 3805 -525 3835
rect -235 3885 -205 3915
rect -235 3805 -205 3835
rect -155 3885 -125 3915
rect 405 4765 435 4795
rect 245 4525 275 4555
rect 1365 5165 1395 5195
rect 1365 5085 1395 5115
rect 1685 5165 1715 5195
rect 1685 5085 1715 5115
rect 2005 5245 2035 5275
rect 2005 5165 2035 5195
rect 2005 5085 2035 5115
rect 2325 5165 2355 5195
rect 2325 5085 2355 5115
rect 2645 5165 2675 5195
rect 2645 5085 2675 5115
rect 2805 5245 2835 5275
rect 2805 5165 2835 5195
rect 2805 5085 2835 5115
rect 2805 5005 2835 5035
rect 3125 5165 3155 5195
rect 3125 5085 3155 5115
rect 3445 5165 3475 5195
rect 3445 5085 3475 5115
rect 3765 5165 3795 5195
rect 3765 5085 3795 5115
rect 4085 5165 4115 5195
rect 4085 5085 4115 5115
rect 4245 5245 4275 5275
rect 4245 5165 4275 5195
rect 4245 5085 4275 5115
rect 4245 5005 4275 5035
rect 4565 5165 4595 5195
rect 4565 5085 4595 5115
rect 650 4925 830 4955
rect 970 4925 1150 4955
rect 1450 4925 1630 4955
rect 1770 4925 1950 4955
rect 2090 4925 2270 4955
rect 2410 4925 2590 4955
rect 2890 4925 3070 4955
rect 3210 4925 3390 4955
rect 3530 4925 3710 4955
rect 3850 4925 4030 4955
rect 4330 4925 4510 4955
rect 565 4285 595 4315
rect 725 4765 755 4795
rect 565 4125 595 4155
rect 1045 4765 1075 4795
rect 885 4525 915 4555
rect 1525 4765 1555 4795
rect 1205 4125 1235 4155
rect 1365 4125 1395 4155
rect 1285 3885 1315 3915
rect -155 3805 -125 3835
rect -795 3725 -765 3755
rect -155 3725 -125 3755
rect 1285 3805 1315 3835
rect 1845 4765 1875 4795
rect 1685 4525 1715 4555
rect 2165 4765 2195 4795
rect 2005 4125 2035 4155
rect 2485 4765 2515 4795
rect 2325 4525 2355 4555
rect 4085 4765 4115 4795
rect 2645 4125 2675 4155
rect 2965 4125 2995 4155
rect 3285 4125 3315 4155
rect 3605 4125 3635 4155
rect 3925 4125 3955 4155
rect 2725 3885 2755 3915
rect 2725 3805 2755 3835
rect 1285 3725 1315 3755
rect 2805 3885 2835 3915
rect 4405 4125 4435 4155
rect 4165 3885 4195 3915
rect 2805 3805 2835 3835
rect 4165 3805 4195 3835
rect 2725 3725 2755 3755
rect 4245 3885 4275 3915
rect 4245 3805 4275 3835
rect 4565 3885 4595 3915
rect 4565 3805 4595 3835
rect 4645 3885 4675 3915
rect 4645 3805 4675 3835
rect 4165 3725 4195 3755
rect 4645 3725 4675 3755
rect -795 3645 -765 3675
rect -470 3405 -290 3435
rect 10 3405 190 3435
rect 330 3405 510 3435
rect 650 3405 830 3435
rect 970 3405 1150 3435
rect 1450 3405 1630 3435
rect 1770 3405 1950 3435
rect 2090 3405 2270 3435
rect 2410 3405 2590 3435
rect 2890 3405 3070 3435
rect 3210 3405 3390 3435
rect 3530 3405 3710 3435
rect 3850 3405 4030 3435
rect 4085 3405 4115 3435
rect -555 3245 -525 3275
rect -555 3165 -525 3195
rect -235 3245 -205 3275
rect -235 3165 -205 3195
rect 565 3325 595 3355
rect 565 3245 595 3275
rect -470 3005 -290 3035
rect 10 3005 190 3035
rect 330 3005 510 3035
rect 2005 3325 2035 3355
rect 2005 3245 2035 3275
rect 650 3005 830 3035
rect 970 3005 1150 3035
rect 1450 3005 1630 3035
rect 1770 3005 1950 3035
rect 2805 3325 2835 3355
rect 4330 3405 4510 3435
rect 2805 3245 2835 3275
rect 2805 3165 2835 3195
rect 2805 3085 2835 3115
rect 2090 3005 2270 3035
rect 2410 3005 2590 3035
rect 2890 3005 3070 3035
rect 3210 3005 3390 3035
rect 3445 3005 3475 3035
rect 2005 2845 2035 2875
rect 2645 2845 2675 2875
rect 565 2605 595 2635
rect 1205 2605 1235 2635
rect -155 2445 -125 2475
rect -155 2285 -125 2315
rect -395 2205 -365 2235
rect -155 2125 -125 2155
rect -555 1965 -525 1995
rect -555 1885 -525 1915
rect -235 1965 -205 1995
rect -235 1885 -205 1915
rect 85 2365 115 2395
rect 405 2365 435 2395
rect 725 2365 755 2395
rect 1045 2365 1075 2395
rect -155 1965 -125 1995
rect -155 1885 -125 1915
rect -75 1965 -45 1995
rect 1285 2445 1315 2475
rect 1285 2285 1315 2315
rect 1285 2125 1315 2155
rect 1525 2205 1555 2235
rect 1845 2205 1875 2235
rect 2165 2205 2195 2235
rect 2485 2205 2515 2235
rect 1285 1965 1315 1995
rect -75 1885 -45 1915
rect 1285 1885 1315 1915
rect -155 1805 -125 1835
rect 1365 1965 1395 1995
rect 2725 2445 2755 2475
rect 2725 2285 2755 2315
rect 2725 2125 2755 2155
rect 2965 2205 2995 2235
rect 3285 2205 3315 2235
rect 2725 1965 2755 1995
rect 1365 1885 1395 1915
rect 2725 1885 2755 1915
rect 1285 1805 1315 1835
rect 2805 1965 2835 1995
rect 3530 3005 3710 3035
rect 3850 3005 4030 3035
rect 4245 3325 4275 3355
rect 4245 3245 4275 3275
rect 4245 3165 4275 3195
rect 4245 3085 4275 3115
rect 4565 3245 4595 3275
rect 4565 3165 4595 3195
rect 4085 3005 4115 3035
rect 4330 3005 4510 3035
rect 4165 2445 4195 2475
rect 4165 2285 4195 2315
rect 3605 2205 3635 2235
rect 3925 2205 3955 2235
rect 4645 2445 4675 2475
rect 4645 2285 4675 2315
rect 4165 2125 4195 2155
rect 4085 1965 4115 1995
rect 2805 1885 2835 1915
rect 4085 1885 4115 1915
rect 4405 2205 4435 2235
rect 4645 2125 4675 2155
rect 4165 1965 4195 1995
rect 4165 1885 4195 1915
rect 2725 1805 2755 1835
rect 4245 1965 4275 1995
rect 4245 1885 4275 1915
rect 4565 1965 4595 1995
rect 4565 1885 4595 1915
rect 4645 1965 4675 1995
rect 4645 1885 4675 1915
rect 4165 1805 4195 1835
rect 4645 1805 4675 1835
rect -470 1485 -290 1515
rect 10 1485 190 1515
rect 330 1485 510 1515
rect 650 1485 830 1515
rect 970 1485 1150 1515
rect 1450 1485 1630 1515
rect 1770 1485 1950 1515
rect 2090 1485 2270 1515
rect 2410 1485 2590 1515
rect 2890 1485 3070 1515
rect 3210 1485 3390 1515
rect 3530 1485 3710 1515
rect 3850 1485 4030 1515
rect 4330 1485 4510 1515
rect -555 1405 -525 1435
rect -555 1325 -525 1355
rect -555 1245 -525 1275
rect -555 1165 -525 1195
rect -235 1405 -205 1435
rect -235 1325 -205 1355
rect -235 1245 -205 1275
rect -235 1165 -205 1195
rect 245 1405 275 1435
rect 245 1325 275 1355
rect -470 1085 -290 1115
rect 10 1085 190 1115
rect -155 845 -125 875
rect -155 685 -125 715
rect -155 525 -125 555
rect -155 365 -125 395
rect -395 285 -365 315
rect -155 205 -125 235
rect -555 45 -525 75
rect -555 -35 -525 -5
rect -235 45 -205 75
rect -235 -35 -205 -5
rect 85 765 115 795
rect 885 1405 915 1435
rect 885 1325 915 1355
rect 330 1085 510 1115
rect 650 1085 830 1115
rect 245 765 275 795
rect 405 765 435 795
rect 725 765 755 795
rect 565 445 595 475
rect -155 45 -125 75
rect -155 -35 -125 -5
rect -75 45 -45 75
rect 2005 1405 2035 1435
rect 2005 1325 2035 1355
rect 970 1085 1150 1115
rect 1450 1085 1630 1115
rect 1770 1085 1950 1115
rect 1285 845 1315 875
rect 885 765 915 795
rect 1045 765 1075 795
rect 1205 765 1235 795
rect 1285 685 1315 715
rect 1285 525 1315 555
rect 1285 365 1315 395
rect 1285 205 1315 235
rect 1525 765 1555 795
rect 1845 765 1875 795
rect 3445 1405 3475 1435
rect 3445 1325 3475 1355
rect 2090 1085 2270 1115
rect 2410 1085 2590 1115
rect 2890 1085 3070 1115
rect 3210 1085 3390 1115
rect 2725 845 2755 875
rect 2725 685 2755 715
rect 2005 605 2035 635
rect 2165 605 2195 635
rect 2005 445 2035 475
rect 1285 45 1315 75
rect -75 -35 -45 -5
rect 1285 -35 1315 -5
rect -155 -115 -125 -85
rect 1365 45 1395 75
rect 2485 605 2515 635
rect 2645 605 2675 635
rect 2725 525 2755 555
rect 2725 365 2755 395
rect 2725 205 2755 235
rect 2965 285 2995 315
rect 3285 285 3315 315
rect 4245 1405 4275 1435
rect 4245 1325 4275 1355
rect 4245 1245 4275 1275
rect 4245 1165 4275 1195
rect 4565 1405 4595 1435
rect 4565 1325 4595 1355
rect 4565 1245 4595 1275
rect 4565 1165 4595 1195
rect 3530 1085 3710 1115
rect 3850 1085 4030 1115
rect 4330 1085 4510 1115
rect 4165 845 4195 875
rect 4165 685 4195 715
rect 4165 525 4195 555
rect 4165 365 4195 395
rect 3445 285 3475 315
rect 3605 285 3635 315
rect 3925 285 3955 315
rect 4085 285 4115 315
rect 2725 45 2755 75
rect 1365 -35 1395 -5
rect 2725 -35 2755 -5
rect 1285 -115 1315 -85
rect 2805 45 2835 75
rect 4645 845 4675 875
rect 4645 685 4675 715
rect 4645 525 4675 555
rect 4645 365 4675 395
rect 4165 205 4195 235
rect 4405 285 4435 315
rect 4645 205 4675 235
rect 4165 45 4195 75
rect 2805 -35 2835 -5
rect 4165 -35 4195 -5
rect 2725 -115 2755 -85
rect 4245 45 4275 75
rect 4245 -35 4275 -5
rect 4565 45 4595 75
rect 4565 -35 4595 -5
rect 4645 45 4675 75
rect 4645 -35 4675 -5
rect 4165 -115 4195 -85
rect 4645 -115 4675 -85
<< metal2 >>
rect -800 5595 4920 5600
rect -800 5565 -795 5595
rect -765 5565 4885 5595
rect 4915 5565 4920 5595
rect -800 5560 4920 5565
rect -880 5515 4840 5520
rect -880 5485 -875 5515
rect -845 5485 4840 5515
rect -880 5480 4840 5485
rect -880 5435 4840 5440
rect -880 5405 -875 5435
rect -845 5405 4840 5435
rect -880 5400 4840 5405
rect -960 5355 1160 5360
rect -960 5325 -955 5355
rect -925 5325 -470 5355
rect -290 5325 10 5355
rect 190 5325 330 5355
rect 510 5325 650 5355
rect 830 5325 970 5355
rect 1150 5325 1160 5355
rect -960 5320 1160 5325
rect 1440 5355 4840 5360
rect 1440 5325 1450 5355
rect 1630 5325 1770 5355
rect 1950 5325 2090 5355
rect 2270 5325 2410 5355
rect 2590 5325 2890 5355
rect 3070 5325 3210 5355
rect 3390 5325 3530 5355
rect 3710 5325 3850 5355
rect 4030 5325 4330 5355
rect 4510 5325 4840 5355
rect 1440 5320 4840 5325
rect -880 5275 4840 5280
rect -880 5245 -875 5275
rect -845 5245 565 5275
rect 595 5245 2005 5275
rect 2035 5245 2805 5275
rect 2835 5245 4245 5275
rect 4275 5245 4840 5275
rect -880 5240 4840 5245
rect -880 5195 4840 5200
rect -880 5165 -875 5195
rect -845 5165 -555 5195
rect -525 5165 -235 5195
rect -205 5165 565 5195
rect 595 5165 1365 5195
rect 1395 5165 1685 5195
rect 1715 5165 2005 5195
rect 2035 5165 2325 5195
rect 2355 5165 2645 5195
rect 2675 5165 2805 5195
rect 2835 5165 3125 5195
rect 3155 5165 3445 5195
rect 3475 5165 3765 5195
rect 3795 5165 4085 5195
rect 4115 5165 4245 5195
rect 4275 5165 4565 5195
rect 4595 5165 4840 5195
rect -880 5160 4840 5165
rect -880 5115 4840 5120
rect -880 5085 -875 5115
rect -845 5085 -555 5115
rect -525 5085 -235 5115
rect -205 5085 1365 5115
rect 1395 5085 1685 5115
rect 1715 5085 2005 5115
rect 2035 5085 2325 5115
rect 2355 5085 2645 5115
rect 2675 5085 2805 5115
rect 2835 5085 3125 5115
rect 3155 5085 3445 5115
rect 3475 5085 3765 5115
rect 3795 5085 4085 5115
rect 4115 5085 4245 5115
rect 4275 5085 4565 5115
rect 4595 5085 4840 5115
rect -880 5080 4840 5085
rect -1200 5035 4840 5040
rect -1200 5005 -1195 5035
rect -1165 5005 -1035 5035
rect -1005 5005 -875 5035
rect -845 5005 2805 5035
rect 2835 5005 4245 5035
rect 4275 5005 4840 5035
rect -1200 5000 4840 5005
rect -1120 4955 1160 4960
rect -1120 4925 -1115 4955
rect -1085 4925 -470 4955
rect -290 4925 10 4955
rect 190 4925 330 4955
rect 510 4925 650 4955
rect 830 4925 970 4955
rect 1150 4925 1160 4955
rect -1120 4920 1160 4925
rect 1440 4955 4840 4960
rect 1440 4925 1450 4955
rect 1630 4925 1770 4955
rect 1950 4925 2090 4955
rect 2270 4925 2410 4955
rect 2590 4925 2890 4955
rect 3070 4925 3210 4955
rect 3390 4925 3530 4955
rect 3710 4925 3850 4955
rect 4030 4925 4330 4955
rect 4510 4925 4840 4955
rect 1440 4920 4840 4925
rect -1520 4875 4840 4880
rect -1520 4845 -1515 4875
rect -1485 4845 -1355 4875
rect -1325 4845 -1195 4875
rect -1165 4845 -1035 4875
rect -1005 4845 -875 4875
rect -845 4845 4840 4875
rect -1520 4840 4840 4845
rect -1440 4795 4840 4800
rect -1440 4765 -1435 4795
rect -1405 4765 85 4795
rect 115 4765 405 4795
rect 435 4765 725 4795
rect 755 4765 1045 4795
rect 1075 4765 1525 4795
rect 1555 4765 1845 4795
rect 1875 4765 2165 4795
rect 2195 4765 2485 4795
rect 2515 4765 2965 4795
rect 2995 4765 3285 4795
rect 3315 4765 3605 4795
rect 3635 4765 3925 4795
rect 3955 4765 4085 4795
rect 4115 4765 4405 4795
rect 4435 4765 4840 4795
rect -1440 4760 4840 4765
rect -1520 4715 4840 4720
rect -1520 4685 -1515 4715
rect -1485 4685 -1355 4715
rect -1325 4685 -1195 4715
rect -1165 4685 -1035 4715
rect -1005 4685 -875 4715
rect -845 4685 4840 4715
rect -1520 4680 4840 4685
rect -1040 4635 4840 4640
rect -1040 4605 -1035 4635
rect -1005 4605 -875 4635
rect -845 4605 4840 4635
rect -1040 4600 4840 4605
rect -960 4555 4840 4560
rect -960 4525 -955 4555
rect -925 4525 245 4555
rect 275 4525 885 4555
rect 915 4525 1685 4555
rect 1715 4525 2325 4555
rect 2355 4525 4840 4555
rect -960 4520 4840 4525
rect -1040 4475 4840 4480
rect -1040 4445 -1035 4475
rect -1005 4445 -875 4475
rect -845 4445 4840 4475
rect -1040 4440 4840 4445
rect -800 4395 5720 4400
rect -800 4365 4885 4395
rect 4915 4365 5045 4395
rect 5075 4365 5205 4395
rect 5235 4365 5365 4395
rect 5395 4365 5525 4395
rect 5555 4365 5685 4395
rect 5715 4365 5720 4395
rect -800 4360 5720 4365
rect -800 4315 5640 4320
rect -800 4285 565 4315
rect 595 4285 5605 4315
rect 5635 4285 5640 4315
rect -800 4280 5640 4285
rect -800 4235 5720 4240
rect -800 4205 4885 4235
rect 4915 4205 5045 4235
rect 5075 4205 5205 4235
rect 5235 4205 5365 4235
rect 5395 4205 5525 4235
rect 5555 4205 5685 4235
rect 5715 4205 5720 4235
rect -800 4200 5720 4205
rect -800 4155 5000 4160
rect -800 4125 -395 4155
rect -365 4125 -75 4155
rect -45 4125 565 4155
rect 595 4125 1205 4155
rect 1235 4125 1365 4155
rect 1395 4125 2005 4155
rect 2035 4125 2645 4155
rect 2675 4125 2965 4155
rect 2995 4125 3285 4155
rect 3315 4125 3605 4155
rect 3635 4125 3925 4155
rect 3955 4125 4405 4155
rect 4435 4125 4965 4155
rect 4995 4125 5000 4155
rect -800 4120 5000 4125
rect -800 4075 5080 4080
rect -800 4045 -795 4075
rect -765 4045 4885 4075
rect 4915 4045 5045 4075
rect 5075 4045 5080 4075
rect -800 4040 5080 4045
rect -800 3995 4920 4000
rect -800 3965 4885 3995
rect 4915 3965 4920 3995
rect -800 3960 4920 3965
rect -800 3915 -80 3920
rect -800 3885 -795 3915
rect -765 3885 -555 3915
rect -525 3885 -235 3915
rect -205 3885 -155 3915
rect -125 3885 -80 3915
rect -800 3880 -80 3885
rect -40 3915 1360 3920
rect -40 3885 1285 3915
rect 1315 3885 1360 3915
rect -40 3880 1360 3885
rect 1400 3915 4920 3920
rect 1400 3885 2725 3915
rect 2755 3885 2805 3915
rect 2835 3885 4165 3915
rect 4195 3885 4245 3915
rect 4275 3885 4565 3915
rect 4595 3885 4645 3915
rect 4675 3885 4885 3915
rect 4915 3885 4920 3915
rect 1400 3880 4920 3885
rect -800 3835 4920 3840
rect -800 3805 -795 3835
rect -765 3805 -555 3835
rect -525 3805 -235 3835
rect -205 3805 -155 3835
rect -125 3805 1285 3835
rect 1315 3805 2725 3835
rect 2755 3805 2805 3835
rect 2835 3805 4165 3835
rect 4195 3805 4245 3835
rect 4275 3805 4565 3835
rect 4595 3805 4645 3835
rect 4675 3805 4885 3835
rect 4915 3805 4920 3835
rect -800 3800 4920 3805
rect -800 3755 4920 3760
rect -800 3725 -795 3755
rect -765 3725 -155 3755
rect -125 3725 1285 3755
rect 1315 3725 2725 3755
rect 2755 3725 4165 3755
rect 4195 3725 4645 3755
rect 4675 3725 4885 3755
rect 4915 3725 4920 3755
rect -800 3720 4920 3725
rect -800 3675 4920 3680
rect -800 3645 -795 3675
rect -765 3645 4885 3675
rect 4915 3645 4920 3675
rect -800 3640 4920 3645
rect -880 3595 4840 3600
rect -880 3565 -875 3595
rect -845 3565 4840 3595
rect -880 3560 4840 3565
rect -1360 3515 4840 3520
rect -1360 3485 -1355 3515
rect -1325 3485 -1195 3515
rect -1165 3485 -1035 3515
rect -1005 3485 -875 3515
rect -845 3485 4840 3515
rect -1360 3480 4840 3485
rect -1280 3435 2600 3440
rect -1280 3405 -1275 3435
rect -1245 3405 -470 3435
rect -290 3405 10 3435
rect 190 3405 330 3435
rect 510 3405 650 3435
rect 830 3405 970 3435
rect 1150 3405 1450 3435
rect 1630 3405 1770 3435
rect 1950 3405 2090 3435
rect 2270 3405 2410 3435
rect 2590 3405 2600 3435
rect -1280 3400 2600 3405
rect 2880 3435 4840 3440
rect 2880 3405 2890 3435
rect 3070 3405 3210 3435
rect 3390 3405 3530 3435
rect 3710 3405 3850 3435
rect 4030 3405 4085 3435
rect 4115 3405 4330 3435
rect 4510 3405 4840 3435
rect 2880 3400 4840 3405
rect -1360 3355 4840 3360
rect -1360 3325 -1355 3355
rect -1325 3325 -1195 3355
rect -1165 3325 -1035 3355
rect -1005 3325 -875 3355
rect -845 3325 565 3355
rect 595 3325 2005 3355
rect 2035 3325 2805 3355
rect 2835 3325 4245 3355
rect 4275 3325 4840 3355
rect -1360 3320 4840 3325
rect -880 3275 4840 3280
rect -880 3245 -875 3275
rect -845 3245 -555 3275
rect -525 3245 -235 3275
rect -205 3245 565 3275
rect 595 3245 2005 3275
rect 2035 3245 2805 3275
rect 2835 3245 4245 3275
rect 4275 3245 4565 3275
rect 4595 3245 4840 3275
rect -880 3240 4840 3245
rect -880 3195 4840 3200
rect -880 3165 -875 3195
rect -845 3165 -555 3195
rect -525 3165 -235 3195
rect -205 3165 2805 3195
rect 2835 3165 4245 3195
rect 4275 3165 4565 3195
rect 4595 3165 4840 3195
rect -880 3160 4840 3165
rect -1200 3115 4840 3120
rect -1200 3085 -1195 3115
rect -1165 3085 -1035 3115
rect -1005 3085 -875 3115
rect -845 3085 2805 3115
rect 2835 3085 4245 3115
rect 4275 3085 4840 3115
rect -1200 3080 4840 3085
rect -1120 3035 4840 3040
rect -1120 3005 -1115 3035
rect -1085 3005 -470 3035
rect -290 3005 10 3035
rect 190 3005 330 3035
rect 510 3005 650 3035
rect 830 3005 970 3035
rect 1150 3005 1450 3035
rect 1630 3005 1770 3035
rect 1950 3005 2090 3035
rect 2270 3005 2410 3035
rect 2590 3005 2890 3035
rect 3070 3005 3210 3035
rect 3390 3005 3445 3035
rect 3475 3005 3530 3035
rect 3710 3005 3850 3035
rect 4030 3005 4085 3035
rect 4115 3005 4330 3035
rect 4510 3005 4840 3035
rect -1120 3000 4840 3005
rect -1200 2955 4840 2960
rect -1200 2925 -1195 2955
rect -1165 2925 -1035 2955
rect -1005 2925 -875 2955
rect -845 2925 4840 2955
rect -1200 2920 4840 2925
rect -960 2875 4840 2880
rect -960 2845 -955 2875
rect -925 2845 2005 2875
rect 2035 2845 2645 2875
rect 2675 2845 4840 2875
rect -960 2840 4840 2845
rect -1040 2795 4840 2800
rect -1040 2765 -1035 2795
rect -1005 2765 -875 2795
rect -845 2765 4840 2795
rect -1040 2760 4840 2765
rect -1360 2715 4840 2720
rect -1360 2685 -1355 2715
rect -1325 2685 -1195 2715
rect -1165 2685 -1035 2715
rect -1005 2685 -875 2715
rect -845 2685 4840 2715
rect -1360 2680 4840 2685
rect -1280 2635 4840 2640
rect -1280 2605 -1275 2635
rect -1245 2605 565 2635
rect 595 2605 1205 2635
rect 1235 2605 4840 2635
rect -1280 2600 4840 2605
rect -1360 2555 4840 2560
rect -1360 2525 -1355 2555
rect -1325 2525 -1195 2555
rect -1165 2525 -1035 2555
rect -1005 2525 -875 2555
rect -845 2525 4840 2555
rect -1360 2520 4840 2525
rect -800 2475 5400 2480
rect -800 2445 -155 2475
rect -125 2445 1285 2475
rect 1315 2445 2725 2475
rect 2755 2445 4165 2475
rect 4195 2445 4645 2475
rect 4675 2445 4885 2475
rect 4915 2445 5045 2475
rect 5075 2445 5205 2475
rect 5235 2445 5365 2475
rect 5395 2445 5400 2475
rect -800 2440 5400 2445
rect -800 2395 5320 2400
rect -800 2365 85 2395
rect 115 2365 405 2395
rect 435 2365 725 2395
rect 755 2365 1045 2395
rect 1075 2365 5285 2395
rect 5315 2365 5320 2395
rect -800 2360 5320 2365
rect -800 2315 5400 2320
rect -800 2285 -155 2315
rect -125 2285 1285 2315
rect 1315 2285 2725 2315
rect 2755 2285 4165 2315
rect 4195 2285 4645 2315
rect 4675 2285 4885 2315
rect 4915 2285 5045 2315
rect 5075 2285 5205 2315
rect 5235 2285 5365 2315
rect 5395 2285 5400 2315
rect -800 2280 5400 2285
rect -800 2235 5000 2240
rect -800 2205 -395 2235
rect -365 2205 1525 2235
rect 1555 2205 1845 2235
rect 1875 2205 2165 2235
rect 2195 2205 2485 2235
rect 2515 2205 2965 2235
rect 2995 2205 3285 2235
rect 3315 2205 3605 2235
rect 3635 2205 3925 2235
rect 3955 2205 4405 2235
rect 4435 2205 4965 2235
rect 4995 2205 5000 2235
rect -800 2200 5000 2205
rect -800 2155 5080 2160
rect -800 2125 -155 2155
rect -125 2125 1285 2155
rect 1315 2125 2725 2155
rect 2755 2125 4165 2155
rect 4195 2125 4645 2155
rect 4675 2125 4885 2155
rect 4915 2125 5045 2155
rect 5075 2125 5080 2155
rect -800 2120 5080 2125
rect -800 2075 4920 2080
rect -800 2045 4885 2075
rect 4915 2045 4920 2075
rect -800 2040 4920 2045
rect -800 1995 4920 2000
rect -800 1965 -555 1995
rect -525 1965 -235 1995
rect -205 1965 -155 1995
rect -125 1965 -75 1995
rect -45 1965 1285 1995
rect 1315 1965 1365 1995
rect 1395 1965 2725 1995
rect 2755 1965 2805 1995
rect 2835 1965 4085 1995
rect 4115 1965 4165 1995
rect 4195 1965 4245 1995
rect 4275 1965 4565 1995
rect 4595 1965 4645 1995
rect 4675 1965 4885 1995
rect 4915 1965 4920 1995
rect -800 1960 4920 1965
rect -800 1915 4920 1920
rect -800 1885 -555 1915
rect -525 1885 -235 1915
rect -205 1885 -155 1915
rect -125 1885 -75 1915
rect -45 1885 1285 1915
rect 1315 1885 1365 1915
rect 1395 1885 2725 1915
rect 2755 1885 2805 1915
rect 2835 1885 4085 1915
rect 4115 1885 4165 1915
rect 4195 1885 4245 1915
rect 4275 1885 4565 1915
rect 4595 1885 4645 1915
rect 4675 1885 4885 1915
rect 4915 1885 4920 1915
rect -800 1880 4920 1885
rect -800 1835 4920 1840
rect -800 1805 -155 1835
rect -125 1805 1285 1835
rect 1315 1805 2725 1835
rect 2755 1805 4165 1835
rect 4195 1805 4645 1835
rect 4675 1805 4885 1835
rect 4915 1805 4920 1835
rect -800 1800 4920 1805
rect -760 1755 4920 1760
rect -760 1725 4885 1755
rect 4915 1725 4920 1755
rect -760 1720 4920 1725
rect -880 1675 4840 1680
rect -880 1645 -875 1675
rect -845 1645 4840 1675
rect -880 1640 4840 1645
rect -1040 1595 4840 1600
rect -1040 1565 -1035 1595
rect -1005 1565 -875 1595
rect -845 1565 4840 1595
rect -1040 1560 4840 1565
rect -960 1515 4840 1520
rect -960 1485 -955 1515
rect -925 1485 -470 1515
rect -290 1485 10 1515
rect 190 1485 330 1515
rect 510 1485 650 1515
rect 830 1485 970 1515
rect 1150 1485 1450 1515
rect 1630 1485 1770 1515
rect 1950 1485 2090 1515
rect 2270 1485 2410 1515
rect 2590 1485 2890 1515
rect 3070 1485 3210 1515
rect 3390 1485 3530 1515
rect 3710 1485 3850 1515
rect 4030 1485 4330 1515
rect 4510 1485 4840 1515
rect -960 1480 4840 1485
rect -1040 1435 4840 1440
rect -1040 1405 -1035 1435
rect -1005 1405 -875 1435
rect -845 1405 -555 1435
rect -525 1405 -235 1435
rect -205 1405 245 1435
rect 275 1405 885 1435
rect 915 1405 2005 1435
rect 2035 1405 3445 1435
rect 3475 1405 4245 1435
rect 4275 1405 4565 1435
rect 4595 1405 4840 1435
rect -1040 1400 4840 1405
rect -880 1355 4840 1360
rect -880 1325 -875 1355
rect -845 1325 -555 1355
rect -525 1325 -235 1355
rect -205 1325 245 1355
rect 275 1325 885 1355
rect 915 1325 2005 1355
rect 2035 1325 3445 1355
rect 3475 1325 4245 1355
rect 4275 1325 4565 1355
rect 4595 1325 4840 1355
rect -880 1320 4840 1325
rect -880 1275 4840 1280
rect -880 1245 -875 1275
rect -845 1245 -555 1275
rect -525 1245 -235 1275
rect -205 1245 4245 1275
rect 4275 1245 4565 1275
rect 4595 1245 4840 1275
rect -880 1240 4840 1245
rect -1200 1195 4840 1200
rect -1200 1165 -1195 1195
rect -1165 1165 -1035 1195
rect -1005 1165 -875 1195
rect -845 1165 -555 1195
rect -525 1165 -235 1195
rect -205 1165 4245 1195
rect 4275 1165 4565 1195
rect 4595 1165 4840 1195
rect -1200 1160 4840 1165
rect -1120 1115 4840 1120
rect -1120 1085 -1115 1115
rect -1085 1085 -470 1115
rect -290 1085 10 1115
rect 190 1085 330 1115
rect 510 1085 650 1115
rect 830 1085 970 1115
rect 1150 1085 1450 1115
rect 1630 1085 1770 1115
rect 1950 1085 2090 1115
rect 2270 1085 2410 1115
rect 2590 1085 2890 1115
rect 3070 1085 3210 1115
rect 3390 1085 3530 1115
rect 3710 1085 3850 1115
rect 4030 1085 4330 1115
rect 4510 1085 4840 1115
rect -1120 1080 4840 1085
rect -1200 1035 4840 1040
rect -1200 1005 -1195 1035
rect -1165 1005 -1035 1035
rect -1005 1005 -875 1035
rect -845 1005 4840 1035
rect -1200 1000 4840 1005
rect -880 955 4840 960
rect -880 925 -875 955
rect -845 925 4840 955
rect -880 920 4840 925
rect -800 875 5560 880
rect -800 845 -155 875
rect -125 845 1285 875
rect 1315 845 2725 875
rect 2755 845 4165 875
rect 4195 845 4645 875
rect 4675 845 4885 875
rect 4915 845 5045 875
rect 5075 845 5205 875
rect 5235 845 5365 875
rect 5395 845 5525 875
rect 5555 845 5560 875
rect -800 840 5560 845
rect -800 795 5480 800
rect -800 765 85 795
rect 115 765 245 795
rect 275 765 405 795
rect 435 765 725 795
rect 755 765 885 795
rect 915 765 1045 795
rect 1075 765 1205 795
rect 1235 765 1525 795
rect 1555 765 1845 795
rect 1875 765 5445 795
rect 5475 765 5480 795
rect -800 760 5480 765
rect -800 715 5560 720
rect -800 685 -155 715
rect -125 685 1285 715
rect 1315 685 2725 715
rect 2755 685 4165 715
rect 4195 685 4645 715
rect 4675 685 4885 715
rect 4915 685 5045 715
rect 5075 685 5205 715
rect 5235 685 5365 715
rect 5395 685 5525 715
rect 5555 685 5560 715
rect -800 680 5560 685
rect -800 635 5320 640
rect -800 605 2005 635
rect 2035 605 2165 635
rect 2195 605 2485 635
rect 2515 605 2645 635
rect 2675 605 5285 635
rect 5315 605 5320 635
rect -800 600 5320 605
rect -800 555 5400 560
rect -800 525 -155 555
rect -125 525 1285 555
rect 1315 525 2725 555
rect 2755 525 4165 555
rect 4195 525 4645 555
rect 4675 525 4885 555
rect 4915 525 5045 555
rect 5075 525 5205 555
rect 5235 525 5365 555
rect 5395 525 5400 555
rect -800 520 5400 525
rect -800 475 5160 480
rect -800 445 565 475
rect 595 445 2005 475
rect 2035 445 5125 475
rect 5155 445 5160 475
rect -800 440 5160 445
rect -800 395 5240 400
rect -800 365 -155 395
rect -125 365 1285 395
rect 1315 365 2725 395
rect 2755 365 4165 395
rect 4195 365 4645 395
rect 4675 365 4885 395
rect 4915 365 5045 395
rect 5075 365 5205 395
rect 5235 365 5240 395
rect -800 360 5240 365
rect -800 315 5000 320
rect -800 285 -395 315
rect -365 285 2965 315
rect 2995 285 3285 315
rect 3315 285 3445 315
rect 3475 285 3605 315
rect 3635 285 3925 315
rect 3955 285 4085 315
rect 4115 285 4405 315
rect 4435 285 4965 315
rect 4995 285 5000 315
rect -800 280 5000 285
rect -800 235 5080 240
rect -800 205 -155 235
rect -125 205 1285 235
rect 1315 205 2725 235
rect 2755 205 4165 235
rect 4195 205 4645 235
rect 4675 205 4885 235
rect 4915 205 5045 235
rect 5075 205 5080 235
rect -800 200 5080 205
rect -800 155 4920 160
rect -800 125 4885 155
rect 4915 125 4920 155
rect -800 120 4920 125
rect -800 75 4920 80
rect -800 45 -555 75
rect -525 45 -235 75
rect -205 45 -155 75
rect -125 45 -75 75
rect -45 45 1285 75
rect 1315 45 1365 75
rect 1395 45 2725 75
rect 2755 45 2805 75
rect 2835 45 4165 75
rect 4195 45 4245 75
rect 4275 45 4565 75
rect 4595 45 4645 75
rect 4675 45 4885 75
rect 4915 45 4920 75
rect -800 40 4920 45
rect -800 -5 4920 0
rect -800 -35 -555 -5
rect -525 -35 -235 -5
rect -205 -35 -155 -5
rect -125 -35 -75 -5
rect -45 -35 1285 -5
rect 1315 -35 1365 -5
rect 1395 -35 2725 -5
rect 2755 -35 2805 -5
rect 2835 -35 4165 -5
rect 4195 -35 4245 -5
rect 4275 -35 4565 -5
rect 4595 -35 4645 -5
rect 4675 -35 4885 -5
rect 4915 -35 4920 -5
rect -800 -40 4920 -35
rect -800 -85 4920 -80
rect -800 -115 -155 -85
rect -125 -115 1285 -85
rect 1315 -115 2725 -85
rect 2755 -115 4165 -85
rect 4195 -115 4645 -85
rect 4675 -115 4885 -85
rect 4915 -115 4920 -85
rect -800 -120 4920 -115
<< via2 >>
rect 4885 5565 4915 5595
rect -875 5485 -845 5515
rect -875 5405 -845 5435
rect -955 5325 -925 5355
rect 1525 5325 1555 5355
rect 1845 5325 1875 5355
rect 2165 5325 2195 5355
rect 2485 5325 2515 5355
rect 2965 5325 2995 5355
rect 3285 5325 3315 5355
rect 3605 5325 3635 5355
rect 3925 5325 3955 5355
rect 4405 5325 4435 5355
rect -875 5245 -845 5275
rect -875 5165 -845 5195
rect -875 5085 -845 5115
rect -1195 5005 -1165 5035
rect -1035 5005 -1005 5035
rect -875 5005 -845 5035
rect -1115 4925 -1085 4955
rect 1525 4925 1555 4955
rect 1845 4925 1875 4955
rect 2165 4925 2195 4955
rect 2485 4925 2515 4955
rect 2965 4925 2995 4955
rect 3285 4925 3315 4955
rect 3605 4925 3635 4955
rect 3925 4925 3955 4955
rect 4405 4925 4435 4955
rect -1515 4845 -1485 4875
rect -1355 4845 -1325 4875
rect -1195 4845 -1165 4875
rect -1035 4845 -1005 4875
rect -875 4845 -845 4875
rect -1435 4765 -1405 4795
rect 1525 4765 1555 4795
rect 1845 4765 1875 4795
rect 2165 4765 2195 4795
rect 2485 4765 2515 4795
rect 2965 4765 2995 4795
rect 3285 4765 3315 4795
rect 3605 4765 3635 4795
rect 3925 4765 3955 4795
rect 4405 4765 4435 4795
rect -1515 4685 -1485 4715
rect -1355 4685 -1325 4715
rect -1195 4685 -1165 4715
rect -1035 4685 -1005 4715
rect -875 4685 -845 4715
rect -1035 4605 -1005 4635
rect -875 4605 -845 4635
rect -955 4525 -925 4555
rect -1035 4445 -1005 4475
rect -875 4445 -845 4475
rect 4885 4365 4915 4395
rect 5045 4365 5075 4395
rect 5205 4365 5235 4395
rect 5365 4365 5395 4395
rect 5525 4365 5555 4395
rect 5685 4365 5715 4395
rect 5605 4285 5635 4315
rect 4885 4205 4915 4235
rect 5045 4205 5075 4235
rect 5205 4205 5235 4235
rect 5365 4205 5395 4235
rect 5525 4205 5555 4235
rect 5685 4205 5715 4235
rect 4965 4125 4995 4155
rect 4885 4045 4915 4075
rect 5045 4045 5075 4075
rect 4885 3965 4915 3995
rect 4885 3885 4915 3915
rect 4885 3805 4915 3835
rect 4885 3725 4915 3755
rect 4885 3645 4915 3675
rect -875 3565 -845 3595
rect -1355 3485 -1325 3515
rect -1195 3485 -1165 3515
rect -1035 3485 -1005 3515
rect -875 3485 -845 3515
rect -1275 3405 -1245 3435
rect -1355 3325 -1325 3355
rect -1195 3325 -1165 3355
rect -1035 3325 -1005 3355
rect -875 3325 -845 3355
rect -875 3245 -845 3275
rect -875 3165 -845 3195
rect -1195 3085 -1165 3115
rect -1035 3085 -1005 3115
rect -875 3085 -845 3115
rect -1115 3005 -1085 3035
rect -1195 2925 -1165 2955
rect -1035 2925 -1005 2955
rect -875 2925 -845 2955
rect -955 2845 -925 2875
rect -1035 2765 -1005 2795
rect -875 2765 -845 2795
rect -1355 2685 -1325 2715
rect -1195 2685 -1165 2715
rect -1035 2685 -1005 2715
rect -875 2685 -845 2715
rect -1275 2605 -1245 2635
rect -1355 2525 -1325 2555
rect -1195 2525 -1165 2555
rect -1035 2525 -1005 2555
rect -875 2525 -845 2555
rect 4885 2445 4915 2475
rect 5045 2445 5075 2475
rect 5205 2445 5235 2475
rect 5365 2445 5395 2475
rect 5285 2365 5315 2395
rect 4885 2285 4915 2315
rect 5045 2285 5075 2315
rect 5205 2285 5235 2315
rect 5365 2285 5395 2315
rect 4965 2205 4995 2235
rect 4885 2125 4915 2155
rect 5045 2125 5075 2155
rect 4885 2045 4915 2075
rect 4885 1965 4915 1995
rect 4885 1885 4915 1915
rect 4885 1805 4915 1835
rect 4885 1725 4915 1755
rect -875 1645 -845 1675
rect -1035 1565 -1005 1595
rect -875 1565 -845 1595
rect -955 1485 -925 1515
rect -1035 1405 -1005 1435
rect -875 1405 -845 1435
rect -875 1325 -845 1355
rect -875 1245 -845 1275
rect -1195 1165 -1165 1195
rect -1035 1165 -1005 1195
rect -875 1165 -845 1195
rect -1115 1085 -1085 1115
rect -1195 1005 -1165 1035
rect -1035 1005 -1005 1035
rect -875 1005 -845 1035
rect -875 925 -845 955
rect 4885 845 4915 875
rect 5045 845 5075 875
rect 5205 845 5235 875
rect 5365 845 5395 875
rect 5525 845 5555 875
rect 5445 765 5475 795
rect 4885 685 4915 715
rect 5045 685 5075 715
rect 5205 685 5235 715
rect 5365 685 5395 715
rect 5525 685 5555 715
rect 5285 605 5315 635
rect 4885 525 4915 555
rect 5045 525 5075 555
rect 5205 525 5235 555
rect 5365 525 5395 555
rect 5125 445 5155 475
rect 4885 365 4915 395
rect 5045 365 5075 395
rect 5205 365 5235 395
rect 4965 285 4995 315
rect 4885 205 4915 235
rect 5045 205 5075 235
rect 4885 125 4915 155
rect 4885 45 4915 75
rect 4885 -35 4915 -5
rect 4885 -115 4915 -85
<< metal3 >>
rect -1520 4875 -1480 5600
rect -1520 4845 -1515 4875
rect -1485 4845 -1480 4875
rect -1520 4715 -1480 4845
rect -1520 4685 -1515 4715
rect -1485 4685 -1480 4715
rect -1520 -120 -1480 4685
rect -1440 4795 -1400 5600
rect -1440 4765 -1435 4795
rect -1405 4765 -1400 4795
rect -1440 -120 -1400 4765
rect -1360 4875 -1320 5600
rect -1360 4845 -1355 4875
rect -1325 4845 -1320 4875
rect -1360 4715 -1320 4845
rect -1360 4685 -1355 4715
rect -1325 4685 -1320 4715
rect -1360 3515 -1320 4685
rect -1360 3485 -1355 3515
rect -1325 3485 -1320 3515
rect -1360 3355 -1320 3485
rect -1360 3325 -1355 3355
rect -1325 3325 -1320 3355
rect -1360 2715 -1320 3325
rect -1360 2685 -1355 2715
rect -1325 2685 -1320 2715
rect -1360 2555 -1320 2685
rect -1360 2525 -1355 2555
rect -1325 2525 -1320 2555
rect -1360 -120 -1320 2525
rect -1280 3435 -1240 5600
rect -1280 3405 -1275 3435
rect -1245 3405 -1240 3435
rect -1280 2635 -1240 3405
rect -1280 2605 -1275 2635
rect -1245 2605 -1240 2635
rect -1280 -120 -1240 2605
rect -1200 5035 -1160 5600
rect -1200 5005 -1195 5035
rect -1165 5005 -1160 5035
rect -1200 4875 -1160 5005
rect -1200 4845 -1195 4875
rect -1165 4845 -1160 4875
rect -1200 4715 -1160 4845
rect -1200 4685 -1195 4715
rect -1165 4685 -1160 4715
rect -1200 3515 -1160 4685
rect -1200 3485 -1195 3515
rect -1165 3485 -1160 3515
rect -1200 3355 -1160 3485
rect -1200 3325 -1195 3355
rect -1165 3325 -1160 3355
rect -1200 3115 -1160 3325
rect -1200 3085 -1195 3115
rect -1165 3085 -1160 3115
rect -1200 2955 -1160 3085
rect -1200 2925 -1195 2955
rect -1165 2925 -1160 2955
rect -1200 2715 -1160 2925
rect -1200 2685 -1195 2715
rect -1165 2685 -1160 2715
rect -1200 2555 -1160 2685
rect -1200 2525 -1195 2555
rect -1165 2525 -1160 2555
rect -1200 1195 -1160 2525
rect -1200 1165 -1195 1195
rect -1165 1165 -1160 1195
rect -1200 1035 -1160 1165
rect -1200 1005 -1195 1035
rect -1165 1005 -1160 1035
rect -1200 -120 -1160 1005
rect -1120 4955 -1080 5600
rect -1120 4925 -1115 4955
rect -1085 4925 -1080 4955
rect -1120 3035 -1080 4925
rect -1120 3005 -1115 3035
rect -1085 3005 -1080 3035
rect -1120 1115 -1080 3005
rect -1120 1085 -1115 1115
rect -1085 1085 -1080 1115
rect -1120 -120 -1080 1085
rect -1040 5035 -1000 5600
rect -1040 5005 -1035 5035
rect -1005 5005 -1000 5035
rect -1040 4875 -1000 5005
rect -1040 4845 -1035 4875
rect -1005 4845 -1000 4875
rect -1040 4715 -1000 4845
rect -1040 4685 -1035 4715
rect -1005 4685 -1000 4715
rect -1040 4635 -1000 4685
rect -1040 4605 -1035 4635
rect -1005 4605 -1000 4635
rect -1040 4475 -1000 4605
rect -1040 4445 -1035 4475
rect -1005 4445 -1000 4475
rect -1040 3515 -1000 4445
rect -1040 3485 -1035 3515
rect -1005 3485 -1000 3515
rect -1040 3355 -1000 3485
rect -1040 3325 -1035 3355
rect -1005 3325 -1000 3355
rect -1040 3115 -1000 3325
rect -1040 3085 -1035 3115
rect -1005 3085 -1000 3115
rect -1040 2955 -1000 3085
rect -1040 2925 -1035 2955
rect -1005 2925 -1000 2955
rect -1040 2795 -1000 2925
rect -1040 2765 -1035 2795
rect -1005 2765 -1000 2795
rect -1040 2715 -1000 2765
rect -1040 2685 -1035 2715
rect -1005 2685 -1000 2715
rect -1040 2555 -1000 2685
rect -1040 2525 -1035 2555
rect -1005 2525 -1000 2555
rect -1040 1595 -1000 2525
rect -1040 1565 -1035 1595
rect -1005 1565 -1000 1595
rect -1040 1435 -1000 1565
rect -1040 1405 -1035 1435
rect -1005 1405 -1000 1435
rect -1040 1195 -1000 1405
rect -1040 1165 -1035 1195
rect -1005 1165 -1000 1195
rect -1040 1035 -1000 1165
rect -1040 1005 -1035 1035
rect -1005 1005 -1000 1035
rect -1040 -120 -1000 1005
rect -960 5355 -920 5600
rect -960 5325 -955 5355
rect -925 5325 -920 5355
rect -960 4555 -920 5325
rect -960 4525 -955 4555
rect -925 4525 -920 4555
rect -960 2875 -920 4525
rect -960 2845 -955 2875
rect -925 2845 -920 2875
rect -960 1515 -920 2845
rect -960 1485 -955 1515
rect -925 1485 -920 1515
rect -960 -120 -920 1485
rect -880 5515 -840 5600
rect -880 5485 -875 5515
rect -845 5485 -840 5515
rect -880 5435 -840 5485
rect -880 5405 -875 5435
rect -845 5405 -840 5435
rect -880 5275 -840 5405
rect 4880 5595 4920 5600
rect 4880 5565 4885 5595
rect 4915 5565 4920 5595
rect -880 5245 -875 5275
rect -845 5245 -840 5275
rect -880 5195 -840 5245
rect -880 5165 -875 5195
rect -845 5165 -840 5195
rect -880 5115 -840 5165
rect -880 5085 -875 5115
rect -845 5085 -840 5115
rect -880 5035 -840 5085
rect -880 5005 -875 5035
rect -845 5005 -840 5035
rect -880 4875 -840 5005
rect -880 4845 -875 4875
rect -845 4845 -840 4875
rect -880 4715 -840 4845
rect 1520 5355 1560 5360
rect 1520 5325 1525 5355
rect 1555 5325 1560 5355
rect 1520 4955 1560 5325
rect 1520 4925 1525 4955
rect 1555 4925 1560 4955
rect 1520 4795 1560 4925
rect 1520 4765 1525 4795
rect 1555 4765 1560 4795
rect 1520 4760 1560 4765
rect 1840 5355 1880 5360
rect 1840 5325 1845 5355
rect 1875 5325 1880 5355
rect 1840 4955 1880 5325
rect 1840 4925 1845 4955
rect 1875 4925 1880 4955
rect 1840 4795 1880 4925
rect 1840 4765 1845 4795
rect 1875 4765 1880 4795
rect 1840 4760 1880 4765
rect 2160 5355 2200 5360
rect 2160 5325 2165 5355
rect 2195 5325 2200 5355
rect 2160 4955 2200 5325
rect 2160 4925 2165 4955
rect 2195 4925 2200 4955
rect 2160 4795 2200 4925
rect 2160 4765 2165 4795
rect 2195 4765 2200 4795
rect 2160 4760 2200 4765
rect 2480 5355 2520 5360
rect 2480 5325 2485 5355
rect 2515 5325 2520 5355
rect 2480 4955 2520 5325
rect 2480 4925 2485 4955
rect 2515 4925 2520 4955
rect 2480 4795 2520 4925
rect 2480 4765 2485 4795
rect 2515 4765 2520 4795
rect 2480 4760 2520 4765
rect 2960 5355 3000 5360
rect 2960 5325 2965 5355
rect 2995 5325 3000 5355
rect 2960 4955 3000 5325
rect 2960 4925 2965 4955
rect 2995 4925 3000 4955
rect 2960 4795 3000 4925
rect 2960 4765 2965 4795
rect 2995 4765 3000 4795
rect 2960 4760 3000 4765
rect 3280 5355 3320 5360
rect 3280 5325 3285 5355
rect 3315 5325 3320 5355
rect 3280 4955 3320 5325
rect 3280 4925 3285 4955
rect 3315 4925 3320 4955
rect 3280 4795 3320 4925
rect 3280 4765 3285 4795
rect 3315 4765 3320 4795
rect 3280 4760 3320 4765
rect 3600 5355 3640 5360
rect 3600 5325 3605 5355
rect 3635 5325 3640 5355
rect 3600 4955 3640 5325
rect 3600 4925 3605 4955
rect 3635 4925 3640 4955
rect 3600 4795 3640 4925
rect 3600 4765 3605 4795
rect 3635 4765 3640 4795
rect 3600 4760 3640 4765
rect 3920 5355 3960 5360
rect 3920 5325 3925 5355
rect 3955 5325 3960 5355
rect 3920 4955 3960 5325
rect 3920 4925 3925 4955
rect 3955 4925 3960 4955
rect 3920 4795 3960 4925
rect 3920 4765 3925 4795
rect 3955 4765 3960 4795
rect 3920 4760 3960 4765
rect 4400 5355 4440 5360
rect 4400 5325 4405 5355
rect 4435 5325 4440 5355
rect 4400 4955 4440 5325
rect 4400 4925 4405 4955
rect 4435 4925 4440 4955
rect 4400 4795 4440 4925
rect 4400 4765 4405 4795
rect 4435 4765 4440 4795
rect 4400 4760 4440 4765
rect -880 4685 -875 4715
rect -845 4685 -840 4715
rect -880 4635 -840 4685
rect -880 4605 -875 4635
rect -845 4605 -840 4635
rect -880 4475 -840 4605
rect -880 4445 -875 4475
rect -845 4445 -840 4475
rect -880 3595 -840 4445
rect -880 3565 -875 3595
rect -845 3565 -840 3595
rect -880 3515 -840 3565
rect -880 3485 -875 3515
rect -845 3485 -840 3515
rect -880 3355 -840 3485
rect -880 3325 -875 3355
rect -845 3325 -840 3355
rect -880 3275 -840 3325
rect -880 3245 -875 3275
rect -845 3245 -840 3275
rect -880 3195 -840 3245
rect -880 3165 -875 3195
rect -845 3165 -840 3195
rect -880 3115 -840 3165
rect -880 3085 -875 3115
rect -845 3085 -840 3115
rect -880 2955 -840 3085
rect -880 2925 -875 2955
rect -845 2925 -840 2955
rect -880 2795 -840 2925
rect -880 2765 -875 2795
rect -845 2765 -840 2795
rect -880 2715 -840 2765
rect -880 2685 -875 2715
rect -845 2685 -840 2715
rect -880 2555 -840 2685
rect -880 2525 -875 2555
rect -845 2525 -840 2555
rect -880 1675 -840 2525
rect -880 1645 -875 1675
rect -845 1645 -840 1675
rect -880 1595 -840 1645
rect -880 1565 -875 1595
rect -845 1565 -840 1595
rect -880 1435 -840 1565
rect -880 1405 -875 1435
rect -845 1405 -840 1435
rect -880 1355 -840 1405
rect -880 1325 -875 1355
rect -845 1325 -840 1355
rect -880 1275 -840 1325
rect -880 1245 -875 1275
rect -845 1245 -840 1275
rect -880 1195 -840 1245
rect -880 1165 -875 1195
rect -845 1165 -840 1195
rect -880 1035 -840 1165
rect -880 1005 -875 1035
rect -845 1005 -840 1035
rect -880 955 -840 1005
rect -880 925 -875 955
rect -845 925 -840 955
rect -880 -120 -840 925
rect 4880 4395 4920 5565
rect 4880 4365 4885 4395
rect 4915 4365 4920 4395
rect 4880 4235 4920 4365
rect 4880 4205 4885 4235
rect 4915 4205 4920 4235
rect 4880 4075 4920 4205
rect 4880 4045 4885 4075
rect 4915 4045 4920 4075
rect 4880 3995 4920 4045
rect 4880 3965 4885 3995
rect 4915 3965 4920 3995
rect 4880 3915 4920 3965
rect 4880 3885 4885 3915
rect 4915 3885 4920 3915
rect 4880 3835 4920 3885
rect 4880 3805 4885 3835
rect 4915 3805 4920 3835
rect 4880 3755 4920 3805
rect 4880 3725 4885 3755
rect 4915 3725 4920 3755
rect 4880 3675 4920 3725
rect 4880 3645 4885 3675
rect 4915 3645 4920 3675
rect 4880 2475 4920 3645
rect 4880 2445 4885 2475
rect 4915 2445 4920 2475
rect 4880 2315 4920 2445
rect 4880 2285 4885 2315
rect 4915 2285 4920 2315
rect 4880 2155 4920 2285
rect 4880 2125 4885 2155
rect 4915 2125 4920 2155
rect 4880 2075 4920 2125
rect 4880 2045 4885 2075
rect 4915 2045 4920 2075
rect 4880 1995 4920 2045
rect 4880 1965 4885 1995
rect 4915 1965 4920 1995
rect 4880 1915 4920 1965
rect 4880 1885 4885 1915
rect 4915 1885 4920 1915
rect 4880 1835 4920 1885
rect 4880 1805 4885 1835
rect 4915 1805 4920 1835
rect 4880 1755 4920 1805
rect 4880 1725 4885 1755
rect 4915 1725 4920 1755
rect 4880 875 4920 1725
rect 4880 845 4885 875
rect 4915 845 4920 875
rect 4880 715 4920 845
rect 4880 685 4885 715
rect 4915 685 4920 715
rect 4880 555 4920 685
rect 4880 525 4885 555
rect 4915 525 4920 555
rect 4880 395 4920 525
rect 4880 365 4885 395
rect 4915 365 4920 395
rect 4880 235 4920 365
rect 4880 205 4885 235
rect 4915 205 4920 235
rect 4880 155 4920 205
rect 4880 125 4885 155
rect 4915 125 4920 155
rect 4880 75 4920 125
rect 4880 45 4885 75
rect 4915 45 4920 75
rect 4880 -5 4920 45
rect 4880 -35 4885 -5
rect 4915 -35 4920 -5
rect 4880 -85 4920 -35
rect 4880 -115 4885 -85
rect 4915 -115 4920 -85
rect 4880 -120 4920 -115
rect 4960 4155 5000 5600
rect 4960 4125 4965 4155
rect 4995 4125 5000 4155
rect 4960 2235 5000 4125
rect 4960 2205 4965 2235
rect 4995 2205 5000 2235
rect 4960 315 5000 2205
rect 4960 285 4965 315
rect 4995 285 5000 315
rect 4960 -120 5000 285
rect 5040 4395 5080 5600
rect 5040 4365 5045 4395
rect 5075 4365 5080 4395
rect 5040 4235 5080 4365
rect 5040 4205 5045 4235
rect 5075 4205 5080 4235
rect 5040 4075 5080 4205
rect 5040 4045 5045 4075
rect 5075 4045 5080 4075
rect 5040 2475 5080 4045
rect 5040 2445 5045 2475
rect 5075 2445 5080 2475
rect 5040 2315 5080 2445
rect 5040 2285 5045 2315
rect 5075 2285 5080 2315
rect 5040 2155 5080 2285
rect 5040 2125 5045 2155
rect 5075 2125 5080 2155
rect 5040 875 5080 2125
rect 5040 845 5045 875
rect 5075 845 5080 875
rect 5040 715 5080 845
rect 5040 685 5045 715
rect 5075 685 5080 715
rect 5040 555 5080 685
rect 5040 525 5045 555
rect 5075 525 5080 555
rect 5040 395 5080 525
rect 5040 365 5045 395
rect 5075 365 5080 395
rect 5040 235 5080 365
rect 5040 205 5045 235
rect 5075 205 5080 235
rect 5040 -120 5080 205
rect 5120 475 5160 5600
rect 5120 445 5125 475
rect 5155 445 5160 475
rect 5120 -120 5160 445
rect 5200 4395 5240 5600
rect 5200 4365 5205 4395
rect 5235 4365 5240 4395
rect 5200 4235 5240 4365
rect 5200 4205 5205 4235
rect 5235 4205 5240 4235
rect 5200 2475 5240 4205
rect 5200 2445 5205 2475
rect 5235 2445 5240 2475
rect 5200 2315 5240 2445
rect 5200 2285 5205 2315
rect 5235 2285 5240 2315
rect 5200 875 5240 2285
rect 5200 845 5205 875
rect 5235 845 5240 875
rect 5200 715 5240 845
rect 5200 685 5205 715
rect 5235 685 5240 715
rect 5200 555 5240 685
rect 5200 525 5205 555
rect 5235 525 5240 555
rect 5200 395 5240 525
rect 5200 365 5205 395
rect 5235 365 5240 395
rect 5200 -120 5240 365
rect 5280 2395 5320 5600
rect 5280 2365 5285 2395
rect 5315 2365 5320 2395
rect 5280 635 5320 2365
rect 5280 605 5285 635
rect 5315 605 5320 635
rect 5280 -120 5320 605
rect 5360 4395 5400 5600
rect 5360 4365 5365 4395
rect 5395 4365 5400 4395
rect 5360 4235 5400 4365
rect 5360 4205 5365 4235
rect 5395 4205 5400 4235
rect 5360 2475 5400 4205
rect 5360 2445 5365 2475
rect 5395 2445 5400 2475
rect 5360 2315 5400 2445
rect 5360 2285 5365 2315
rect 5395 2285 5400 2315
rect 5360 875 5400 2285
rect 5360 845 5365 875
rect 5395 845 5400 875
rect 5360 715 5400 845
rect 5360 685 5365 715
rect 5395 685 5400 715
rect 5360 555 5400 685
rect 5360 525 5365 555
rect 5395 525 5400 555
rect 5360 -120 5400 525
rect 5440 795 5480 5600
rect 5440 765 5445 795
rect 5475 765 5480 795
rect 5440 -120 5480 765
rect 5520 4395 5560 5600
rect 5520 4365 5525 4395
rect 5555 4365 5560 4395
rect 5520 4235 5560 4365
rect 5520 4205 5525 4235
rect 5555 4205 5560 4235
rect 5520 875 5560 4205
rect 5520 845 5525 875
rect 5555 845 5560 875
rect 5520 715 5560 845
rect 5520 685 5525 715
rect 5555 685 5560 715
rect 5520 -120 5560 685
rect 5600 4315 5640 5600
rect 5600 4285 5605 4315
rect 5635 4285 5640 4315
rect 5600 -120 5640 4285
rect 5680 4395 5720 5600
rect 5680 4365 5685 4395
rect 5715 4365 5720 4395
rect 5680 4235 5720 4365
rect 5680 4205 5685 4235
rect 5715 4205 5720 4235
rect 5680 -120 5720 4205
<< labels >>
rlabel metal3 4960 5560 5000 5600 0 n
rlabel metal3 5120 5560 5160 5600 0 z
rlabel metal3 5280 5560 5320 5600 0 y
rlabel metal3 5440 5560 5480 5600 0 x
port 4 nsew
rlabel metal3 5600 5560 5640 5600 0 io
port 1 nsew
rlabel metal3 -960 5560 -920 5600 0 p1
rlabel metal3 -1120 5560 -1080 5600 0 p2
rlabel metal3 -1280 5560 -1240 5600 0 p0
rlabel metal3 -1440 5560 -1400 5600 0 s
rlabel metal3 -1520 5560 -1480 5600 0 vdda
port 2 nsew
rlabel metal3 5680 5560 5720 5600 0 vssa
port 3 nsew
<< end >>
