magic
tech sky130A
timestamp 1641007606
<< nwell >>
rect -200 480 10520 920
rect -240 -1200 10480 -760
rect -240 -1920 10480 -1480
rect -200 -3600 10520 -3160
<< pmoslvt >>
rect 0 660 200 760
rect 320 660 520 760
rect 640 660 840 760
rect 960 660 1160 760
rect 1280 660 1480 760
rect 1600 660 1800 760
rect 1920 660 2120 760
rect 2240 660 2440 760
rect 2560 660 2760 760
rect 2880 660 3080 760
rect 3200 660 3400 760
rect 3520 660 3720 760
rect 3840 660 4040 760
rect 4160 660 4360 760
rect 4480 660 4680 760
rect 4800 660 5000 760
rect 5280 660 5480 760
rect 5600 660 5800 760
rect 5920 660 6120 760
rect 6240 660 6440 760
rect 6560 660 6760 760
rect 6880 660 7080 760
rect 7200 660 7400 760
rect 7520 660 7720 760
rect 7840 660 8040 760
rect 8160 660 8360 760
rect 8480 660 8680 760
rect 8800 660 9000 760
rect 9120 660 9320 760
rect 9440 660 9640 760
rect 9760 660 9960 760
rect 10080 660 10280 760
rect 0 -1040 200 -940
rect 320 -1040 520 -940
rect 640 -1040 840 -940
rect 960 -1040 1160 -940
rect 1280 -1040 1480 -940
rect 1600 -1040 1800 -940
rect 1920 -1040 2120 -940
rect 2240 -1040 2440 -940
rect 2560 -1040 2760 -940
rect 2880 -1040 3080 -940
rect 3200 -1040 3400 -940
rect 3520 -1040 3720 -940
rect 3840 -1040 4040 -940
rect 4160 -1040 4360 -940
rect 4480 -1040 4680 -940
rect 4800 -1040 5000 -940
rect 5280 -1040 5480 -940
rect 5600 -1040 5800 -940
rect 5920 -1040 6120 -940
rect 6240 -1040 6440 -940
rect 6560 -1040 6760 -940
rect 6880 -1040 7080 -940
rect 7200 -1040 7400 -940
rect 7520 -1040 7720 -940
rect 7840 -1040 8040 -940
rect 8160 -1040 8360 -940
rect 8480 -1040 8680 -940
rect 8800 -1040 9000 -940
rect 9120 -1040 9320 -940
rect 9440 -1040 9640 -940
rect 9760 -1040 9960 -940
rect 10080 -1040 10280 -940
rect 0 -1740 200 -1640
rect 320 -1740 520 -1640
rect 640 -1740 840 -1640
rect 960 -1740 1160 -1640
rect 1280 -1740 1480 -1640
rect 1600 -1740 1800 -1640
rect 1920 -1740 2120 -1640
rect 2240 -1740 2440 -1640
rect 2560 -1740 2760 -1640
rect 2880 -1740 3080 -1640
rect 3200 -1740 3400 -1640
rect 3520 -1740 3720 -1640
rect 3840 -1740 4040 -1640
rect 4160 -1740 4360 -1640
rect 4480 -1740 4680 -1640
rect 4800 -1740 5000 -1640
rect 5280 -1740 5480 -1640
rect 5600 -1740 5800 -1640
rect 5920 -1740 6120 -1640
rect 6240 -1740 6440 -1640
rect 6560 -1740 6760 -1640
rect 6880 -1740 7080 -1640
rect 7200 -1740 7400 -1640
rect 7520 -1740 7720 -1640
rect 7840 -1740 8040 -1640
rect 8160 -1740 8360 -1640
rect 8480 -1740 8680 -1640
rect 8800 -1740 9000 -1640
rect 9120 -1740 9320 -1640
rect 9440 -1740 9640 -1640
rect 9760 -1740 9960 -1640
rect 10080 -1740 10280 -1640
rect 0 -3440 200 -3340
rect 320 -3440 520 -3340
rect 640 -3440 840 -3340
rect 960 -3440 1160 -3340
rect 1280 -3440 1480 -3340
rect 1600 -3440 1800 -3340
rect 1920 -3440 2120 -3340
rect 2240 -3440 2440 -3340
rect 2560 -3440 2760 -3340
rect 2880 -3440 3080 -3340
rect 3200 -3440 3400 -3340
rect 3520 -3440 3720 -3340
rect 3840 -3440 4040 -3340
rect 4160 -3440 4360 -3340
rect 4480 -3440 4680 -3340
rect 4800 -3440 5000 -3340
rect 5280 -3440 5480 -3340
rect 5600 -3440 5800 -3340
rect 5920 -3440 6120 -3340
rect 6240 -3440 6440 -3340
rect 6560 -3440 6760 -3340
rect 6880 -3440 7080 -3340
rect 7200 -3440 7400 -3340
rect 7520 -3440 7720 -3340
rect 7840 -3440 8040 -3340
rect 8160 -3440 8360 -3340
rect 8480 -3440 8680 -3340
rect 8800 -3440 9000 -3340
rect 9120 -3440 9320 -3340
rect 9440 -3440 9640 -3340
rect 9760 -3440 9960 -3340
rect 10080 -3440 10280 -3340
<< nmoslvt >>
rect 0 0 200 100
rect 320 0 520 100
rect 640 0 840 100
rect 960 0 1160 100
rect 1280 0 1480 100
rect 1600 0 1800 100
rect 1920 0 2120 100
rect 2240 0 2440 100
rect 2560 0 2760 100
rect 2880 0 3080 100
rect 3200 0 3400 100
rect 3520 0 3720 100
rect 3840 0 4040 100
rect 4160 0 4360 100
rect 4480 0 4680 100
rect 4800 0 5000 100
rect 5280 0 5480 100
rect 5600 0 5800 100
rect 5920 0 6120 100
rect 6240 0 6440 100
rect 6560 0 6760 100
rect 6880 0 7080 100
rect 7200 0 7400 100
rect 7520 0 7720 100
rect 7840 0 8040 100
rect 8160 0 8360 100
rect 8480 0 8680 100
rect 8800 0 9000 100
rect 9120 0 9320 100
rect 9440 0 9640 100
rect 9760 0 9960 100
rect 10080 0 10280 100
rect 0 -380 200 -280
rect 320 -380 520 -280
rect 640 -380 840 -280
rect 960 -380 1160 -280
rect 1280 -380 1480 -280
rect 1600 -380 1800 -280
rect 1920 -380 2120 -280
rect 2240 -380 2440 -280
rect 2560 -380 2760 -280
rect 2880 -380 3080 -280
rect 3200 -380 3400 -280
rect 3520 -380 3720 -280
rect 3840 -380 4040 -280
rect 4160 -380 4360 -280
rect 4480 -380 4680 -280
rect 4800 -380 5000 -280
rect 5280 -380 5480 -280
rect 5600 -380 5800 -280
rect 5920 -380 6120 -280
rect 6240 -380 6440 -280
rect 6560 -380 6760 -280
rect 6880 -380 7080 -280
rect 7200 -380 7400 -280
rect 7520 -380 7720 -280
rect 7840 -380 8040 -280
rect 8160 -380 8360 -280
rect 8480 -380 8680 -280
rect 8800 -380 9000 -280
rect 9120 -380 9320 -280
rect 9440 -380 9640 -280
rect 9760 -380 9960 -280
rect 10080 -380 10280 -280
rect 0 -2400 200 -2300
rect 320 -2400 520 -2300
rect 640 -2400 840 -2300
rect 960 -2400 1160 -2300
rect 1280 -2400 1480 -2300
rect 1600 -2400 1800 -2300
rect 1920 -2400 2120 -2300
rect 2240 -2400 2440 -2300
rect 2560 -2400 2760 -2300
rect 2880 -2400 3080 -2300
rect 3200 -2400 3400 -2300
rect 3520 -2400 3720 -2300
rect 3840 -2400 4040 -2300
rect 4160 -2400 4360 -2300
rect 4480 -2400 4680 -2300
rect 4800 -2400 5000 -2300
rect 5280 -2400 5480 -2300
rect 5600 -2400 5800 -2300
rect 5920 -2400 6120 -2300
rect 6240 -2400 6440 -2300
rect 6560 -2400 6760 -2300
rect 6880 -2400 7080 -2300
rect 7200 -2400 7400 -2300
rect 7520 -2400 7720 -2300
rect 7840 -2400 8040 -2300
rect 8160 -2400 8360 -2300
rect 8480 -2400 8680 -2300
rect 8800 -2400 9000 -2300
rect 9120 -2400 9320 -2300
rect 9440 -2400 9640 -2300
rect 9760 -2400 9960 -2300
rect 10080 -2400 10280 -2300
rect 0 -2780 200 -2680
rect 320 -2780 520 -2680
rect 640 -2780 840 -2680
rect 960 -2780 1160 -2680
rect 1280 -2780 1480 -2680
rect 1600 -2780 1800 -2680
rect 1920 -2780 2120 -2680
rect 2240 -2780 2440 -2680
rect 2560 -2780 2760 -2680
rect 2880 -2780 3080 -2680
rect 3200 -2780 3400 -2680
rect 3520 -2780 3720 -2680
rect 3840 -2780 4040 -2680
rect 4160 -2780 4360 -2680
rect 4480 -2780 4680 -2680
rect 4800 -2780 5000 -2680
rect 5280 -2780 5480 -2680
rect 5600 -2780 5800 -2680
rect 5920 -2780 6120 -2680
rect 6240 -2780 6440 -2680
rect 6560 -2780 6760 -2680
rect 6880 -2780 7080 -2680
rect 7200 -2780 7400 -2680
rect 7520 -2780 7720 -2680
rect 7840 -2780 8040 -2680
rect 8160 -2780 8360 -2680
rect 8480 -2780 8680 -2680
rect 8800 -2780 9000 -2680
rect 9120 -2780 9320 -2680
rect 9440 -2780 9640 -2680
rect 9760 -2780 9960 -2680
rect 10080 -2780 10280 -2680
<< ndiff >>
rect -80 90 0 100
rect -80 10 -75 90
rect -45 10 0 90
rect -80 0 0 10
rect 200 90 320 100
rect 200 10 245 90
rect 275 10 320 90
rect 200 0 320 10
rect 520 90 640 100
rect 520 10 565 90
rect 595 10 640 90
rect 520 0 640 10
rect 840 90 960 100
rect 840 10 885 90
rect 915 10 960 90
rect 840 0 960 10
rect 1160 90 1280 100
rect 1160 10 1205 90
rect 1235 10 1280 90
rect 1160 0 1280 10
rect 1480 90 1600 100
rect 1480 10 1525 90
rect 1555 10 1600 90
rect 1480 0 1600 10
rect 1800 90 1920 100
rect 1800 10 1845 90
rect 1875 10 1920 90
rect 1800 0 1920 10
rect 2120 90 2240 100
rect 2120 10 2165 90
rect 2195 10 2240 90
rect 2120 0 2240 10
rect 2440 90 2560 100
rect 2440 10 2485 90
rect 2515 10 2560 90
rect 2440 0 2560 10
rect 2760 90 2880 100
rect 2760 10 2805 90
rect 2835 10 2880 90
rect 2760 0 2880 10
rect 3080 90 3200 100
rect 3080 10 3125 90
rect 3155 10 3200 90
rect 3080 0 3200 10
rect 3400 90 3520 100
rect 3400 10 3445 90
rect 3475 10 3520 90
rect 3400 0 3520 10
rect 3720 90 3840 100
rect 3720 10 3765 90
rect 3795 10 3840 90
rect 3720 0 3840 10
rect 4040 90 4160 100
rect 4040 10 4085 90
rect 4115 10 4160 90
rect 4040 0 4160 10
rect 4360 90 4480 100
rect 4360 10 4405 90
rect 4435 10 4480 90
rect 4360 0 4480 10
rect 4680 90 4800 100
rect 4680 10 4725 90
rect 4755 10 4800 90
rect 4680 0 4800 10
rect 5000 90 5080 100
rect 5000 10 5045 90
rect 5075 10 5080 90
rect 5000 0 5080 10
rect 5200 90 5280 100
rect 5200 10 5205 90
rect 5235 10 5280 90
rect 5200 0 5280 10
rect 5480 90 5600 100
rect 5480 10 5525 90
rect 5555 10 5600 90
rect 5480 0 5600 10
rect 5800 90 5920 100
rect 5800 10 5845 90
rect 5875 10 5920 90
rect 5800 0 5920 10
rect 6120 90 6240 100
rect 6120 10 6165 90
rect 6195 10 6240 90
rect 6120 0 6240 10
rect 6440 90 6560 100
rect 6440 10 6485 90
rect 6515 10 6560 90
rect 6440 0 6560 10
rect 6760 90 6880 100
rect 6760 10 6805 90
rect 6835 10 6880 90
rect 6760 0 6880 10
rect 7080 90 7200 100
rect 7080 10 7125 90
rect 7155 10 7200 90
rect 7080 0 7200 10
rect 7400 90 7520 100
rect 7400 10 7445 90
rect 7475 10 7520 90
rect 7400 0 7520 10
rect 7720 90 7840 100
rect 7720 10 7765 90
rect 7795 10 7840 90
rect 7720 0 7840 10
rect 8040 90 8160 100
rect 8040 10 8085 90
rect 8115 10 8160 90
rect 8040 0 8160 10
rect 8360 90 8480 100
rect 8360 10 8405 90
rect 8435 10 8480 90
rect 8360 0 8480 10
rect 8680 90 8800 100
rect 8680 10 8725 90
rect 8755 10 8800 90
rect 8680 0 8800 10
rect 9000 90 9120 100
rect 9000 10 9045 90
rect 9075 10 9120 90
rect 9000 0 9120 10
rect 9320 90 9440 100
rect 9320 10 9365 90
rect 9395 10 9440 90
rect 9320 0 9440 10
rect 9640 90 9760 100
rect 9640 10 9685 90
rect 9715 10 9760 90
rect 9640 0 9760 10
rect 9960 90 10080 100
rect 9960 10 10005 90
rect 10035 10 10080 90
rect 9960 0 10080 10
rect 10280 90 10360 100
rect 10280 10 10325 90
rect 10355 10 10360 90
rect 10280 0 10360 10
rect -80 -290 0 -280
rect -80 -370 -75 -290
rect -45 -370 0 -290
rect -80 -380 0 -370
rect 200 -290 320 -280
rect 200 -370 245 -290
rect 275 -370 320 -290
rect 200 -380 320 -370
rect 520 -290 640 -280
rect 520 -370 565 -290
rect 595 -370 640 -290
rect 520 -380 640 -370
rect 840 -290 960 -280
rect 840 -370 885 -290
rect 915 -370 960 -290
rect 840 -380 960 -370
rect 1160 -290 1280 -280
rect 1160 -370 1205 -290
rect 1235 -370 1280 -290
rect 1160 -380 1280 -370
rect 1480 -290 1600 -280
rect 1480 -370 1525 -290
rect 1555 -370 1600 -290
rect 1480 -380 1600 -370
rect 1800 -290 1920 -280
rect 1800 -370 1845 -290
rect 1875 -370 1920 -290
rect 1800 -380 1920 -370
rect 2120 -290 2240 -280
rect 2120 -370 2165 -290
rect 2195 -370 2240 -290
rect 2120 -380 2240 -370
rect 2440 -290 2560 -280
rect 2440 -370 2485 -290
rect 2515 -370 2560 -290
rect 2440 -380 2560 -370
rect 2760 -290 2880 -280
rect 2760 -370 2805 -290
rect 2835 -370 2880 -290
rect 2760 -380 2880 -370
rect 3080 -290 3200 -280
rect 3080 -370 3125 -290
rect 3155 -370 3200 -290
rect 3080 -380 3200 -370
rect 3400 -290 3520 -280
rect 3400 -370 3445 -290
rect 3475 -370 3520 -290
rect 3400 -380 3520 -370
rect 3720 -290 3840 -280
rect 3720 -370 3765 -290
rect 3795 -370 3840 -290
rect 3720 -380 3840 -370
rect 4040 -290 4160 -280
rect 4040 -370 4085 -290
rect 4115 -370 4160 -290
rect 4040 -380 4160 -370
rect 4360 -290 4480 -280
rect 4360 -370 4405 -290
rect 4435 -370 4480 -290
rect 4360 -380 4480 -370
rect 4680 -290 4800 -280
rect 4680 -370 4725 -290
rect 4755 -370 4800 -290
rect 4680 -380 4800 -370
rect 5000 -290 5080 -280
rect 5000 -370 5045 -290
rect 5075 -370 5080 -290
rect 5000 -380 5080 -370
rect 5200 -290 5280 -280
rect 5200 -370 5205 -290
rect 5235 -370 5280 -290
rect 5200 -380 5280 -370
rect 5480 -290 5600 -280
rect 5480 -370 5525 -290
rect 5555 -370 5600 -290
rect 5480 -380 5600 -370
rect 5800 -290 5920 -280
rect 5800 -370 5845 -290
rect 5875 -370 5920 -290
rect 5800 -380 5920 -370
rect 6120 -290 6240 -280
rect 6120 -370 6165 -290
rect 6195 -370 6240 -290
rect 6120 -380 6240 -370
rect 6440 -290 6560 -280
rect 6440 -370 6485 -290
rect 6515 -370 6560 -290
rect 6440 -380 6560 -370
rect 6760 -290 6880 -280
rect 6760 -370 6805 -290
rect 6835 -370 6880 -290
rect 6760 -380 6880 -370
rect 7080 -290 7200 -280
rect 7080 -370 7125 -290
rect 7155 -370 7200 -290
rect 7080 -380 7200 -370
rect 7400 -290 7520 -280
rect 7400 -370 7445 -290
rect 7475 -370 7520 -290
rect 7400 -380 7520 -370
rect 7720 -290 7840 -280
rect 7720 -370 7765 -290
rect 7795 -370 7840 -290
rect 7720 -380 7840 -370
rect 8040 -290 8160 -280
rect 8040 -370 8085 -290
rect 8115 -370 8160 -290
rect 8040 -380 8160 -370
rect 8360 -290 8480 -280
rect 8360 -370 8405 -290
rect 8435 -370 8480 -290
rect 8360 -380 8480 -370
rect 8680 -290 8800 -280
rect 8680 -370 8725 -290
rect 8755 -370 8800 -290
rect 8680 -380 8800 -370
rect 9000 -290 9120 -280
rect 9000 -370 9045 -290
rect 9075 -370 9120 -290
rect 9000 -380 9120 -370
rect 9320 -290 9440 -280
rect 9320 -370 9365 -290
rect 9395 -370 9440 -290
rect 9320 -380 9440 -370
rect 9640 -290 9760 -280
rect 9640 -370 9685 -290
rect 9715 -370 9760 -290
rect 9640 -380 9760 -370
rect 9960 -290 10080 -280
rect 9960 -370 10005 -290
rect 10035 -370 10080 -290
rect 9960 -380 10080 -370
rect 10280 -290 10360 -280
rect 10280 -370 10325 -290
rect 10355 -370 10360 -290
rect 10280 -380 10360 -370
rect -80 -2310 0 -2300
rect -80 -2390 -75 -2310
rect -45 -2390 0 -2310
rect -80 -2400 0 -2390
rect 200 -2310 320 -2300
rect 200 -2390 245 -2310
rect 275 -2390 320 -2310
rect 200 -2400 320 -2390
rect 520 -2310 640 -2300
rect 520 -2390 565 -2310
rect 595 -2390 640 -2310
rect 520 -2400 640 -2390
rect 840 -2310 960 -2300
rect 840 -2390 885 -2310
rect 915 -2390 960 -2310
rect 840 -2400 960 -2390
rect 1160 -2310 1280 -2300
rect 1160 -2390 1205 -2310
rect 1235 -2390 1280 -2310
rect 1160 -2400 1280 -2390
rect 1480 -2310 1600 -2300
rect 1480 -2390 1525 -2310
rect 1555 -2390 1600 -2310
rect 1480 -2400 1600 -2390
rect 1800 -2310 1920 -2300
rect 1800 -2390 1845 -2310
rect 1875 -2390 1920 -2310
rect 1800 -2400 1920 -2390
rect 2120 -2310 2240 -2300
rect 2120 -2390 2165 -2310
rect 2195 -2390 2240 -2310
rect 2120 -2400 2240 -2390
rect 2440 -2310 2560 -2300
rect 2440 -2390 2485 -2310
rect 2515 -2390 2560 -2310
rect 2440 -2400 2560 -2390
rect 2760 -2310 2880 -2300
rect 2760 -2390 2805 -2310
rect 2835 -2390 2880 -2310
rect 2760 -2400 2880 -2390
rect 3080 -2310 3200 -2300
rect 3080 -2390 3125 -2310
rect 3155 -2390 3200 -2310
rect 3080 -2400 3200 -2390
rect 3400 -2310 3520 -2300
rect 3400 -2390 3445 -2310
rect 3475 -2390 3520 -2310
rect 3400 -2400 3520 -2390
rect 3720 -2310 3840 -2300
rect 3720 -2390 3765 -2310
rect 3795 -2390 3840 -2310
rect 3720 -2400 3840 -2390
rect 4040 -2310 4160 -2300
rect 4040 -2390 4085 -2310
rect 4115 -2390 4160 -2310
rect 4040 -2400 4160 -2390
rect 4360 -2310 4480 -2300
rect 4360 -2390 4405 -2310
rect 4435 -2390 4480 -2310
rect 4360 -2400 4480 -2390
rect 4680 -2310 4800 -2300
rect 4680 -2390 4725 -2310
rect 4755 -2390 4800 -2310
rect 4680 -2400 4800 -2390
rect 5000 -2310 5080 -2300
rect 5000 -2390 5045 -2310
rect 5075 -2390 5080 -2310
rect 5000 -2400 5080 -2390
rect 5200 -2310 5280 -2300
rect 5200 -2390 5205 -2310
rect 5235 -2390 5280 -2310
rect 5200 -2400 5280 -2390
rect 5480 -2310 5600 -2300
rect 5480 -2390 5525 -2310
rect 5555 -2390 5600 -2310
rect 5480 -2400 5600 -2390
rect 5800 -2310 5920 -2300
rect 5800 -2390 5845 -2310
rect 5875 -2390 5920 -2310
rect 5800 -2400 5920 -2390
rect 6120 -2310 6240 -2300
rect 6120 -2390 6165 -2310
rect 6195 -2390 6240 -2310
rect 6120 -2400 6240 -2390
rect 6440 -2310 6560 -2300
rect 6440 -2390 6485 -2310
rect 6515 -2390 6560 -2310
rect 6440 -2400 6560 -2390
rect 6760 -2310 6880 -2300
rect 6760 -2390 6805 -2310
rect 6835 -2390 6880 -2310
rect 6760 -2400 6880 -2390
rect 7080 -2310 7200 -2300
rect 7080 -2390 7125 -2310
rect 7155 -2390 7200 -2310
rect 7080 -2400 7200 -2390
rect 7400 -2310 7520 -2300
rect 7400 -2390 7445 -2310
rect 7475 -2390 7520 -2310
rect 7400 -2400 7520 -2390
rect 7720 -2310 7840 -2300
rect 7720 -2390 7765 -2310
rect 7795 -2390 7840 -2310
rect 7720 -2400 7840 -2390
rect 8040 -2310 8160 -2300
rect 8040 -2390 8085 -2310
rect 8115 -2390 8160 -2310
rect 8040 -2400 8160 -2390
rect 8360 -2310 8480 -2300
rect 8360 -2390 8405 -2310
rect 8435 -2390 8480 -2310
rect 8360 -2400 8480 -2390
rect 8680 -2310 8800 -2300
rect 8680 -2390 8725 -2310
rect 8755 -2390 8800 -2310
rect 8680 -2400 8800 -2390
rect 9000 -2310 9120 -2300
rect 9000 -2390 9045 -2310
rect 9075 -2390 9120 -2310
rect 9000 -2400 9120 -2390
rect 9320 -2310 9440 -2300
rect 9320 -2390 9365 -2310
rect 9395 -2390 9440 -2310
rect 9320 -2400 9440 -2390
rect 9640 -2310 9760 -2300
rect 9640 -2390 9685 -2310
rect 9715 -2390 9760 -2310
rect 9640 -2400 9760 -2390
rect 9960 -2310 10080 -2300
rect 9960 -2390 10005 -2310
rect 10035 -2390 10080 -2310
rect 9960 -2400 10080 -2390
rect 10280 -2310 10360 -2300
rect 10280 -2390 10325 -2310
rect 10355 -2390 10360 -2310
rect 10280 -2400 10360 -2390
rect -80 -2690 0 -2680
rect -80 -2770 -75 -2690
rect -45 -2770 0 -2690
rect -80 -2780 0 -2770
rect 200 -2690 320 -2680
rect 200 -2770 245 -2690
rect 275 -2770 320 -2690
rect 200 -2780 320 -2770
rect 520 -2690 640 -2680
rect 520 -2770 565 -2690
rect 595 -2770 640 -2690
rect 520 -2780 640 -2770
rect 840 -2690 960 -2680
rect 840 -2770 885 -2690
rect 915 -2770 960 -2690
rect 840 -2780 960 -2770
rect 1160 -2690 1280 -2680
rect 1160 -2770 1205 -2690
rect 1235 -2770 1280 -2690
rect 1160 -2780 1280 -2770
rect 1480 -2690 1600 -2680
rect 1480 -2770 1525 -2690
rect 1555 -2770 1600 -2690
rect 1480 -2780 1600 -2770
rect 1800 -2690 1920 -2680
rect 1800 -2770 1845 -2690
rect 1875 -2770 1920 -2690
rect 1800 -2780 1920 -2770
rect 2120 -2690 2240 -2680
rect 2120 -2770 2165 -2690
rect 2195 -2770 2240 -2690
rect 2120 -2780 2240 -2770
rect 2440 -2690 2560 -2680
rect 2440 -2770 2485 -2690
rect 2515 -2770 2560 -2690
rect 2440 -2780 2560 -2770
rect 2760 -2690 2880 -2680
rect 2760 -2770 2805 -2690
rect 2835 -2770 2880 -2690
rect 2760 -2780 2880 -2770
rect 3080 -2690 3200 -2680
rect 3080 -2770 3125 -2690
rect 3155 -2770 3200 -2690
rect 3080 -2780 3200 -2770
rect 3400 -2690 3520 -2680
rect 3400 -2770 3445 -2690
rect 3475 -2770 3520 -2690
rect 3400 -2780 3520 -2770
rect 3720 -2690 3840 -2680
rect 3720 -2770 3765 -2690
rect 3795 -2770 3840 -2690
rect 3720 -2780 3840 -2770
rect 4040 -2690 4160 -2680
rect 4040 -2770 4085 -2690
rect 4115 -2770 4160 -2690
rect 4040 -2780 4160 -2770
rect 4360 -2690 4480 -2680
rect 4360 -2770 4405 -2690
rect 4435 -2770 4480 -2690
rect 4360 -2780 4480 -2770
rect 4680 -2690 4800 -2680
rect 4680 -2770 4725 -2690
rect 4755 -2770 4800 -2690
rect 4680 -2780 4800 -2770
rect 5000 -2690 5080 -2680
rect 5000 -2770 5045 -2690
rect 5075 -2770 5080 -2690
rect 5000 -2780 5080 -2770
rect 5200 -2690 5280 -2680
rect 5200 -2770 5205 -2690
rect 5235 -2770 5280 -2690
rect 5200 -2780 5280 -2770
rect 5480 -2690 5600 -2680
rect 5480 -2770 5525 -2690
rect 5555 -2770 5600 -2690
rect 5480 -2780 5600 -2770
rect 5800 -2690 5920 -2680
rect 5800 -2770 5845 -2690
rect 5875 -2770 5920 -2690
rect 5800 -2780 5920 -2770
rect 6120 -2690 6240 -2680
rect 6120 -2770 6165 -2690
rect 6195 -2770 6240 -2690
rect 6120 -2780 6240 -2770
rect 6440 -2690 6560 -2680
rect 6440 -2770 6485 -2690
rect 6515 -2770 6560 -2690
rect 6440 -2780 6560 -2770
rect 6760 -2690 6880 -2680
rect 6760 -2770 6805 -2690
rect 6835 -2770 6880 -2690
rect 6760 -2780 6880 -2770
rect 7080 -2690 7200 -2680
rect 7080 -2770 7125 -2690
rect 7155 -2770 7200 -2690
rect 7080 -2780 7200 -2770
rect 7400 -2690 7520 -2680
rect 7400 -2770 7445 -2690
rect 7475 -2770 7520 -2690
rect 7400 -2780 7520 -2770
rect 7720 -2690 7840 -2680
rect 7720 -2770 7765 -2690
rect 7795 -2770 7840 -2690
rect 7720 -2780 7840 -2770
rect 8040 -2690 8160 -2680
rect 8040 -2770 8085 -2690
rect 8115 -2770 8160 -2690
rect 8040 -2780 8160 -2770
rect 8360 -2690 8480 -2680
rect 8360 -2770 8405 -2690
rect 8435 -2770 8480 -2690
rect 8360 -2780 8480 -2770
rect 8680 -2690 8800 -2680
rect 8680 -2770 8725 -2690
rect 8755 -2770 8800 -2690
rect 8680 -2780 8800 -2770
rect 9000 -2690 9120 -2680
rect 9000 -2770 9045 -2690
rect 9075 -2770 9120 -2690
rect 9000 -2780 9120 -2770
rect 9320 -2690 9440 -2680
rect 9320 -2770 9365 -2690
rect 9395 -2770 9440 -2690
rect 9320 -2780 9440 -2770
rect 9640 -2690 9760 -2680
rect 9640 -2770 9685 -2690
rect 9715 -2770 9760 -2690
rect 9640 -2780 9760 -2770
rect 9960 -2690 10080 -2680
rect 9960 -2770 10005 -2690
rect 10035 -2770 10080 -2690
rect 9960 -2780 10080 -2770
rect 10280 -2690 10360 -2680
rect 10280 -2770 10325 -2690
rect 10355 -2770 10360 -2690
rect 10280 -2780 10360 -2770
<< pdiff >>
rect -80 750 0 760
rect -80 670 -75 750
rect -45 670 0 750
rect -80 660 0 670
rect 200 750 320 760
rect 200 670 245 750
rect 275 670 320 750
rect 200 660 320 670
rect 520 750 640 760
rect 520 670 565 750
rect 595 670 640 750
rect 520 660 640 670
rect 840 750 960 760
rect 840 670 885 750
rect 915 670 960 750
rect 840 660 960 670
rect 1160 750 1280 760
rect 1160 670 1205 750
rect 1235 670 1280 750
rect 1160 660 1280 670
rect 1480 750 1600 760
rect 1480 670 1525 750
rect 1555 670 1600 750
rect 1480 660 1600 670
rect 1800 750 1920 760
rect 1800 670 1845 750
rect 1875 670 1920 750
rect 1800 660 1920 670
rect 2120 750 2240 760
rect 2120 670 2165 750
rect 2195 670 2240 750
rect 2120 660 2240 670
rect 2440 750 2560 760
rect 2440 670 2485 750
rect 2515 670 2560 750
rect 2440 660 2560 670
rect 2760 750 2880 760
rect 2760 670 2805 750
rect 2835 670 2880 750
rect 2760 660 2880 670
rect 3080 750 3200 760
rect 3080 670 3125 750
rect 3155 670 3200 750
rect 3080 660 3200 670
rect 3400 750 3520 760
rect 3400 670 3445 750
rect 3475 670 3520 750
rect 3400 660 3520 670
rect 3720 750 3840 760
rect 3720 670 3765 750
rect 3795 670 3840 750
rect 3720 660 3840 670
rect 4040 750 4160 760
rect 4040 670 4085 750
rect 4115 670 4160 750
rect 4040 660 4160 670
rect 4360 750 4480 760
rect 4360 670 4405 750
rect 4435 670 4480 750
rect 4360 660 4480 670
rect 4680 750 4800 760
rect 4680 670 4725 750
rect 4755 670 4800 750
rect 4680 660 4800 670
rect 5000 750 5080 760
rect 5000 670 5045 750
rect 5075 670 5080 750
rect 5000 660 5080 670
rect 5200 750 5280 760
rect 5200 670 5205 750
rect 5235 670 5280 750
rect 5200 660 5280 670
rect 5480 750 5600 760
rect 5480 670 5525 750
rect 5555 670 5600 750
rect 5480 660 5600 670
rect 5800 750 5920 760
rect 5800 670 5845 750
rect 5875 670 5920 750
rect 5800 660 5920 670
rect 6120 750 6240 760
rect 6120 670 6165 750
rect 6195 670 6240 750
rect 6120 660 6240 670
rect 6440 750 6560 760
rect 6440 670 6485 750
rect 6515 670 6560 750
rect 6440 660 6560 670
rect 6760 750 6880 760
rect 6760 670 6805 750
rect 6835 670 6880 750
rect 6760 660 6880 670
rect 7080 750 7200 760
rect 7080 670 7125 750
rect 7155 670 7200 750
rect 7080 660 7200 670
rect 7400 750 7520 760
rect 7400 670 7445 750
rect 7475 670 7520 750
rect 7400 660 7520 670
rect 7720 750 7840 760
rect 7720 670 7765 750
rect 7795 670 7840 750
rect 7720 660 7840 670
rect 8040 750 8160 760
rect 8040 670 8085 750
rect 8115 670 8160 750
rect 8040 660 8160 670
rect 8360 750 8480 760
rect 8360 670 8405 750
rect 8435 670 8480 750
rect 8360 660 8480 670
rect 8680 750 8800 760
rect 8680 670 8725 750
rect 8755 670 8800 750
rect 8680 660 8800 670
rect 9000 750 9120 760
rect 9000 670 9045 750
rect 9075 670 9120 750
rect 9000 660 9120 670
rect 9320 750 9440 760
rect 9320 670 9365 750
rect 9395 670 9440 750
rect 9320 660 9440 670
rect 9640 750 9760 760
rect 9640 670 9685 750
rect 9715 670 9760 750
rect 9640 660 9760 670
rect 9960 750 10080 760
rect 9960 670 10005 750
rect 10035 670 10080 750
rect 9960 660 10080 670
rect 10280 750 10360 760
rect 10280 670 10325 750
rect 10355 670 10360 750
rect 10280 660 10360 670
rect -80 -950 0 -940
rect -80 -1030 -75 -950
rect -45 -1030 0 -950
rect -80 -1040 0 -1030
rect 200 -950 320 -940
rect 200 -1030 245 -950
rect 275 -1030 320 -950
rect 200 -1040 320 -1030
rect 520 -950 640 -940
rect 520 -1030 565 -950
rect 595 -1030 640 -950
rect 520 -1040 640 -1030
rect 840 -950 960 -940
rect 840 -1030 885 -950
rect 915 -1030 960 -950
rect 840 -1040 960 -1030
rect 1160 -950 1280 -940
rect 1160 -1030 1205 -950
rect 1235 -1030 1280 -950
rect 1160 -1040 1280 -1030
rect 1480 -950 1600 -940
rect 1480 -1030 1525 -950
rect 1555 -1030 1600 -950
rect 1480 -1040 1600 -1030
rect 1800 -950 1920 -940
rect 1800 -1030 1845 -950
rect 1875 -1030 1920 -950
rect 1800 -1040 1920 -1030
rect 2120 -950 2240 -940
rect 2120 -1030 2165 -950
rect 2195 -1030 2240 -950
rect 2120 -1040 2240 -1030
rect 2440 -950 2560 -940
rect 2440 -1030 2485 -950
rect 2515 -1030 2560 -950
rect 2440 -1040 2560 -1030
rect 2760 -950 2880 -940
rect 2760 -1030 2805 -950
rect 2835 -1030 2880 -950
rect 2760 -1040 2880 -1030
rect 3080 -950 3200 -940
rect 3080 -1030 3125 -950
rect 3155 -1030 3200 -950
rect 3080 -1040 3200 -1030
rect 3400 -950 3520 -940
rect 3400 -1030 3445 -950
rect 3475 -1030 3520 -950
rect 3400 -1040 3520 -1030
rect 3720 -950 3840 -940
rect 3720 -1030 3765 -950
rect 3795 -1030 3840 -950
rect 3720 -1040 3840 -1030
rect 4040 -950 4160 -940
rect 4040 -1030 4085 -950
rect 4115 -1030 4160 -950
rect 4040 -1040 4160 -1030
rect 4360 -950 4480 -940
rect 4360 -1030 4405 -950
rect 4435 -1030 4480 -950
rect 4360 -1040 4480 -1030
rect 4680 -950 4800 -940
rect 4680 -1030 4725 -950
rect 4755 -1030 4800 -950
rect 4680 -1040 4800 -1030
rect 5000 -950 5080 -940
rect 5000 -1030 5045 -950
rect 5075 -1030 5080 -950
rect 5000 -1040 5080 -1030
rect 5200 -950 5280 -940
rect 5200 -1030 5205 -950
rect 5235 -1030 5280 -950
rect 5200 -1040 5280 -1030
rect 5480 -950 5600 -940
rect 5480 -1030 5525 -950
rect 5555 -1030 5600 -950
rect 5480 -1040 5600 -1030
rect 5800 -950 5920 -940
rect 5800 -1030 5845 -950
rect 5875 -1030 5920 -950
rect 5800 -1040 5920 -1030
rect 6120 -950 6240 -940
rect 6120 -1030 6165 -950
rect 6195 -1030 6240 -950
rect 6120 -1040 6240 -1030
rect 6440 -950 6560 -940
rect 6440 -1030 6485 -950
rect 6515 -1030 6560 -950
rect 6440 -1040 6560 -1030
rect 6760 -950 6880 -940
rect 6760 -1030 6805 -950
rect 6835 -1030 6880 -950
rect 6760 -1040 6880 -1030
rect 7080 -950 7200 -940
rect 7080 -1030 7125 -950
rect 7155 -1030 7200 -950
rect 7080 -1040 7200 -1030
rect 7400 -950 7520 -940
rect 7400 -1030 7445 -950
rect 7475 -1030 7520 -950
rect 7400 -1040 7520 -1030
rect 7720 -950 7840 -940
rect 7720 -1030 7765 -950
rect 7795 -1030 7840 -950
rect 7720 -1040 7840 -1030
rect 8040 -950 8160 -940
rect 8040 -1030 8085 -950
rect 8115 -1030 8160 -950
rect 8040 -1040 8160 -1030
rect 8360 -950 8480 -940
rect 8360 -1030 8405 -950
rect 8435 -1030 8480 -950
rect 8360 -1040 8480 -1030
rect 8680 -950 8800 -940
rect 8680 -1030 8725 -950
rect 8755 -1030 8800 -950
rect 8680 -1040 8800 -1030
rect 9000 -950 9120 -940
rect 9000 -1030 9045 -950
rect 9075 -1030 9120 -950
rect 9000 -1040 9120 -1030
rect 9320 -950 9440 -940
rect 9320 -1030 9365 -950
rect 9395 -1030 9440 -950
rect 9320 -1040 9440 -1030
rect 9640 -950 9760 -940
rect 9640 -1030 9685 -950
rect 9715 -1030 9760 -950
rect 9640 -1040 9760 -1030
rect 9960 -950 10080 -940
rect 9960 -1030 10005 -950
rect 10035 -1030 10080 -950
rect 9960 -1040 10080 -1030
rect 10280 -950 10360 -940
rect 10280 -1030 10325 -950
rect 10355 -1030 10360 -950
rect 10280 -1040 10360 -1030
rect -80 -1650 0 -1640
rect -80 -1730 -75 -1650
rect -45 -1730 0 -1650
rect -80 -1740 0 -1730
rect 200 -1650 320 -1640
rect 200 -1730 245 -1650
rect 275 -1730 320 -1650
rect 200 -1740 320 -1730
rect 520 -1650 640 -1640
rect 520 -1730 565 -1650
rect 595 -1730 640 -1650
rect 520 -1740 640 -1730
rect 840 -1650 960 -1640
rect 840 -1730 885 -1650
rect 915 -1730 960 -1650
rect 840 -1740 960 -1730
rect 1160 -1650 1280 -1640
rect 1160 -1730 1205 -1650
rect 1235 -1730 1280 -1650
rect 1160 -1740 1280 -1730
rect 1480 -1650 1600 -1640
rect 1480 -1730 1525 -1650
rect 1555 -1730 1600 -1650
rect 1480 -1740 1600 -1730
rect 1800 -1650 1920 -1640
rect 1800 -1730 1845 -1650
rect 1875 -1730 1920 -1650
rect 1800 -1740 1920 -1730
rect 2120 -1650 2240 -1640
rect 2120 -1730 2165 -1650
rect 2195 -1730 2240 -1650
rect 2120 -1740 2240 -1730
rect 2440 -1650 2560 -1640
rect 2440 -1730 2485 -1650
rect 2515 -1730 2560 -1650
rect 2440 -1740 2560 -1730
rect 2760 -1650 2880 -1640
rect 2760 -1730 2805 -1650
rect 2835 -1730 2880 -1650
rect 2760 -1740 2880 -1730
rect 3080 -1650 3200 -1640
rect 3080 -1730 3125 -1650
rect 3155 -1730 3200 -1650
rect 3080 -1740 3200 -1730
rect 3400 -1650 3520 -1640
rect 3400 -1730 3445 -1650
rect 3475 -1730 3520 -1650
rect 3400 -1740 3520 -1730
rect 3720 -1650 3840 -1640
rect 3720 -1730 3765 -1650
rect 3795 -1730 3840 -1650
rect 3720 -1740 3840 -1730
rect 4040 -1650 4160 -1640
rect 4040 -1730 4085 -1650
rect 4115 -1730 4160 -1650
rect 4040 -1740 4160 -1730
rect 4360 -1650 4480 -1640
rect 4360 -1730 4405 -1650
rect 4435 -1730 4480 -1650
rect 4360 -1740 4480 -1730
rect 4680 -1650 4800 -1640
rect 4680 -1730 4725 -1650
rect 4755 -1730 4800 -1650
rect 4680 -1740 4800 -1730
rect 5000 -1650 5080 -1640
rect 5000 -1730 5045 -1650
rect 5075 -1730 5080 -1650
rect 5000 -1740 5080 -1730
rect 5200 -1650 5280 -1640
rect 5200 -1730 5205 -1650
rect 5235 -1730 5280 -1650
rect 5200 -1740 5280 -1730
rect 5480 -1650 5600 -1640
rect 5480 -1730 5525 -1650
rect 5555 -1730 5600 -1650
rect 5480 -1740 5600 -1730
rect 5800 -1650 5920 -1640
rect 5800 -1730 5845 -1650
rect 5875 -1730 5920 -1650
rect 5800 -1740 5920 -1730
rect 6120 -1650 6240 -1640
rect 6120 -1730 6165 -1650
rect 6195 -1730 6240 -1650
rect 6120 -1740 6240 -1730
rect 6440 -1650 6560 -1640
rect 6440 -1730 6485 -1650
rect 6515 -1730 6560 -1650
rect 6440 -1740 6560 -1730
rect 6760 -1650 6880 -1640
rect 6760 -1730 6805 -1650
rect 6835 -1730 6880 -1650
rect 6760 -1740 6880 -1730
rect 7080 -1650 7200 -1640
rect 7080 -1730 7125 -1650
rect 7155 -1730 7200 -1650
rect 7080 -1740 7200 -1730
rect 7400 -1650 7520 -1640
rect 7400 -1730 7445 -1650
rect 7475 -1730 7520 -1650
rect 7400 -1740 7520 -1730
rect 7720 -1650 7840 -1640
rect 7720 -1730 7765 -1650
rect 7795 -1730 7840 -1650
rect 7720 -1740 7840 -1730
rect 8040 -1650 8160 -1640
rect 8040 -1730 8085 -1650
rect 8115 -1730 8160 -1650
rect 8040 -1740 8160 -1730
rect 8360 -1650 8480 -1640
rect 8360 -1730 8405 -1650
rect 8435 -1730 8480 -1650
rect 8360 -1740 8480 -1730
rect 8680 -1650 8800 -1640
rect 8680 -1730 8725 -1650
rect 8755 -1730 8800 -1650
rect 8680 -1740 8800 -1730
rect 9000 -1650 9120 -1640
rect 9000 -1730 9045 -1650
rect 9075 -1730 9120 -1650
rect 9000 -1740 9120 -1730
rect 9320 -1650 9440 -1640
rect 9320 -1730 9365 -1650
rect 9395 -1730 9440 -1650
rect 9320 -1740 9440 -1730
rect 9640 -1650 9760 -1640
rect 9640 -1730 9685 -1650
rect 9715 -1730 9760 -1650
rect 9640 -1740 9760 -1730
rect 9960 -1650 10080 -1640
rect 9960 -1730 10005 -1650
rect 10035 -1730 10080 -1650
rect 9960 -1740 10080 -1730
rect 10280 -1650 10360 -1640
rect 10280 -1730 10325 -1650
rect 10355 -1730 10360 -1650
rect 10280 -1740 10360 -1730
rect -80 -3350 0 -3340
rect -80 -3430 -75 -3350
rect -45 -3430 0 -3350
rect -80 -3440 0 -3430
rect 200 -3350 320 -3340
rect 200 -3430 245 -3350
rect 275 -3430 320 -3350
rect 200 -3440 320 -3430
rect 520 -3350 640 -3340
rect 520 -3430 565 -3350
rect 595 -3430 640 -3350
rect 520 -3440 640 -3430
rect 840 -3350 960 -3340
rect 840 -3430 885 -3350
rect 915 -3430 960 -3350
rect 840 -3440 960 -3430
rect 1160 -3350 1280 -3340
rect 1160 -3430 1205 -3350
rect 1235 -3430 1280 -3350
rect 1160 -3440 1280 -3430
rect 1480 -3350 1600 -3340
rect 1480 -3430 1525 -3350
rect 1555 -3430 1600 -3350
rect 1480 -3440 1600 -3430
rect 1800 -3350 1920 -3340
rect 1800 -3430 1845 -3350
rect 1875 -3430 1920 -3350
rect 1800 -3440 1920 -3430
rect 2120 -3350 2240 -3340
rect 2120 -3430 2165 -3350
rect 2195 -3430 2240 -3350
rect 2120 -3440 2240 -3430
rect 2440 -3350 2560 -3340
rect 2440 -3430 2485 -3350
rect 2515 -3430 2560 -3350
rect 2440 -3440 2560 -3430
rect 2760 -3350 2880 -3340
rect 2760 -3430 2805 -3350
rect 2835 -3430 2880 -3350
rect 2760 -3440 2880 -3430
rect 3080 -3350 3200 -3340
rect 3080 -3430 3125 -3350
rect 3155 -3430 3200 -3350
rect 3080 -3440 3200 -3430
rect 3400 -3350 3520 -3340
rect 3400 -3430 3445 -3350
rect 3475 -3430 3520 -3350
rect 3400 -3440 3520 -3430
rect 3720 -3350 3840 -3340
rect 3720 -3430 3765 -3350
rect 3795 -3430 3840 -3350
rect 3720 -3440 3840 -3430
rect 4040 -3350 4160 -3340
rect 4040 -3430 4085 -3350
rect 4115 -3430 4160 -3350
rect 4040 -3440 4160 -3430
rect 4360 -3350 4480 -3340
rect 4360 -3430 4405 -3350
rect 4435 -3430 4480 -3350
rect 4360 -3440 4480 -3430
rect 4680 -3350 4800 -3340
rect 4680 -3430 4725 -3350
rect 4755 -3430 4800 -3350
rect 4680 -3440 4800 -3430
rect 5000 -3350 5080 -3340
rect 5000 -3430 5045 -3350
rect 5075 -3430 5080 -3350
rect 5000 -3440 5080 -3430
rect 5200 -3350 5280 -3340
rect 5200 -3430 5205 -3350
rect 5235 -3430 5280 -3350
rect 5200 -3440 5280 -3430
rect 5480 -3350 5600 -3340
rect 5480 -3430 5525 -3350
rect 5555 -3430 5600 -3350
rect 5480 -3440 5600 -3430
rect 5800 -3350 5920 -3340
rect 5800 -3430 5845 -3350
rect 5875 -3430 5920 -3350
rect 5800 -3440 5920 -3430
rect 6120 -3350 6240 -3340
rect 6120 -3430 6165 -3350
rect 6195 -3430 6240 -3350
rect 6120 -3440 6240 -3430
rect 6440 -3350 6560 -3340
rect 6440 -3430 6485 -3350
rect 6515 -3430 6560 -3350
rect 6440 -3440 6560 -3430
rect 6760 -3350 6880 -3340
rect 6760 -3430 6805 -3350
rect 6835 -3430 6880 -3350
rect 6760 -3440 6880 -3430
rect 7080 -3350 7200 -3340
rect 7080 -3430 7125 -3350
rect 7155 -3430 7200 -3350
rect 7080 -3440 7200 -3430
rect 7400 -3350 7520 -3340
rect 7400 -3430 7445 -3350
rect 7475 -3430 7520 -3350
rect 7400 -3440 7520 -3430
rect 7720 -3350 7840 -3340
rect 7720 -3430 7765 -3350
rect 7795 -3430 7840 -3350
rect 7720 -3440 7840 -3430
rect 8040 -3350 8160 -3340
rect 8040 -3430 8085 -3350
rect 8115 -3430 8160 -3350
rect 8040 -3440 8160 -3430
rect 8360 -3350 8480 -3340
rect 8360 -3430 8405 -3350
rect 8435 -3430 8480 -3350
rect 8360 -3440 8480 -3430
rect 8680 -3350 8800 -3340
rect 8680 -3430 8725 -3350
rect 8755 -3430 8800 -3350
rect 8680 -3440 8800 -3430
rect 9000 -3350 9120 -3340
rect 9000 -3430 9045 -3350
rect 9075 -3430 9120 -3350
rect 9000 -3440 9120 -3430
rect 9320 -3350 9440 -3340
rect 9320 -3430 9365 -3350
rect 9395 -3430 9440 -3350
rect 9320 -3440 9440 -3430
rect 9640 -3350 9760 -3340
rect 9640 -3430 9685 -3350
rect 9715 -3430 9760 -3350
rect 9640 -3440 9760 -3430
rect 9960 -3350 10080 -3340
rect 9960 -3430 10005 -3350
rect 10035 -3430 10080 -3350
rect 9960 -3440 10080 -3430
rect 10280 -3350 10360 -3340
rect 10280 -3430 10325 -3350
rect 10355 -3430 10360 -3350
rect 10280 -3440 10360 -3430
<< ndiffc >>
rect -75 10 -45 90
rect 245 10 275 90
rect 565 10 595 90
rect 885 10 915 90
rect 1205 10 1235 90
rect 1525 10 1555 90
rect 1845 10 1875 90
rect 2165 10 2195 90
rect 2485 10 2515 90
rect 2805 10 2835 90
rect 3125 10 3155 90
rect 3445 10 3475 90
rect 3765 10 3795 90
rect 4085 10 4115 90
rect 4405 10 4435 90
rect 4725 10 4755 90
rect 5045 10 5075 90
rect 5205 10 5235 90
rect 5525 10 5555 90
rect 5845 10 5875 90
rect 6165 10 6195 90
rect 6485 10 6515 90
rect 6805 10 6835 90
rect 7125 10 7155 90
rect 7445 10 7475 90
rect 7765 10 7795 90
rect 8085 10 8115 90
rect 8405 10 8435 90
rect 8725 10 8755 90
rect 9045 10 9075 90
rect 9365 10 9395 90
rect 9685 10 9715 90
rect 10005 10 10035 90
rect 10325 10 10355 90
rect -75 -370 -45 -290
rect 245 -370 275 -290
rect 565 -370 595 -290
rect 885 -370 915 -290
rect 1205 -370 1235 -290
rect 1525 -370 1555 -290
rect 1845 -370 1875 -290
rect 2165 -370 2195 -290
rect 2485 -370 2515 -290
rect 2805 -370 2835 -290
rect 3125 -370 3155 -290
rect 3445 -370 3475 -290
rect 3765 -370 3795 -290
rect 4085 -370 4115 -290
rect 4405 -370 4435 -290
rect 4725 -370 4755 -290
rect 5045 -370 5075 -290
rect 5205 -370 5235 -290
rect 5525 -370 5555 -290
rect 5845 -370 5875 -290
rect 6165 -370 6195 -290
rect 6485 -370 6515 -290
rect 6805 -370 6835 -290
rect 7125 -370 7155 -290
rect 7445 -370 7475 -290
rect 7765 -370 7795 -290
rect 8085 -370 8115 -290
rect 8405 -370 8435 -290
rect 8725 -370 8755 -290
rect 9045 -370 9075 -290
rect 9365 -370 9395 -290
rect 9685 -370 9715 -290
rect 10005 -370 10035 -290
rect 10325 -370 10355 -290
rect -75 -2390 -45 -2310
rect 245 -2390 275 -2310
rect 565 -2390 595 -2310
rect 885 -2390 915 -2310
rect 1205 -2390 1235 -2310
rect 1525 -2390 1555 -2310
rect 1845 -2390 1875 -2310
rect 2165 -2390 2195 -2310
rect 2485 -2390 2515 -2310
rect 2805 -2390 2835 -2310
rect 3125 -2390 3155 -2310
rect 3445 -2390 3475 -2310
rect 3765 -2390 3795 -2310
rect 4085 -2390 4115 -2310
rect 4405 -2390 4435 -2310
rect 4725 -2390 4755 -2310
rect 5045 -2390 5075 -2310
rect 5205 -2390 5235 -2310
rect 5525 -2390 5555 -2310
rect 5845 -2390 5875 -2310
rect 6165 -2390 6195 -2310
rect 6485 -2390 6515 -2310
rect 6805 -2390 6835 -2310
rect 7125 -2390 7155 -2310
rect 7445 -2390 7475 -2310
rect 7765 -2390 7795 -2310
rect 8085 -2390 8115 -2310
rect 8405 -2390 8435 -2310
rect 8725 -2390 8755 -2310
rect 9045 -2390 9075 -2310
rect 9365 -2390 9395 -2310
rect 9685 -2390 9715 -2310
rect 10005 -2390 10035 -2310
rect 10325 -2390 10355 -2310
rect -75 -2770 -45 -2690
rect 245 -2770 275 -2690
rect 565 -2770 595 -2690
rect 885 -2770 915 -2690
rect 1205 -2770 1235 -2690
rect 1525 -2770 1555 -2690
rect 1845 -2770 1875 -2690
rect 2165 -2770 2195 -2690
rect 2485 -2770 2515 -2690
rect 2805 -2770 2835 -2690
rect 3125 -2770 3155 -2690
rect 3445 -2770 3475 -2690
rect 3765 -2770 3795 -2690
rect 4085 -2770 4115 -2690
rect 4405 -2770 4435 -2690
rect 4725 -2770 4755 -2690
rect 5045 -2770 5075 -2690
rect 5205 -2770 5235 -2690
rect 5525 -2770 5555 -2690
rect 5845 -2770 5875 -2690
rect 6165 -2770 6195 -2690
rect 6485 -2770 6515 -2690
rect 6805 -2770 6835 -2690
rect 7125 -2770 7155 -2690
rect 7445 -2770 7475 -2690
rect 7765 -2770 7795 -2690
rect 8085 -2770 8115 -2690
rect 8405 -2770 8435 -2690
rect 8725 -2770 8755 -2690
rect 9045 -2770 9075 -2690
rect 9365 -2770 9395 -2690
rect 9685 -2770 9715 -2690
rect 10005 -2770 10035 -2690
rect 10325 -2770 10355 -2690
<< pdiffc >>
rect -75 670 -45 750
rect 245 670 275 750
rect 565 670 595 750
rect 885 670 915 750
rect 1205 670 1235 750
rect 1525 670 1555 750
rect 1845 670 1875 750
rect 2165 670 2195 750
rect 2485 670 2515 750
rect 2805 670 2835 750
rect 3125 670 3155 750
rect 3445 670 3475 750
rect 3765 670 3795 750
rect 4085 670 4115 750
rect 4405 670 4435 750
rect 4725 670 4755 750
rect 5045 670 5075 750
rect 5205 670 5235 750
rect 5525 670 5555 750
rect 5845 670 5875 750
rect 6165 670 6195 750
rect 6485 670 6515 750
rect 6805 670 6835 750
rect 7125 670 7155 750
rect 7445 670 7475 750
rect 7765 670 7795 750
rect 8085 670 8115 750
rect 8405 670 8435 750
rect 8725 670 8755 750
rect 9045 670 9075 750
rect 9365 670 9395 750
rect 9685 670 9715 750
rect 10005 670 10035 750
rect 10325 670 10355 750
rect -75 -1030 -45 -950
rect 245 -1030 275 -950
rect 565 -1030 595 -950
rect 885 -1030 915 -950
rect 1205 -1030 1235 -950
rect 1525 -1030 1555 -950
rect 1845 -1030 1875 -950
rect 2165 -1030 2195 -950
rect 2485 -1030 2515 -950
rect 2805 -1030 2835 -950
rect 3125 -1030 3155 -950
rect 3445 -1030 3475 -950
rect 3765 -1030 3795 -950
rect 4085 -1030 4115 -950
rect 4405 -1030 4435 -950
rect 4725 -1030 4755 -950
rect 5045 -1030 5075 -950
rect 5205 -1030 5235 -950
rect 5525 -1030 5555 -950
rect 5845 -1030 5875 -950
rect 6165 -1030 6195 -950
rect 6485 -1030 6515 -950
rect 6805 -1030 6835 -950
rect 7125 -1030 7155 -950
rect 7445 -1030 7475 -950
rect 7765 -1030 7795 -950
rect 8085 -1030 8115 -950
rect 8405 -1030 8435 -950
rect 8725 -1030 8755 -950
rect 9045 -1030 9075 -950
rect 9365 -1030 9395 -950
rect 9685 -1030 9715 -950
rect 10005 -1030 10035 -950
rect 10325 -1030 10355 -950
rect -75 -1730 -45 -1650
rect 245 -1730 275 -1650
rect 565 -1730 595 -1650
rect 885 -1730 915 -1650
rect 1205 -1730 1235 -1650
rect 1525 -1730 1555 -1650
rect 1845 -1730 1875 -1650
rect 2165 -1730 2195 -1650
rect 2485 -1730 2515 -1650
rect 2805 -1730 2835 -1650
rect 3125 -1730 3155 -1650
rect 3445 -1730 3475 -1650
rect 3765 -1730 3795 -1650
rect 4085 -1730 4115 -1650
rect 4405 -1730 4435 -1650
rect 4725 -1730 4755 -1650
rect 5045 -1730 5075 -1650
rect 5205 -1730 5235 -1650
rect 5525 -1730 5555 -1650
rect 5845 -1730 5875 -1650
rect 6165 -1730 6195 -1650
rect 6485 -1730 6515 -1650
rect 6805 -1730 6835 -1650
rect 7125 -1730 7155 -1650
rect 7445 -1730 7475 -1650
rect 7765 -1730 7795 -1650
rect 8085 -1730 8115 -1650
rect 8405 -1730 8435 -1650
rect 8725 -1730 8755 -1650
rect 9045 -1730 9075 -1650
rect 9365 -1730 9395 -1650
rect 9685 -1730 9715 -1650
rect 10005 -1730 10035 -1650
rect 10325 -1730 10355 -1650
rect -75 -3430 -45 -3350
rect 245 -3430 275 -3350
rect 565 -3430 595 -3350
rect 885 -3430 915 -3350
rect 1205 -3430 1235 -3350
rect 1525 -3430 1555 -3350
rect 1845 -3430 1875 -3350
rect 2165 -3430 2195 -3350
rect 2485 -3430 2515 -3350
rect 2805 -3430 2835 -3350
rect 3125 -3430 3155 -3350
rect 3445 -3430 3475 -3350
rect 3765 -3430 3795 -3350
rect 4085 -3430 4115 -3350
rect 4405 -3430 4435 -3350
rect 4725 -3430 4755 -3350
rect 5045 -3430 5075 -3350
rect 5205 -3430 5235 -3350
rect 5525 -3430 5555 -3350
rect 5845 -3430 5875 -3350
rect 6165 -3430 6195 -3350
rect 6485 -3430 6515 -3350
rect 6805 -3430 6835 -3350
rect 7125 -3430 7155 -3350
rect 7445 -3430 7475 -3350
rect 7765 -3430 7795 -3350
rect 8085 -3430 8115 -3350
rect 8405 -3430 8435 -3350
rect 8725 -3430 8755 -3350
rect 9045 -3430 9075 -3350
rect 9365 -3430 9395 -3350
rect 9685 -3430 9715 -3350
rect 10005 -3430 10035 -3350
rect 10325 -3430 10355 -3350
<< psubdiff >>
rect -320 1000 -40 1040
rect 240 1000 280 1040
rect 560 1000 600 1040
rect 880 1000 920 1040
rect 1200 1000 1240 1040
rect 1520 1000 1560 1040
rect 1840 1000 1880 1040
rect 2160 1000 2200 1040
rect 2480 1000 2520 1040
rect 2800 1000 2840 1040
rect 3120 1000 3160 1040
rect 3440 1000 3480 1040
rect 3760 1000 3800 1040
rect 4080 1000 4120 1040
rect 4400 1000 4440 1040
rect 4720 1000 4760 1040
rect 5040 1000 5240 1040
rect 5520 1000 5560 1040
rect 5840 1000 5880 1040
rect 6160 1000 6200 1040
rect 6480 1000 6520 1040
rect 6800 1000 6840 1040
rect 7120 1000 7160 1040
rect 7440 1000 7480 1040
rect 7760 1000 7800 1040
rect 8080 1000 8120 1040
rect 8400 1000 8440 1040
rect 8720 1000 8760 1040
rect 9040 1000 9080 1040
rect 9360 1000 9400 1040
rect 9680 1000 9720 1040
rect 10000 1000 10040 1040
rect 10320 1000 10600 1040
rect -320 960 -280 1000
rect 10560 960 10600 1000
rect -280 360 -40 400
rect 240 360 280 400
rect 560 360 600 400
rect 880 360 920 400
rect 1200 360 1240 400
rect 1520 360 1560 400
rect 1840 360 1880 400
rect 2160 360 2200 400
rect 2480 360 2520 400
rect 2800 360 2840 400
rect 3120 360 3160 400
rect 3440 360 3480 400
rect 3760 360 3800 400
rect 4080 360 4120 400
rect 4400 360 4440 400
rect 4720 360 4760 400
rect 5040 360 5240 400
rect 5520 360 5560 400
rect 5840 360 5880 400
rect 6160 360 6200 400
rect 6480 360 6520 400
rect 6800 360 6840 400
rect 7120 360 7160 400
rect 7440 360 7480 400
rect 7760 360 7800 400
rect 8080 360 8120 400
rect 8400 360 8440 400
rect 8720 360 8760 400
rect 9040 360 9080 400
rect 9360 360 9400 400
rect 9680 360 9720 400
rect 10000 360 10040 400
rect 10320 360 10560 400
rect -320 -80 -280 -40
rect -160 200 -40 240
rect 240 200 280 240
rect 560 200 600 240
rect 880 200 920 240
rect 1200 200 1240 240
rect 1520 200 1560 240
rect 1840 200 1880 240
rect 2160 200 2200 240
rect 2480 200 2520 240
rect 2800 200 2840 240
rect 3120 200 3160 240
rect 3440 200 3480 240
rect 3760 200 3800 240
rect 4080 200 4120 240
rect 4400 200 4440 240
rect 4720 200 4760 240
rect 5040 200 5240 240
rect 5520 200 5560 240
rect 5840 200 5880 240
rect 6160 200 6200 240
rect 6480 200 6520 240
rect 6800 200 6840 240
rect 7120 200 7160 240
rect 7440 200 7480 240
rect 7760 200 7800 240
rect 8080 200 8120 240
rect 8400 200 8440 240
rect 8720 200 8760 240
rect 9040 200 9080 240
rect 9360 200 9400 240
rect 9680 200 9720 240
rect 10000 200 10040 240
rect 10320 200 10480 240
rect -160 160 -120 200
rect 5120 160 5160 200
rect 10400 160 10440 200
rect -160 -80 -120 -40
rect 5120 -80 5160 -40
rect 10400 -80 10440 -40
rect 10560 -80 10600 -40
rect -320 -120 -40 -80
rect 240 -120 280 -80
rect 560 -120 600 -80
rect 880 -120 920 -80
rect 1200 -120 1240 -80
rect 1520 -120 1560 -80
rect 1840 -120 1880 -80
rect 2160 -120 2200 -80
rect 2480 -120 2520 -80
rect 2800 -120 2840 -80
rect 3120 -120 3160 -80
rect 3440 -120 3480 -80
rect 3760 -120 3800 -80
rect 4080 -120 4120 -80
rect 4400 -120 4440 -80
rect 4720 -120 4760 -80
rect 5040 -120 5240 -80
rect 5520 -120 5560 -80
rect 5840 -120 5880 -80
rect 6160 -120 6200 -80
rect 6480 -120 6520 -80
rect 6800 -120 6840 -80
rect 7120 -120 7160 -80
rect 7440 -120 7480 -80
rect 7760 -120 7800 -80
rect 8080 -120 8120 -80
rect 8400 -120 8440 -80
rect 8720 -120 8760 -80
rect 9040 -120 9080 -80
rect 9360 -120 9400 -80
rect 9680 -120 9720 -80
rect 10000 -120 10040 -80
rect 10320 -120 10600 -80
rect -320 -200 -40 -160
rect 240 -200 280 -160
rect 560 -200 600 -160
rect 880 -200 920 -160
rect 1200 -200 1240 -160
rect 1520 -200 1560 -160
rect 1840 -200 1880 -160
rect 2160 -200 2200 -160
rect 2480 -200 2520 -160
rect 2800 -200 2840 -160
rect 3120 -200 3160 -160
rect 3440 -200 3480 -160
rect 3760 -200 3800 -160
rect 4080 -200 4120 -160
rect 4400 -200 4440 -160
rect 4720 -200 4760 -160
rect 5040 -200 5240 -160
rect 5520 -200 5560 -160
rect 5840 -200 5880 -160
rect 6160 -200 6200 -160
rect 6480 -200 6520 -160
rect 6800 -200 6840 -160
rect 7120 -200 7160 -160
rect 7440 -200 7480 -160
rect 7760 -200 7800 -160
rect 8080 -200 8120 -160
rect 8400 -200 8440 -160
rect 8720 -200 8760 -160
rect 9040 -200 9080 -160
rect 9360 -200 9400 -160
rect 9680 -200 9720 -160
rect 10000 -200 10040 -160
rect 10320 -200 10600 -160
rect -320 -240 -280 -200
rect -160 -240 -120 -200
rect 5120 -240 5160 -200
rect 10400 -240 10440 -200
rect -160 -480 -120 -440
rect 5120 -480 5160 -440
rect 10400 -480 10440 -440
rect -200 -520 -40 -480
rect 240 -520 280 -480
rect 560 -520 600 -480
rect 880 -520 920 -480
rect 1200 -520 1240 -480
rect 1520 -520 1560 -480
rect 1840 -520 1880 -480
rect 2160 -520 2200 -480
rect 2480 -520 2520 -480
rect 2800 -520 2840 -480
rect 3120 -520 3160 -480
rect 3440 -520 3480 -480
rect 3760 -520 3800 -480
rect 4080 -520 4120 -480
rect 4400 -520 4440 -480
rect 4720 -520 4760 -480
rect 5040 -520 5240 -480
rect 5520 -520 5560 -480
rect 5840 -520 5880 -480
rect 6160 -520 6200 -480
rect 6480 -520 6520 -480
rect 6800 -520 6840 -480
rect 7120 -520 7160 -480
rect 7440 -520 7480 -480
rect 7760 -520 7800 -480
rect 8080 -520 8120 -480
rect 8400 -520 8440 -480
rect 8720 -520 8760 -480
rect 9040 -520 9080 -480
rect 9360 -520 9400 -480
rect 9680 -520 9720 -480
rect 10000 -520 10040 -480
rect 10320 -520 10440 -480
rect 10560 -240 10600 -200
rect -280 -680 -40 -640
rect 240 -680 280 -640
rect 560 -680 600 -640
rect 880 -680 920 -640
rect 1200 -680 1240 -640
rect 1520 -680 1560 -640
rect 1840 -680 1880 -640
rect 2160 -680 2200 -640
rect 2480 -680 2520 -640
rect 2800 -680 2840 -640
rect 3120 -680 3160 -640
rect 3440 -680 3480 -640
rect 3760 -680 3800 -640
rect 4080 -680 4120 -640
rect 4400 -680 4440 -640
rect 4720 -680 4760 -640
rect 5040 -680 5240 -640
rect 5520 -680 5560 -640
rect 5840 -680 5880 -640
rect 6160 -680 6200 -640
rect 6480 -680 6520 -640
rect 6800 -680 6840 -640
rect 7120 -680 7160 -640
rect 7440 -680 7480 -640
rect 7760 -680 7800 -640
rect 8080 -680 8120 -640
rect 8400 -680 8440 -640
rect 8720 -680 8760 -640
rect 9040 -680 9080 -640
rect 9360 -680 9400 -640
rect 9680 -680 9720 -640
rect 10000 -680 10040 -640
rect 10320 -680 10560 -640
rect -320 -1280 -280 -1240
rect 10560 -1280 10600 -1240
rect -320 -1320 -40 -1280
rect 240 -1320 280 -1280
rect 560 -1320 600 -1280
rect 880 -1320 920 -1280
rect 1200 -1320 1240 -1280
rect 1520 -1320 1560 -1280
rect 1840 -1320 1880 -1280
rect 2160 -1320 2200 -1280
rect 2480 -1320 2520 -1280
rect 2800 -1320 2840 -1280
rect 3120 -1320 3160 -1280
rect 3440 -1320 3480 -1280
rect 3760 -1320 3800 -1280
rect 4080 -1320 4120 -1280
rect 4400 -1320 4440 -1280
rect 4720 -1320 4760 -1280
rect 5040 -1320 5240 -1280
rect 5520 -1320 5560 -1280
rect 5840 -1320 5880 -1280
rect 6160 -1320 6200 -1280
rect 6480 -1320 6520 -1280
rect 6800 -1320 6840 -1280
rect 7120 -1320 7160 -1280
rect 7440 -1320 7480 -1280
rect 7760 -1320 7800 -1280
rect 8080 -1320 8120 -1280
rect 8400 -1320 8440 -1280
rect 8720 -1320 8760 -1280
rect 9040 -1320 9080 -1280
rect 9360 -1320 9400 -1280
rect 9680 -1320 9720 -1280
rect 10000 -1320 10040 -1280
rect 10320 -1320 10600 -1280
rect -320 -1400 -40 -1360
rect 240 -1400 280 -1360
rect 560 -1400 600 -1360
rect 880 -1400 920 -1360
rect 1200 -1400 1240 -1360
rect 1520 -1400 1560 -1360
rect 1840 -1400 1880 -1360
rect 2160 -1400 2200 -1360
rect 2480 -1400 2520 -1360
rect 2800 -1400 2840 -1360
rect 3120 -1400 3160 -1360
rect 3440 -1400 3480 -1360
rect 3760 -1400 3800 -1360
rect 4080 -1400 4120 -1360
rect 4400 -1400 4440 -1360
rect 4720 -1400 4760 -1360
rect 5040 -1400 5240 -1360
rect 5520 -1400 5560 -1360
rect 5840 -1400 5880 -1360
rect 6160 -1400 6200 -1360
rect 6480 -1400 6520 -1360
rect 6800 -1400 6840 -1360
rect 7120 -1400 7160 -1360
rect 7440 -1400 7480 -1360
rect 7760 -1400 7800 -1360
rect 8080 -1400 8120 -1360
rect 8400 -1400 8440 -1360
rect 8720 -1400 8760 -1360
rect 9040 -1400 9080 -1360
rect 9360 -1400 9400 -1360
rect 9680 -1400 9720 -1360
rect 10000 -1400 10040 -1360
rect 10320 -1400 10600 -1360
rect -320 -1440 -280 -1400
rect 10560 -1440 10600 -1400
rect -280 -2040 -40 -2000
rect 240 -2040 280 -2000
rect 560 -2040 600 -2000
rect 880 -2040 920 -2000
rect 1200 -2040 1240 -2000
rect 1520 -2040 1560 -2000
rect 1840 -2040 1880 -2000
rect 2160 -2040 2200 -2000
rect 2480 -2040 2520 -2000
rect 2800 -2040 2840 -2000
rect 3120 -2040 3160 -2000
rect 3440 -2040 3480 -2000
rect 3760 -2040 3800 -2000
rect 4080 -2040 4120 -2000
rect 4400 -2040 4440 -2000
rect 4720 -2040 4760 -2000
rect 5040 -2040 5240 -2000
rect 5520 -2040 5560 -2000
rect 5840 -2040 5880 -2000
rect 6160 -2040 6200 -2000
rect 6480 -2040 6520 -2000
rect 6800 -2040 6840 -2000
rect 7120 -2040 7160 -2000
rect 7440 -2040 7480 -2000
rect 7760 -2040 7800 -2000
rect 8080 -2040 8120 -2000
rect 8400 -2040 8440 -2000
rect 8720 -2040 8760 -2000
rect 9040 -2040 9080 -2000
rect 9360 -2040 9400 -2000
rect 9680 -2040 9720 -2000
rect 10000 -2040 10040 -2000
rect 10320 -2040 10560 -2000
rect -200 -2200 -40 -2160
rect 240 -2200 280 -2160
rect 560 -2200 600 -2160
rect 880 -2200 920 -2160
rect 1200 -2200 1240 -2160
rect 1520 -2200 1560 -2160
rect 1840 -2200 1880 -2160
rect 2160 -2200 2200 -2160
rect 2480 -2200 2520 -2160
rect 2800 -2200 2840 -2160
rect 3120 -2200 3160 -2160
rect 3440 -2200 3480 -2160
rect 3760 -2200 3800 -2160
rect 4080 -2200 4120 -2160
rect 4400 -2200 4440 -2160
rect 4720 -2200 4760 -2160
rect 5040 -2200 5240 -2160
rect 5520 -2200 5560 -2160
rect 5840 -2200 5880 -2160
rect 6160 -2200 6200 -2160
rect 6480 -2200 6520 -2160
rect 6800 -2200 6840 -2160
rect 7120 -2200 7160 -2160
rect 7440 -2200 7480 -2160
rect 7760 -2200 7800 -2160
rect 8080 -2200 8120 -2160
rect 8400 -2200 8440 -2160
rect 8720 -2200 8760 -2160
rect 9040 -2200 9080 -2160
rect 9360 -2200 9400 -2160
rect 9680 -2200 9720 -2160
rect 10000 -2200 10040 -2160
rect 10320 -2200 10440 -2160
rect -320 -2480 -280 -2440
rect -160 -2240 -120 -2200
rect 5120 -2240 5160 -2200
rect 10400 -2240 10440 -2200
rect -160 -2480 -120 -2440
rect 5120 -2480 5160 -2440
rect 10400 -2480 10440 -2440
rect 10560 -2480 10600 -2440
rect -320 -2520 -40 -2480
rect 240 -2520 280 -2480
rect 560 -2520 600 -2480
rect 880 -2520 920 -2480
rect 1200 -2520 1240 -2480
rect 1520 -2520 1560 -2480
rect 1840 -2520 1880 -2480
rect 2160 -2520 2200 -2480
rect 2480 -2520 2520 -2480
rect 2800 -2520 2840 -2480
rect 3120 -2520 3160 -2480
rect 3440 -2520 3480 -2480
rect 3760 -2520 3800 -2480
rect 4080 -2520 4120 -2480
rect 4400 -2520 4440 -2480
rect 4720 -2520 4760 -2480
rect 5040 -2520 5240 -2480
rect 5520 -2520 5560 -2480
rect 5840 -2520 5880 -2480
rect 6160 -2520 6200 -2480
rect 6480 -2520 6520 -2480
rect 6800 -2520 6840 -2480
rect 7120 -2520 7160 -2480
rect 7440 -2520 7480 -2480
rect 7760 -2520 7800 -2480
rect 8080 -2520 8120 -2480
rect 8400 -2520 8440 -2480
rect 8720 -2520 8760 -2480
rect 9040 -2520 9080 -2480
rect 9360 -2520 9400 -2480
rect 9680 -2520 9720 -2480
rect 10000 -2520 10040 -2480
rect 10320 -2520 10600 -2480
rect -320 -2600 -40 -2560
rect 240 -2600 280 -2560
rect 560 -2600 600 -2560
rect 880 -2600 920 -2560
rect 1200 -2600 1240 -2560
rect 1520 -2600 1560 -2560
rect 1840 -2600 1880 -2560
rect 2160 -2600 2200 -2560
rect 2480 -2600 2520 -2560
rect 2800 -2600 2840 -2560
rect 3120 -2600 3160 -2560
rect 3440 -2600 3480 -2560
rect 3760 -2600 3800 -2560
rect 4080 -2600 4120 -2560
rect 4400 -2600 4440 -2560
rect 4720 -2600 4760 -2560
rect 5040 -2600 5240 -2560
rect 5520 -2600 5560 -2560
rect 5840 -2600 5880 -2560
rect 6160 -2600 6200 -2560
rect 6480 -2600 6520 -2560
rect 6800 -2600 6840 -2560
rect 7120 -2600 7160 -2560
rect 7440 -2600 7480 -2560
rect 7760 -2600 7800 -2560
rect 8080 -2600 8120 -2560
rect 8400 -2600 8440 -2560
rect 8720 -2600 8760 -2560
rect 9040 -2600 9080 -2560
rect 9360 -2600 9400 -2560
rect 9680 -2600 9720 -2560
rect 10000 -2600 10040 -2560
rect 10320 -2600 10600 -2560
rect -320 -2640 -280 -2600
rect -160 -2640 -120 -2600
rect 5120 -2640 5160 -2600
rect 10400 -2640 10440 -2600
rect -160 -2880 -120 -2840
rect 5120 -2880 5160 -2840
rect 10400 -2880 10440 -2840
rect 10560 -2640 10600 -2600
rect -160 -2920 -40 -2880
rect 240 -2920 280 -2880
rect 560 -2920 600 -2880
rect 880 -2920 920 -2880
rect 1200 -2920 1240 -2880
rect 1520 -2920 1560 -2880
rect 1840 -2920 1880 -2880
rect 2160 -2920 2200 -2880
rect 2480 -2920 2520 -2880
rect 2800 -2920 2840 -2880
rect 3120 -2920 3160 -2880
rect 3440 -2920 3480 -2880
rect 3760 -2920 3800 -2880
rect 4080 -2920 4120 -2880
rect 4400 -2920 4440 -2880
rect 4720 -2920 4760 -2880
rect 5040 -2920 5240 -2880
rect 5520 -2920 5560 -2880
rect 5840 -2920 5880 -2880
rect 6160 -2920 6200 -2880
rect 6480 -2920 6520 -2880
rect 6800 -2920 6840 -2880
rect 7120 -2920 7160 -2880
rect 7440 -2920 7480 -2880
rect 7760 -2920 7800 -2880
rect 8080 -2920 8120 -2880
rect 8400 -2920 8440 -2880
rect 8720 -2920 8760 -2880
rect 9040 -2920 9080 -2880
rect 9360 -2920 9400 -2880
rect 9680 -2920 9720 -2880
rect 10000 -2920 10040 -2880
rect 10320 -2920 10480 -2880
rect -280 -3080 -40 -3040
rect 240 -3080 280 -3040
rect 560 -3080 600 -3040
rect 880 -3080 920 -3040
rect 1200 -3080 1240 -3040
rect 1520 -3080 1560 -3040
rect 1840 -3080 1880 -3040
rect 2160 -3080 2200 -3040
rect 2480 -3080 2520 -3040
rect 2800 -3080 2840 -3040
rect 3120 -3080 3160 -3040
rect 3440 -3080 3480 -3040
rect 3760 -3080 3800 -3040
rect 4080 -3080 4120 -3040
rect 4400 -3080 4440 -3040
rect 4720 -3080 4760 -3040
rect 5040 -3080 5240 -3040
rect 5520 -3080 5560 -3040
rect 5840 -3080 5880 -3040
rect 6160 -3080 6200 -3040
rect 6480 -3080 6520 -3040
rect 6800 -3080 6840 -3040
rect 7120 -3080 7160 -3040
rect 7440 -3080 7480 -3040
rect 7760 -3080 7800 -3040
rect 8080 -3080 8120 -3040
rect 8400 -3080 8440 -3040
rect 8720 -3080 8760 -3040
rect 9040 -3080 9080 -3040
rect 9360 -3080 9400 -3040
rect 9680 -3080 9720 -3040
rect 10000 -3080 10040 -3040
rect 10320 -3080 10560 -3040
rect -320 -3680 -280 -3640
rect 10560 -3680 10600 -3640
rect -320 -3720 -40 -3680
rect 240 -3720 280 -3680
rect 560 -3720 600 -3680
rect 880 -3720 920 -3680
rect 1200 -3720 1240 -3680
rect 1520 -3720 1560 -3680
rect 1840 -3720 1880 -3680
rect 2160 -3720 2200 -3680
rect 2480 -3720 2520 -3680
rect 2800 -3720 2840 -3680
rect 3120 -3720 3160 -3680
rect 3440 -3720 3480 -3680
rect 3760 -3720 3800 -3680
rect 4080 -3720 4120 -3680
rect 4400 -3720 4440 -3680
rect 4720 -3720 4760 -3680
rect 5040 -3720 5240 -3680
rect 5520 -3720 5560 -3680
rect 5840 -3720 5880 -3680
rect 6160 -3720 6200 -3680
rect 6480 -3720 6520 -3680
rect 6800 -3720 6840 -3680
rect 7120 -3720 7160 -3680
rect 7440 -3720 7480 -3680
rect 7760 -3720 7800 -3680
rect 8080 -3720 8120 -3680
rect 8400 -3720 8440 -3680
rect 8720 -3720 8760 -3680
rect 9040 -3720 9080 -3680
rect 9360 -3720 9400 -3680
rect 9680 -3720 9720 -3680
rect 10000 -3720 10040 -3680
rect 10320 -3720 10600 -3680
<< nsubdiff >>
rect -160 840 -40 880
rect 240 840 280 880
rect 560 840 600 880
rect 880 840 920 880
rect 1200 840 1240 880
rect 1520 840 1560 880
rect 1840 840 1880 880
rect 2160 840 2200 880
rect 2480 840 2520 880
rect 2800 840 2840 880
rect 3120 840 3160 880
rect 3440 840 3480 880
rect 3760 840 3800 880
rect 4080 840 4120 880
rect 4400 840 4440 880
rect 4720 840 4760 880
rect 5040 840 5240 880
rect 5520 840 5560 880
rect 5840 840 5880 880
rect 6160 840 6200 880
rect 6480 840 6520 880
rect 6800 840 6840 880
rect 7120 840 7160 880
rect 7440 840 7480 880
rect 7760 840 7800 880
rect 8080 840 8120 880
rect 8400 840 8440 880
rect 8720 840 8760 880
rect 9040 840 9080 880
rect 9360 840 9400 880
rect 9680 840 9720 880
rect 10000 840 10040 880
rect 10320 840 10480 880
rect -160 800 -120 840
rect 5120 800 5160 840
rect 10400 800 10440 840
rect -160 560 -120 600
rect 5120 560 5160 600
rect 10400 560 10440 600
rect -160 520 -40 560
rect 240 520 280 560
rect 560 520 600 560
rect 880 520 920 560
rect 1200 520 1240 560
rect 1520 520 1560 560
rect 1840 520 1880 560
rect 2160 520 2200 560
rect 2480 520 2520 560
rect 2800 520 2840 560
rect 3120 520 3160 560
rect 3440 520 3480 560
rect 3760 520 3800 560
rect 4080 520 4120 560
rect 4400 520 4440 560
rect 4720 520 4760 560
rect 5040 520 5240 560
rect 5520 520 5560 560
rect 5840 520 5880 560
rect 6160 520 6200 560
rect 6480 520 6520 560
rect 6800 520 6840 560
rect 7120 520 7160 560
rect 7440 520 7480 560
rect 7760 520 7800 560
rect 8080 520 8120 560
rect 8400 520 8440 560
rect 8720 520 8760 560
rect 9040 520 9080 560
rect 9360 520 9400 560
rect 9680 520 9720 560
rect 10000 520 10040 560
rect 10320 520 10480 560
rect -200 -840 -40 -800
rect 240 -840 280 -800
rect 560 -840 600 -800
rect 880 -840 920 -800
rect 1200 -840 1240 -800
rect 1520 -840 1560 -800
rect 1840 -840 1880 -800
rect 2160 -840 2200 -800
rect 2480 -840 2520 -800
rect 2800 -840 2840 -800
rect 3120 -840 3160 -800
rect 3440 -840 3480 -800
rect 3760 -840 3800 -800
rect 4080 -840 4120 -800
rect 4400 -840 4440 -800
rect 4720 -840 4760 -800
rect 5040 -840 5240 -800
rect 5520 -840 5560 -800
rect 5840 -840 5880 -800
rect 6160 -840 6200 -800
rect 6480 -840 6520 -800
rect 6800 -840 6840 -800
rect 7120 -840 7160 -800
rect 7440 -840 7480 -800
rect 7760 -840 7800 -800
rect 8080 -840 8120 -800
rect 8400 -840 8440 -800
rect 8720 -840 8760 -800
rect 9040 -840 9080 -800
rect 9360 -840 9400 -800
rect 9680 -840 9720 -800
rect 10000 -840 10040 -800
rect 10320 -840 10440 -800
rect -160 -880 -120 -840
rect 5120 -880 5160 -840
rect 10400 -880 10440 -840
rect -160 -1120 -120 -1080
rect 5120 -1120 5160 -1080
rect 10400 -1120 10440 -1080
rect -200 -1160 -40 -1120
rect 240 -1160 280 -1120
rect 560 -1160 600 -1120
rect 880 -1160 920 -1120
rect 1200 -1160 1240 -1120
rect 1520 -1160 1560 -1120
rect 1840 -1160 1880 -1120
rect 2160 -1160 2200 -1120
rect 2480 -1160 2520 -1120
rect 2800 -1160 2840 -1120
rect 3120 -1160 3160 -1120
rect 3440 -1160 3480 -1120
rect 3760 -1160 3800 -1120
rect 4080 -1160 4120 -1120
rect 4400 -1160 4440 -1120
rect 4720 -1160 4760 -1120
rect 5040 -1160 5240 -1120
rect 5520 -1160 5560 -1120
rect 5840 -1160 5880 -1120
rect 6160 -1160 6200 -1120
rect 6480 -1160 6520 -1120
rect 6800 -1160 6840 -1120
rect 7120 -1160 7160 -1120
rect 7440 -1160 7480 -1120
rect 7760 -1160 7800 -1120
rect 8080 -1160 8120 -1120
rect 8400 -1160 8440 -1120
rect 8720 -1160 8760 -1120
rect 9040 -1160 9080 -1120
rect 9360 -1160 9400 -1120
rect 9680 -1160 9720 -1120
rect 10000 -1160 10040 -1120
rect 10320 -1160 10440 -1120
rect -200 -1560 -40 -1520
rect 240 -1560 280 -1520
rect 560 -1560 600 -1520
rect 880 -1560 920 -1520
rect 1200 -1560 1240 -1520
rect 1520 -1560 1560 -1520
rect 1840 -1560 1880 -1520
rect 2160 -1560 2200 -1520
rect 2480 -1560 2520 -1520
rect 2800 -1560 2840 -1520
rect 3120 -1560 3160 -1520
rect 3440 -1560 3480 -1520
rect 3760 -1560 3800 -1520
rect 4080 -1560 4120 -1520
rect 4400 -1560 4440 -1520
rect 4720 -1560 4760 -1520
rect 5040 -1560 5240 -1520
rect 5520 -1560 5560 -1520
rect 5840 -1560 5880 -1520
rect 6160 -1560 6200 -1520
rect 6480 -1560 6520 -1520
rect 6800 -1560 6840 -1520
rect 7120 -1560 7160 -1520
rect 7440 -1560 7480 -1520
rect 7760 -1560 7800 -1520
rect 8080 -1560 8120 -1520
rect 8400 -1560 8440 -1520
rect 8720 -1560 8760 -1520
rect 9040 -1560 9080 -1520
rect 9360 -1560 9400 -1520
rect 9680 -1560 9720 -1520
rect 10000 -1560 10040 -1520
rect 10320 -1560 10440 -1520
rect -160 -1600 -120 -1560
rect 5120 -1600 5160 -1560
rect 10400 -1600 10440 -1560
rect -160 -1840 -120 -1800
rect 5120 -1840 5160 -1800
rect 10400 -1840 10440 -1800
rect -200 -1880 -40 -1840
rect 240 -1880 280 -1840
rect 560 -1880 600 -1840
rect 880 -1880 920 -1840
rect 1200 -1880 1240 -1840
rect 1520 -1880 1560 -1840
rect 1840 -1880 1880 -1840
rect 2160 -1880 2200 -1840
rect 2480 -1880 2520 -1840
rect 2800 -1880 2840 -1840
rect 3120 -1880 3160 -1840
rect 3440 -1880 3480 -1840
rect 3760 -1880 3800 -1840
rect 4080 -1880 4120 -1840
rect 4400 -1880 4440 -1840
rect 4720 -1880 4760 -1840
rect 5040 -1880 5240 -1840
rect 5520 -1880 5560 -1840
rect 5840 -1880 5880 -1840
rect 6160 -1880 6200 -1840
rect 6480 -1880 6520 -1840
rect 6800 -1880 6840 -1840
rect 7120 -1880 7160 -1840
rect 7440 -1880 7480 -1840
rect 7760 -1880 7800 -1840
rect 8080 -1880 8120 -1840
rect 8400 -1880 8440 -1840
rect 8720 -1880 8760 -1840
rect 9040 -1880 9080 -1840
rect 9360 -1880 9400 -1840
rect 9680 -1880 9720 -1840
rect 10000 -1880 10040 -1840
rect 10320 -1880 10440 -1840
rect -160 -3240 -40 -3200
rect 240 -3240 280 -3200
rect 560 -3240 600 -3200
rect 880 -3240 920 -3200
rect 1200 -3240 1240 -3200
rect 1520 -3240 1560 -3200
rect 1840 -3240 1880 -3200
rect 2160 -3240 2200 -3200
rect 2480 -3240 2520 -3200
rect 2800 -3240 2840 -3200
rect 3120 -3240 3160 -3200
rect 3440 -3240 3480 -3200
rect 3760 -3240 3800 -3200
rect 4080 -3240 4120 -3200
rect 4400 -3240 4440 -3200
rect 4720 -3240 4760 -3200
rect 5040 -3240 5240 -3200
rect 5520 -3240 5560 -3200
rect 5840 -3240 5880 -3200
rect 6160 -3240 6200 -3200
rect 6480 -3240 6520 -3200
rect 6800 -3240 6840 -3200
rect 7120 -3240 7160 -3200
rect 7440 -3240 7480 -3200
rect 7760 -3240 7800 -3200
rect 8080 -3240 8120 -3200
rect 8400 -3240 8440 -3200
rect 8720 -3240 8760 -3200
rect 9040 -3240 9080 -3200
rect 9360 -3240 9400 -3200
rect 9680 -3240 9720 -3200
rect 10000 -3240 10040 -3200
rect 10320 -3240 10480 -3200
rect -160 -3280 -120 -3240
rect 5120 -3280 5160 -3240
rect 10400 -3280 10440 -3240
rect -160 -3520 -120 -3480
rect 5120 -3520 5160 -3480
rect 10400 -3520 10440 -3480
rect -160 -3560 -40 -3520
rect 240 -3560 280 -3520
rect 560 -3560 600 -3520
rect 880 -3560 920 -3520
rect 1200 -3560 1240 -3520
rect 1520 -3560 1560 -3520
rect 1840 -3560 1880 -3520
rect 2160 -3560 2200 -3520
rect 2480 -3560 2520 -3520
rect 2800 -3560 2840 -3520
rect 3120 -3560 3160 -3520
rect 3440 -3560 3480 -3520
rect 3760 -3560 3800 -3520
rect 4080 -3560 4120 -3520
rect 4400 -3560 4440 -3520
rect 4720 -3560 4760 -3520
rect 5040 -3560 5240 -3520
rect 5520 -3560 5560 -3520
rect 5840 -3560 5880 -3520
rect 6160 -3560 6200 -3520
rect 6480 -3560 6520 -3520
rect 6800 -3560 6840 -3520
rect 7120 -3560 7160 -3520
rect 7440 -3560 7480 -3520
rect 7760 -3560 7800 -3520
rect 8080 -3560 8120 -3520
rect 8400 -3560 8440 -3520
rect 8720 -3560 8760 -3520
rect 9040 -3560 9080 -3520
rect 9360 -3560 9400 -3520
rect 9680 -3560 9720 -3520
rect 10000 -3560 10040 -3520
rect 10320 -3560 10480 -3520
<< psubdiffcont >>
rect -40 1000 240 1040
rect 280 1000 560 1040
rect 600 1000 880 1040
rect 920 1000 1200 1040
rect 1240 1000 1520 1040
rect 1560 1000 1840 1040
rect 1880 1000 2160 1040
rect 2200 1000 2480 1040
rect 2520 1000 2800 1040
rect 2840 1000 3120 1040
rect 3160 1000 3440 1040
rect 3480 1000 3760 1040
rect 3800 1000 4080 1040
rect 4120 1000 4400 1040
rect 4440 1000 4720 1040
rect 4760 1000 5040 1040
rect 5240 1000 5520 1040
rect 5560 1000 5840 1040
rect 5880 1000 6160 1040
rect 6200 1000 6480 1040
rect 6520 1000 6800 1040
rect 6840 1000 7120 1040
rect 7160 1000 7440 1040
rect 7480 1000 7760 1040
rect 7800 1000 8080 1040
rect 8120 1000 8400 1040
rect 8440 1000 8720 1040
rect 8760 1000 9040 1040
rect 9080 1000 9360 1040
rect 9400 1000 9680 1040
rect 9720 1000 10000 1040
rect 10040 1000 10320 1040
rect -320 -40 -280 960
rect -40 360 240 400
rect 280 360 560 400
rect 600 360 880 400
rect 920 360 1200 400
rect 1240 360 1520 400
rect 1560 360 1840 400
rect 1880 360 2160 400
rect 2200 360 2480 400
rect 2520 360 2800 400
rect 2840 360 3120 400
rect 3160 360 3440 400
rect 3480 360 3760 400
rect 3800 360 4080 400
rect 4120 360 4400 400
rect 4440 360 4720 400
rect 4760 360 5040 400
rect 5240 360 5520 400
rect 5560 360 5840 400
rect 5880 360 6160 400
rect 6200 360 6480 400
rect 6520 360 6800 400
rect 6840 360 7120 400
rect 7160 360 7440 400
rect 7480 360 7760 400
rect 7800 360 8080 400
rect 8120 360 8400 400
rect 8440 360 8720 400
rect 8760 360 9040 400
rect 9080 360 9360 400
rect 9400 360 9680 400
rect 9720 360 10000 400
rect 10040 360 10320 400
rect -40 200 240 240
rect 280 200 560 240
rect 600 200 880 240
rect 920 200 1200 240
rect 1240 200 1520 240
rect 1560 200 1840 240
rect 1880 200 2160 240
rect 2200 200 2480 240
rect 2520 200 2800 240
rect 2840 200 3120 240
rect 3160 200 3440 240
rect 3480 200 3760 240
rect 3800 200 4080 240
rect 4120 200 4400 240
rect 4440 200 4720 240
rect 4760 200 5040 240
rect 5240 200 5520 240
rect 5560 200 5840 240
rect 5880 200 6160 240
rect 6200 200 6480 240
rect 6520 200 6800 240
rect 6840 200 7120 240
rect 7160 200 7440 240
rect 7480 200 7760 240
rect 7800 200 8080 240
rect 8120 200 8400 240
rect 8440 200 8720 240
rect 8760 200 9040 240
rect 9080 200 9360 240
rect 9400 200 9680 240
rect 9720 200 10000 240
rect 10040 200 10320 240
rect -160 -40 -120 160
rect 5120 -40 5160 160
rect 10400 -40 10440 160
rect 10560 -40 10600 960
rect -40 -120 240 -80
rect 280 -120 560 -80
rect 600 -120 880 -80
rect 920 -120 1200 -80
rect 1240 -120 1520 -80
rect 1560 -120 1840 -80
rect 1880 -120 2160 -80
rect 2200 -120 2480 -80
rect 2520 -120 2800 -80
rect 2840 -120 3120 -80
rect 3160 -120 3440 -80
rect 3480 -120 3760 -80
rect 3800 -120 4080 -80
rect 4120 -120 4400 -80
rect 4440 -120 4720 -80
rect 4760 -120 5040 -80
rect 5240 -120 5520 -80
rect 5560 -120 5840 -80
rect 5880 -120 6160 -80
rect 6200 -120 6480 -80
rect 6520 -120 6800 -80
rect 6840 -120 7120 -80
rect 7160 -120 7440 -80
rect 7480 -120 7760 -80
rect 7800 -120 8080 -80
rect 8120 -120 8400 -80
rect 8440 -120 8720 -80
rect 8760 -120 9040 -80
rect 9080 -120 9360 -80
rect 9400 -120 9680 -80
rect 9720 -120 10000 -80
rect 10040 -120 10320 -80
rect -40 -200 240 -160
rect 280 -200 560 -160
rect 600 -200 880 -160
rect 920 -200 1200 -160
rect 1240 -200 1520 -160
rect 1560 -200 1840 -160
rect 1880 -200 2160 -160
rect 2200 -200 2480 -160
rect 2520 -200 2800 -160
rect 2840 -200 3120 -160
rect 3160 -200 3440 -160
rect 3480 -200 3760 -160
rect 3800 -200 4080 -160
rect 4120 -200 4400 -160
rect 4440 -200 4720 -160
rect 4760 -200 5040 -160
rect 5240 -200 5520 -160
rect 5560 -200 5840 -160
rect 5880 -200 6160 -160
rect 6200 -200 6480 -160
rect 6520 -200 6800 -160
rect 6840 -200 7120 -160
rect 7160 -200 7440 -160
rect 7480 -200 7760 -160
rect 7800 -200 8080 -160
rect 8120 -200 8400 -160
rect 8440 -200 8720 -160
rect 8760 -200 9040 -160
rect 9080 -200 9360 -160
rect 9400 -200 9680 -160
rect 9720 -200 10000 -160
rect 10040 -200 10320 -160
rect -320 -1240 -280 -240
rect -160 -440 -120 -240
rect 5120 -440 5160 -240
rect 10400 -440 10440 -240
rect -40 -520 240 -480
rect 280 -520 560 -480
rect 600 -520 880 -480
rect 920 -520 1200 -480
rect 1240 -520 1520 -480
rect 1560 -520 1840 -480
rect 1880 -520 2160 -480
rect 2200 -520 2480 -480
rect 2520 -520 2800 -480
rect 2840 -520 3120 -480
rect 3160 -520 3440 -480
rect 3480 -520 3760 -480
rect 3800 -520 4080 -480
rect 4120 -520 4400 -480
rect 4440 -520 4720 -480
rect 4760 -520 5040 -480
rect 5240 -520 5520 -480
rect 5560 -520 5840 -480
rect 5880 -520 6160 -480
rect 6200 -520 6480 -480
rect 6520 -520 6800 -480
rect 6840 -520 7120 -480
rect 7160 -520 7440 -480
rect 7480 -520 7760 -480
rect 7800 -520 8080 -480
rect 8120 -520 8400 -480
rect 8440 -520 8720 -480
rect 8760 -520 9040 -480
rect 9080 -520 9360 -480
rect 9400 -520 9680 -480
rect 9720 -520 10000 -480
rect 10040 -520 10320 -480
rect -40 -680 240 -640
rect 280 -680 560 -640
rect 600 -680 880 -640
rect 920 -680 1200 -640
rect 1240 -680 1520 -640
rect 1560 -680 1840 -640
rect 1880 -680 2160 -640
rect 2200 -680 2480 -640
rect 2520 -680 2800 -640
rect 2840 -680 3120 -640
rect 3160 -680 3440 -640
rect 3480 -680 3760 -640
rect 3800 -680 4080 -640
rect 4120 -680 4400 -640
rect 4440 -680 4720 -640
rect 4760 -680 5040 -640
rect 5240 -680 5520 -640
rect 5560 -680 5840 -640
rect 5880 -680 6160 -640
rect 6200 -680 6480 -640
rect 6520 -680 6800 -640
rect 6840 -680 7120 -640
rect 7160 -680 7440 -640
rect 7480 -680 7760 -640
rect 7800 -680 8080 -640
rect 8120 -680 8400 -640
rect 8440 -680 8720 -640
rect 8760 -680 9040 -640
rect 9080 -680 9360 -640
rect 9400 -680 9680 -640
rect 9720 -680 10000 -640
rect 10040 -680 10320 -640
rect 10560 -1240 10600 -240
rect -40 -1320 240 -1280
rect 280 -1320 560 -1280
rect 600 -1320 880 -1280
rect 920 -1320 1200 -1280
rect 1240 -1320 1520 -1280
rect 1560 -1320 1840 -1280
rect 1880 -1320 2160 -1280
rect 2200 -1320 2480 -1280
rect 2520 -1320 2800 -1280
rect 2840 -1320 3120 -1280
rect 3160 -1320 3440 -1280
rect 3480 -1320 3760 -1280
rect 3800 -1320 4080 -1280
rect 4120 -1320 4400 -1280
rect 4440 -1320 4720 -1280
rect 4760 -1320 5040 -1280
rect 5240 -1320 5520 -1280
rect 5560 -1320 5840 -1280
rect 5880 -1320 6160 -1280
rect 6200 -1320 6480 -1280
rect 6520 -1320 6800 -1280
rect 6840 -1320 7120 -1280
rect 7160 -1320 7440 -1280
rect 7480 -1320 7760 -1280
rect 7800 -1320 8080 -1280
rect 8120 -1320 8400 -1280
rect 8440 -1320 8720 -1280
rect 8760 -1320 9040 -1280
rect 9080 -1320 9360 -1280
rect 9400 -1320 9680 -1280
rect 9720 -1320 10000 -1280
rect 10040 -1320 10320 -1280
rect -40 -1400 240 -1360
rect 280 -1400 560 -1360
rect 600 -1400 880 -1360
rect 920 -1400 1200 -1360
rect 1240 -1400 1520 -1360
rect 1560 -1400 1840 -1360
rect 1880 -1400 2160 -1360
rect 2200 -1400 2480 -1360
rect 2520 -1400 2800 -1360
rect 2840 -1400 3120 -1360
rect 3160 -1400 3440 -1360
rect 3480 -1400 3760 -1360
rect 3800 -1400 4080 -1360
rect 4120 -1400 4400 -1360
rect 4440 -1400 4720 -1360
rect 4760 -1400 5040 -1360
rect 5240 -1400 5520 -1360
rect 5560 -1400 5840 -1360
rect 5880 -1400 6160 -1360
rect 6200 -1400 6480 -1360
rect 6520 -1400 6800 -1360
rect 6840 -1400 7120 -1360
rect 7160 -1400 7440 -1360
rect 7480 -1400 7760 -1360
rect 7800 -1400 8080 -1360
rect 8120 -1400 8400 -1360
rect 8440 -1400 8720 -1360
rect 8760 -1400 9040 -1360
rect 9080 -1400 9360 -1360
rect 9400 -1400 9680 -1360
rect 9720 -1400 10000 -1360
rect 10040 -1400 10320 -1360
rect -320 -2440 -280 -1440
rect -40 -2040 240 -2000
rect 280 -2040 560 -2000
rect 600 -2040 880 -2000
rect 920 -2040 1200 -2000
rect 1240 -2040 1520 -2000
rect 1560 -2040 1840 -2000
rect 1880 -2040 2160 -2000
rect 2200 -2040 2480 -2000
rect 2520 -2040 2800 -2000
rect 2840 -2040 3120 -2000
rect 3160 -2040 3440 -2000
rect 3480 -2040 3760 -2000
rect 3800 -2040 4080 -2000
rect 4120 -2040 4400 -2000
rect 4440 -2040 4720 -2000
rect 4760 -2040 5040 -2000
rect 5240 -2040 5520 -2000
rect 5560 -2040 5840 -2000
rect 5880 -2040 6160 -2000
rect 6200 -2040 6480 -2000
rect 6520 -2040 6800 -2000
rect 6840 -2040 7120 -2000
rect 7160 -2040 7440 -2000
rect 7480 -2040 7760 -2000
rect 7800 -2040 8080 -2000
rect 8120 -2040 8400 -2000
rect 8440 -2040 8720 -2000
rect 8760 -2040 9040 -2000
rect 9080 -2040 9360 -2000
rect 9400 -2040 9680 -2000
rect 9720 -2040 10000 -2000
rect 10040 -2040 10320 -2000
rect -40 -2200 240 -2160
rect 280 -2200 560 -2160
rect 600 -2200 880 -2160
rect 920 -2200 1200 -2160
rect 1240 -2200 1520 -2160
rect 1560 -2200 1840 -2160
rect 1880 -2200 2160 -2160
rect 2200 -2200 2480 -2160
rect 2520 -2200 2800 -2160
rect 2840 -2200 3120 -2160
rect 3160 -2200 3440 -2160
rect 3480 -2200 3760 -2160
rect 3800 -2200 4080 -2160
rect 4120 -2200 4400 -2160
rect 4440 -2200 4720 -2160
rect 4760 -2200 5040 -2160
rect 5240 -2200 5520 -2160
rect 5560 -2200 5840 -2160
rect 5880 -2200 6160 -2160
rect 6200 -2200 6480 -2160
rect 6520 -2200 6800 -2160
rect 6840 -2200 7120 -2160
rect 7160 -2200 7440 -2160
rect 7480 -2200 7760 -2160
rect 7800 -2200 8080 -2160
rect 8120 -2200 8400 -2160
rect 8440 -2200 8720 -2160
rect 8760 -2200 9040 -2160
rect 9080 -2200 9360 -2160
rect 9400 -2200 9680 -2160
rect 9720 -2200 10000 -2160
rect 10040 -2200 10320 -2160
rect -160 -2440 -120 -2240
rect 5120 -2440 5160 -2240
rect 10400 -2440 10440 -2240
rect 10560 -2440 10600 -1440
rect -40 -2520 240 -2480
rect 280 -2520 560 -2480
rect 600 -2520 880 -2480
rect 920 -2520 1200 -2480
rect 1240 -2520 1520 -2480
rect 1560 -2520 1840 -2480
rect 1880 -2520 2160 -2480
rect 2200 -2520 2480 -2480
rect 2520 -2520 2800 -2480
rect 2840 -2520 3120 -2480
rect 3160 -2520 3440 -2480
rect 3480 -2520 3760 -2480
rect 3800 -2520 4080 -2480
rect 4120 -2520 4400 -2480
rect 4440 -2520 4720 -2480
rect 4760 -2520 5040 -2480
rect 5240 -2520 5520 -2480
rect 5560 -2520 5840 -2480
rect 5880 -2520 6160 -2480
rect 6200 -2520 6480 -2480
rect 6520 -2520 6800 -2480
rect 6840 -2520 7120 -2480
rect 7160 -2520 7440 -2480
rect 7480 -2520 7760 -2480
rect 7800 -2520 8080 -2480
rect 8120 -2520 8400 -2480
rect 8440 -2520 8720 -2480
rect 8760 -2520 9040 -2480
rect 9080 -2520 9360 -2480
rect 9400 -2520 9680 -2480
rect 9720 -2520 10000 -2480
rect 10040 -2520 10320 -2480
rect -40 -2600 240 -2560
rect 280 -2600 560 -2560
rect 600 -2600 880 -2560
rect 920 -2600 1200 -2560
rect 1240 -2600 1520 -2560
rect 1560 -2600 1840 -2560
rect 1880 -2600 2160 -2560
rect 2200 -2600 2480 -2560
rect 2520 -2600 2800 -2560
rect 2840 -2600 3120 -2560
rect 3160 -2600 3440 -2560
rect 3480 -2600 3760 -2560
rect 3800 -2600 4080 -2560
rect 4120 -2600 4400 -2560
rect 4440 -2600 4720 -2560
rect 4760 -2600 5040 -2560
rect 5240 -2600 5520 -2560
rect 5560 -2600 5840 -2560
rect 5880 -2600 6160 -2560
rect 6200 -2600 6480 -2560
rect 6520 -2600 6800 -2560
rect 6840 -2600 7120 -2560
rect 7160 -2600 7440 -2560
rect 7480 -2600 7760 -2560
rect 7800 -2600 8080 -2560
rect 8120 -2600 8400 -2560
rect 8440 -2600 8720 -2560
rect 8760 -2600 9040 -2560
rect 9080 -2600 9360 -2560
rect 9400 -2600 9680 -2560
rect 9720 -2600 10000 -2560
rect 10040 -2600 10320 -2560
rect -320 -3640 -280 -2640
rect -160 -2840 -120 -2640
rect 5120 -2840 5160 -2640
rect 10400 -2840 10440 -2640
rect -40 -2920 240 -2880
rect 280 -2920 560 -2880
rect 600 -2920 880 -2880
rect 920 -2920 1200 -2880
rect 1240 -2920 1520 -2880
rect 1560 -2920 1840 -2880
rect 1880 -2920 2160 -2880
rect 2200 -2920 2480 -2880
rect 2520 -2920 2800 -2880
rect 2840 -2920 3120 -2880
rect 3160 -2920 3440 -2880
rect 3480 -2920 3760 -2880
rect 3800 -2920 4080 -2880
rect 4120 -2920 4400 -2880
rect 4440 -2920 4720 -2880
rect 4760 -2920 5040 -2880
rect 5240 -2920 5520 -2880
rect 5560 -2920 5840 -2880
rect 5880 -2920 6160 -2880
rect 6200 -2920 6480 -2880
rect 6520 -2920 6800 -2880
rect 6840 -2920 7120 -2880
rect 7160 -2920 7440 -2880
rect 7480 -2920 7760 -2880
rect 7800 -2920 8080 -2880
rect 8120 -2920 8400 -2880
rect 8440 -2920 8720 -2880
rect 8760 -2920 9040 -2880
rect 9080 -2920 9360 -2880
rect 9400 -2920 9680 -2880
rect 9720 -2920 10000 -2880
rect 10040 -2920 10320 -2880
rect -40 -3080 240 -3040
rect 280 -3080 560 -3040
rect 600 -3080 880 -3040
rect 920 -3080 1200 -3040
rect 1240 -3080 1520 -3040
rect 1560 -3080 1840 -3040
rect 1880 -3080 2160 -3040
rect 2200 -3080 2480 -3040
rect 2520 -3080 2800 -3040
rect 2840 -3080 3120 -3040
rect 3160 -3080 3440 -3040
rect 3480 -3080 3760 -3040
rect 3800 -3080 4080 -3040
rect 4120 -3080 4400 -3040
rect 4440 -3080 4720 -3040
rect 4760 -3080 5040 -3040
rect 5240 -3080 5520 -3040
rect 5560 -3080 5840 -3040
rect 5880 -3080 6160 -3040
rect 6200 -3080 6480 -3040
rect 6520 -3080 6800 -3040
rect 6840 -3080 7120 -3040
rect 7160 -3080 7440 -3040
rect 7480 -3080 7760 -3040
rect 7800 -3080 8080 -3040
rect 8120 -3080 8400 -3040
rect 8440 -3080 8720 -3040
rect 8760 -3080 9040 -3040
rect 9080 -3080 9360 -3040
rect 9400 -3080 9680 -3040
rect 9720 -3080 10000 -3040
rect 10040 -3080 10320 -3040
rect 10560 -3640 10600 -2640
rect -40 -3720 240 -3680
rect 280 -3720 560 -3680
rect 600 -3720 880 -3680
rect 920 -3720 1200 -3680
rect 1240 -3720 1520 -3680
rect 1560 -3720 1840 -3680
rect 1880 -3720 2160 -3680
rect 2200 -3720 2480 -3680
rect 2520 -3720 2800 -3680
rect 2840 -3720 3120 -3680
rect 3160 -3720 3440 -3680
rect 3480 -3720 3760 -3680
rect 3800 -3720 4080 -3680
rect 4120 -3720 4400 -3680
rect 4440 -3720 4720 -3680
rect 4760 -3720 5040 -3680
rect 5240 -3720 5520 -3680
rect 5560 -3720 5840 -3680
rect 5880 -3720 6160 -3680
rect 6200 -3720 6480 -3680
rect 6520 -3720 6800 -3680
rect 6840 -3720 7120 -3680
rect 7160 -3720 7440 -3680
rect 7480 -3720 7760 -3680
rect 7800 -3720 8080 -3680
rect 8120 -3720 8400 -3680
rect 8440 -3720 8720 -3680
rect 8760 -3720 9040 -3680
rect 9080 -3720 9360 -3680
rect 9400 -3720 9680 -3680
rect 9720 -3720 10000 -3680
rect 10040 -3720 10320 -3680
<< nsubdiffcont >>
rect -40 840 240 880
rect 280 840 560 880
rect 600 840 880 880
rect 920 840 1200 880
rect 1240 840 1520 880
rect 1560 840 1840 880
rect 1880 840 2160 880
rect 2200 840 2480 880
rect 2520 840 2800 880
rect 2840 840 3120 880
rect 3160 840 3440 880
rect 3480 840 3760 880
rect 3800 840 4080 880
rect 4120 840 4400 880
rect 4440 840 4720 880
rect 4760 840 5040 880
rect 5240 840 5520 880
rect 5560 840 5840 880
rect 5880 840 6160 880
rect 6200 840 6480 880
rect 6520 840 6800 880
rect 6840 840 7120 880
rect 7160 840 7440 880
rect 7480 840 7760 880
rect 7800 840 8080 880
rect 8120 840 8400 880
rect 8440 840 8720 880
rect 8760 840 9040 880
rect 9080 840 9360 880
rect 9400 840 9680 880
rect 9720 840 10000 880
rect 10040 840 10320 880
rect -160 600 -120 800
rect 5120 600 5160 800
rect 10400 600 10440 800
rect -40 520 240 560
rect 280 520 560 560
rect 600 520 880 560
rect 920 520 1200 560
rect 1240 520 1520 560
rect 1560 520 1840 560
rect 1880 520 2160 560
rect 2200 520 2480 560
rect 2520 520 2800 560
rect 2840 520 3120 560
rect 3160 520 3440 560
rect 3480 520 3760 560
rect 3800 520 4080 560
rect 4120 520 4400 560
rect 4440 520 4720 560
rect 4760 520 5040 560
rect 5240 520 5520 560
rect 5560 520 5840 560
rect 5880 520 6160 560
rect 6200 520 6480 560
rect 6520 520 6800 560
rect 6840 520 7120 560
rect 7160 520 7440 560
rect 7480 520 7760 560
rect 7800 520 8080 560
rect 8120 520 8400 560
rect 8440 520 8720 560
rect 8760 520 9040 560
rect 9080 520 9360 560
rect 9400 520 9680 560
rect 9720 520 10000 560
rect 10040 520 10320 560
rect -40 -840 240 -800
rect 280 -840 560 -800
rect 600 -840 880 -800
rect 920 -840 1200 -800
rect 1240 -840 1520 -800
rect 1560 -840 1840 -800
rect 1880 -840 2160 -800
rect 2200 -840 2480 -800
rect 2520 -840 2800 -800
rect 2840 -840 3120 -800
rect 3160 -840 3440 -800
rect 3480 -840 3760 -800
rect 3800 -840 4080 -800
rect 4120 -840 4400 -800
rect 4440 -840 4720 -800
rect 4760 -840 5040 -800
rect 5240 -840 5520 -800
rect 5560 -840 5840 -800
rect 5880 -840 6160 -800
rect 6200 -840 6480 -800
rect 6520 -840 6800 -800
rect 6840 -840 7120 -800
rect 7160 -840 7440 -800
rect 7480 -840 7760 -800
rect 7800 -840 8080 -800
rect 8120 -840 8400 -800
rect 8440 -840 8720 -800
rect 8760 -840 9040 -800
rect 9080 -840 9360 -800
rect 9400 -840 9680 -800
rect 9720 -840 10000 -800
rect 10040 -840 10320 -800
rect -160 -1080 -120 -880
rect 5120 -1080 5160 -880
rect 10400 -1080 10440 -880
rect -40 -1160 240 -1120
rect 280 -1160 560 -1120
rect 600 -1160 880 -1120
rect 920 -1160 1200 -1120
rect 1240 -1160 1520 -1120
rect 1560 -1160 1840 -1120
rect 1880 -1160 2160 -1120
rect 2200 -1160 2480 -1120
rect 2520 -1160 2800 -1120
rect 2840 -1160 3120 -1120
rect 3160 -1160 3440 -1120
rect 3480 -1160 3760 -1120
rect 3800 -1160 4080 -1120
rect 4120 -1160 4400 -1120
rect 4440 -1160 4720 -1120
rect 4760 -1160 5040 -1120
rect 5240 -1160 5520 -1120
rect 5560 -1160 5840 -1120
rect 5880 -1160 6160 -1120
rect 6200 -1160 6480 -1120
rect 6520 -1160 6800 -1120
rect 6840 -1160 7120 -1120
rect 7160 -1160 7440 -1120
rect 7480 -1160 7760 -1120
rect 7800 -1160 8080 -1120
rect 8120 -1160 8400 -1120
rect 8440 -1160 8720 -1120
rect 8760 -1160 9040 -1120
rect 9080 -1160 9360 -1120
rect 9400 -1160 9680 -1120
rect 9720 -1160 10000 -1120
rect 10040 -1160 10320 -1120
rect -40 -1560 240 -1520
rect 280 -1560 560 -1520
rect 600 -1560 880 -1520
rect 920 -1560 1200 -1520
rect 1240 -1560 1520 -1520
rect 1560 -1560 1840 -1520
rect 1880 -1560 2160 -1520
rect 2200 -1560 2480 -1520
rect 2520 -1560 2800 -1520
rect 2840 -1560 3120 -1520
rect 3160 -1560 3440 -1520
rect 3480 -1560 3760 -1520
rect 3800 -1560 4080 -1520
rect 4120 -1560 4400 -1520
rect 4440 -1560 4720 -1520
rect 4760 -1560 5040 -1520
rect 5240 -1560 5520 -1520
rect 5560 -1560 5840 -1520
rect 5880 -1560 6160 -1520
rect 6200 -1560 6480 -1520
rect 6520 -1560 6800 -1520
rect 6840 -1560 7120 -1520
rect 7160 -1560 7440 -1520
rect 7480 -1560 7760 -1520
rect 7800 -1560 8080 -1520
rect 8120 -1560 8400 -1520
rect 8440 -1560 8720 -1520
rect 8760 -1560 9040 -1520
rect 9080 -1560 9360 -1520
rect 9400 -1560 9680 -1520
rect 9720 -1560 10000 -1520
rect 10040 -1560 10320 -1520
rect -160 -1800 -120 -1600
rect 5120 -1800 5160 -1600
rect 10400 -1800 10440 -1600
rect -40 -1880 240 -1840
rect 280 -1880 560 -1840
rect 600 -1880 880 -1840
rect 920 -1880 1200 -1840
rect 1240 -1880 1520 -1840
rect 1560 -1880 1840 -1840
rect 1880 -1880 2160 -1840
rect 2200 -1880 2480 -1840
rect 2520 -1880 2800 -1840
rect 2840 -1880 3120 -1840
rect 3160 -1880 3440 -1840
rect 3480 -1880 3760 -1840
rect 3800 -1880 4080 -1840
rect 4120 -1880 4400 -1840
rect 4440 -1880 4720 -1840
rect 4760 -1880 5040 -1840
rect 5240 -1880 5520 -1840
rect 5560 -1880 5840 -1840
rect 5880 -1880 6160 -1840
rect 6200 -1880 6480 -1840
rect 6520 -1880 6800 -1840
rect 6840 -1880 7120 -1840
rect 7160 -1880 7440 -1840
rect 7480 -1880 7760 -1840
rect 7800 -1880 8080 -1840
rect 8120 -1880 8400 -1840
rect 8440 -1880 8720 -1840
rect 8760 -1880 9040 -1840
rect 9080 -1880 9360 -1840
rect 9400 -1880 9680 -1840
rect 9720 -1880 10000 -1840
rect 10040 -1880 10320 -1840
rect -40 -3240 240 -3200
rect 280 -3240 560 -3200
rect 600 -3240 880 -3200
rect 920 -3240 1200 -3200
rect 1240 -3240 1520 -3200
rect 1560 -3240 1840 -3200
rect 1880 -3240 2160 -3200
rect 2200 -3240 2480 -3200
rect 2520 -3240 2800 -3200
rect 2840 -3240 3120 -3200
rect 3160 -3240 3440 -3200
rect 3480 -3240 3760 -3200
rect 3800 -3240 4080 -3200
rect 4120 -3240 4400 -3200
rect 4440 -3240 4720 -3200
rect 4760 -3240 5040 -3200
rect 5240 -3240 5520 -3200
rect 5560 -3240 5840 -3200
rect 5880 -3240 6160 -3200
rect 6200 -3240 6480 -3200
rect 6520 -3240 6800 -3200
rect 6840 -3240 7120 -3200
rect 7160 -3240 7440 -3200
rect 7480 -3240 7760 -3200
rect 7800 -3240 8080 -3200
rect 8120 -3240 8400 -3200
rect 8440 -3240 8720 -3200
rect 8760 -3240 9040 -3200
rect 9080 -3240 9360 -3200
rect 9400 -3240 9680 -3200
rect 9720 -3240 10000 -3200
rect 10040 -3240 10320 -3200
rect -160 -3480 -120 -3280
rect 5120 -3480 5160 -3280
rect 10400 -3480 10440 -3280
rect -40 -3560 240 -3520
rect 280 -3560 560 -3520
rect 600 -3560 880 -3520
rect 920 -3560 1200 -3520
rect 1240 -3560 1520 -3520
rect 1560 -3560 1840 -3520
rect 1880 -3560 2160 -3520
rect 2200 -3560 2480 -3520
rect 2520 -3560 2800 -3520
rect 2840 -3560 3120 -3520
rect 3160 -3560 3440 -3520
rect 3480 -3560 3760 -3520
rect 3800 -3560 4080 -3520
rect 4120 -3560 4400 -3520
rect 4440 -3560 4720 -3520
rect 4760 -3560 5040 -3520
rect 5240 -3560 5520 -3520
rect 5560 -3560 5840 -3520
rect 5880 -3560 6160 -3520
rect 6200 -3560 6480 -3520
rect 6520 -3560 6800 -3520
rect 6840 -3560 7120 -3520
rect 7160 -3560 7440 -3520
rect 7480 -3560 7760 -3520
rect 7800 -3560 8080 -3520
rect 8120 -3560 8400 -3520
rect 8440 -3560 8720 -3520
rect 8760 -3560 9040 -3520
rect 9080 -3560 9360 -3520
rect 9400 -3560 9680 -3520
rect 9720 -3560 10000 -3520
rect 10040 -3560 10320 -3520
<< poly >>
rect 0 760 200 780
rect 320 760 520 780
rect 640 760 840 780
rect 960 760 1160 780
rect 1280 760 1480 780
rect 1600 760 1800 780
rect 1920 760 2120 780
rect 2240 760 2440 780
rect 2560 760 2760 780
rect 2880 760 3080 780
rect 3200 760 3400 780
rect 3520 760 3720 780
rect 3840 760 4040 780
rect 4160 760 4360 780
rect 4480 760 4680 780
rect 4800 760 5000 780
rect 0 635 200 660
rect 0 605 10 635
rect 190 605 200 635
rect 0 600 200 605
rect 320 635 520 660
rect 320 605 330 635
rect 510 605 520 635
rect 320 600 520 605
rect 640 635 840 660
rect 640 605 650 635
rect 830 605 840 635
rect 640 600 840 605
rect 960 635 1160 660
rect 960 605 970 635
rect 1150 605 1160 635
rect 960 600 1160 605
rect 1280 635 1480 660
rect 1280 605 1290 635
rect 1470 605 1480 635
rect 1280 600 1480 605
rect 1600 635 1800 660
rect 1600 605 1610 635
rect 1790 605 1800 635
rect 1600 600 1800 605
rect 1920 635 2120 660
rect 1920 605 1930 635
rect 2110 605 2120 635
rect 1920 600 2120 605
rect 2240 635 2440 660
rect 2240 605 2250 635
rect 2430 605 2440 635
rect 2240 600 2440 605
rect 2560 635 2760 660
rect 2560 605 2570 635
rect 2750 605 2760 635
rect 2560 600 2760 605
rect 2880 635 3080 660
rect 2880 605 2890 635
rect 3070 605 3080 635
rect 2880 600 3080 605
rect 3200 635 3400 660
rect 3200 605 3210 635
rect 3390 605 3400 635
rect 3200 600 3400 605
rect 3520 635 3720 660
rect 3520 605 3530 635
rect 3710 605 3720 635
rect 3520 600 3720 605
rect 3840 635 4040 660
rect 3840 605 3850 635
rect 4030 605 4040 635
rect 3840 600 4040 605
rect 4160 635 4360 660
rect 4160 605 4170 635
rect 4350 605 4360 635
rect 4160 600 4360 605
rect 4480 635 4680 660
rect 4480 605 4490 635
rect 4670 605 4680 635
rect 4480 600 4680 605
rect 4800 635 5000 660
rect 4800 605 4810 635
rect 4990 605 5000 635
rect 4800 600 5000 605
rect 5280 760 5480 780
rect 5600 760 5800 780
rect 5920 760 6120 780
rect 6240 760 6440 780
rect 6560 760 6760 780
rect 6880 760 7080 780
rect 7200 760 7400 780
rect 7520 760 7720 780
rect 7840 760 8040 780
rect 8160 760 8360 780
rect 8480 760 8680 780
rect 8800 760 9000 780
rect 9120 760 9320 780
rect 9440 760 9640 780
rect 9760 760 9960 780
rect 10080 760 10280 780
rect 5280 635 5480 660
rect 5280 605 5290 635
rect 5470 605 5480 635
rect 5280 600 5480 605
rect 5600 635 5800 660
rect 5600 605 5610 635
rect 5790 605 5800 635
rect 5600 600 5800 605
rect 5920 635 6120 660
rect 5920 605 5930 635
rect 6110 605 6120 635
rect 5920 600 6120 605
rect 6240 635 6440 660
rect 6240 605 6250 635
rect 6430 605 6440 635
rect 6240 600 6440 605
rect 6560 635 6760 660
rect 6560 605 6570 635
rect 6750 605 6760 635
rect 6560 600 6760 605
rect 6880 635 7080 660
rect 6880 605 6890 635
rect 7070 605 7080 635
rect 6880 600 7080 605
rect 7200 635 7400 660
rect 7200 605 7210 635
rect 7390 605 7400 635
rect 7200 600 7400 605
rect 7520 635 7720 660
rect 7520 605 7530 635
rect 7710 605 7720 635
rect 7520 600 7720 605
rect 7840 635 8040 660
rect 7840 605 7850 635
rect 8030 605 8040 635
rect 7840 600 8040 605
rect 8160 635 8360 660
rect 8160 605 8170 635
rect 8350 605 8360 635
rect 8160 600 8360 605
rect 8480 635 8680 660
rect 8480 605 8490 635
rect 8670 605 8680 635
rect 8480 600 8680 605
rect 8800 635 9000 660
rect 8800 605 8810 635
rect 8990 605 9000 635
rect 8800 600 9000 605
rect 9120 635 9320 660
rect 9120 605 9130 635
rect 9310 605 9320 635
rect 9120 600 9320 605
rect 9440 635 9640 660
rect 9440 605 9450 635
rect 9630 605 9640 635
rect 9440 600 9640 605
rect 9760 635 9960 660
rect 9760 605 9770 635
rect 9950 605 9960 635
rect 9760 600 9960 605
rect 10080 635 10280 660
rect 10080 605 10090 635
rect 10270 605 10280 635
rect 10080 600 10280 605
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 100 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 100 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 100 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 100 1160 125
rect 1280 155 1480 160
rect 1280 125 1290 155
rect 1470 125 1480 155
rect 1280 100 1480 125
rect 1600 155 1800 160
rect 1600 125 1610 155
rect 1790 125 1800 155
rect 1600 100 1800 125
rect 1920 155 2120 160
rect 1920 125 1930 155
rect 2110 125 2120 155
rect 1920 100 2120 125
rect 2240 155 2440 160
rect 2240 125 2250 155
rect 2430 125 2440 155
rect 2240 100 2440 125
rect 2560 155 2760 160
rect 2560 125 2570 155
rect 2750 125 2760 155
rect 2560 100 2760 125
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 100 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 100 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 100 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 100 4040 125
rect 4160 155 4360 160
rect 4160 125 4170 155
rect 4350 125 4360 155
rect 4160 100 4360 125
rect 4480 155 4680 160
rect 4480 125 4490 155
rect 4670 125 4680 155
rect 4480 100 4680 125
rect 4800 155 5000 160
rect 4800 125 4810 155
rect 4990 125 5000 155
rect 4800 100 5000 125
rect 0 -20 200 0
rect 320 -20 520 0
rect 640 -20 840 0
rect 960 -20 1160 0
rect 1280 -20 1480 0
rect 1600 -20 1800 0
rect 1920 -20 2120 0
rect 2240 -20 2440 0
rect 2560 -20 2760 0
rect 2880 -20 3080 0
rect 3200 -20 3400 0
rect 3520 -20 3720 0
rect 3840 -20 4040 0
rect 4160 -20 4360 0
rect 4480 -20 4680 0
rect 4800 -20 5000 0
rect 5280 155 5480 160
rect 5280 125 5290 155
rect 5470 125 5480 155
rect 5280 100 5480 125
rect 5600 155 5800 160
rect 5600 125 5610 155
rect 5790 125 5800 155
rect 5600 100 5800 125
rect 5920 155 6120 160
rect 5920 125 5930 155
rect 6110 125 6120 155
rect 5920 100 6120 125
rect 6240 155 6440 160
rect 6240 125 6250 155
rect 6430 125 6440 155
rect 6240 100 6440 125
rect 6560 155 6760 160
rect 6560 125 6570 155
rect 6750 125 6760 155
rect 6560 100 6760 125
rect 6880 155 7080 160
rect 6880 125 6890 155
rect 7070 125 7080 155
rect 6880 100 7080 125
rect 7200 155 7400 160
rect 7200 125 7210 155
rect 7390 125 7400 155
rect 7200 100 7400 125
rect 7520 155 7720 160
rect 7520 125 7530 155
rect 7710 125 7720 155
rect 7520 100 7720 125
rect 7840 155 8040 160
rect 7840 125 7850 155
rect 8030 125 8040 155
rect 7840 100 8040 125
rect 8160 155 8360 160
rect 8160 125 8170 155
rect 8350 125 8360 155
rect 8160 100 8360 125
rect 8480 155 8680 160
rect 8480 125 8490 155
rect 8670 125 8680 155
rect 8480 100 8680 125
rect 8800 155 9000 160
rect 8800 125 8810 155
rect 8990 125 9000 155
rect 8800 100 9000 125
rect 9120 155 9320 160
rect 9120 125 9130 155
rect 9310 125 9320 155
rect 9120 100 9320 125
rect 9440 155 9640 160
rect 9440 125 9450 155
rect 9630 125 9640 155
rect 9440 100 9640 125
rect 9760 155 9960 160
rect 9760 125 9770 155
rect 9950 125 9960 155
rect 9760 100 9960 125
rect 10080 155 10280 160
rect 10080 125 10090 155
rect 10270 125 10280 155
rect 10080 100 10280 125
rect 5280 -20 5480 0
rect 5600 -20 5800 0
rect 5920 -20 6120 0
rect 6240 -20 6440 0
rect 6560 -20 6760 0
rect 6880 -20 7080 0
rect 7200 -20 7400 0
rect 7520 -20 7720 0
rect 7840 -20 8040 0
rect 8160 -20 8360 0
rect 8480 -20 8680 0
rect 8800 -20 9000 0
rect 9120 -20 9320 0
rect 9440 -20 9640 0
rect 9760 -20 9960 0
rect 10080 -20 10280 0
rect 0 -280 200 -260
rect 320 -280 520 -260
rect 640 -280 840 -260
rect 960 -280 1160 -260
rect 1280 -280 1480 -260
rect 1600 -280 1800 -260
rect 1920 -280 2120 -260
rect 2240 -280 2440 -260
rect 2560 -280 2760 -260
rect 2880 -280 3080 -260
rect 3200 -280 3400 -260
rect 3520 -280 3720 -260
rect 3840 -280 4040 -260
rect 4160 -280 4360 -260
rect 4480 -280 4680 -260
rect 4800 -280 5000 -260
rect 0 -405 200 -380
rect 0 -435 10 -405
rect 190 -435 200 -405
rect 0 -440 200 -435
rect 320 -405 520 -380
rect 320 -435 330 -405
rect 510 -435 520 -405
rect 320 -440 520 -435
rect 640 -405 840 -380
rect 640 -435 650 -405
rect 830 -435 840 -405
rect 640 -440 840 -435
rect 960 -405 1160 -380
rect 960 -435 970 -405
rect 1150 -435 1160 -405
rect 960 -440 1160 -435
rect 1280 -405 1480 -380
rect 1280 -435 1290 -405
rect 1470 -435 1480 -405
rect 1280 -440 1480 -435
rect 1600 -405 1800 -380
rect 1600 -435 1610 -405
rect 1790 -435 1800 -405
rect 1600 -440 1800 -435
rect 1920 -405 2120 -380
rect 1920 -435 1930 -405
rect 2110 -435 2120 -405
rect 1920 -440 2120 -435
rect 2240 -405 2440 -380
rect 2240 -435 2250 -405
rect 2430 -435 2440 -405
rect 2240 -440 2440 -435
rect 2560 -405 2760 -380
rect 2560 -435 2570 -405
rect 2750 -435 2760 -405
rect 2560 -440 2760 -435
rect 2880 -405 3080 -380
rect 2880 -435 2890 -405
rect 3070 -435 3080 -405
rect 2880 -440 3080 -435
rect 3200 -405 3400 -380
rect 3200 -435 3210 -405
rect 3390 -435 3400 -405
rect 3200 -440 3400 -435
rect 3520 -405 3720 -380
rect 3520 -435 3530 -405
rect 3710 -435 3720 -405
rect 3520 -440 3720 -435
rect 3840 -405 4040 -380
rect 3840 -435 3850 -405
rect 4030 -435 4040 -405
rect 3840 -440 4040 -435
rect 4160 -405 4360 -380
rect 4160 -435 4170 -405
rect 4350 -435 4360 -405
rect 4160 -440 4360 -435
rect 4480 -405 4680 -380
rect 4480 -435 4490 -405
rect 4670 -435 4680 -405
rect 4480 -440 4680 -435
rect 4800 -405 5000 -380
rect 4800 -435 4810 -405
rect 4990 -435 5000 -405
rect 4800 -440 5000 -435
rect 5280 -280 5480 -260
rect 5600 -280 5800 -260
rect 5920 -280 6120 -260
rect 6240 -280 6440 -260
rect 6560 -280 6760 -260
rect 6880 -280 7080 -260
rect 7200 -280 7400 -260
rect 7520 -280 7720 -260
rect 7840 -280 8040 -260
rect 8160 -280 8360 -260
rect 8480 -280 8680 -260
rect 8800 -280 9000 -260
rect 9120 -280 9320 -260
rect 9440 -280 9640 -260
rect 9760 -280 9960 -260
rect 10080 -280 10280 -260
rect 5280 -405 5480 -380
rect 5280 -435 5290 -405
rect 5470 -435 5480 -405
rect 5280 -440 5480 -435
rect 5600 -405 5800 -380
rect 5600 -435 5610 -405
rect 5790 -435 5800 -405
rect 5600 -440 5800 -435
rect 5920 -405 6120 -380
rect 5920 -435 5930 -405
rect 6110 -435 6120 -405
rect 5920 -440 6120 -435
rect 6240 -405 6440 -380
rect 6240 -435 6250 -405
rect 6430 -435 6440 -405
rect 6240 -440 6440 -435
rect 6560 -405 6760 -380
rect 6560 -435 6570 -405
rect 6750 -435 6760 -405
rect 6560 -440 6760 -435
rect 6880 -405 7080 -380
rect 6880 -435 6890 -405
rect 7070 -435 7080 -405
rect 6880 -440 7080 -435
rect 7200 -405 7400 -380
rect 7200 -435 7210 -405
rect 7390 -435 7400 -405
rect 7200 -440 7400 -435
rect 7520 -405 7720 -380
rect 7520 -435 7530 -405
rect 7710 -435 7720 -405
rect 7520 -440 7720 -435
rect 7840 -405 8040 -380
rect 7840 -435 7850 -405
rect 8030 -435 8040 -405
rect 7840 -440 8040 -435
rect 8160 -405 8360 -380
rect 8160 -435 8170 -405
rect 8350 -435 8360 -405
rect 8160 -440 8360 -435
rect 8480 -405 8680 -380
rect 8480 -435 8490 -405
rect 8670 -435 8680 -405
rect 8480 -440 8680 -435
rect 8800 -405 9000 -380
rect 8800 -435 8810 -405
rect 8990 -435 9000 -405
rect 8800 -440 9000 -435
rect 9120 -405 9320 -380
rect 9120 -435 9130 -405
rect 9310 -435 9320 -405
rect 9120 -440 9320 -435
rect 9440 -405 9640 -380
rect 9440 -435 9450 -405
rect 9630 -435 9640 -405
rect 9440 -440 9640 -435
rect 9760 -405 9960 -380
rect 9760 -435 9770 -405
rect 9950 -435 9960 -405
rect 9760 -440 9960 -435
rect 10080 -405 10280 -380
rect 10080 -435 10090 -405
rect 10270 -435 10280 -405
rect 10080 -440 10280 -435
rect 0 -885 200 -880
rect 0 -915 10 -885
rect 190 -915 200 -885
rect 0 -940 200 -915
rect 320 -885 520 -880
rect 320 -915 330 -885
rect 510 -915 520 -885
rect 320 -940 520 -915
rect 640 -885 840 -880
rect 640 -915 650 -885
rect 830 -915 840 -885
rect 640 -940 840 -915
rect 960 -885 1160 -880
rect 960 -915 970 -885
rect 1150 -915 1160 -885
rect 960 -940 1160 -915
rect 1280 -885 1480 -880
rect 1280 -915 1290 -885
rect 1470 -915 1480 -885
rect 1280 -940 1480 -915
rect 1600 -885 1800 -880
rect 1600 -915 1610 -885
rect 1790 -915 1800 -885
rect 1600 -940 1800 -915
rect 1920 -885 2120 -880
rect 1920 -915 1930 -885
rect 2110 -915 2120 -885
rect 1920 -940 2120 -915
rect 2240 -885 2440 -880
rect 2240 -915 2250 -885
rect 2430 -915 2440 -885
rect 2240 -940 2440 -915
rect 2560 -885 2760 -880
rect 2560 -915 2570 -885
rect 2750 -915 2760 -885
rect 2560 -940 2760 -915
rect 2880 -885 3080 -880
rect 2880 -915 2890 -885
rect 3070 -915 3080 -885
rect 2880 -940 3080 -915
rect 3200 -885 3400 -880
rect 3200 -915 3210 -885
rect 3390 -915 3400 -885
rect 3200 -940 3400 -915
rect 3520 -885 3720 -880
rect 3520 -915 3530 -885
rect 3710 -915 3720 -885
rect 3520 -940 3720 -915
rect 3840 -885 4040 -880
rect 3840 -915 3850 -885
rect 4030 -915 4040 -885
rect 3840 -940 4040 -915
rect 4160 -885 4360 -880
rect 4160 -915 4170 -885
rect 4350 -915 4360 -885
rect 4160 -940 4360 -915
rect 4480 -885 4680 -880
rect 4480 -915 4490 -885
rect 4670 -915 4680 -885
rect 4480 -940 4680 -915
rect 4800 -885 5000 -880
rect 4800 -915 4810 -885
rect 4990 -915 5000 -885
rect 4800 -940 5000 -915
rect 0 -1060 200 -1040
rect 320 -1060 520 -1040
rect 640 -1060 840 -1040
rect 960 -1060 1160 -1040
rect 1280 -1060 1480 -1040
rect 1600 -1060 1800 -1040
rect 1920 -1060 2120 -1040
rect 2240 -1060 2440 -1040
rect 2560 -1060 2760 -1040
rect 2880 -1060 3080 -1040
rect 3200 -1060 3400 -1040
rect 3520 -1060 3720 -1040
rect 3840 -1060 4040 -1040
rect 4160 -1060 4360 -1040
rect 4480 -1060 4680 -1040
rect 4800 -1060 5000 -1040
rect 5280 -885 5480 -880
rect 5280 -915 5290 -885
rect 5470 -915 5480 -885
rect 5280 -940 5480 -915
rect 5600 -885 5800 -880
rect 5600 -915 5610 -885
rect 5790 -915 5800 -885
rect 5600 -940 5800 -915
rect 5920 -885 6120 -880
rect 5920 -915 5930 -885
rect 6110 -915 6120 -885
rect 5920 -940 6120 -915
rect 6240 -885 6440 -880
rect 6240 -915 6250 -885
rect 6430 -915 6440 -885
rect 6240 -940 6440 -915
rect 6560 -885 6760 -880
rect 6560 -915 6570 -885
rect 6750 -915 6760 -885
rect 6560 -940 6760 -915
rect 6880 -885 7080 -880
rect 6880 -915 6890 -885
rect 7070 -915 7080 -885
rect 6880 -940 7080 -915
rect 7200 -885 7400 -880
rect 7200 -915 7210 -885
rect 7390 -915 7400 -885
rect 7200 -940 7400 -915
rect 7520 -885 7720 -880
rect 7520 -915 7530 -885
rect 7710 -915 7720 -885
rect 7520 -940 7720 -915
rect 7840 -885 8040 -880
rect 7840 -915 7850 -885
rect 8030 -915 8040 -885
rect 7840 -940 8040 -915
rect 8160 -885 8360 -880
rect 8160 -915 8170 -885
rect 8350 -915 8360 -885
rect 8160 -940 8360 -915
rect 8480 -885 8680 -880
rect 8480 -915 8490 -885
rect 8670 -915 8680 -885
rect 8480 -940 8680 -915
rect 8800 -885 9000 -880
rect 8800 -915 8810 -885
rect 8990 -915 9000 -885
rect 8800 -940 9000 -915
rect 9120 -885 9320 -880
rect 9120 -915 9130 -885
rect 9310 -915 9320 -885
rect 9120 -940 9320 -915
rect 9440 -885 9640 -880
rect 9440 -915 9450 -885
rect 9630 -915 9640 -885
rect 9440 -940 9640 -915
rect 9760 -885 9960 -880
rect 9760 -915 9770 -885
rect 9950 -915 9960 -885
rect 9760 -940 9960 -915
rect 10080 -885 10280 -880
rect 10080 -915 10090 -885
rect 10270 -915 10280 -885
rect 10080 -940 10280 -915
rect 5280 -1060 5480 -1040
rect 5600 -1060 5800 -1040
rect 5920 -1060 6120 -1040
rect 6240 -1060 6440 -1040
rect 6560 -1060 6760 -1040
rect 6880 -1060 7080 -1040
rect 7200 -1060 7400 -1040
rect 7520 -1060 7720 -1040
rect 7840 -1060 8040 -1040
rect 8160 -1060 8360 -1040
rect 8480 -1060 8680 -1040
rect 8800 -1060 9000 -1040
rect 9120 -1060 9320 -1040
rect 9440 -1060 9640 -1040
rect 9760 -1060 9960 -1040
rect 10080 -1060 10280 -1040
rect 0 -1640 200 -1620
rect 320 -1640 520 -1620
rect 640 -1640 840 -1620
rect 960 -1640 1160 -1620
rect 1280 -1640 1480 -1620
rect 1600 -1640 1800 -1620
rect 1920 -1640 2120 -1620
rect 2240 -1640 2440 -1620
rect 2560 -1640 2760 -1620
rect 2880 -1640 3080 -1620
rect 3200 -1640 3400 -1620
rect 3520 -1640 3720 -1620
rect 3840 -1640 4040 -1620
rect 4160 -1640 4360 -1620
rect 4480 -1640 4680 -1620
rect 4800 -1640 5000 -1620
rect 0 -1765 200 -1740
rect 0 -1795 10 -1765
rect 190 -1795 200 -1765
rect 0 -1800 200 -1795
rect 320 -1765 520 -1740
rect 320 -1795 330 -1765
rect 510 -1795 520 -1765
rect 320 -1800 520 -1795
rect 640 -1765 840 -1740
rect 640 -1795 650 -1765
rect 830 -1795 840 -1765
rect 640 -1800 840 -1795
rect 960 -1765 1160 -1740
rect 960 -1795 970 -1765
rect 1150 -1795 1160 -1765
rect 960 -1800 1160 -1795
rect 1280 -1765 1480 -1740
rect 1280 -1795 1290 -1765
rect 1470 -1795 1480 -1765
rect 1280 -1800 1480 -1795
rect 1600 -1765 1800 -1740
rect 1600 -1795 1610 -1765
rect 1790 -1795 1800 -1765
rect 1600 -1800 1800 -1795
rect 1920 -1765 2120 -1740
rect 1920 -1795 1930 -1765
rect 2110 -1795 2120 -1765
rect 1920 -1800 2120 -1795
rect 2240 -1765 2440 -1740
rect 2240 -1795 2250 -1765
rect 2430 -1795 2440 -1765
rect 2240 -1800 2440 -1795
rect 2560 -1765 2760 -1740
rect 2560 -1795 2570 -1765
rect 2750 -1795 2760 -1765
rect 2560 -1800 2760 -1795
rect 2880 -1765 3080 -1740
rect 2880 -1795 2890 -1765
rect 3070 -1795 3080 -1765
rect 2880 -1800 3080 -1795
rect 3200 -1765 3400 -1740
rect 3200 -1795 3210 -1765
rect 3390 -1795 3400 -1765
rect 3200 -1800 3400 -1795
rect 3520 -1765 3720 -1740
rect 3520 -1795 3530 -1765
rect 3710 -1795 3720 -1765
rect 3520 -1800 3720 -1795
rect 3840 -1765 4040 -1740
rect 3840 -1795 3850 -1765
rect 4030 -1795 4040 -1765
rect 3840 -1800 4040 -1795
rect 4160 -1765 4360 -1740
rect 4160 -1795 4170 -1765
rect 4350 -1795 4360 -1765
rect 4160 -1800 4360 -1795
rect 4480 -1765 4680 -1740
rect 4480 -1795 4490 -1765
rect 4670 -1795 4680 -1765
rect 4480 -1800 4680 -1795
rect 4800 -1765 5000 -1740
rect 4800 -1795 4810 -1765
rect 4990 -1795 5000 -1765
rect 4800 -1800 5000 -1795
rect 5280 -1640 5480 -1620
rect 5600 -1640 5800 -1620
rect 5920 -1640 6120 -1620
rect 6240 -1640 6440 -1620
rect 6560 -1640 6760 -1620
rect 6880 -1640 7080 -1620
rect 7200 -1640 7400 -1620
rect 7520 -1640 7720 -1620
rect 7840 -1640 8040 -1620
rect 8160 -1640 8360 -1620
rect 8480 -1640 8680 -1620
rect 8800 -1640 9000 -1620
rect 9120 -1640 9320 -1620
rect 9440 -1640 9640 -1620
rect 9760 -1640 9960 -1620
rect 10080 -1640 10280 -1620
rect 5280 -1765 5480 -1740
rect 5280 -1795 5290 -1765
rect 5470 -1795 5480 -1765
rect 5280 -1800 5480 -1795
rect 5600 -1765 5800 -1740
rect 5600 -1795 5610 -1765
rect 5790 -1795 5800 -1765
rect 5600 -1800 5800 -1795
rect 5920 -1765 6120 -1740
rect 5920 -1795 5930 -1765
rect 6110 -1795 6120 -1765
rect 5920 -1800 6120 -1795
rect 6240 -1765 6440 -1740
rect 6240 -1795 6250 -1765
rect 6430 -1795 6440 -1765
rect 6240 -1800 6440 -1795
rect 6560 -1765 6760 -1740
rect 6560 -1795 6570 -1765
rect 6750 -1795 6760 -1765
rect 6560 -1800 6760 -1795
rect 6880 -1765 7080 -1740
rect 6880 -1795 6890 -1765
rect 7070 -1795 7080 -1765
rect 6880 -1800 7080 -1795
rect 7200 -1765 7400 -1740
rect 7200 -1795 7210 -1765
rect 7390 -1795 7400 -1765
rect 7200 -1800 7400 -1795
rect 7520 -1765 7720 -1740
rect 7520 -1795 7530 -1765
rect 7710 -1795 7720 -1765
rect 7520 -1800 7720 -1795
rect 7840 -1765 8040 -1740
rect 7840 -1795 7850 -1765
rect 8030 -1795 8040 -1765
rect 7840 -1800 8040 -1795
rect 8160 -1765 8360 -1740
rect 8160 -1795 8170 -1765
rect 8350 -1795 8360 -1765
rect 8160 -1800 8360 -1795
rect 8480 -1765 8680 -1740
rect 8480 -1795 8490 -1765
rect 8670 -1795 8680 -1765
rect 8480 -1800 8680 -1795
rect 8800 -1765 9000 -1740
rect 8800 -1795 8810 -1765
rect 8990 -1795 9000 -1765
rect 8800 -1800 9000 -1795
rect 9120 -1765 9320 -1740
rect 9120 -1795 9130 -1765
rect 9310 -1795 9320 -1765
rect 9120 -1800 9320 -1795
rect 9440 -1765 9640 -1740
rect 9440 -1795 9450 -1765
rect 9630 -1795 9640 -1765
rect 9440 -1800 9640 -1795
rect 9760 -1765 9960 -1740
rect 9760 -1795 9770 -1765
rect 9950 -1795 9960 -1765
rect 9760 -1800 9960 -1795
rect 10080 -1765 10280 -1740
rect 10080 -1795 10090 -1765
rect 10270 -1795 10280 -1765
rect 10080 -1800 10280 -1795
rect 0 -2245 200 -2240
rect 0 -2275 10 -2245
rect 190 -2275 200 -2245
rect 0 -2300 200 -2275
rect 320 -2245 520 -2240
rect 320 -2275 330 -2245
rect 510 -2275 520 -2245
rect 320 -2300 520 -2275
rect 640 -2245 840 -2240
rect 640 -2275 650 -2245
rect 830 -2275 840 -2245
rect 640 -2300 840 -2275
rect 960 -2245 1160 -2240
rect 960 -2275 970 -2245
rect 1150 -2275 1160 -2245
rect 960 -2300 1160 -2275
rect 1280 -2245 1480 -2240
rect 1280 -2275 1290 -2245
rect 1470 -2275 1480 -2245
rect 1280 -2300 1480 -2275
rect 1600 -2245 1800 -2240
rect 1600 -2275 1610 -2245
rect 1790 -2275 1800 -2245
rect 1600 -2300 1800 -2275
rect 1920 -2245 2120 -2240
rect 1920 -2275 1930 -2245
rect 2110 -2275 2120 -2245
rect 1920 -2300 2120 -2275
rect 2240 -2245 2440 -2240
rect 2240 -2275 2250 -2245
rect 2430 -2275 2440 -2245
rect 2240 -2300 2440 -2275
rect 2560 -2245 2760 -2240
rect 2560 -2275 2570 -2245
rect 2750 -2275 2760 -2245
rect 2560 -2300 2760 -2275
rect 2880 -2245 3080 -2240
rect 2880 -2275 2890 -2245
rect 3070 -2275 3080 -2245
rect 2880 -2300 3080 -2275
rect 3200 -2245 3400 -2240
rect 3200 -2275 3210 -2245
rect 3390 -2275 3400 -2245
rect 3200 -2300 3400 -2275
rect 3520 -2245 3720 -2240
rect 3520 -2275 3530 -2245
rect 3710 -2275 3720 -2245
rect 3520 -2300 3720 -2275
rect 3840 -2245 4040 -2240
rect 3840 -2275 3850 -2245
rect 4030 -2275 4040 -2245
rect 3840 -2300 4040 -2275
rect 4160 -2245 4360 -2240
rect 4160 -2275 4170 -2245
rect 4350 -2275 4360 -2245
rect 4160 -2300 4360 -2275
rect 4480 -2245 4680 -2240
rect 4480 -2275 4490 -2245
rect 4670 -2275 4680 -2245
rect 4480 -2300 4680 -2275
rect 4800 -2245 5000 -2240
rect 4800 -2275 4810 -2245
rect 4990 -2275 5000 -2245
rect 4800 -2300 5000 -2275
rect 0 -2420 200 -2400
rect 320 -2420 520 -2400
rect 640 -2420 840 -2400
rect 960 -2420 1160 -2400
rect 1280 -2420 1480 -2400
rect 1600 -2420 1800 -2400
rect 1920 -2420 2120 -2400
rect 2240 -2420 2440 -2400
rect 2560 -2420 2760 -2400
rect 2880 -2420 3080 -2400
rect 3200 -2420 3400 -2400
rect 3520 -2420 3720 -2400
rect 3840 -2420 4040 -2400
rect 4160 -2420 4360 -2400
rect 4480 -2420 4680 -2400
rect 4800 -2420 5000 -2400
rect 5280 -2245 5480 -2240
rect 5280 -2275 5290 -2245
rect 5470 -2275 5480 -2245
rect 5280 -2300 5480 -2275
rect 5600 -2245 5800 -2240
rect 5600 -2275 5610 -2245
rect 5790 -2275 5800 -2245
rect 5600 -2300 5800 -2275
rect 5920 -2245 6120 -2240
rect 5920 -2275 5930 -2245
rect 6110 -2275 6120 -2245
rect 5920 -2300 6120 -2275
rect 6240 -2245 6440 -2240
rect 6240 -2275 6250 -2245
rect 6430 -2275 6440 -2245
rect 6240 -2300 6440 -2275
rect 6560 -2245 6760 -2240
rect 6560 -2275 6570 -2245
rect 6750 -2275 6760 -2245
rect 6560 -2300 6760 -2275
rect 6880 -2245 7080 -2240
rect 6880 -2275 6890 -2245
rect 7070 -2275 7080 -2245
rect 6880 -2300 7080 -2275
rect 7200 -2245 7400 -2240
rect 7200 -2275 7210 -2245
rect 7390 -2275 7400 -2245
rect 7200 -2300 7400 -2275
rect 7520 -2245 7720 -2240
rect 7520 -2275 7530 -2245
rect 7710 -2275 7720 -2245
rect 7520 -2300 7720 -2275
rect 7840 -2245 8040 -2240
rect 7840 -2275 7850 -2245
rect 8030 -2275 8040 -2245
rect 7840 -2300 8040 -2275
rect 8160 -2245 8360 -2240
rect 8160 -2275 8170 -2245
rect 8350 -2275 8360 -2245
rect 8160 -2300 8360 -2275
rect 8480 -2245 8680 -2240
rect 8480 -2275 8490 -2245
rect 8670 -2275 8680 -2245
rect 8480 -2300 8680 -2275
rect 8800 -2245 9000 -2240
rect 8800 -2275 8810 -2245
rect 8990 -2275 9000 -2245
rect 8800 -2300 9000 -2275
rect 9120 -2245 9320 -2240
rect 9120 -2275 9130 -2245
rect 9310 -2275 9320 -2245
rect 9120 -2300 9320 -2275
rect 9440 -2245 9640 -2240
rect 9440 -2275 9450 -2245
rect 9630 -2275 9640 -2245
rect 9440 -2300 9640 -2275
rect 9760 -2245 9960 -2240
rect 9760 -2275 9770 -2245
rect 9950 -2275 9960 -2245
rect 9760 -2300 9960 -2275
rect 10080 -2245 10280 -2240
rect 10080 -2275 10090 -2245
rect 10270 -2275 10280 -2245
rect 10080 -2300 10280 -2275
rect 5280 -2420 5480 -2400
rect 5600 -2420 5800 -2400
rect 5920 -2420 6120 -2400
rect 6240 -2420 6440 -2400
rect 6560 -2420 6760 -2400
rect 6880 -2420 7080 -2400
rect 7200 -2420 7400 -2400
rect 7520 -2420 7720 -2400
rect 7840 -2420 8040 -2400
rect 8160 -2420 8360 -2400
rect 8480 -2420 8680 -2400
rect 8800 -2420 9000 -2400
rect 9120 -2420 9320 -2400
rect 9440 -2420 9640 -2400
rect 9760 -2420 9960 -2400
rect 10080 -2420 10280 -2400
rect 0 -2680 200 -2660
rect 320 -2680 520 -2660
rect 640 -2680 840 -2660
rect 960 -2680 1160 -2660
rect 1280 -2680 1480 -2660
rect 1600 -2680 1800 -2660
rect 1920 -2680 2120 -2660
rect 2240 -2680 2440 -2660
rect 2560 -2680 2760 -2660
rect 2880 -2680 3080 -2660
rect 3200 -2680 3400 -2660
rect 3520 -2680 3720 -2660
rect 3840 -2680 4040 -2660
rect 4160 -2680 4360 -2660
rect 4480 -2680 4680 -2660
rect 4800 -2680 5000 -2660
rect 0 -2805 200 -2780
rect 0 -2835 10 -2805
rect 190 -2835 200 -2805
rect 0 -2840 200 -2835
rect 320 -2805 520 -2780
rect 320 -2835 330 -2805
rect 510 -2835 520 -2805
rect 320 -2840 520 -2835
rect 640 -2805 840 -2780
rect 640 -2835 650 -2805
rect 830 -2835 840 -2805
rect 640 -2840 840 -2835
rect 960 -2805 1160 -2780
rect 960 -2835 970 -2805
rect 1150 -2835 1160 -2805
rect 960 -2840 1160 -2835
rect 1280 -2805 1480 -2780
rect 1280 -2835 1290 -2805
rect 1470 -2835 1480 -2805
rect 1280 -2840 1480 -2835
rect 1600 -2805 1800 -2780
rect 1600 -2835 1610 -2805
rect 1790 -2835 1800 -2805
rect 1600 -2840 1800 -2835
rect 1920 -2805 2120 -2780
rect 1920 -2835 1930 -2805
rect 2110 -2835 2120 -2805
rect 1920 -2840 2120 -2835
rect 2240 -2805 2440 -2780
rect 2240 -2835 2250 -2805
rect 2430 -2835 2440 -2805
rect 2240 -2840 2440 -2835
rect 2560 -2805 2760 -2780
rect 2560 -2835 2570 -2805
rect 2750 -2835 2760 -2805
rect 2560 -2840 2760 -2835
rect 2880 -2805 3080 -2780
rect 2880 -2835 2890 -2805
rect 3070 -2835 3080 -2805
rect 2880 -2840 3080 -2835
rect 3200 -2805 3400 -2780
rect 3200 -2835 3210 -2805
rect 3390 -2835 3400 -2805
rect 3200 -2840 3400 -2835
rect 3520 -2805 3720 -2780
rect 3520 -2835 3530 -2805
rect 3710 -2835 3720 -2805
rect 3520 -2840 3720 -2835
rect 3840 -2805 4040 -2780
rect 3840 -2835 3850 -2805
rect 4030 -2835 4040 -2805
rect 3840 -2840 4040 -2835
rect 4160 -2805 4360 -2780
rect 4160 -2835 4170 -2805
rect 4350 -2835 4360 -2805
rect 4160 -2840 4360 -2835
rect 4480 -2805 4680 -2780
rect 4480 -2835 4490 -2805
rect 4670 -2835 4680 -2805
rect 4480 -2840 4680 -2835
rect 4800 -2805 5000 -2780
rect 4800 -2835 4810 -2805
rect 4990 -2835 5000 -2805
rect 4800 -2840 5000 -2835
rect 5280 -2680 5480 -2660
rect 5600 -2680 5800 -2660
rect 5920 -2680 6120 -2660
rect 6240 -2680 6440 -2660
rect 6560 -2680 6760 -2660
rect 6880 -2680 7080 -2660
rect 7200 -2680 7400 -2660
rect 7520 -2680 7720 -2660
rect 7840 -2680 8040 -2660
rect 8160 -2680 8360 -2660
rect 8480 -2680 8680 -2660
rect 8800 -2680 9000 -2660
rect 9120 -2680 9320 -2660
rect 9440 -2680 9640 -2660
rect 9760 -2680 9960 -2660
rect 10080 -2680 10280 -2660
rect 5280 -2805 5480 -2780
rect 5280 -2835 5290 -2805
rect 5470 -2835 5480 -2805
rect 5280 -2840 5480 -2835
rect 5600 -2805 5800 -2780
rect 5600 -2835 5610 -2805
rect 5790 -2835 5800 -2805
rect 5600 -2840 5800 -2835
rect 5920 -2805 6120 -2780
rect 5920 -2835 5930 -2805
rect 6110 -2835 6120 -2805
rect 5920 -2840 6120 -2835
rect 6240 -2805 6440 -2780
rect 6240 -2835 6250 -2805
rect 6430 -2835 6440 -2805
rect 6240 -2840 6440 -2835
rect 6560 -2805 6760 -2780
rect 6560 -2835 6570 -2805
rect 6750 -2835 6760 -2805
rect 6560 -2840 6760 -2835
rect 6880 -2805 7080 -2780
rect 6880 -2835 6890 -2805
rect 7070 -2835 7080 -2805
rect 6880 -2840 7080 -2835
rect 7200 -2805 7400 -2780
rect 7200 -2835 7210 -2805
rect 7390 -2835 7400 -2805
rect 7200 -2840 7400 -2835
rect 7520 -2805 7720 -2780
rect 7520 -2835 7530 -2805
rect 7710 -2835 7720 -2805
rect 7520 -2840 7720 -2835
rect 7840 -2805 8040 -2780
rect 7840 -2835 7850 -2805
rect 8030 -2835 8040 -2805
rect 7840 -2840 8040 -2835
rect 8160 -2805 8360 -2780
rect 8160 -2835 8170 -2805
rect 8350 -2835 8360 -2805
rect 8160 -2840 8360 -2835
rect 8480 -2805 8680 -2780
rect 8480 -2835 8490 -2805
rect 8670 -2835 8680 -2805
rect 8480 -2840 8680 -2835
rect 8800 -2805 9000 -2780
rect 8800 -2835 8810 -2805
rect 8990 -2835 9000 -2805
rect 8800 -2840 9000 -2835
rect 9120 -2805 9320 -2780
rect 9120 -2835 9130 -2805
rect 9310 -2835 9320 -2805
rect 9120 -2840 9320 -2835
rect 9440 -2805 9640 -2780
rect 9440 -2835 9450 -2805
rect 9630 -2835 9640 -2805
rect 9440 -2840 9640 -2835
rect 9760 -2805 9960 -2780
rect 9760 -2835 9770 -2805
rect 9950 -2835 9960 -2805
rect 9760 -2840 9960 -2835
rect 10080 -2805 10280 -2780
rect 10080 -2835 10090 -2805
rect 10270 -2835 10280 -2805
rect 10080 -2840 10280 -2835
rect 0 -3285 200 -3280
rect 0 -3315 10 -3285
rect 190 -3315 200 -3285
rect 0 -3340 200 -3315
rect 320 -3285 520 -3280
rect 320 -3315 330 -3285
rect 510 -3315 520 -3285
rect 320 -3340 520 -3315
rect 640 -3285 840 -3280
rect 640 -3315 650 -3285
rect 830 -3315 840 -3285
rect 640 -3340 840 -3315
rect 960 -3285 1160 -3280
rect 960 -3315 970 -3285
rect 1150 -3315 1160 -3285
rect 960 -3340 1160 -3315
rect 1280 -3285 1480 -3280
rect 1280 -3315 1290 -3285
rect 1470 -3315 1480 -3285
rect 1280 -3340 1480 -3315
rect 1600 -3285 1800 -3280
rect 1600 -3315 1610 -3285
rect 1790 -3315 1800 -3285
rect 1600 -3340 1800 -3315
rect 1920 -3285 2120 -3280
rect 1920 -3315 1930 -3285
rect 2110 -3315 2120 -3285
rect 1920 -3340 2120 -3315
rect 2240 -3285 2440 -3280
rect 2240 -3315 2250 -3285
rect 2430 -3315 2440 -3285
rect 2240 -3340 2440 -3315
rect 2560 -3285 2760 -3280
rect 2560 -3315 2570 -3285
rect 2750 -3315 2760 -3285
rect 2560 -3340 2760 -3315
rect 2880 -3285 3080 -3280
rect 2880 -3315 2890 -3285
rect 3070 -3315 3080 -3285
rect 2880 -3340 3080 -3315
rect 3200 -3285 3400 -3280
rect 3200 -3315 3210 -3285
rect 3390 -3315 3400 -3285
rect 3200 -3340 3400 -3315
rect 3520 -3285 3720 -3280
rect 3520 -3315 3530 -3285
rect 3710 -3315 3720 -3285
rect 3520 -3340 3720 -3315
rect 3840 -3285 4040 -3280
rect 3840 -3315 3850 -3285
rect 4030 -3315 4040 -3285
rect 3840 -3340 4040 -3315
rect 4160 -3285 4360 -3280
rect 4160 -3315 4170 -3285
rect 4350 -3315 4360 -3285
rect 4160 -3340 4360 -3315
rect 4480 -3285 4680 -3280
rect 4480 -3315 4490 -3285
rect 4670 -3315 4680 -3285
rect 4480 -3340 4680 -3315
rect 4800 -3285 5000 -3280
rect 4800 -3315 4810 -3285
rect 4990 -3315 5000 -3285
rect 4800 -3340 5000 -3315
rect 0 -3460 200 -3440
rect 320 -3460 520 -3440
rect 640 -3460 840 -3440
rect 960 -3460 1160 -3440
rect 1280 -3460 1480 -3440
rect 1600 -3460 1800 -3440
rect 1920 -3460 2120 -3440
rect 2240 -3460 2440 -3440
rect 2560 -3460 2760 -3440
rect 2880 -3460 3080 -3440
rect 3200 -3460 3400 -3440
rect 3520 -3460 3720 -3440
rect 3840 -3460 4040 -3440
rect 4160 -3460 4360 -3440
rect 4480 -3460 4680 -3440
rect 4800 -3460 5000 -3440
rect 5280 -3285 5480 -3280
rect 5280 -3315 5290 -3285
rect 5470 -3315 5480 -3285
rect 5280 -3340 5480 -3315
rect 5600 -3285 5800 -3280
rect 5600 -3315 5610 -3285
rect 5790 -3315 5800 -3285
rect 5600 -3340 5800 -3315
rect 5920 -3285 6120 -3280
rect 5920 -3315 5930 -3285
rect 6110 -3315 6120 -3285
rect 5920 -3340 6120 -3315
rect 6240 -3285 6440 -3280
rect 6240 -3315 6250 -3285
rect 6430 -3315 6440 -3285
rect 6240 -3340 6440 -3315
rect 6560 -3285 6760 -3280
rect 6560 -3315 6570 -3285
rect 6750 -3315 6760 -3285
rect 6560 -3340 6760 -3315
rect 6880 -3285 7080 -3280
rect 6880 -3315 6890 -3285
rect 7070 -3315 7080 -3285
rect 6880 -3340 7080 -3315
rect 7200 -3285 7400 -3280
rect 7200 -3315 7210 -3285
rect 7390 -3315 7400 -3285
rect 7200 -3340 7400 -3315
rect 7520 -3285 7720 -3280
rect 7520 -3315 7530 -3285
rect 7710 -3315 7720 -3285
rect 7520 -3340 7720 -3315
rect 7840 -3285 8040 -3280
rect 7840 -3315 7850 -3285
rect 8030 -3315 8040 -3285
rect 7840 -3340 8040 -3315
rect 8160 -3285 8360 -3280
rect 8160 -3315 8170 -3285
rect 8350 -3315 8360 -3285
rect 8160 -3340 8360 -3315
rect 8480 -3285 8680 -3280
rect 8480 -3315 8490 -3285
rect 8670 -3315 8680 -3285
rect 8480 -3340 8680 -3315
rect 8800 -3285 9000 -3280
rect 8800 -3315 8810 -3285
rect 8990 -3315 9000 -3285
rect 8800 -3340 9000 -3315
rect 9120 -3285 9320 -3280
rect 9120 -3315 9130 -3285
rect 9310 -3315 9320 -3285
rect 9120 -3340 9320 -3315
rect 9440 -3285 9640 -3280
rect 9440 -3315 9450 -3285
rect 9630 -3315 9640 -3285
rect 9440 -3340 9640 -3315
rect 9760 -3285 9960 -3280
rect 9760 -3315 9770 -3285
rect 9950 -3315 9960 -3285
rect 9760 -3340 9960 -3315
rect 10080 -3285 10280 -3280
rect 10080 -3315 10090 -3285
rect 10270 -3315 10280 -3285
rect 10080 -3340 10280 -3315
rect 5280 -3460 5480 -3440
rect 5600 -3460 5800 -3440
rect 5920 -3460 6120 -3440
rect 6240 -3460 6440 -3440
rect 6560 -3460 6760 -3440
rect 6880 -3460 7080 -3440
rect 7200 -3460 7400 -3440
rect 7520 -3460 7720 -3440
rect 7840 -3460 8040 -3440
rect 8160 -3460 8360 -3440
rect 8480 -3460 8680 -3440
rect 8800 -3460 9000 -3440
rect 9120 -3460 9320 -3440
rect 9440 -3460 9640 -3440
rect 9760 -3460 9960 -3440
rect 10080 -3460 10280 -3440
<< polycont >>
rect 10 605 190 635
rect 330 605 510 635
rect 650 605 830 635
rect 970 605 1150 635
rect 1290 605 1470 635
rect 1610 605 1790 635
rect 1930 605 2110 635
rect 2250 605 2430 635
rect 2570 605 2750 635
rect 2890 605 3070 635
rect 3210 605 3390 635
rect 3530 605 3710 635
rect 3850 605 4030 635
rect 4170 605 4350 635
rect 4490 605 4670 635
rect 4810 605 4990 635
rect 5290 605 5470 635
rect 5610 605 5790 635
rect 5930 605 6110 635
rect 6250 605 6430 635
rect 6570 605 6750 635
rect 6890 605 7070 635
rect 7210 605 7390 635
rect 7530 605 7710 635
rect 7850 605 8030 635
rect 8170 605 8350 635
rect 8490 605 8670 635
rect 8810 605 8990 635
rect 9130 605 9310 635
rect 9450 605 9630 635
rect 9770 605 9950 635
rect 10090 605 10270 635
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect 1290 125 1470 155
rect 1610 125 1790 155
rect 1930 125 2110 155
rect 2250 125 2430 155
rect 2570 125 2750 155
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3850 125 4030 155
rect 4170 125 4350 155
rect 4490 125 4670 155
rect 4810 125 4990 155
rect 5290 125 5470 155
rect 5610 125 5790 155
rect 5930 125 6110 155
rect 6250 125 6430 155
rect 6570 125 6750 155
rect 6890 125 7070 155
rect 7210 125 7390 155
rect 7530 125 7710 155
rect 7850 125 8030 155
rect 8170 125 8350 155
rect 8490 125 8670 155
rect 8810 125 8990 155
rect 9130 125 9310 155
rect 9450 125 9630 155
rect 9770 125 9950 155
rect 10090 125 10270 155
rect 10 -435 190 -405
rect 330 -435 510 -405
rect 650 -435 830 -405
rect 970 -435 1150 -405
rect 1290 -435 1470 -405
rect 1610 -435 1790 -405
rect 1930 -435 2110 -405
rect 2250 -435 2430 -405
rect 2570 -435 2750 -405
rect 2890 -435 3070 -405
rect 3210 -435 3390 -405
rect 3530 -435 3710 -405
rect 3850 -435 4030 -405
rect 4170 -435 4350 -405
rect 4490 -435 4670 -405
rect 4810 -435 4990 -405
rect 5290 -435 5470 -405
rect 5610 -435 5790 -405
rect 5930 -435 6110 -405
rect 6250 -435 6430 -405
rect 6570 -435 6750 -405
rect 6890 -435 7070 -405
rect 7210 -435 7390 -405
rect 7530 -435 7710 -405
rect 7850 -435 8030 -405
rect 8170 -435 8350 -405
rect 8490 -435 8670 -405
rect 8810 -435 8990 -405
rect 9130 -435 9310 -405
rect 9450 -435 9630 -405
rect 9770 -435 9950 -405
rect 10090 -435 10270 -405
rect 10 -915 190 -885
rect 330 -915 510 -885
rect 650 -915 830 -885
rect 970 -915 1150 -885
rect 1290 -915 1470 -885
rect 1610 -915 1790 -885
rect 1930 -915 2110 -885
rect 2250 -915 2430 -885
rect 2570 -915 2750 -885
rect 2890 -915 3070 -885
rect 3210 -915 3390 -885
rect 3530 -915 3710 -885
rect 3850 -915 4030 -885
rect 4170 -915 4350 -885
rect 4490 -915 4670 -885
rect 4810 -915 4990 -885
rect 5290 -915 5470 -885
rect 5610 -915 5790 -885
rect 5930 -915 6110 -885
rect 6250 -915 6430 -885
rect 6570 -915 6750 -885
rect 6890 -915 7070 -885
rect 7210 -915 7390 -885
rect 7530 -915 7710 -885
rect 7850 -915 8030 -885
rect 8170 -915 8350 -885
rect 8490 -915 8670 -885
rect 8810 -915 8990 -885
rect 9130 -915 9310 -885
rect 9450 -915 9630 -885
rect 9770 -915 9950 -885
rect 10090 -915 10270 -885
rect 10 -1795 190 -1765
rect 330 -1795 510 -1765
rect 650 -1795 830 -1765
rect 970 -1795 1150 -1765
rect 1290 -1795 1470 -1765
rect 1610 -1795 1790 -1765
rect 1930 -1795 2110 -1765
rect 2250 -1795 2430 -1765
rect 2570 -1795 2750 -1765
rect 2890 -1795 3070 -1765
rect 3210 -1795 3390 -1765
rect 3530 -1795 3710 -1765
rect 3850 -1795 4030 -1765
rect 4170 -1795 4350 -1765
rect 4490 -1795 4670 -1765
rect 4810 -1795 4990 -1765
rect 5290 -1795 5470 -1765
rect 5610 -1795 5790 -1765
rect 5930 -1795 6110 -1765
rect 6250 -1795 6430 -1765
rect 6570 -1795 6750 -1765
rect 6890 -1795 7070 -1765
rect 7210 -1795 7390 -1765
rect 7530 -1795 7710 -1765
rect 7850 -1795 8030 -1765
rect 8170 -1795 8350 -1765
rect 8490 -1795 8670 -1765
rect 8810 -1795 8990 -1765
rect 9130 -1795 9310 -1765
rect 9450 -1795 9630 -1765
rect 9770 -1795 9950 -1765
rect 10090 -1795 10270 -1765
rect 10 -2275 190 -2245
rect 330 -2275 510 -2245
rect 650 -2275 830 -2245
rect 970 -2275 1150 -2245
rect 1290 -2275 1470 -2245
rect 1610 -2275 1790 -2245
rect 1930 -2275 2110 -2245
rect 2250 -2275 2430 -2245
rect 2570 -2275 2750 -2245
rect 2890 -2275 3070 -2245
rect 3210 -2275 3390 -2245
rect 3530 -2275 3710 -2245
rect 3850 -2275 4030 -2245
rect 4170 -2275 4350 -2245
rect 4490 -2275 4670 -2245
rect 4810 -2275 4990 -2245
rect 5290 -2275 5470 -2245
rect 5610 -2275 5790 -2245
rect 5930 -2275 6110 -2245
rect 6250 -2275 6430 -2245
rect 6570 -2275 6750 -2245
rect 6890 -2275 7070 -2245
rect 7210 -2275 7390 -2245
rect 7530 -2275 7710 -2245
rect 7850 -2275 8030 -2245
rect 8170 -2275 8350 -2245
rect 8490 -2275 8670 -2245
rect 8810 -2275 8990 -2245
rect 9130 -2275 9310 -2245
rect 9450 -2275 9630 -2245
rect 9770 -2275 9950 -2245
rect 10090 -2275 10270 -2245
rect 10 -2835 190 -2805
rect 330 -2835 510 -2805
rect 650 -2835 830 -2805
rect 970 -2835 1150 -2805
rect 1290 -2835 1470 -2805
rect 1610 -2835 1790 -2805
rect 1930 -2835 2110 -2805
rect 2250 -2835 2430 -2805
rect 2570 -2835 2750 -2805
rect 2890 -2835 3070 -2805
rect 3210 -2835 3390 -2805
rect 3530 -2835 3710 -2805
rect 3850 -2835 4030 -2805
rect 4170 -2835 4350 -2805
rect 4490 -2835 4670 -2805
rect 4810 -2835 4990 -2805
rect 5290 -2835 5470 -2805
rect 5610 -2835 5790 -2805
rect 5930 -2835 6110 -2805
rect 6250 -2835 6430 -2805
rect 6570 -2835 6750 -2805
rect 6890 -2835 7070 -2805
rect 7210 -2835 7390 -2805
rect 7530 -2835 7710 -2805
rect 7850 -2835 8030 -2805
rect 8170 -2835 8350 -2805
rect 8490 -2835 8670 -2805
rect 8810 -2835 8990 -2805
rect 9130 -2835 9310 -2805
rect 9450 -2835 9630 -2805
rect 9770 -2835 9950 -2805
rect 10090 -2835 10270 -2805
rect 10 -3315 190 -3285
rect 330 -3315 510 -3285
rect 650 -3315 830 -3285
rect 970 -3315 1150 -3285
rect 1290 -3315 1470 -3285
rect 1610 -3315 1790 -3285
rect 1930 -3315 2110 -3285
rect 2250 -3315 2430 -3285
rect 2570 -3315 2750 -3285
rect 2890 -3315 3070 -3285
rect 3210 -3315 3390 -3285
rect 3530 -3315 3710 -3285
rect 3850 -3315 4030 -3285
rect 4170 -3315 4350 -3285
rect 4490 -3315 4670 -3285
rect 4810 -3315 4990 -3285
rect 5290 -3315 5470 -3285
rect 5610 -3315 5790 -3285
rect 5930 -3315 6110 -3285
rect 6250 -3315 6430 -3285
rect 6570 -3315 6750 -3285
rect 6890 -3315 7070 -3285
rect 7210 -3315 7390 -3285
rect 7530 -3315 7710 -3285
rect 7850 -3315 8030 -3285
rect 8170 -3315 8350 -3285
rect 8490 -3315 8670 -3285
rect 8810 -3315 8990 -3285
rect 9130 -3315 9310 -3285
rect 9450 -3315 9630 -3285
rect 9770 -3315 9950 -3285
rect 10090 -3315 10270 -3285
<< locali >>
rect -320 1000 -40 1040
rect 240 1000 280 1040
rect 560 1000 600 1040
rect 880 1000 920 1040
rect 1200 1000 1240 1040
rect 1520 1000 1560 1040
rect 1840 1000 1880 1040
rect 2160 1000 2200 1040
rect 2480 1000 2520 1040
rect 2800 1000 2840 1040
rect 3120 1000 3160 1040
rect 3440 1000 3480 1040
rect 3760 1000 3800 1040
rect 4080 1000 4120 1040
rect 4400 1000 4440 1040
rect 4720 1000 4760 1040
rect 5040 1000 5240 1040
rect 5520 1000 5560 1040
rect 5840 1000 5880 1040
rect 6160 1000 6200 1040
rect 6480 1000 6520 1040
rect 6800 1000 6840 1040
rect 7120 1000 7160 1040
rect 7440 1000 7480 1040
rect 7760 1000 7800 1040
rect 8080 1000 8120 1040
rect 8400 1000 8440 1040
rect 8720 1000 8760 1040
rect 9040 1000 9080 1040
rect 9360 1000 9400 1040
rect 9680 1000 9720 1040
rect 10000 1000 10040 1040
rect 10320 1000 10600 1040
rect -320 960 -280 1000
rect 10560 960 10600 1000
rect -160 840 -40 880
rect 240 840 280 880
rect 560 840 600 880
rect 880 840 920 880
rect 1200 840 1240 880
rect 1520 840 1560 880
rect 1840 840 1880 880
rect 2160 840 2200 880
rect 2480 840 2520 880
rect 2800 840 2840 880
rect 3120 840 3160 880
rect 3440 840 3480 880
rect 3760 840 3800 880
rect 4080 840 4120 880
rect 4400 840 4440 880
rect 4720 840 4760 880
rect 5040 840 5240 880
rect 5520 840 5560 880
rect -160 800 -120 840
rect -160 560 -120 600
rect -80 750 -40 840
rect 5120 800 5160 840
rect -80 670 -75 750
rect -45 670 -40 750
rect -80 560 -40 670
rect 240 750 280 760
rect 240 670 245 750
rect 275 670 280 750
rect 240 660 280 670
rect 560 750 600 760
rect 560 670 565 750
rect 595 670 600 750
rect 560 660 600 670
rect 880 750 920 760
rect 880 670 885 750
rect 915 670 920 750
rect 880 660 920 670
rect 1200 750 1240 760
rect 1200 670 1205 750
rect 1235 670 1240 750
rect 1200 660 1240 670
rect 1520 750 1560 760
rect 1520 670 1525 750
rect 1555 670 1560 750
rect 1520 660 1560 670
rect 1840 750 1880 760
rect 1840 670 1845 750
rect 1875 670 1880 750
rect 1840 660 1880 670
rect 2160 750 2200 760
rect 2160 670 2165 750
rect 2195 670 2200 750
rect 2160 660 2200 670
rect 2480 750 2520 760
rect 2480 670 2485 750
rect 2515 670 2520 750
rect 2480 660 2520 670
rect 2800 750 2840 760
rect 2800 670 2805 750
rect 2835 670 2840 750
rect 2800 660 2840 670
rect 3120 750 3160 760
rect 3120 670 3125 750
rect 3155 670 3160 750
rect 3120 660 3160 670
rect 3440 750 3480 760
rect 3440 670 3445 750
rect 3475 670 3480 750
rect 3440 660 3480 670
rect 3760 750 3800 760
rect 3760 670 3765 750
rect 3795 670 3800 750
rect 3760 660 3800 670
rect 4080 750 4120 760
rect 4080 670 4085 750
rect 4115 670 4120 750
rect 4080 660 4120 670
rect 4400 750 4440 760
rect 4400 670 4405 750
rect 4435 670 4440 750
rect 4400 660 4440 670
rect 4720 750 4760 760
rect 4720 670 4725 750
rect 4755 670 4760 750
rect 4720 660 4760 670
rect 5040 750 5080 760
rect 5040 670 5045 750
rect 5075 670 5080 750
rect 5040 660 5080 670
rect 0 635 200 640
rect 0 605 10 635
rect 190 605 200 635
rect 0 600 200 605
rect 320 635 520 640
rect 320 605 330 635
rect 510 605 520 635
rect 320 600 520 605
rect 640 635 840 640
rect 640 605 650 635
rect 830 605 840 635
rect 640 600 840 605
rect 960 635 1160 640
rect 960 605 970 635
rect 1150 605 1160 635
rect 960 600 1160 605
rect 1280 635 1480 640
rect 1280 605 1290 635
rect 1470 605 1480 635
rect 1280 600 1480 605
rect 1600 635 1800 640
rect 1600 605 1610 635
rect 1790 605 1800 635
rect 1600 600 1800 605
rect 1920 635 2120 640
rect 1920 605 1930 635
rect 2110 605 2120 635
rect 1920 600 2120 605
rect 2240 635 2440 640
rect 2240 605 2250 635
rect 2430 605 2440 635
rect 2240 600 2440 605
rect 2560 635 2760 640
rect 2560 605 2570 635
rect 2750 605 2760 635
rect 2560 600 2760 605
rect 2880 635 3080 640
rect 2880 605 2890 635
rect 3070 605 3080 635
rect 2880 600 3080 605
rect 3200 635 3400 640
rect 3200 605 3210 635
rect 3390 605 3400 635
rect 3200 600 3400 605
rect 3520 635 3720 640
rect 3520 605 3530 635
rect 3710 605 3720 635
rect 3520 600 3720 605
rect 3840 635 4040 640
rect 3840 605 3850 635
rect 4030 605 4040 635
rect 3840 600 4040 605
rect 4160 635 4360 640
rect 4160 605 4170 635
rect 4350 605 4360 635
rect 4160 600 4360 605
rect 4480 635 4680 640
rect 4480 605 4490 635
rect 4670 605 4680 635
rect 4480 600 4680 605
rect 4800 635 5000 640
rect 4800 605 4810 635
rect 4990 605 5000 635
rect 4800 600 5000 605
rect 5120 560 5160 600
rect 5200 750 5240 840
rect 5200 670 5205 750
rect 5235 670 5240 750
rect 5200 560 5240 670
rect 5520 750 5560 760
rect 5520 670 5525 750
rect 5555 670 5560 750
rect 5520 660 5560 670
rect 5840 750 5880 880
rect 6160 840 6200 880
rect 5840 670 5845 750
rect 5875 670 5880 750
rect 5280 635 5480 640
rect 5280 605 5290 635
rect 5470 605 5480 635
rect 5280 600 5480 605
rect 5600 635 5800 640
rect 5600 605 5610 635
rect 5790 605 5800 635
rect 5600 600 5800 605
rect -160 520 -40 560
rect 240 520 280 560
rect 560 520 600 560
rect 880 520 920 560
rect 1200 520 1240 560
rect 1520 520 1560 560
rect 1840 520 1880 560
rect 2160 520 2200 560
rect 2480 520 2520 560
rect 2800 520 2840 560
rect 3120 520 3160 560
rect 3440 520 3480 560
rect 3760 520 3800 560
rect 4080 520 4120 560
rect 4400 520 4440 560
rect 4720 520 4760 560
rect 5040 520 5240 560
rect 5520 520 5560 560
rect 5840 520 5880 670
rect 6160 750 6200 760
rect 6160 670 6165 750
rect 6195 670 6200 750
rect 6160 660 6200 670
rect 6480 750 6520 880
rect 6800 840 6840 880
rect 6480 670 6485 750
rect 6515 670 6520 750
rect 5920 635 6120 640
rect 5920 605 5930 635
rect 6110 605 6120 635
rect 5920 600 6120 605
rect 6240 635 6440 640
rect 6240 605 6250 635
rect 6430 605 6440 635
rect 6240 600 6440 605
rect 6160 520 6200 560
rect 6480 520 6520 670
rect 6800 750 6840 760
rect 6800 670 6805 750
rect 6835 670 6840 750
rect 6800 660 6840 670
rect 7120 750 7160 880
rect 7440 840 7480 880
rect 7120 670 7125 750
rect 7155 670 7160 750
rect 6560 635 6760 640
rect 6560 605 6570 635
rect 6750 605 6760 635
rect 6560 600 6760 605
rect 6880 635 7080 640
rect 6880 605 6890 635
rect 7070 605 7080 635
rect 6880 600 7080 605
rect 6800 520 6840 560
rect 7120 520 7160 670
rect 7440 750 7480 760
rect 7440 670 7445 750
rect 7475 670 7480 750
rect 7440 660 7480 670
rect 7760 750 7800 880
rect 8080 840 8120 880
rect 7760 670 7765 750
rect 7795 670 7800 750
rect 7200 635 7400 640
rect 7200 605 7210 635
rect 7390 605 7400 635
rect 7200 600 7400 605
rect 7520 635 7720 640
rect 7520 605 7530 635
rect 7710 605 7720 635
rect 7520 600 7720 605
rect 7440 520 7480 560
rect 7760 520 7800 670
rect 8080 750 8120 760
rect 8080 670 8085 750
rect 8115 670 8120 750
rect 8080 660 8120 670
rect 8400 750 8440 880
rect 8720 840 8760 880
rect 8400 670 8405 750
rect 8435 670 8440 750
rect 7840 635 8040 640
rect 7840 605 7850 635
rect 8030 605 8040 635
rect 7840 600 8040 605
rect 8160 635 8360 640
rect 8160 605 8170 635
rect 8350 605 8360 635
rect 8160 600 8360 605
rect 8080 520 8120 560
rect 8400 520 8440 670
rect 8720 750 8760 760
rect 8720 670 8725 750
rect 8755 670 8760 750
rect 8720 660 8760 670
rect 9040 750 9080 880
rect 9360 840 9400 880
rect 9040 670 9045 750
rect 9075 670 9080 750
rect 8480 635 8680 640
rect 8480 605 8490 635
rect 8670 605 8680 635
rect 8480 600 8680 605
rect 8800 635 9000 640
rect 8800 605 8810 635
rect 8990 605 9000 635
rect 8800 600 9000 605
rect 8720 520 8760 560
rect 9040 520 9080 670
rect 9360 750 9400 760
rect 9360 670 9365 750
rect 9395 670 9400 750
rect 9360 660 9400 670
rect 9680 750 9720 880
rect 10000 840 10040 880
rect 10320 840 10480 880
rect 9680 670 9685 750
rect 9715 670 9720 750
rect 9120 635 9320 640
rect 9120 605 9130 635
rect 9310 605 9320 635
rect 9120 600 9320 605
rect 9440 635 9640 640
rect 9440 605 9450 635
rect 9630 605 9640 635
rect 9440 600 9640 605
rect 9360 520 9400 560
rect 9680 520 9720 670
rect 10000 750 10040 760
rect 10000 670 10005 750
rect 10035 670 10040 750
rect 10000 660 10040 670
rect 10320 750 10360 840
rect 10320 670 10325 750
rect 10355 670 10360 750
rect 9760 635 9960 640
rect 9760 605 9770 635
rect 9950 605 9960 635
rect 9760 600 9960 605
rect 10080 635 10280 640
rect 10080 605 10090 635
rect 10270 605 10280 635
rect 10080 600 10280 605
rect 10320 560 10360 670
rect 10400 800 10440 840
rect 10400 560 10440 600
rect 10000 520 10040 560
rect 10320 520 10480 560
rect -280 360 -40 400
rect 240 360 280 400
rect 560 360 600 400
rect 880 360 920 400
rect 1200 360 1240 400
rect 1520 360 1560 400
rect 1840 360 1880 400
rect 2160 360 2200 400
rect 2480 360 2520 400
rect 2800 360 2840 400
rect 3120 360 3160 400
rect 3440 360 3480 400
rect 3760 360 3800 400
rect 4080 360 4120 400
rect 4400 360 4440 400
rect 4720 360 4760 400
rect 5040 360 5240 400
rect 5520 360 5560 400
rect 5840 360 5880 400
rect 6160 360 6200 400
rect 6480 360 6520 400
rect 6800 360 6840 400
rect 7120 360 7160 400
rect 7440 360 7480 400
rect 7760 360 7800 400
rect 8080 360 8120 400
rect 8400 360 8440 400
rect 8720 360 8760 400
rect 9040 360 9080 400
rect 9360 360 9400 400
rect 9680 360 9720 400
rect 10000 360 10040 400
rect 10320 360 10560 400
rect -320 -80 -280 -40
rect -160 200 -40 240
rect 240 200 280 240
rect 560 200 600 240
rect 880 200 920 240
rect 1200 200 1240 240
rect 1520 200 1560 240
rect 1840 200 1880 240
rect 2160 200 2200 240
rect -160 160 -120 200
rect -160 -80 -120 -40
rect -80 90 -40 200
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 120 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 120 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 120 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 120 1160 125
rect 1280 155 1480 160
rect 1280 125 1290 155
rect 1470 125 1480 155
rect 1280 120 1480 125
rect 1600 155 1800 160
rect 1600 125 1610 155
rect 1790 125 1800 155
rect 1600 120 1800 125
rect 1920 155 2120 160
rect 1920 125 1930 155
rect 2110 125 2120 155
rect 1920 120 2120 125
rect 2240 155 2440 160
rect 2240 125 2250 155
rect 2430 125 2440 155
rect 2240 120 2440 125
rect -80 10 -75 90
rect -45 10 -40 90
rect -80 -80 -40 10
rect 240 90 280 100
rect 240 10 245 90
rect 275 10 280 90
rect 240 0 280 10
rect 560 90 600 100
rect 560 10 565 90
rect 595 10 600 90
rect 560 0 600 10
rect 880 90 920 100
rect 880 10 885 90
rect 915 10 920 90
rect 880 0 920 10
rect 1200 90 1240 100
rect 1200 10 1205 90
rect 1235 10 1240 90
rect 1200 0 1240 10
rect 1520 90 1560 100
rect 1520 10 1525 90
rect 1555 10 1560 90
rect 1520 0 1560 10
rect 1840 90 1880 100
rect 1840 10 1845 90
rect 1875 10 1880 90
rect 1840 0 1880 10
rect 2160 90 2200 100
rect 2160 10 2165 90
rect 2195 10 2200 90
rect 2160 0 2200 10
rect 2480 90 2520 240
rect 2800 200 2840 240
rect 3120 200 3160 240
rect 3440 200 3480 240
rect 3760 200 3800 240
rect 4080 200 4120 240
rect 4400 200 4440 240
rect 4720 200 4760 240
rect 5040 200 5240 240
rect 5520 200 5560 240
rect 5840 200 5880 240
rect 6160 200 6200 240
rect 6480 200 6520 240
rect 6800 200 6840 240
rect 7120 200 7160 240
rect 7440 200 7480 240
rect 2560 155 2760 160
rect 2560 125 2570 155
rect 2750 125 2760 155
rect 2560 120 2760 125
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 120 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 120 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 120 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 120 4040 125
rect 4160 155 4360 160
rect 4160 125 4170 155
rect 4350 125 4360 155
rect 4160 120 4360 125
rect 4480 155 4680 160
rect 4480 125 4490 155
rect 4670 125 4680 155
rect 4480 120 4680 125
rect 4800 155 5000 160
rect 4800 125 4810 155
rect 4990 125 5000 155
rect 4800 120 5000 125
rect 2480 10 2485 90
rect 2515 10 2520 90
rect -320 -120 -40 -80
rect 240 -120 280 -80
rect 560 -120 600 -80
rect 880 -120 920 -80
rect 1200 -120 1240 -80
rect 1520 -120 1560 -80
rect 1840 -120 1880 -80
rect 2160 -120 2200 -80
rect 2480 -120 2520 10
rect 2800 90 2840 100
rect 2800 10 2805 90
rect 2835 10 2840 90
rect 2800 0 2840 10
rect 3120 90 3160 100
rect 3120 10 3125 90
rect 3155 10 3160 90
rect 3120 0 3160 10
rect 3440 90 3480 100
rect 3440 10 3445 90
rect 3475 10 3480 90
rect 3440 0 3480 10
rect 3760 90 3800 100
rect 3760 10 3765 90
rect 3795 10 3800 90
rect 3760 0 3800 10
rect 4080 90 4120 100
rect 4080 10 4085 90
rect 4115 10 4120 90
rect 4080 0 4120 10
rect 4400 90 4440 100
rect 4400 10 4405 90
rect 4435 10 4440 90
rect 4400 0 4440 10
rect 4720 90 4760 100
rect 4720 10 4725 90
rect 4755 10 4760 90
rect 4720 0 4760 10
rect 5040 90 5080 200
rect 5040 10 5045 90
rect 5075 10 5080 90
rect 5040 -80 5080 10
rect 5120 160 5160 200
rect 5120 -80 5160 -40
rect 5200 90 5240 200
rect 5280 155 5480 160
rect 5280 125 5290 155
rect 5470 125 5480 155
rect 5280 120 5480 125
rect 5600 155 5800 160
rect 5600 125 5610 155
rect 5790 125 5800 155
rect 5600 120 5800 125
rect 5920 155 6120 160
rect 5920 125 5930 155
rect 6110 125 6120 155
rect 5920 120 6120 125
rect 6240 155 6440 160
rect 6240 125 6250 155
rect 6430 125 6440 155
rect 6240 120 6440 125
rect 6560 155 6760 160
rect 6560 125 6570 155
rect 6750 125 6760 155
rect 6560 120 6760 125
rect 6880 155 7080 160
rect 6880 125 6890 155
rect 7070 125 7080 155
rect 6880 120 7080 125
rect 7200 155 7400 160
rect 7200 125 7210 155
rect 7390 125 7400 155
rect 7200 120 7400 125
rect 7520 155 7720 160
rect 7520 125 7530 155
rect 7710 125 7720 155
rect 7520 120 7720 125
rect 5200 10 5205 90
rect 5235 10 5240 90
rect 5200 -80 5240 10
rect 5520 90 5560 100
rect 5520 10 5525 90
rect 5555 10 5560 90
rect 5520 0 5560 10
rect 5840 90 5880 100
rect 5840 10 5845 90
rect 5875 10 5880 90
rect 5840 0 5880 10
rect 6160 90 6200 100
rect 6160 10 6165 90
rect 6195 10 6200 90
rect 6160 0 6200 10
rect 6480 90 6520 100
rect 6480 10 6485 90
rect 6515 10 6520 90
rect 6480 0 6520 10
rect 6800 90 6840 100
rect 6800 10 6805 90
rect 6835 10 6840 90
rect 6800 0 6840 10
rect 7120 90 7160 100
rect 7120 10 7125 90
rect 7155 10 7160 90
rect 7120 0 7160 10
rect 7440 90 7480 100
rect 7440 10 7445 90
rect 7475 10 7480 90
rect 7440 0 7480 10
rect 7760 90 7800 240
rect 8080 200 8120 240
rect 8400 200 8440 240
rect 8720 200 8760 240
rect 9040 200 9080 240
rect 9360 200 9400 240
rect 9680 200 9720 240
rect 10000 200 10040 240
rect 10320 200 10480 240
rect 7840 155 8040 160
rect 7840 125 7850 155
rect 8030 125 8040 155
rect 7840 120 8040 125
rect 8160 155 8360 160
rect 8160 125 8170 155
rect 8350 125 8360 155
rect 8160 120 8360 125
rect 8480 155 8680 160
rect 8480 125 8490 155
rect 8670 125 8680 155
rect 8480 120 8680 125
rect 8800 155 9000 160
rect 8800 125 8810 155
rect 8990 125 9000 155
rect 8800 120 9000 125
rect 9120 155 9320 160
rect 9120 125 9130 155
rect 9310 125 9320 155
rect 9120 120 9320 125
rect 9440 155 9640 160
rect 9440 125 9450 155
rect 9630 125 9640 155
rect 9440 120 9640 125
rect 9760 155 9960 160
rect 9760 125 9770 155
rect 9950 125 9960 155
rect 9760 120 9960 125
rect 10080 155 10280 160
rect 10080 125 10090 155
rect 10270 125 10280 155
rect 10080 120 10280 125
rect 7760 10 7765 90
rect 7795 10 7800 90
rect 2800 -120 2840 -80
rect 3120 -120 3160 -80
rect 3440 -120 3480 -80
rect 3760 -120 3800 -80
rect 4080 -120 4120 -80
rect 4400 -120 4440 -80
rect 4720 -120 4760 -80
rect 5040 -120 5240 -80
rect 5520 -120 5560 -80
rect 5840 -120 5880 -80
rect 6160 -120 6200 -80
rect 6480 -120 6520 -80
rect 6800 -120 6840 -80
rect 7120 -120 7160 -80
rect 7440 -120 7480 -80
rect 7760 -120 7800 10
rect 8080 90 8120 100
rect 8080 10 8085 90
rect 8115 10 8120 90
rect 8080 0 8120 10
rect 8400 90 8440 100
rect 8400 10 8405 90
rect 8435 10 8440 90
rect 8400 0 8440 10
rect 8720 90 8760 100
rect 8720 10 8725 90
rect 8755 10 8760 90
rect 8720 0 8760 10
rect 9040 90 9080 100
rect 9040 10 9045 90
rect 9075 10 9080 90
rect 9040 0 9080 10
rect 9360 90 9400 100
rect 9360 10 9365 90
rect 9395 10 9400 90
rect 9360 0 9400 10
rect 9680 90 9720 100
rect 9680 10 9685 90
rect 9715 10 9720 90
rect 9680 0 9720 10
rect 10000 90 10040 100
rect 10000 10 10005 90
rect 10035 10 10040 90
rect 10000 0 10040 10
rect 10320 90 10360 200
rect 10320 10 10325 90
rect 10355 10 10360 90
rect 10320 -80 10360 10
rect 10400 160 10440 200
rect 10400 -80 10440 -40
rect 10560 -80 10600 -40
rect 8080 -120 8120 -80
rect 8400 -120 8440 -80
rect 8720 -120 8760 -80
rect 9040 -120 9080 -80
rect 9360 -120 9400 -80
rect 9680 -120 9720 -80
rect 10000 -120 10040 -80
rect 10320 -120 10600 -80
rect -320 -200 -40 -160
rect 240 -200 280 -160
rect 560 -200 600 -160
rect 880 -200 920 -160
rect 1200 -200 1240 -160
rect 1520 -200 1560 -160
rect 1840 -200 1880 -160
rect 2160 -200 2200 -160
rect -320 -240 -280 -200
rect -160 -240 -120 -200
rect -160 -480 -120 -440
rect -80 -290 -40 -200
rect -80 -370 -75 -290
rect -45 -370 -40 -290
rect -80 -480 -40 -370
rect 240 -290 280 -280
rect 240 -370 245 -290
rect 275 -370 280 -290
rect 240 -380 280 -370
rect 560 -290 600 -280
rect 560 -370 565 -290
rect 595 -370 600 -290
rect 560 -380 600 -370
rect 880 -290 920 -280
rect 880 -370 885 -290
rect 915 -370 920 -290
rect 880 -380 920 -370
rect 1200 -290 1240 -280
rect 1200 -370 1205 -290
rect 1235 -370 1240 -290
rect 1200 -380 1240 -370
rect 1520 -290 1560 -280
rect 1520 -370 1525 -290
rect 1555 -370 1560 -290
rect 1520 -380 1560 -370
rect 1840 -290 1880 -280
rect 1840 -370 1845 -290
rect 1875 -370 1880 -290
rect 1840 -380 1880 -370
rect 2160 -290 2200 -280
rect 2160 -370 2165 -290
rect 2195 -370 2200 -290
rect 2160 -380 2200 -370
rect 2480 -290 2520 -160
rect 2800 -200 2840 -160
rect 3120 -200 3160 -160
rect 3440 -200 3480 -160
rect 3760 -200 3800 -160
rect 4080 -200 4120 -160
rect 4400 -200 4440 -160
rect 4720 -200 4760 -160
rect 5040 -200 5240 -160
rect 5520 -200 5560 -160
rect 5840 -200 5880 -160
rect 6160 -200 6200 -160
rect 6480 -200 6520 -160
rect 6800 -200 6840 -160
rect 7120 -200 7160 -160
rect 7440 -200 7480 -160
rect 2480 -370 2485 -290
rect 2515 -370 2520 -290
rect 0 -405 200 -400
rect 0 -435 10 -405
rect 190 -435 200 -405
rect 0 -440 200 -435
rect 320 -405 520 -400
rect 320 -435 330 -405
rect 510 -435 520 -405
rect 320 -440 520 -435
rect 640 -405 840 -400
rect 640 -435 650 -405
rect 830 -435 840 -405
rect 640 -440 840 -435
rect 960 -405 1160 -400
rect 960 -435 970 -405
rect 1150 -435 1160 -405
rect 960 -440 1160 -435
rect 1280 -405 1480 -400
rect 1280 -435 1290 -405
rect 1470 -435 1480 -405
rect 1280 -440 1480 -435
rect 1600 -405 1800 -400
rect 1600 -435 1610 -405
rect 1790 -435 1800 -405
rect 1600 -440 1800 -435
rect 1920 -405 2120 -400
rect 1920 -435 1930 -405
rect 2110 -435 2120 -405
rect 1920 -440 2120 -435
rect 2240 -405 2440 -400
rect 2240 -435 2250 -405
rect 2430 -435 2440 -405
rect 2240 -440 2440 -435
rect -200 -520 -40 -480
rect 240 -520 280 -480
rect 560 -520 600 -480
rect 880 -520 920 -480
rect 1200 -520 1240 -480
rect 1520 -520 1560 -480
rect 1840 -520 1880 -480
rect 2160 -520 2200 -480
rect 2480 -520 2520 -370
rect 2800 -290 2840 -280
rect 2800 -370 2805 -290
rect 2835 -370 2840 -290
rect 2800 -380 2840 -370
rect 3120 -290 3160 -280
rect 3120 -370 3125 -290
rect 3155 -370 3160 -290
rect 3120 -380 3160 -370
rect 3440 -290 3480 -280
rect 3440 -370 3445 -290
rect 3475 -370 3480 -290
rect 3440 -380 3480 -370
rect 3760 -290 3800 -280
rect 3760 -370 3765 -290
rect 3795 -370 3800 -290
rect 3760 -380 3800 -370
rect 4080 -290 4120 -280
rect 4080 -370 4085 -290
rect 4115 -370 4120 -290
rect 4080 -380 4120 -370
rect 4400 -290 4440 -280
rect 4400 -370 4405 -290
rect 4435 -370 4440 -290
rect 4400 -380 4440 -370
rect 4720 -290 4760 -280
rect 4720 -370 4725 -290
rect 4755 -370 4760 -290
rect 4720 -380 4760 -370
rect 5040 -290 5080 -200
rect 5040 -370 5045 -290
rect 5075 -370 5080 -290
rect 2560 -405 2760 -400
rect 2560 -435 2570 -405
rect 2750 -435 2760 -405
rect 2560 -440 2760 -435
rect 2880 -405 3080 -400
rect 2880 -435 2890 -405
rect 3070 -435 3080 -405
rect 2880 -440 3080 -435
rect 3200 -405 3400 -400
rect 3200 -435 3210 -405
rect 3390 -435 3400 -405
rect 3200 -440 3400 -435
rect 3520 -405 3720 -400
rect 3520 -435 3530 -405
rect 3710 -435 3720 -405
rect 3520 -440 3720 -435
rect 3840 -405 4040 -400
rect 3840 -435 3850 -405
rect 4030 -435 4040 -405
rect 3840 -440 4040 -435
rect 4160 -405 4360 -400
rect 4160 -435 4170 -405
rect 4350 -435 4360 -405
rect 4160 -440 4360 -435
rect 4480 -405 4680 -400
rect 4480 -435 4490 -405
rect 4670 -435 4680 -405
rect 4480 -440 4680 -435
rect 4800 -405 5000 -400
rect 4800 -435 4810 -405
rect 4990 -435 5000 -405
rect 4800 -440 5000 -435
rect 5040 -480 5080 -370
rect 5120 -240 5160 -200
rect 5120 -480 5160 -440
rect 5200 -290 5240 -200
rect 5200 -370 5205 -290
rect 5235 -370 5240 -290
rect 5200 -480 5240 -370
rect 5520 -290 5560 -280
rect 5520 -370 5525 -290
rect 5555 -370 5560 -290
rect 5520 -380 5560 -370
rect 5840 -290 5880 -280
rect 5840 -370 5845 -290
rect 5875 -370 5880 -290
rect 5840 -380 5880 -370
rect 6160 -290 6200 -280
rect 6160 -370 6165 -290
rect 6195 -370 6200 -290
rect 6160 -380 6200 -370
rect 6480 -290 6520 -280
rect 6480 -370 6485 -290
rect 6515 -370 6520 -290
rect 6480 -380 6520 -370
rect 6800 -290 6840 -280
rect 6800 -370 6805 -290
rect 6835 -370 6840 -290
rect 6800 -380 6840 -370
rect 7120 -290 7160 -280
rect 7120 -370 7125 -290
rect 7155 -370 7160 -290
rect 7120 -380 7160 -370
rect 7440 -290 7480 -280
rect 7440 -370 7445 -290
rect 7475 -370 7480 -290
rect 7440 -380 7480 -370
rect 7760 -290 7800 -160
rect 8080 -200 8120 -160
rect 8400 -200 8440 -160
rect 8720 -200 8760 -160
rect 9040 -200 9080 -160
rect 9360 -200 9400 -160
rect 9680 -200 9720 -160
rect 10000 -200 10040 -160
rect 10320 -200 10600 -160
rect 7760 -370 7765 -290
rect 7795 -370 7800 -290
rect 5280 -405 5480 -400
rect 5280 -435 5290 -405
rect 5470 -435 5480 -405
rect 5280 -440 5480 -435
rect 5600 -405 5800 -400
rect 5600 -435 5610 -405
rect 5790 -435 5800 -405
rect 5600 -440 5800 -435
rect 5920 -405 6120 -400
rect 5920 -435 5930 -405
rect 6110 -435 6120 -405
rect 5920 -440 6120 -435
rect 6240 -405 6440 -400
rect 6240 -435 6250 -405
rect 6430 -435 6440 -405
rect 6240 -440 6440 -435
rect 6560 -405 6760 -400
rect 6560 -435 6570 -405
rect 6750 -435 6760 -405
rect 6560 -440 6760 -435
rect 6880 -405 7080 -400
rect 6880 -435 6890 -405
rect 7070 -435 7080 -405
rect 6880 -440 7080 -435
rect 7200 -405 7400 -400
rect 7200 -435 7210 -405
rect 7390 -435 7400 -405
rect 7200 -440 7400 -435
rect 7520 -405 7720 -400
rect 7520 -435 7530 -405
rect 7710 -435 7720 -405
rect 7520 -440 7720 -435
rect 2800 -520 2840 -480
rect 3120 -520 3160 -480
rect 3440 -520 3480 -480
rect 3760 -520 3800 -480
rect 4080 -520 4120 -480
rect 4400 -520 4440 -480
rect 4720 -520 4760 -480
rect 5040 -520 5240 -480
rect 5520 -520 5560 -480
rect 5840 -520 5880 -480
rect 6160 -520 6200 -480
rect 6480 -520 6520 -480
rect 6800 -520 6840 -480
rect 7120 -520 7160 -480
rect 7440 -520 7480 -480
rect 7760 -520 7800 -370
rect 8080 -290 8120 -280
rect 8080 -370 8085 -290
rect 8115 -370 8120 -290
rect 8080 -380 8120 -370
rect 8400 -290 8440 -280
rect 8400 -370 8405 -290
rect 8435 -370 8440 -290
rect 8400 -380 8440 -370
rect 8720 -290 8760 -280
rect 8720 -370 8725 -290
rect 8755 -370 8760 -290
rect 8720 -380 8760 -370
rect 9040 -290 9080 -280
rect 9040 -370 9045 -290
rect 9075 -370 9080 -290
rect 9040 -380 9080 -370
rect 9360 -290 9400 -280
rect 9360 -370 9365 -290
rect 9395 -370 9400 -290
rect 9360 -380 9400 -370
rect 9680 -290 9720 -280
rect 9680 -370 9685 -290
rect 9715 -370 9720 -290
rect 9680 -380 9720 -370
rect 10000 -290 10040 -280
rect 10000 -370 10005 -290
rect 10035 -370 10040 -290
rect 10000 -380 10040 -370
rect 10320 -290 10360 -200
rect 10320 -370 10325 -290
rect 10355 -370 10360 -290
rect 7840 -405 8040 -400
rect 7840 -435 7850 -405
rect 8030 -435 8040 -405
rect 7840 -440 8040 -435
rect 8160 -405 8360 -400
rect 8160 -435 8170 -405
rect 8350 -435 8360 -405
rect 8160 -440 8360 -435
rect 8480 -405 8680 -400
rect 8480 -435 8490 -405
rect 8670 -435 8680 -405
rect 8480 -440 8680 -435
rect 8800 -405 9000 -400
rect 8800 -435 8810 -405
rect 8990 -435 9000 -405
rect 8800 -440 9000 -435
rect 9120 -405 9320 -400
rect 9120 -435 9130 -405
rect 9310 -435 9320 -405
rect 9120 -440 9320 -435
rect 9440 -405 9640 -400
rect 9440 -435 9450 -405
rect 9630 -435 9640 -405
rect 9440 -440 9640 -435
rect 9760 -405 9960 -400
rect 9760 -435 9770 -405
rect 9950 -435 9960 -405
rect 9760 -440 9960 -435
rect 10080 -405 10280 -400
rect 10080 -435 10090 -405
rect 10270 -435 10280 -405
rect 10080 -440 10280 -435
rect 10320 -480 10360 -370
rect 10400 -240 10440 -200
rect 10400 -480 10440 -440
rect 8080 -520 8120 -480
rect 8400 -520 8440 -480
rect 8720 -520 8760 -480
rect 9040 -520 9080 -480
rect 9360 -520 9400 -480
rect 9680 -520 9720 -480
rect 10000 -520 10040 -480
rect 10320 -520 10440 -480
rect 10560 -240 10600 -200
rect -280 -680 -40 -640
rect 240 -680 280 -640
rect 560 -680 600 -640
rect 880 -680 920 -640
rect 1200 -680 1240 -640
rect 1520 -680 1560 -640
rect 1840 -680 1880 -640
rect 2160 -680 2200 -640
rect 2480 -680 2520 -640
rect 2800 -680 2840 -640
rect 3120 -680 3160 -640
rect 3440 -680 3480 -640
rect 3760 -680 3800 -640
rect 4080 -680 4120 -640
rect 4400 -680 4440 -640
rect 4720 -680 4760 -640
rect 5040 -680 5240 -640
rect 5520 -680 5560 -640
rect 5840 -680 5880 -640
rect 6160 -680 6200 -640
rect 6480 -680 6520 -640
rect 6800 -680 6840 -640
rect 7120 -680 7160 -640
rect 7440 -680 7480 -640
rect 7760 -680 7800 -640
rect 8080 -680 8120 -640
rect 8400 -680 8440 -640
rect 8720 -680 8760 -640
rect 9040 -680 9080 -640
rect 9360 -680 9400 -640
rect 9680 -680 9720 -640
rect 10000 -680 10040 -640
rect 10320 -680 10560 -640
rect -200 -840 -40 -800
rect 240 -840 280 -800
rect -160 -880 -120 -840
rect -160 -1120 -120 -1080
rect -80 -950 -40 -840
rect 0 -885 200 -880
rect 0 -915 10 -885
rect 190 -915 200 -885
rect 0 -920 200 -915
rect 320 -885 520 -880
rect 320 -915 330 -885
rect 510 -915 520 -885
rect 320 -920 520 -915
rect -80 -1030 -75 -950
rect -45 -1030 -40 -950
rect -80 -1120 -40 -1030
rect 240 -950 280 -940
rect 240 -1030 245 -950
rect 275 -1030 280 -950
rect 240 -1040 280 -1030
rect 560 -950 600 -800
rect 880 -840 920 -800
rect 640 -885 840 -880
rect 640 -915 650 -885
rect 830 -915 840 -885
rect 640 -920 840 -915
rect 960 -885 1160 -880
rect 960 -915 970 -885
rect 1150 -915 1160 -885
rect 960 -920 1160 -915
rect 560 -1030 565 -950
rect 595 -1030 600 -950
rect -200 -1160 -40 -1120
rect 240 -1160 280 -1120
rect 560 -1160 600 -1030
rect 880 -950 920 -940
rect 880 -1030 885 -950
rect 915 -1030 920 -950
rect 880 -1040 920 -1030
rect 1200 -950 1240 -800
rect 1520 -840 1560 -800
rect 1280 -885 1480 -880
rect 1280 -915 1290 -885
rect 1470 -915 1480 -885
rect 1280 -920 1480 -915
rect 1600 -885 1800 -880
rect 1600 -915 1610 -885
rect 1790 -915 1800 -885
rect 1600 -920 1800 -915
rect 1200 -1030 1205 -950
rect 1235 -1030 1240 -950
rect 880 -1160 920 -1120
rect 1200 -1160 1240 -1030
rect 1520 -950 1560 -940
rect 1520 -1030 1525 -950
rect 1555 -1030 1560 -950
rect 1520 -1040 1560 -1030
rect 1840 -950 1880 -800
rect 2160 -840 2200 -800
rect 1920 -885 2120 -880
rect 1920 -915 1930 -885
rect 2110 -915 2120 -885
rect 1920 -920 2120 -915
rect 2240 -885 2440 -880
rect 2240 -915 2250 -885
rect 2430 -915 2440 -885
rect 2240 -920 2440 -915
rect 1840 -1030 1845 -950
rect 1875 -1030 1880 -950
rect 1520 -1160 1560 -1120
rect 1840 -1160 1880 -1030
rect 2160 -950 2200 -940
rect 2160 -1030 2165 -950
rect 2195 -1030 2200 -950
rect 2160 -1040 2200 -1030
rect 2480 -950 2520 -800
rect 2800 -840 2840 -800
rect 2560 -885 2760 -880
rect 2560 -915 2570 -885
rect 2750 -915 2760 -885
rect 2560 -920 2760 -915
rect 2880 -885 3080 -880
rect 2880 -915 2890 -885
rect 3070 -915 3080 -885
rect 2880 -920 3080 -915
rect 2480 -1030 2485 -950
rect 2515 -1030 2520 -950
rect 2160 -1160 2200 -1120
rect 2480 -1160 2520 -1030
rect 2800 -950 2840 -940
rect 2800 -1030 2805 -950
rect 2835 -1030 2840 -950
rect 2800 -1040 2840 -1030
rect 3120 -950 3160 -800
rect 3440 -840 3480 -800
rect 3200 -885 3400 -880
rect 3200 -915 3210 -885
rect 3390 -915 3400 -885
rect 3200 -920 3400 -915
rect 3520 -885 3720 -880
rect 3520 -915 3530 -885
rect 3710 -915 3720 -885
rect 3520 -920 3720 -915
rect 3120 -1030 3125 -950
rect 3155 -1030 3160 -950
rect 2800 -1160 2840 -1120
rect 3120 -1160 3160 -1030
rect 3440 -950 3480 -940
rect 3440 -1030 3445 -950
rect 3475 -1030 3480 -950
rect 3440 -1040 3480 -1030
rect 3760 -950 3800 -800
rect 4080 -840 4120 -800
rect 3840 -885 4040 -880
rect 3840 -915 3850 -885
rect 4030 -915 4040 -885
rect 3840 -920 4040 -915
rect 4160 -885 4360 -880
rect 4160 -915 4170 -885
rect 4350 -915 4360 -885
rect 4160 -920 4360 -915
rect 3760 -1030 3765 -950
rect 3795 -1030 3800 -950
rect 3440 -1160 3480 -1120
rect 3760 -1160 3800 -1030
rect 4080 -950 4120 -940
rect 4080 -1030 4085 -950
rect 4115 -1030 4120 -950
rect 4080 -1040 4120 -1030
rect 4400 -950 4440 -800
rect 4720 -840 4760 -800
rect 5040 -840 5240 -800
rect 5520 -840 5560 -800
rect 5840 -840 5880 -800
rect 6160 -840 6200 -800
rect 6480 -840 6520 -800
rect 6800 -840 6840 -800
rect 7120 -840 7160 -800
rect 7440 -840 7480 -800
rect 7760 -840 7800 -800
rect 8080 -840 8120 -800
rect 8400 -840 8440 -800
rect 8720 -840 8760 -800
rect 9040 -840 9080 -800
rect 9360 -840 9400 -800
rect 9680 -840 9720 -800
rect 10000 -840 10040 -800
rect 10320 -840 10440 -800
rect 4480 -885 4680 -880
rect 4480 -915 4490 -885
rect 4670 -915 4680 -885
rect 4480 -920 4680 -915
rect 4800 -885 5000 -880
rect 4800 -915 4810 -885
rect 4990 -915 5000 -885
rect 4800 -920 5000 -915
rect 4400 -1030 4405 -950
rect 4435 -1030 4440 -950
rect 4080 -1160 4120 -1120
rect 4400 -1160 4440 -1030
rect 4720 -950 4760 -940
rect 4720 -1030 4725 -950
rect 4755 -1030 4760 -950
rect 4720 -1040 4760 -1030
rect 5040 -950 5080 -840
rect 5040 -1030 5045 -950
rect 5075 -1030 5080 -950
rect 5040 -1120 5080 -1030
rect 5120 -880 5160 -840
rect 5280 -885 5480 -880
rect 5280 -915 5290 -885
rect 5470 -915 5480 -885
rect 5280 -920 5480 -915
rect 5600 -885 5800 -880
rect 5600 -915 5610 -885
rect 5790 -915 5800 -885
rect 5600 -920 5800 -915
rect 5920 -885 6120 -880
rect 5920 -915 5930 -885
rect 6110 -915 6120 -885
rect 5920 -920 6120 -915
rect 6240 -885 6440 -880
rect 6240 -915 6250 -885
rect 6430 -915 6440 -885
rect 6240 -920 6440 -915
rect 6560 -885 6760 -880
rect 6560 -915 6570 -885
rect 6750 -915 6760 -885
rect 6560 -920 6760 -915
rect 6880 -885 7080 -880
rect 6880 -915 6890 -885
rect 7070 -915 7080 -885
rect 6880 -920 7080 -915
rect 7200 -885 7400 -880
rect 7200 -915 7210 -885
rect 7390 -915 7400 -885
rect 7200 -920 7400 -915
rect 7520 -885 7720 -880
rect 7520 -915 7530 -885
rect 7710 -915 7720 -885
rect 7520 -920 7720 -915
rect 7840 -885 8040 -880
rect 7840 -915 7850 -885
rect 8030 -915 8040 -885
rect 7840 -920 8040 -915
rect 8160 -885 8360 -880
rect 8160 -915 8170 -885
rect 8350 -915 8360 -885
rect 8160 -920 8360 -915
rect 8480 -885 8680 -880
rect 8480 -915 8490 -885
rect 8670 -915 8680 -885
rect 8480 -920 8680 -915
rect 8800 -885 9000 -880
rect 8800 -915 8810 -885
rect 8990 -915 9000 -885
rect 8800 -920 9000 -915
rect 9120 -885 9320 -880
rect 9120 -915 9130 -885
rect 9310 -915 9320 -885
rect 9120 -920 9320 -915
rect 9440 -885 9640 -880
rect 9440 -915 9450 -885
rect 9630 -915 9640 -885
rect 9440 -920 9640 -915
rect 9760 -885 9960 -880
rect 9760 -915 9770 -885
rect 9950 -915 9960 -885
rect 9760 -920 9960 -915
rect 10080 -885 10280 -880
rect 10080 -915 10090 -885
rect 10270 -915 10280 -885
rect 10080 -920 10280 -915
rect 5200 -950 5240 -940
rect 5200 -1030 5205 -950
rect 5235 -1030 5240 -950
rect 5200 -1040 5240 -1030
rect 5520 -950 5560 -940
rect 5520 -1030 5525 -950
rect 5555 -1030 5560 -950
rect 5520 -1040 5560 -1030
rect 5840 -950 5880 -940
rect 5840 -1030 5845 -950
rect 5875 -1030 5880 -950
rect 5840 -1040 5880 -1030
rect 6160 -950 6200 -940
rect 6160 -1030 6165 -950
rect 6195 -1030 6200 -950
rect 6160 -1040 6200 -1030
rect 6480 -950 6520 -940
rect 6480 -1030 6485 -950
rect 6515 -1030 6520 -950
rect 6480 -1040 6520 -1030
rect 6800 -950 6840 -940
rect 6800 -1030 6805 -950
rect 6835 -1030 6840 -950
rect 6800 -1040 6840 -1030
rect 7120 -950 7160 -940
rect 7120 -1030 7125 -950
rect 7155 -1030 7160 -950
rect 7120 -1040 7160 -1030
rect 7440 -950 7480 -940
rect 7440 -1030 7445 -950
rect 7475 -1030 7480 -950
rect 7440 -1040 7480 -1030
rect 7760 -950 7800 -940
rect 7760 -1030 7765 -950
rect 7795 -1030 7800 -950
rect 7760 -1040 7800 -1030
rect 8080 -950 8120 -940
rect 8080 -1030 8085 -950
rect 8115 -1030 8120 -950
rect 8080 -1040 8120 -1030
rect 8400 -950 8440 -940
rect 8400 -1030 8405 -950
rect 8435 -1030 8440 -950
rect 8400 -1040 8440 -1030
rect 8720 -950 8760 -940
rect 8720 -1030 8725 -950
rect 8755 -1030 8760 -950
rect 8720 -1040 8760 -1030
rect 9040 -950 9080 -940
rect 9040 -1030 9045 -950
rect 9075 -1030 9080 -950
rect 9040 -1040 9080 -1030
rect 9360 -950 9400 -940
rect 9360 -1030 9365 -950
rect 9395 -1030 9400 -950
rect 9360 -1040 9400 -1030
rect 9680 -950 9720 -940
rect 9680 -1030 9685 -950
rect 9715 -1030 9720 -950
rect 9680 -1040 9720 -1030
rect 10000 -950 10040 -940
rect 10000 -1030 10005 -950
rect 10035 -1030 10040 -950
rect 10000 -1040 10040 -1030
rect 10320 -950 10360 -840
rect 10320 -1030 10325 -950
rect 10355 -1030 10360 -950
rect 5120 -1120 5160 -1080
rect 10320 -1120 10360 -1030
rect 10400 -880 10440 -840
rect 10400 -1120 10440 -1080
rect 4720 -1160 4760 -1120
rect 5040 -1160 5240 -1120
rect 5520 -1160 5560 -1120
rect 5840 -1160 5880 -1120
rect 6160 -1160 6200 -1120
rect 6480 -1160 6520 -1120
rect 6800 -1160 6840 -1120
rect 7120 -1160 7160 -1120
rect 7440 -1160 7480 -1120
rect 7760 -1160 7800 -1120
rect 8080 -1160 8120 -1120
rect 8400 -1160 8440 -1120
rect 8720 -1160 8760 -1120
rect 9040 -1160 9080 -1120
rect 9360 -1160 9400 -1120
rect 9680 -1160 9720 -1120
rect 10000 -1160 10040 -1120
rect 10320 -1160 10440 -1120
rect -320 -1280 -280 -1240
rect 10560 -1280 10600 -1240
rect -320 -1320 -40 -1280
rect 240 -1320 280 -1280
rect 560 -1320 600 -1280
rect 880 -1320 920 -1280
rect 1200 -1320 1240 -1280
rect 1520 -1320 1560 -1280
rect 1840 -1320 1880 -1280
rect 2160 -1320 2200 -1280
rect 2480 -1320 2520 -1280
rect 2800 -1320 2840 -1280
rect 3120 -1320 3160 -1280
rect 3440 -1320 3480 -1280
rect 3760 -1320 3800 -1280
rect 4080 -1320 4120 -1280
rect 4400 -1320 4440 -1280
rect 4720 -1320 4760 -1280
rect 5040 -1320 5240 -1280
rect 5520 -1320 5560 -1280
rect 5840 -1320 5880 -1280
rect 6160 -1320 6200 -1280
rect 6480 -1320 6520 -1280
rect 6800 -1320 6840 -1280
rect 7120 -1320 7160 -1280
rect 7440 -1320 7480 -1280
rect 7760 -1320 7800 -1280
rect 8080 -1320 8120 -1280
rect 8400 -1320 8440 -1280
rect 8720 -1320 8760 -1280
rect 9040 -1320 9080 -1280
rect 9360 -1320 9400 -1280
rect 9680 -1320 9720 -1280
rect 10000 -1320 10040 -1280
rect 10320 -1320 10600 -1280
rect -320 -1400 -40 -1360
rect 240 -1400 280 -1360
rect 560 -1400 600 -1360
rect 880 -1400 920 -1360
rect 1200 -1400 1240 -1360
rect 1520 -1400 1560 -1360
rect 1840 -1400 1880 -1360
rect 2160 -1400 2200 -1360
rect 2480 -1400 2520 -1360
rect 2800 -1400 2840 -1360
rect 3120 -1400 3160 -1360
rect 3440 -1400 3480 -1360
rect 3760 -1400 3800 -1360
rect 4080 -1400 4120 -1360
rect 4400 -1400 4440 -1360
rect 4720 -1400 4760 -1360
rect 5040 -1400 5240 -1360
rect 5520 -1400 5560 -1360
rect 5840 -1400 5880 -1360
rect 6160 -1400 6200 -1360
rect 6480 -1400 6520 -1360
rect 6800 -1400 6840 -1360
rect 7120 -1400 7160 -1360
rect 7440 -1400 7480 -1360
rect 7760 -1400 7800 -1360
rect 8080 -1400 8120 -1360
rect 8400 -1400 8440 -1360
rect 8720 -1400 8760 -1360
rect 9040 -1400 9080 -1360
rect 9360 -1400 9400 -1360
rect 9680 -1400 9720 -1360
rect 10000 -1400 10040 -1360
rect 10320 -1400 10600 -1360
rect -320 -1440 -280 -1400
rect 10560 -1440 10600 -1400
rect -200 -1560 -40 -1520
rect 240 -1560 280 -1520
rect -160 -1600 -120 -1560
rect -160 -1840 -120 -1800
rect -80 -1650 -40 -1560
rect -80 -1730 -75 -1650
rect -45 -1730 -40 -1650
rect -80 -1840 -40 -1730
rect 240 -1650 280 -1640
rect 240 -1730 245 -1650
rect 275 -1730 280 -1650
rect 240 -1740 280 -1730
rect 560 -1650 600 -1520
rect 880 -1560 920 -1520
rect 560 -1730 565 -1650
rect 595 -1730 600 -1650
rect 0 -1765 200 -1760
rect 0 -1795 10 -1765
rect 190 -1795 200 -1765
rect 0 -1800 200 -1795
rect 320 -1765 520 -1760
rect 320 -1795 330 -1765
rect 510 -1795 520 -1765
rect 320 -1800 520 -1795
rect -200 -1880 -40 -1840
rect 240 -1880 280 -1840
rect 560 -1880 600 -1730
rect 880 -1650 920 -1640
rect 880 -1730 885 -1650
rect 915 -1730 920 -1650
rect 880 -1740 920 -1730
rect 1200 -1650 1240 -1520
rect 1520 -1560 1560 -1520
rect 1200 -1730 1205 -1650
rect 1235 -1730 1240 -1650
rect 640 -1765 840 -1760
rect 640 -1795 650 -1765
rect 830 -1795 840 -1765
rect 640 -1800 840 -1795
rect 960 -1765 1160 -1760
rect 960 -1795 970 -1765
rect 1150 -1795 1160 -1765
rect 960 -1800 1160 -1795
rect 880 -1880 920 -1840
rect 1200 -1880 1240 -1730
rect 1520 -1650 1560 -1640
rect 1520 -1730 1525 -1650
rect 1555 -1730 1560 -1650
rect 1520 -1740 1560 -1730
rect 1840 -1650 1880 -1520
rect 2160 -1560 2200 -1520
rect 1840 -1730 1845 -1650
rect 1875 -1730 1880 -1650
rect 1280 -1765 1480 -1760
rect 1280 -1795 1290 -1765
rect 1470 -1795 1480 -1765
rect 1280 -1800 1480 -1795
rect 1600 -1765 1800 -1760
rect 1600 -1795 1610 -1765
rect 1790 -1795 1800 -1765
rect 1600 -1800 1800 -1795
rect 1520 -1880 1560 -1840
rect 1840 -1880 1880 -1730
rect 2160 -1650 2200 -1640
rect 2160 -1730 2165 -1650
rect 2195 -1730 2200 -1650
rect 2160 -1740 2200 -1730
rect 2480 -1650 2520 -1520
rect 2800 -1560 2840 -1520
rect 2480 -1730 2485 -1650
rect 2515 -1730 2520 -1650
rect 1920 -1765 2120 -1760
rect 1920 -1795 1930 -1765
rect 2110 -1795 2120 -1765
rect 1920 -1800 2120 -1795
rect 2240 -1765 2440 -1760
rect 2240 -1795 2250 -1765
rect 2430 -1795 2440 -1765
rect 2240 -1800 2440 -1795
rect 2160 -1880 2200 -1840
rect 2480 -1880 2520 -1730
rect 2800 -1650 2840 -1640
rect 2800 -1730 2805 -1650
rect 2835 -1730 2840 -1650
rect 2800 -1740 2840 -1730
rect 3120 -1650 3160 -1520
rect 3440 -1560 3480 -1520
rect 3120 -1730 3125 -1650
rect 3155 -1730 3160 -1650
rect 2560 -1765 2760 -1760
rect 2560 -1795 2570 -1765
rect 2750 -1795 2760 -1765
rect 2560 -1800 2760 -1795
rect 2880 -1765 3080 -1760
rect 2880 -1795 2890 -1765
rect 3070 -1795 3080 -1765
rect 2880 -1800 3080 -1795
rect 2800 -1880 2840 -1840
rect 3120 -1880 3160 -1730
rect 3440 -1650 3480 -1640
rect 3440 -1730 3445 -1650
rect 3475 -1730 3480 -1650
rect 3440 -1740 3480 -1730
rect 3760 -1650 3800 -1520
rect 4080 -1560 4120 -1520
rect 3760 -1730 3765 -1650
rect 3795 -1730 3800 -1650
rect 3200 -1765 3400 -1760
rect 3200 -1795 3210 -1765
rect 3390 -1795 3400 -1765
rect 3200 -1800 3400 -1795
rect 3520 -1765 3720 -1760
rect 3520 -1795 3530 -1765
rect 3710 -1795 3720 -1765
rect 3520 -1800 3720 -1795
rect 3440 -1880 3480 -1840
rect 3760 -1880 3800 -1730
rect 4080 -1650 4120 -1640
rect 4080 -1730 4085 -1650
rect 4115 -1730 4120 -1650
rect 4080 -1740 4120 -1730
rect 4400 -1650 4440 -1520
rect 4720 -1560 4760 -1520
rect 5040 -1560 5240 -1520
rect 5520 -1560 5560 -1520
rect 5840 -1560 5880 -1520
rect 6160 -1560 6200 -1520
rect 6480 -1560 6520 -1520
rect 6800 -1560 6840 -1520
rect 7120 -1560 7160 -1520
rect 7440 -1560 7480 -1520
rect 7760 -1560 7800 -1520
rect 8080 -1560 8120 -1520
rect 8400 -1560 8440 -1520
rect 8720 -1560 8760 -1520
rect 9040 -1560 9080 -1520
rect 9360 -1560 9400 -1520
rect 9680 -1560 9720 -1520
rect 10000 -1560 10040 -1520
rect 10320 -1560 10440 -1520
rect 4400 -1730 4405 -1650
rect 4435 -1730 4440 -1650
rect 3840 -1765 4040 -1760
rect 3840 -1795 3850 -1765
rect 4030 -1795 4040 -1765
rect 3840 -1800 4040 -1795
rect 4160 -1765 4360 -1760
rect 4160 -1795 4170 -1765
rect 4350 -1795 4360 -1765
rect 4160 -1800 4360 -1795
rect 4080 -1880 4120 -1840
rect 4400 -1880 4440 -1730
rect 4720 -1650 4760 -1640
rect 4720 -1730 4725 -1650
rect 4755 -1730 4760 -1650
rect 4720 -1740 4760 -1730
rect 5040 -1650 5080 -1560
rect 5040 -1730 5045 -1650
rect 5075 -1730 5080 -1650
rect 4480 -1765 4680 -1760
rect 4480 -1795 4490 -1765
rect 4670 -1795 4680 -1765
rect 4480 -1800 4680 -1795
rect 4800 -1765 5000 -1760
rect 4800 -1795 4810 -1765
rect 4990 -1795 5000 -1765
rect 4800 -1800 5000 -1795
rect 5040 -1840 5080 -1730
rect 5120 -1600 5160 -1560
rect 5200 -1650 5240 -1640
rect 5200 -1730 5205 -1650
rect 5235 -1730 5240 -1650
rect 5200 -1740 5240 -1730
rect 5520 -1650 5560 -1640
rect 5520 -1730 5525 -1650
rect 5555 -1730 5560 -1650
rect 5520 -1740 5560 -1730
rect 5840 -1650 5880 -1640
rect 5840 -1730 5845 -1650
rect 5875 -1730 5880 -1650
rect 5840 -1740 5880 -1730
rect 6160 -1650 6200 -1640
rect 6160 -1730 6165 -1650
rect 6195 -1730 6200 -1650
rect 6160 -1740 6200 -1730
rect 6480 -1650 6520 -1640
rect 6480 -1730 6485 -1650
rect 6515 -1730 6520 -1650
rect 6480 -1740 6520 -1730
rect 6800 -1650 6840 -1640
rect 6800 -1730 6805 -1650
rect 6835 -1730 6840 -1650
rect 6800 -1740 6840 -1730
rect 7120 -1650 7160 -1640
rect 7120 -1730 7125 -1650
rect 7155 -1730 7160 -1650
rect 7120 -1740 7160 -1730
rect 7440 -1650 7480 -1640
rect 7440 -1730 7445 -1650
rect 7475 -1730 7480 -1650
rect 7440 -1740 7480 -1730
rect 7760 -1650 7800 -1640
rect 7760 -1730 7765 -1650
rect 7795 -1730 7800 -1650
rect 7760 -1740 7800 -1730
rect 8080 -1650 8120 -1640
rect 8080 -1730 8085 -1650
rect 8115 -1730 8120 -1650
rect 8080 -1740 8120 -1730
rect 8400 -1650 8440 -1640
rect 8400 -1730 8405 -1650
rect 8435 -1730 8440 -1650
rect 8400 -1740 8440 -1730
rect 8720 -1650 8760 -1640
rect 8720 -1730 8725 -1650
rect 8755 -1730 8760 -1650
rect 8720 -1740 8760 -1730
rect 9040 -1650 9080 -1640
rect 9040 -1730 9045 -1650
rect 9075 -1730 9080 -1650
rect 9040 -1740 9080 -1730
rect 9360 -1650 9400 -1640
rect 9360 -1730 9365 -1650
rect 9395 -1730 9400 -1650
rect 9360 -1740 9400 -1730
rect 9680 -1650 9720 -1640
rect 9680 -1730 9685 -1650
rect 9715 -1730 9720 -1650
rect 9680 -1740 9720 -1730
rect 10000 -1650 10040 -1640
rect 10000 -1730 10005 -1650
rect 10035 -1730 10040 -1650
rect 10000 -1740 10040 -1730
rect 10320 -1650 10360 -1560
rect 10320 -1730 10325 -1650
rect 10355 -1730 10360 -1650
rect 5280 -1765 5480 -1760
rect 5280 -1795 5290 -1765
rect 5470 -1795 5480 -1765
rect 5280 -1800 5480 -1795
rect 5600 -1765 5800 -1760
rect 5600 -1795 5610 -1765
rect 5790 -1795 5800 -1765
rect 5600 -1800 5800 -1795
rect 5920 -1765 6120 -1760
rect 5920 -1795 5930 -1765
rect 6110 -1795 6120 -1765
rect 5920 -1800 6120 -1795
rect 6240 -1765 6440 -1760
rect 6240 -1795 6250 -1765
rect 6430 -1795 6440 -1765
rect 6240 -1800 6440 -1795
rect 6560 -1765 6760 -1760
rect 6560 -1795 6570 -1765
rect 6750 -1795 6760 -1765
rect 6560 -1800 6760 -1795
rect 6880 -1765 7080 -1760
rect 6880 -1795 6890 -1765
rect 7070 -1795 7080 -1765
rect 6880 -1800 7080 -1795
rect 7200 -1765 7400 -1760
rect 7200 -1795 7210 -1765
rect 7390 -1795 7400 -1765
rect 7200 -1800 7400 -1795
rect 7520 -1765 7720 -1760
rect 7520 -1795 7530 -1765
rect 7710 -1795 7720 -1765
rect 7520 -1800 7720 -1795
rect 7840 -1765 8040 -1760
rect 7840 -1795 7850 -1765
rect 8030 -1795 8040 -1765
rect 7840 -1800 8040 -1795
rect 8160 -1765 8360 -1760
rect 8160 -1795 8170 -1765
rect 8350 -1795 8360 -1765
rect 8160 -1800 8360 -1795
rect 8480 -1765 8680 -1760
rect 8480 -1795 8490 -1765
rect 8670 -1795 8680 -1765
rect 8480 -1800 8680 -1795
rect 8800 -1765 9000 -1760
rect 8800 -1795 8810 -1765
rect 8990 -1795 9000 -1765
rect 8800 -1800 9000 -1795
rect 9120 -1765 9320 -1760
rect 9120 -1795 9130 -1765
rect 9310 -1795 9320 -1765
rect 9120 -1800 9320 -1795
rect 9440 -1765 9640 -1760
rect 9440 -1795 9450 -1765
rect 9630 -1795 9640 -1765
rect 9440 -1800 9640 -1795
rect 9760 -1765 9960 -1760
rect 9760 -1795 9770 -1765
rect 9950 -1795 9960 -1765
rect 9760 -1800 9960 -1795
rect 10080 -1765 10280 -1760
rect 10080 -1795 10090 -1765
rect 10270 -1795 10280 -1765
rect 10080 -1800 10280 -1795
rect 5120 -1840 5160 -1800
rect 10320 -1840 10360 -1730
rect 10400 -1600 10440 -1560
rect 10400 -1840 10440 -1800
rect 4720 -1880 4760 -1840
rect 5040 -1880 5240 -1840
rect 5520 -1880 5560 -1840
rect 5840 -1880 5880 -1840
rect 6160 -1880 6200 -1840
rect 6480 -1880 6520 -1840
rect 6800 -1880 6840 -1840
rect 7120 -1880 7160 -1840
rect 7440 -1880 7480 -1840
rect 7760 -1880 7800 -1840
rect 8080 -1880 8120 -1840
rect 8400 -1880 8440 -1840
rect 8720 -1880 8760 -1840
rect 9040 -1880 9080 -1840
rect 9360 -1880 9400 -1840
rect 9680 -1880 9720 -1840
rect 10000 -1880 10040 -1840
rect 10320 -1880 10440 -1840
rect -280 -2040 -40 -2000
rect 240 -2040 280 -2000
rect 560 -2040 600 -2000
rect 880 -2040 920 -2000
rect 1200 -2040 1240 -2000
rect 1520 -2040 1560 -2000
rect 1840 -2040 1880 -2000
rect 2160 -2040 2200 -2000
rect 2480 -2040 2520 -2000
rect 2800 -2040 2840 -2000
rect 3120 -2040 3160 -2000
rect 3440 -2040 3480 -2000
rect 3760 -2040 3800 -2000
rect 4080 -2040 4120 -2000
rect 4400 -2040 4440 -2000
rect 4720 -2040 4760 -2000
rect 5040 -2040 5240 -2000
rect 5520 -2040 5560 -2000
rect 5840 -2040 5880 -2000
rect 6160 -2040 6200 -2000
rect 6480 -2040 6520 -2000
rect 6800 -2040 6840 -2000
rect 7120 -2040 7160 -2000
rect 7440 -2040 7480 -2000
rect 7760 -2040 7800 -2000
rect 8080 -2040 8120 -2000
rect 8400 -2040 8440 -2000
rect 8720 -2040 8760 -2000
rect 9040 -2040 9080 -2000
rect 9360 -2040 9400 -2000
rect 9680 -2040 9720 -2000
rect 10000 -2040 10040 -2000
rect 10320 -2040 10560 -2000
rect -200 -2200 -40 -2160
rect 240 -2200 280 -2160
rect 560 -2200 600 -2160
rect 880 -2200 920 -2160
rect 1200 -2200 1240 -2160
rect 1520 -2200 1560 -2160
rect 1840 -2200 1880 -2160
rect 2160 -2200 2200 -2160
rect -320 -2480 -280 -2440
rect -160 -2240 -120 -2200
rect -160 -2480 -120 -2440
rect -80 -2310 -40 -2200
rect 0 -2245 200 -2240
rect 0 -2275 10 -2245
rect 190 -2275 200 -2245
rect 0 -2280 200 -2275
rect 320 -2245 520 -2240
rect 320 -2275 330 -2245
rect 510 -2275 520 -2245
rect 320 -2280 520 -2275
rect 640 -2245 840 -2240
rect 640 -2275 650 -2245
rect 830 -2275 840 -2245
rect 640 -2280 840 -2275
rect 960 -2245 1160 -2240
rect 960 -2275 970 -2245
rect 1150 -2275 1160 -2245
rect 960 -2280 1160 -2275
rect 1280 -2245 1480 -2240
rect 1280 -2275 1290 -2245
rect 1470 -2275 1480 -2245
rect 1280 -2280 1480 -2275
rect 1600 -2245 1800 -2240
rect 1600 -2275 1610 -2245
rect 1790 -2275 1800 -2245
rect 1600 -2280 1800 -2275
rect 1920 -2245 2120 -2240
rect 1920 -2275 1930 -2245
rect 2110 -2275 2120 -2245
rect 1920 -2280 2120 -2275
rect 2240 -2245 2440 -2240
rect 2240 -2275 2250 -2245
rect 2430 -2275 2440 -2245
rect 2240 -2280 2440 -2275
rect -80 -2390 -75 -2310
rect -45 -2390 -40 -2310
rect -80 -2480 -40 -2390
rect 240 -2310 280 -2300
rect 240 -2390 245 -2310
rect 275 -2390 280 -2310
rect 240 -2400 280 -2390
rect 560 -2310 600 -2300
rect 560 -2390 565 -2310
rect 595 -2390 600 -2310
rect 560 -2400 600 -2390
rect 880 -2310 920 -2300
rect 880 -2390 885 -2310
rect 915 -2390 920 -2310
rect 880 -2400 920 -2390
rect 1200 -2310 1240 -2300
rect 1200 -2390 1205 -2310
rect 1235 -2390 1240 -2310
rect 1200 -2400 1240 -2390
rect 1520 -2310 1560 -2300
rect 1520 -2390 1525 -2310
rect 1555 -2390 1560 -2310
rect 1520 -2400 1560 -2390
rect 1840 -2310 1880 -2300
rect 1840 -2390 1845 -2310
rect 1875 -2390 1880 -2310
rect 1840 -2400 1880 -2390
rect 2160 -2310 2200 -2300
rect 2160 -2390 2165 -2310
rect 2195 -2390 2200 -2310
rect 2160 -2400 2200 -2390
rect 2480 -2310 2520 -2160
rect 2800 -2200 2840 -2160
rect 3120 -2200 3160 -2160
rect 3440 -2200 3480 -2160
rect 3760 -2200 3800 -2160
rect 4080 -2200 4120 -2160
rect 4400 -2200 4440 -2160
rect 4720 -2200 4760 -2160
rect 5040 -2200 5240 -2160
rect 5520 -2200 5560 -2160
rect 5840 -2200 5880 -2160
rect 6160 -2200 6200 -2160
rect 6480 -2200 6520 -2160
rect 6800 -2200 6840 -2160
rect 7120 -2200 7160 -2160
rect 7440 -2200 7480 -2160
rect 2560 -2245 2760 -2240
rect 2560 -2275 2570 -2245
rect 2750 -2275 2760 -2245
rect 2560 -2280 2760 -2275
rect 2880 -2245 3080 -2240
rect 2880 -2275 2890 -2245
rect 3070 -2275 3080 -2245
rect 2880 -2280 3080 -2275
rect 3200 -2245 3400 -2240
rect 3200 -2275 3210 -2245
rect 3390 -2275 3400 -2245
rect 3200 -2280 3400 -2275
rect 3520 -2245 3720 -2240
rect 3520 -2275 3530 -2245
rect 3710 -2275 3720 -2245
rect 3520 -2280 3720 -2275
rect 3840 -2245 4040 -2240
rect 3840 -2275 3850 -2245
rect 4030 -2275 4040 -2245
rect 3840 -2280 4040 -2275
rect 4160 -2245 4360 -2240
rect 4160 -2275 4170 -2245
rect 4350 -2275 4360 -2245
rect 4160 -2280 4360 -2275
rect 4480 -2245 4680 -2240
rect 4480 -2275 4490 -2245
rect 4670 -2275 4680 -2245
rect 4480 -2280 4680 -2275
rect 4800 -2245 5000 -2240
rect 4800 -2275 4810 -2245
rect 4990 -2275 5000 -2245
rect 4800 -2280 5000 -2275
rect 2480 -2390 2485 -2310
rect 2515 -2390 2520 -2310
rect -320 -2520 -40 -2480
rect 240 -2520 280 -2480
rect 560 -2520 600 -2480
rect 880 -2520 920 -2480
rect 1200 -2520 1240 -2480
rect 1520 -2520 1560 -2480
rect 1840 -2520 1880 -2480
rect 2160 -2520 2200 -2480
rect 2480 -2520 2520 -2390
rect 2800 -2310 2840 -2300
rect 2800 -2390 2805 -2310
rect 2835 -2390 2840 -2310
rect 2800 -2400 2840 -2390
rect 3120 -2310 3160 -2300
rect 3120 -2390 3125 -2310
rect 3155 -2390 3160 -2310
rect 3120 -2400 3160 -2390
rect 3440 -2310 3480 -2300
rect 3440 -2390 3445 -2310
rect 3475 -2390 3480 -2310
rect 3440 -2400 3480 -2390
rect 3760 -2310 3800 -2300
rect 3760 -2390 3765 -2310
rect 3795 -2390 3800 -2310
rect 3760 -2400 3800 -2390
rect 4080 -2310 4120 -2300
rect 4080 -2390 4085 -2310
rect 4115 -2390 4120 -2310
rect 4080 -2400 4120 -2390
rect 4400 -2310 4440 -2300
rect 4400 -2390 4405 -2310
rect 4435 -2390 4440 -2310
rect 4400 -2400 4440 -2390
rect 4720 -2310 4760 -2300
rect 4720 -2390 4725 -2310
rect 4755 -2390 4760 -2310
rect 4720 -2400 4760 -2390
rect 5040 -2310 5080 -2200
rect 5040 -2390 5045 -2310
rect 5075 -2390 5080 -2310
rect 5040 -2480 5080 -2390
rect 5120 -2240 5160 -2200
rect 5120 -2480 5160 -2440
rect 5200 -2310 5240 -2200
rect 5280 -2245 5480 -2240
rect 5280 -2275 5290 -2245
rect 5470 -2275 5480 -2245
rect 5280 -2280 5480 -2275
rect 5600 -2245 5800 -2240
rect 5600 -2275 5610 -2245
rect 5790 -2275 5800 -2245
rect 5600 -2280 5800 -2275
rect 5920 -2245 6120 -2240
rect 5920 -2275 5930 -2245
rect 6110 -2275 6120 -2245
rect 5920 -2280 6120 -2275
rect 6240 -2245 6440 -2240
rect 6240 -2275 6250 -2245
rect 6430 -2275 6440 -2245
rect 6240 -2280 6440 -2275
rect 6560 -2245 6760 -2240
rect 6560 -2275 6570 -2245
rect 6750 -2275 6760 -2245
rect 6560 -2280 6760 -2275
rect 6880 -2245 7080 -2240
rect 6880 -2275 6890 -2245
rect 7070 -2275 7080 -2245
rect 6880 -2280 7080 -2275
rect 7200 -2245 7400 -2240
rect 7200 -2275 7210 -2245
rect 7390 -2275 7400 -2245
rect 7200 -2280 7400 -2275
rect 7520 -2245 7720 -2240
rect 7520 -2275 7530 -2245
rect 7710 -2275 7720 -2245
rect 7520 -2280 7720 -2275
rect 5200 -2390 5205 -2310
rect 5235 -2390 5240 -2310
rect 5200 -2480 5240 -2390
rect 5520 -2310 5560 -2300
rect 5520 -2390 5525 -2310
rect 5555 -2390 5560 -2310
rect 5520 -2400 5560 -2390
rect 5840 -2310 5880 -2300
rect 5840 -2390 5845 -2310
rect 5875 -2390 5880 -2310
rect 5840 -2400 5880 -2390
rect 6160 -2310 6200 -2300
rect 6160 -2390 6165 -2310
rect 6195 -2390 6200 -2310
rect 6160 -2400 6200 -2390
rect 6480 -2310 6520 -2300
rect 6480 -2390 6485 -2310
rect 6515 -2390 6520 -2310
rect 6480 -2400 6520 -2390
rect 6800 -2310 6840 -2300
rect 6800 -2390 6805 -2310
rect 6835 -2390 6840 -2310
rect 6800 -2400 6840 -2390
rect 7120 -2310 7160 -2300
rect 7120 -2390 7125 -2310
rect 7155 -2390 7160 -2310
rect 7120 -2400 7160 -2390
rect 7440 -2310 7480 -2300
rect 7440 -2390 7445 -2310
rect 7475 -2390 7480 -2310
rect 7440 -2400 7480 -2390
rect 7760 -2310 7800 -2160
rect 8080 -2200 8120 -2160
rect 8400 -2200 8440 -2160
rect 8720 -2200 8760 -2160
rect 9040 -2200 9080 -2160
rect 9360 -2200 9400 -2160
rect 9680 -2200 9720 -2160
rect 10000 -2200 10040 -2160
rect 10320 -2200 10440 -2160
rect 7840 -2245 8040 -2240
rect 7840 -2275 7850 -2245
rect 8030 -2275 8040 -2245
rect 7840 -2280 8040 -2275
rect 8160 -2245 8360 -2240
rect 8160 -2275 8170 -2245
rect 8350 -2275 8360 -2245
rect 8160 -2280 8360 -2275
rect 8480 -2245 8680 -2240
rect 8480 -2275 8490 -2245
rect 8670 -2275 8680 -2245
rect 8480 -2280 8680 -2275
rect 8800 -2245 9000 -2240
rect 8800 -2275 8810 -2245
rect 8990 -2275 9000 -2245
rect 8800 -2280 9000 -2275
rect 9120 -2245 9320 -2240
rect 9120 -2275 9130 -2245
rect 9310 -2275 9320 -2245
rect 9120 -2280 9320 -2275
rect 9440 -2245 9640 -2240
rect 9440 -2275 9450 -2245
rect 9630 -2275 9640 -2245
rect 9440 -2280 9640 -2275
rect 9760 -2245 9960 -2240
rect 9760 -2275 9770 -2245
rect 9950 -2275 9960 -2245
rect 9760 -2280 9960 -2275
rect 10080 -2245 10280 -2240
rect 10080 -2275 10090 -2245
rect 10270 -2275 10280 -2245
rect 10080 -2280 10280 -2275
rect 7760 -2390 7765 -2310
rect 7795 -2390 7800 -2310
rect 2800 -2520 2840 -2480
rect 3120 -2520 3160 -2480
rect 3440 -2520 3480 -2480
rect 3760 -2520 3800 -2480
rect 4080 -2520 4120 -2480
rect 4400 -2520 4440 -2480
rect 4720 -2520 4760 -2480
rect 5040 -2520 5240 -2480
rect 5520 -2520 5560 -2480
rect 5840 -2520 5880 -2480
rect 6160 -2520 6200 -2480
rect 6480 -2520 6520 -2480
rect 6800 -2520 6840 -2480
rect 7120 -2520 7160 -2480
rect 7440 -2520 7480 -2480
rect 7760 -2520 7800 -2390
rect 8080 -2310 8120 -2300
rect 8080 -2390 8085 -2310
rect 8115 -2390 8120 -2310
rect 8080 -2400 8120 -2390
rect 8400 -2310 8440 -2300
rect 8400 -2390 8405 -2310
rect 8435 -2390 8440 -2310
rect 8400 -2400 8440 -2390
rect 8720 -2310 8760 -2300
rect 8720 -2390 8725 -2310
rect 8755 -2390 8760 -2310
rect 8720 -2400 8760 -2390
rect 9040 -2310 9080 -2300
rect 9040 -2390 9045 -2310
rect 9075 -2390 9080 -2310
rect 9040 -2400 9080 -2390
rect 9360 -2310 9400 -2300
rect 9360 -2390 9365 -2310
rect 9395 -2390 9400 -2310
rect 9360 -2400 9400 -2390
rect 9680 -2310 9720 -2300
rect 9680 -2390 9685 -2310
rect 9715 -2390 9720 -2310
rect 9680 -2400 9720 -2390
rect 10000 -2310 10040 -2300
rect 10000 -2390 10005 -2310
rect 10035 -2390 10040 -2310
rect 10000 -2400 10040 -2390
rect 10320 -2310 10360 -2200
rect 10320 -2390 10325 -2310
rect 10355 -2390 10360 -2310
rect 10320 -2480 10360 -2390
rect 10400 -2240 10440 -2200
rect 10400 -2480 10440 -2440
rect 10560 -2480 10600 -2440
rect 8080 -2520 8120 -2480
rect 8400 -2520 8440 -2480
rect 8720 -2520 8760 -2480
rect 9040 -2520 9080 -2480
rect 9360 -2520 9400 -2480
rect 9680 -2520 9720 -2480
rect 10000 -2520 10040 -2480
rect 10320 -2520 10600 -2480
rect -320 -2600 -40 -2560
rect 240 -2600 280 -2560
rect 560 -2600 600 -2560
rect 880 -2600 920 -2560
rect 1200 -2600 1240 -2560
rect 1520 -2600 1560 -2560
rect 1840 -2600 1880 -2560
rect 2160 -2600 2200 -2560
rect -320 -2640 -280 -2600
rect -160 -2640 -120 -2600
rect -160 -2880 -120 -2840
rect -80 -2690 -40 -2600
rect -80 -2770 -75 -2690
rect -45 -2770 -40 -2690
rect -80 -2880 -40 -2770
rect 240 -2690 280 -2680
rect 240 -2770 245 -2690
rect 275 -2770 280 -2690
rect 240 -2780 280 -2770
rect 560 -2690 600 -2680
rect 560 -2770 565 -2690
rect 595 -2770 600 -2690
rect 560 -2780 600 -2770
rect 880 -2690 920 -2680
rect 880 -2770 885 -2690
rect 915 -2770 920 -2690
rect 880 -2780 920 -2770
rect 1200 -2690 1240 -2680
rect 1200 -2770 1205 -2690
rect 1235 -2770 1240 -2690
rect 1200 -2780 1240 -2770
rect 1520 -2690 1560 -2680
rect 1520 -2770 1525 -2690
rect 1555 -2770 1560 -2690
rect 1520 -2780 1560 -2770
rect 1840 -2690 1880 -2680
rect 1840 -2770 1845 -2690
rect 1875 -2770 1880 -2690
rect 1840 -2780 1880 -2770
rect 2160 -2690 2200 -2680
rect 2160 -2770 2165 -2690
rect 2195 -2770 2200 -2690
rect 2160 -2780 2200 -2770
rect 2480 -2690 2520 -2560
rect 2800 -2600 2840 -2560
rect 3120 -2600 3160 -2560
rect 3440 -2600 3480 -2560
rect 3760 -2600 3800 -2560
rect 4080 -2600 4120 -2560
rect 4400 -2600 4440 -2560
rect 4720 -2600 4760 -2560
rect 5040 -2600 5240 -2560
rect 5520 -2600 5560 -2560
rect 5840 -2600 5880 -2560
rect 6160 -2600 6200 -2560
rect 6480 -2600 6520 -2560
rect 6800 -2600 6840 -2560
rect 7120 -2600 7160 -2560
rect 7440 -2600 7480 -2560
rect 2480 -2770 2485 -2690
rect 2515 -2770 2520 -2690
rect 0 -2805 200 -2800
rect 0 -2835 10 -2805
rect 190 -2835 200 -2805
rect 0 -2840 200 -2835
rect 320 -2805 520 -2800
rect 320 -2835 330 -2805
rect 510 -2835 520 -2805
rect 320 -2840 520 -2835
rect 640 -2805 840 -2800
rect 640 -2835 650 -2805
rect 830 -2835 840 -2805
rect 640 -2840 840 -2835
rect 960 -2805 1160 -2800
rect 960 -2835 970 -2805
rect 1150 -2835 1160 -2805
rect 960 -2840 1160 -2835
rect 1280 -2805 1480 -2800
rect 1280 -2835 1290 -2805
rect 1470 -2835 1480 -2805
rect 1280 -2840 1480 -2835
rect 1600 -2805 1800 -2800
rect 1600 -2835 1610 -2805
rect 1790 -2835 1800 -2805
rect 1600 -2840 1800 -2835
rect 1920 -2805 2120 -2800
rect 1920 -2835 1930 -2805
rect 2110 -2835 2120 -2805
rect 1920 -2840 2120 -2835
rect 2240 -2805 2440 -2800
rect 2240 -2835 2250 -2805
rect 2430 -2835 2440 -2805
rect 2240 -2840 2440 -2835
rect -160 -2920 -40 -2880
rect 240 -2920 280 -2880
rect 560 -2920 600 -2880
rect 880 -2920 920 -2880
rect 1200 -2920 1240 -2880
rect 1520 -2920 1560 -2880
rect 1840 -2920 1880 -2880
rect 2160 -2920 2200 -2880
rect 2480 -2920 2520 -2770
rect 2800 -2690 2840 -2680
rect 2800 -2770 2805 -2690
rect 2835 -2770 2840 -2690
rect 2800 -2780 2840 -2770
rect 3120 -2690 3160 -2680
rect 3120 -2770 3125 -2690
rect 3155 -2770 3160 -2690
rect 3120 -2780 3160 -2770
rect 3440 -2690 3480 -2680
rect 3440 -2770 3445 -2690
rect 3475 -2770 3480 -2690
rect 3440 -2780 3480 -2770
rect 3760 -2690 3800 -2680
rect 3760 -2770 3765 -2690
rect 3795 -2770 3800 -2690
rect 3760 -2780 3800 -2770
rect 4080 -2690 4120 -2680
rect 4080 -2770 4085 -2690
rect 4115 -2770 4120 -2690
rect 4080 -2780 4120 -2770
rect 4400 -2690 4440 -2680
rect 4400 -2770 4405 -2690
rect 4435 -2770 4440 -2690
rect 4400 -2780 4440 -2770
rect 4720 -2690 4760 -2680
rect 4720 -2770 4725 -2690
rect 4755 -2770 4760 -2690
rect 4720 -2780 4760 -2770
rect 5040 -2690 5080 -2600
rect 5040 -2770 5045 -2690
rect 5075 -2770 5080 -2690
rect 2560 -2805 2760 -2800
rect 2560 -2835 2570 -2805
rect 2750 -2835 2760 -2805
rect 2560 -2840 2760 -2835
rect 2880 -2805 3080 -2800
rect 2880 -2835 2890 -2805
rect 3070 -2835 3080 -2805
rect 2880 -2840 3080 -2835
rect 3200 -2805 3400 -2800
rect 3200 -2835 3210 -2805
rect 3390 -2835 3400 -2805
rect 3200 -2840 3400 -2835
rect 3520 -2805 3720 -2800
rect 3520 -2835 3530 -2805
rect 3710 -2835 3720 -2805
rect 3520 -2840 3720 -2835
rect 3840 -2805 4040 -2800
rect 3840 -2835 3850 -2805
rect 4030 -2835 4040 -2805
rect 3840 -2840 4040 -2835
rect 4160 -2805 4360 -2800
rect 4160 -2835 4170 -2805
rect 4350 -2835 4360 -2805
rect 4160 -2840 4360 -2835
rect 4480 -2805 4680 -2800
rect 4480 -2835 4490 -2805
rect 4670 -2835 4680 -2805
rect 4480 -2840 4680 -2835
rect 4800 -2805 5000 -2800
rect 4800 -2835 4810 -2805
rect 4990 -2835 5000 -2805
rect 4800 -2840 5000 -2835
rect 5040 -2880 5080 -2770
rect 5120 -2640 5160 -2600
rect 5120 -2880 5160 -2840
rect 5200 -2690 5240 -2600
rect 5200 -2770 5205 -2690
rect 5235 -2770 5240 -2690
rect 5200 -2880 5240 -2770
rect 5520 -2690 5560 -2680
rect 5520 -2770 5525 -2690
rect 5555 -2770 5560 -2690
rect 5520 -2780 5560 -2770
rect 5840 -2690 5880 -2680
rect 5840 -2770 5845 -2690
rect 5875 -2770 5880 -2690
rect 5840 -2780 5880 -2770
rect 6160 -2690 6200 -2680
rect 6160 -2770 6165 -2690
rect 6195 -2770 6200 -2690
rect 6160 -2780 6200 -2770
rect 6480 -2690 6520 -2680
rect 6480 -2770 6485 -2690
rect 6515 -2770 6520 -2690
rect 6480 -2780 6520 -2770
rect 6800 -2690 6840 -2680
rect 6800 -2770 6805 -2690
rect 6835 -2770 6840 -2690
rect 6800 -2780 6840 -2770
rect 7120 -2690 7160 -2680
rect 7120 -2770 7125 -2690
rect 7155 -2770 7160 -2690
rect 7120 -2780 7160 -2770
rect 7440 -2690 7480 -2680
rect 7440 -2770 7445 -2690
rect 7475 -2770 7480 -2690
rect 7440 -2780 7480 -2770
rect 7760 -2690 7800 -2560
rect 8080 -2600 8120 -2560
rect 8400 -2600 8440 -2560
rect 8720 -2600 8760 -2560
rect 9040 -2600 9080 -2560
rect 9360 -2600 9400 -2560
rect 9680 -2600 9720 -2560
rect 10000 -2600 10040 -2560
rect 10320 -2600 10600 -2560
rect 7760 -2770 7765 -2690
rect 7795 -2770 7800 -2690
rect 5280 -2805 5480 -2800
rect 5280 -2835 5290 -2805
rect 5470 -2835 5480 -2805
rect 5280 -2840 5480 -2835
rect 5600 -2805 5800 -2800
rect 5600 -2835 5610 -2805
rect 5790 -2835 5800 -2805
rect 5600 -2840 5800 -2835
rect 5920 -2805 6120 -2800
rect 5920 -2835 5930 -2805
rect 6110 -2835 6120 -2805
rect 5920 -2840 6120 -2835
rect 6240 -2805 6440 -2800
rect 6240 -2835 6250 -2805
rect 6430 -2835 6440 -2805
rect 6240 -2840 6440 -2835
rect 6560 -2805 6760 -2800
rect 6560 -2835 6570 -2805
rect 6750 -2835 6760 -2805
rect 6560 -2840 6760 -2835
rect 6880 -2805 7080 -2800
rect 6880 -2835 6890 -2805
rect 7070 -2835 7080 -2805
rect 6880 -2840 7080 -2835
rect 7200 -2805 7400 -2800
rect 7200 -2835 7210 -2805
rect 7390 -2835 7400 -2805
rect 7200 -2840 7400 -2835
rect 7520 -2805 7720 -2800
rect 7520 -2835 7530 -2805
rect 7710 -2835 7720 -2805
rect 7520 -2840 7720 -2835
rect 2800 -2920 2840 -2880
rect 3120 -2920 3160 -2880
rect 3440 -2920 3480 -2880
rect 3760 -2920 3800 -2880
rect 4080 -2920 4120 -2880
rect 4400 -2920 4440 -2880
rect 4720 -2920 4760 -2880
rect 5040 -2920 5240 -2880
rect 5520 -2920 5560 -2880
rect 5840 -2920 5880 -2880
rect 6160 -2920 6200 -2880
rect 6480 -2920 6520 -2880
rect 6800 -2920 6840 -2880
rect 7120 -2920 7160 -2880
rect 7440 -2920 7480 -2880
rect 7760 -2920 7800 -2770
rect 8080 -2690 8120 -2680
rect 8080 -2770 8085 -2690
rect 8115 -2770 8120 -2690
rect 8080 -2780 8120 -2770
rect 8400 -2690 8440 -2680
rect 8400 -2770 8405 -2690
rect 8435 -2770 8440 -2690
rect 8400 -2780 8440 -2770
rect 8720 -2690 8760 -2680
rect 8720 -2770 8725 -2690
rect 8755 -2770 8760 -2690
rect 8720 -2780 8760 -2770
rect 9040 -2690 9080 -2680
rect 9040 -2770 9045 -2690
rect 9075 -2770 9080 -2690
rect 9040 -2780 9080 -2770
rect 9360 -2690 9400 -2680
rect 9360 -2770 9365 -2690
rect 9395 -2770 9400 -2690
rect 9360 -2780 9400 -2770
rect 9680 -2690 9720 -2680
rect 9680 -2770 9685 -2690
rect 9715 -2770 9720 -2690
rect 9680 -2780 9720 -2770
rect 10000 -2690 10040 -2680
rect 10000 -2770 10005 -2690
rect 10035 -2770 10040 -2690
rect 10000 -2780 10040 -2770
rect 10320 -2690 10360 -2600
rect 10320 -2770 10325 -2690
rect 10355 -2770 10360 -2690
rect 7840 -2805 8040 -2800
rect 7840 -2835 7850 -2805
rect 8030 -2835 8040 -2805
rect 7840 -2840 8040 -2835
rect 8160 -2805 8360 -2800
rect 8160 -2835 8170 -2805
rect 8350 -2835 8360 -2805
rect 8160 -2840 8360 -2835
rect 8480 -2805 8680 -2800
rect 8480 -2835 8490 -2805
rect 8670 -2835 8680 -2805
rect 8480 -2840 8680 -2835
rect 8800 -2805 9000 -2800
rect 8800 -2835 8810 -2805
rect 8990 -2835 9000 -2805
rect 8800 -2840 9000 -2835
rect 9120 -2805 9320 -2800
rect 9120 -2835 9130 -2805
rect 9310 -2835 9320 -2805
rect 9120 -2840 9320 -2835
rect 9440 -2805 9640 -2800
rect 9440 -2835 9450 -2805
rect 9630 -2835 9640 -2805
rect 9440 -2840 9640 -2835
rect 9760 -2805 9960 -2800
rect 9760 -2835 9770 -2805
rect 9950 -2835 9960 -2805
rect 9760 -2840 9960 -2835
rect 10080 -2805 10280 -2800
rect 10080 -2835 10090 -2805
rect 10270 -2835 10280 -2805
rect 10080 -2840 10280 -2835
rect 10320 -2880 10360 -2770
rect 10400 -2640 10440 -2600
rect 10400 -2880 10440 -2840
rect 10560 -2640 10600 -2600
rect 8080 -2920 8120 -2880
rect 8400 -2920 8440 -2880
rect 8720 -2920 8760 -2880
rect 9040 -2920 9080 -2880
rect 9360 -2920 9400 -2880
rect 9680 -2920 9720 -2880
rect 10000 -2920 10040 -2880
rect 10320 -2920 10480 -2880
rect -280 -3080 -40 -3040
rect 240 -3080 280 -3040
rect 560 -3080 600 -3040
rect 880 -3080 920 -3040
rect 1200 -3080 1240 -3040
rect 1520 -3080 1560 -3040
rect 1840 -3080 1880 -3040
rect 2160 -3080 2200 -3040
rect 2480 -3080 2520 -3040
rect 2800 -3080 2840 -3040
rect 3120 -3080 3160 -3040
rect 3440 -3080 3480 -3040
rect 3760 -3080 3800 -3040
rect 4080 -3080 4120 -3040
rect 4400 -3080 4440 -3040
rect 4720 -3080 4760 -3040
rect 5040 -3080 5240 -3040
rect 5520 -3080 5560 -3040
rect 5840 -3080 5880 -3040
rect 6160 -3080 6200 -3040
rect 6480 -3080 6520 -3040
rect 6800 -3080 6840 -3040
rect 7120 -3080 7160 -3040
rect 7440 -3080 7480 -3040
rect 7760 -3080 7800 -3040
rect 8080 -3080 8120 -3040
rect 8400 -3080 8440 -3040
rect 8720 -3080 8760 -3040
rect 9040 -3080 9080 -3040
rect 9360 -3080 9400 -3040
rect 9680 -3080 9720 -3040
rect 10000 -3080 10040 -3040
rect 10320 -3080 10560 -3040
rect -160 -3240 -40 -3200
rect 240 -3240 280 -3200
rect 560 -3240 600 -3200
rect 880 -3240 920 -3200
rect 1200 -3240 1240 -3200
rect 1520 -3240 1560 -3200
rect 1840 -3240 1880 -3200
rect 2160 -3240 2200 -3200
rect 2480 -3240 2520 -3200
rect 2800 -3240 2840 -3200
rect 3120 -3240 3160 -3200
rect 3440 -3240 3480 -3200
rect 3760 -3240 3800 -3200
rect 4080 -3240 4120 -3200
rect 4400 -3240 4440 -3200
rect 4720 -3240 4760 -3200
rect 5040 -3240 5240 -3200
rect 5520 -3240 5560 -3200
rect -160 -3280 -120 -3240
rect -160 -3520 -120 -3480
rect -80 -3350 -40 -3240
rect 5120 -3280 5160 -3240
rect 0 -3285 200 -3280
rect 0 -3315 10 -3285
rect 190 -3315 200 -3285
rect 0 -3320 200 -3315
rect 320 -3285 520 -3280
rect 320 -3315 330 -3285
rect 510 -3315 520 -3285
rect 320 -3320 520 -3315
rect 640 -3285 840 -3280
rect 640 -3315 650 -3285
rect 830 -3315 840 -3285
rect 640 -3320 840 -3315
rect 960 -3285 1160 -3280
rect 960 -3315 970 -3285
rect 1150 -3315 1160 -3285
rect 960 -3320 1160 -3315
rect 1280 -3285 1480 -3280
rect 1280 -3315 1290 -3285
rect 1470 -3315 1480 -3285
rect 1280 -3320 1480 -3315
rect 1600 -3285 1800 -3280
rect 1600 -3315 1610 -3285
rect 1790 -3315 1800 -3285
rect 1600 -3320 1800 -3315
rect 1920 -3285 2120 -3280
rect 1920 -3315 1930 -3285
rect 2110 -3315 2120 -3285
rect 1920 -3320 2120 -3315
rect 2240 -3285 2440 -3280
rect 2240 -3315 2250 -3285
rect 2430 -3315 2440 -3285
rect 2240 -3320 2440 -3315
rect 2560 -3285 2760 -3280
rect 2560 -3315 2570 -3285
rect 2750 -3315 2760 -3285
rect 2560 -3320 2760 -3315
rect 2880 -3285 3080 -3280
rect 2880 -3315 2890 -3285
rect 3070 -3315 3080 -3285
rect 2880 -3320 3080 -3315
rect 3200 -3285 3400 -3280
rect 3200 -3315 3210 -3285
rect 3390 -3315 3400 -3285
rect 3200 -3320 3400 -3315
rect 3520 -3285 3720 -3280
rect 3520 -3315 3530 -3285
rect 3710 -3315 3720 -3285
rect 3520 -3320 3720 -3315
rect 3840 -3285 4040 -3280
rect 3840 -3315 3850 -3285
rect 4030 -3315 4040 -3285
rect 3840 -3320 4040 -3315
rect 4160 -3285 4360 -3280
rect 4160 -3315 4170 -3285
rect 4350 -3315 4360 -3285
rect 4160 -3320 4360 -3315
rect 4480 -3285 4680 -3280
rect 4480 -3315 4490 -3285
rect 4670 -3315 4680 -3285
rect 4480 -3320 4680 -3315
rect 4800 -3285 5000 -3280
rect 4800 -3315 4810 -3285
rect 4990 -3315 5000 -3285
rect 4800 -3320 5000 -3315
rect -80 -3430 -75 -3350
rect -45 -3430 -40 -3350
rect -80 -3520 -40 -3430
rect 240 -3350 280 -3340
rect 240 -3430 245 -3350
rect 275 -3430 280 -3350
rect 240 -3440 280 -3430
rect 560 -3350 600 -3340
rect 560 -3430 565 -3350
rect 595 -3430 600 -3350
rect 560 -3440 600 -3430
rect 880 -3350 920 -3340
rect 880 -3430 885 -3350
rect 915 -3430 920 -3350
rect 880 -3440 920 -3430
rect 1200 -3350 1240 -3340
rect 1200 -3430 1205 -3350
rect 1235 -3430 1240 -3350
rect 1200 -3440 1240 -3430
rect 1520 -3350 1560 -3340
rect 1520 -3430 1525 -3350
rect 1555 -3430 1560 -3350
rect 1520 -3440 1560 -3430
rect 1840 -3350 1880 -3340
rect 1840 -3430 1845 -3350
rect 1875 -3430 1880 -3350
rect 1840 -3440 1880 -3430
rect 2160 -3350 2200 -3340
rect 2160 -3430 2165 -3350
rect 2195 -3430 2200 -3350
rect 2160 -3440 2200 -3430
rect 2480 -3350 2520 -3340
rect 2480 -3430 2485 -3350
rect 2515 -3430 2520 -3350
rect 2480 -3440 2520 -3430
rect 2800 -3350 2840 -3340
rect 2800 -3430 2805 -3350
rect 2835 -3430 2840 -3350
rect 2800 -3440 2840 -3430
rect 3120 -3350 3160 -3340
rect 3120 -3430 3125 -3350
rect 3155 -3430 3160 -3350
rect 3120 -3440 3160 -3430
rect 3440 -3350 3480 -3340
rect 3440 -3430 3445 -3350
rect 3475 -3430 3480 -3350
rect 3440 -3440 3480 -3430
rect 3760 -3350 3800 -3340
rect 3760 -3430 3765 -3350
rect 3795 -3430 3800 -3350
rect 3760 -3440 3800 -3430
rect 4080 -3350 4120 -3340
rect 4080 -3430 4085 -3350
rect 4115 -3430 4120 -3350
rect 4080 -3440 4120 -3430
rect 4400 -3350 4440 -3340
rect 4400 -3430 4405 -3350
rect 4435 -3430 4440 -3350
rect 4400 -3440 4440 -3430
rect 4720 -3350 4760 -3340
rect 4720 -3430 4725 -3350
rect 4755 -3430 4760 -3350
rect 4720 -3440 4760 -3430
rect 5040 -3350 5080 -3340
rect 5040 -3430 5045 -3350
rect 5075 -3430 5080 -3350
rect 5040 -3440 5080 -3430
rect 5120 -3520 5160 -3480
rect 5200 -3350 5240 -3240
rect 5280 -3285 5480 -3280
rect 5280 -3315 5290 -3285
rect 5470 -3315 5480 -3285
rect 5280 -3320 5480 -3315
rect 5600 -3285 5800 -3280
rect 5600 -3315 5610 -3285
rect 5790 -3315 5800 -3285
rect 5600 -3320 5800 -3315
rect 5200 -3430 5205 -3350
rect 5235 -3430 5240 -3350
rect 5200 -3520 5240 -3430
rect 5520 -3350 5560 -3340
rect 5520 -3430 5525 -3350
rect 5555 -3430 5560 -3350
rect 5520 -3440 5560 -3430
rect 5840 -3350 5880 -3200
rect 6160 -3240 6200 -3200
rect 5920 -3285 6120 -3280
rect 5920 -3315 5930 -3285
rect 6110 -3315 6120 -3285
rect 5920 -3320 6120 -3315
rect 6240 -3285 6440 -3280
rect 6240 -3315 6250 -3285
rect 6430 -3315 6440 -3285
rect 6240 -3320 6440 -3315
rect 5840 -3430 5845 -3350
rect 5875 -3430 5880 -3350
rect -160 -3560 -40 -3520
rect 240 -3560 280 -3520
rect 560 -3560 600 -3520
rect 880 -3560 920 -3520
rect 1200 -3560 1240 -3520
rect 1520 -3560 1560 -3520
rect 1840 -3560 1880 -3520
rect 2160 -3560 2200 -3520
rect 2480 -3560 2520 -3520
rect 2800 -3560 2840 -3520
rect 3120 -3560 3160 -3520
rect 3440 -3560 3480 -3520
rect 3760 -3560 3800 -3520
rect 4080 -3560 4120 -3520
rect 4400 -3560 4440 -3520
rect 4720 -3560 4760 -3520
rect 5040 -3560 5240 -3520
rect 5520 -3560 5560 -3520
rect 5840 -3560 5880 -3430
rect 6160 -3350 6200 -3340
rect 6160 -3430 6165 -3350
rect 6195 -3430 6200 -3350
rect 6160 -3440 6200 -3430
rect 6480 -3350 6520 -3200
rect 6800 -3240 6840 -3200
rect 6560 -3285 6760 -3280
rect 6560 -3315 6570 -3285
rect 6750 -3315 6760 -3285
rect 6560 -3320 6760 -3315
rect 6880 -3285 7080 -3280
rect 6880 -3315 6890 -3285
rect 7070 -3315 7080 -3285
rect 6880 -3320 7080 -3315
rect 6480 -3430 6485 -3350
rect 6515 -3430 6520 -3350
rect 6160 -3560 6200 -3520
rect 6480 -3560 6520 -3430
rect 6800 -3350 6840 -3340
rect 6800 -3430 6805 -3350
rect 6835 -3430 6840 -3350
rect 6800 -3440 6840 -3430
rect 7120 -3350 7160 -3200
rect 7440 -3240 7480 -3200
rect 7200 -3285 7400 -3280
rect 7200 -3315 7210 -3285
rect 7390 -3315 7400 -3285
rect 7200 -3320 7400 -3315
rect 7520 -3285 7720 -3280
rect 7520 -3315 7530 -3285
rect 7710 -3315 7720 -3285
rect 7520 -3320 7720 -3315
rect 7120 -3430 7125 -3350
rect 7155 -3430 7160 -3350
rect 6800 -3560 6840 -3520
rect 7120 -3560 7160 -3430
rect 7440 -3350 7480 -3340
rect 7440 -3430 7445 -3350
rect 7475 -3430 7480 -3350
rect 7440 -3440 7480 -3430
rect 7760 -3350 7800 -3200
rect 8080 -3240 8120 -3200
rect 7840 -3285 8040 -3280
rect 7840 -3315 7850 -3285
rect 8030 -3315 8040 -3285
rect 7840 -3320 8040 -3315
rect 8160 -3285 8360 -3280
rect 8160 -3315 8170 -3285
rect 8350 -3315 8360 -3285
rect 8160 -3320 8360 -3315
rect 7760 -3430 7765 -3350
rect 7795 -3430 7800 -3350
rect 7440 -3560 7480 -3520
rect 7760 -3560 7800 -3430
rect 8080 -3350 8120 -3340
rect 8080 -3430 8085 -3350
rect 8115 -3430 8120 -3350
rect 8080 -3440 8120 -3430
rect 8400 -3350 8440 -3200
rect 8720 -3240 8760 -3200
rect 8480 -3285 8680 -3280
rect 8480 -3315 8490 -3285
rect 8670 -3315 8680 -3285
rect 8480 -3320 8680 -3315
rect 8800 -3285 9000 -3280
rect 8800 -3315 8810 -3285
rect 8990 -3315 9000 -3285
rect 8800 -3320 9000 -3315
rect 8400 -3430 8405 -3350
rect 8435 -3430 8440 -3350
rect 8080 -3560 8120 -3520
rect 8400 -3560 8440 -3430
rect 8720 -3350 8760 -3340
rect 8720 -3430 8725 -3350
rect 8755 -3430 8760 -3350
rect 8720 -3440 8760 -3430
rect 9040 -3350 9080 -3200
rect 9360 -3240 9400 -3200
rect 9120 -3285 9320 -3280
rect 9120 -3315 9130 -3285
rect 9310 -3315 9320 -3285
rect 9120 -3320 9320 -3315
rect 9440 -3285 9640 -3280
rect 9440 -3315 9450 -3285
rect 9630 -3315 9640 -3285
rect 9440 -3320 9640 -3315
rect 9040 -3430 9045 -3350
rect 9075 -3430 9080 -3350
rect 8720 -3560 8760 -3520
rect 9040 -3560 9080 -3430
rect 9360 -3350 9400 -3340
rect 9360 -3430 9365 -3350
rect 9395 -3430 9400 -3350
rect 9360 -3440 9400 -3430
rect 9680 -3350 9720 -3200
rect 10000 -3240 10040 -3200
rect 10320 -3240 10480 -3200
rect 9760 -3285 9960 -3280
rect 9760 -3315 9770 -3285
rect 9950 -3315 9960 -3285
rect 9760 -3320 9960 -3315
rect 10080 -3285 10280 -3280
rect 10080 -3315 10090 -3285
rect 10270 -3315 10280 -3285
rect 10080 -3320 10280 -3315
rect 9680 -3430 9685 -3350
rect 9715 -3430 9720 -3350
rect 9360 -3560 9400 -3520
rect 9680 -3560 9720 -3430
rect 10000 -3350 10040 -3340
rect 10000 -3430 10005 -3350
rect 10035 -3430 10040 -3350
rect 10000 -3440 10040 -3430
rect 10320 -3350 10360 -3240
rect 10320 -3430 10325 -3350
rect 10355 -3430 10360 -3350
rect 10320 -3520 10360 -3430
rect 10400 -3280 10440 -3240
rect 10400 -3520 10440 -3480
rect 10000 -3560 10040 -3520
rect 10320 -3560 10480 -3520
rect -320 -3680 -280 -3640
rect 10560 -3680 10600 -3640
rect -320 -3720 -40 -3680
rect 240 -3720 280 -3680
rect 560 -3720 600 -3680
rect 880 -3720 920 -3680
rect 1200 -3720 1240 -3680
rect 1520 -3720 1560 -3680
rect 1840 -3720 1880 -3680
rect 2160 -3720 2200 -3680
rect 2480 -3720 2520 -3680
rect 2800 -3720 2840 -3680
rect 3120 -3720 3160 -3680
rect 3440 -3720 3480 -3680
rect 3760 -3720 3800 -3680
rect 4080 -3720 4120 -3680
rect 4400 -3720 4440 -3680
rect 4720 -3720 4760 -3680
rect 5040 -3720 5240 -3680
rect 5520 -3720 5560 -3680
rect 5840 -3720 5880 -3680
rect 6160 -3720 6200 -3680
rect 6480 -3720 6520 -3680
rect 6800 -3720 6840 -3680
rect 7120 -3720 7160 -3680
rect 7440 -3720 7480 -3680
rect 7760 -3720 7800 -3680
rect 8080 -3720 8120 -3680
rect 8400 -3720 8440 -3680
rect 8720 -3720 8760 -3680
rect 9040 -3720 9080 -3680
rect 9360 -3720 9400 -3680
rect 9680 -3720 9720 -3680
rect 10000 -3720 10040 -3680
rect 10320 -3720 10600 -3680
<< viali >>
rect -75 670 -45 750
rect 245 670 275 750
rect 565 670 595 750
rect 885 670 915 750
rect 1205 670 1235 750
rect 1525 670 1555 750
rect 1845 670 1875 750
rect 2165 670 2195 750
rect 2485 670 2515 750
rect 2805 670 2835 750
rect 3125 670 3155 750
rect 3445 670 3475 750
rect 3765 670 3795 750
rect 4085 670 4115 750
rect 4405 670 4435 750
rect 4725 670 4755 750
rect 5045 670 5075 750
rect 10 605 190 635
rect 330 605 510 635
rect 650 605 830 635
rect 970 605 1150 635
rect 1290 605 1470 635
rect 1610 605 1790 635
rect 1930 605 2110 635
rect 2250 605 2430 635
rect 2570 605 2750 635
rect 2890 605 3070 635
rect 3210 605 3390 635
rect 3530 605 3710 635
rect 3850 605 4030 635
rect 4170 605 4350 635
rect 4490 605 4670 635
rect 4810 605 4990 635
rect 5205 670 5235 750
rect 5525 670 5555 750
rect 5845 670 5875 750
rect 5290 605 5470 635
rect 5610 605 5790 635
rect 6165 670 6195 750
rect 6485 670 6515 750
rect 5930 605 6110 635
rect 6250 605 6430 635
rect 6805 670 6835 750
rect 7125 670 7155 750
rect 6570 605 6750 635
rect 6890 605 7070 635
rect 7445 670 7475 750
rect 7765 670 7795 750
rect 7210 605 7390 635
rect 7530 605 7710 635
rect 8085 670 8115 750
rect 8405 670 8435 750
rect 7850 605 8030 635
rect 8170 605 8350 635
rect 8725 670 8755 750
rect 9045 670 9075 750
rect 8490 605 8670 635
rect 8810 605 8990 635
rect 9365 670 9395 750
rect 9685 670 9715 750
rect 9130 605 9310 635
rect 9450 605 9630 635
rect 10005 670 10035 750
rect 10325 670 10355 750
rect 9770 605 9950 635
rect 10090 605 10270 635
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect 1290 125 1470 155
rect 1610 125 1790 155
rect 1930 125 2110 155
rect 2250 125 2430 155
rect -75 10 -45 90
rect 245 10 275 90
rect 565 10 595 90
rect 885 10 915 90
rect 1205 10 1235 90
rect 1525 10 1555 90
rect 1845 10 1875 90
rect 2165 10 2195 90
rect 2570 125 2750 155
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3850 125 4030 155
rect 4170 125 4350 155
rect 4490 125 4670 155
rect 4810 125 4990 155
rect 2485 10 2515 90
rect 2805 10 2835 90
rect 3125 10 3155 90
rect 3445 10 3475 90
rect 3765 10 3795 90
rect 4085 10 4115 90
rect 4405 10 4435 90
rect 4725 10 4755 90
rect 5045 10 5075 90
rect 5290 125 5470 155
rect 5610 125 5790 155
rect 5930 125 6110 155
rect 6250 125 6430 155
rect 6570 125 6750 155
rect 6890 125 7070 155
rect 7210 125 7390 155
rect 7530 125 7710 155
rect 5205 10 5235 90
rect 5525 10 5555 90
rect 5845 10 5875 90
rect 6165 10 6195 90
rect 6485 10 6515 90
rect 6805 10 6835 90
rect 7125 10 7155 90
rect 7445 10 7475 90
rect 7850 125 8030 155
rect 8170 125 8350 155
rect 8490 125 8670 155
rect 8810 125 8990 155
rect 9130 125 9310 155
rect 9450 125 9630 155
rect 9770 125 9950 155
rect 10090 125 10270 155
rect 7765 10 7795 90
rect 8085 10 8115 90
rect 8405 10 8435 90
rect 8725 10 8755 90
rect 9045 10 9075 90
rect 9365 10 9395 90
rect 9685 10 9715 90
rect 10005 10 10035 90
rect 10325 10 10355 90
rect -75 -370 -45 -290
rect 245 -370 275 -290
rect 565 -370 595 -290
rect 885 -370 915 -290
rect 1205 -370 1235 -290
rect 1525 -370 1555 -290
rect 1845 -370 1875 -290
rect 2165 -370 2195 -290
rect 2485 -370 2515 -290
rect 10 -435 190 -405
rect 330 -435 510 -405
rect 650 -435 830 -405
rect 970 -435 1150 -405
rect 1290 -435 1470 -405
rect 1610 -435 1790 -405
rect 1930 -435 2110 -405
rect 2250 -435 2430 -405
rect 2805 -370 2835 -290
rect 3125 -370 3155 -290
rect 3445 -370 3475 -290
rect 3765 -370 3795 -290
rect 4085 -370 4115 -290
rect 4405 -370 4435 -290
rect 4725 -370 4755 -290
rect 5045 -370 5075 -290
rect 2570 -435 2750 -405
rect 2890 -435 3070 -405
rect 3210 -435 3390 -405
rect 3530 -435 3710 -405
rect 3850 -435 4030 -405
rect 4170 -435 4350 -405
rect 4490 -435 4670 -405
rect 4810 -435 4990 -405
rect 5205 -370 5235 -290
rect 5525 -370 5555 -290
rect 5845 -370 5875 -290
rect 6165 -370 6195 -290
rect 6485 -370 6515 -290
rect 6805 -370 6835 -290
rect 7125 -370 7155 -290
rect 7445 -370 7475 -290
rect 7765 -370 7795 -290
rect 5290 -435 5470 -405
rect 5610 -435 5790 -405
rect 5930 -435 6110 -405
rect 6250 -435 6430 -405
rect 6570 -435 6750 -405
rect 6890 -435 7070 -405
rect 7210 -435 7390 -405
rect 7530 -435 7710 -405
rect 8085 -370 8115 -290
rect 8405 -370 8435 -290
rect 8725 -370 8755 -290
rect 9045 -370 9075 -290
rect 9365 -370 9395 -290
rect 9685 -370 9715 -290
rect 10005 -370 10035 -290
rect 10325 -370 10355 -290
rect 7850 -435 8030 -405
rect 8170 -435 8350 -405
rect 8490 -435 8670 -405
rect 8810 -435 8990 -405
rect 9130 -435 9310 -405
rect 9450 -435 9630 -405
rect 9770 -435 9950 -405
rect 10090 -435 10270 -405
rect 10 -915 190 -885
rect 330 -915 510 -885
rect -75 -1030 -45 -950
rect 245 -1030 275 -950
rect 650 -915 830 -885
rect 970 -915 1150 -885
rect 565 -1030 595 -950
rect 885 -1030 915 -950
rect 1290 -915 1470 -885
rect 1610 -915 1790 -885
rect 1205 -1030 1235 -950
rect 1525 -1030 1555 -950
rect 1930 -915 2110 -885
rect 2250 -915 2430 -885
rect 1845 -1030 1875 -950
rect 2165 -1030 2195 -950
rect 2570 -915 2750 -885
rect 2890 -915 3070 -885
rect 2485 -1030 2515 -950
rect 2805 -1030 2835 -950
rect 3210 -915 3390 -885
rect 3530 -915 3710 -885
rect 3125 -1030 3155 -950
rect 3445 -1030 3475 -950
rect 3850 -915 4030 -885
rect 4170 -915 4350 -885
rect 3765 -1030 3795 -950
rect 4085 -1030 4115 -950
rect 4490 -915 4670 -885
rect 4810 -915 4990 -885
rect 4405 -1030 4435 -950
rect 4725 -1030 4755 -950
rect 5045 -1030 5075 -950
rect 5290 -915 5470 -885
rect 5610 -915 5790 -885
rect 5930 -915 6110 -885
rect 6250 -915 6430 -885
rect 6570 -915 6750 -885
rect 6890 -915 7070 -885
rect 7210 -915 7390 -885
rect 7530 -915 7710 -885
rect 7850 -915 8030 -885
rect 8170 -915 8350 -885
rect 8490 -915 8670 -885
rect 8810 -915 8990 -885
rect 9130 -915 9310 -885
rect 9450 -915 9630 -885
rect 9770 -915 9950 -885
rect 10090 -915 10270 -885
rect 5205 -1030 5235 -950
rect 5525 -1030 5555 -950
rect 5845 -1030 5875 -950
rect 6165 -1030 6195 -950
rect 6485 -1030 6515 -950
rect 6805 -1030 6835 -950
rect 7125 -1030 7155 -950
rect 7445 -1030 7475 -950
rect 7765 -1030 7795 -950
rect 8085 -1030 8115 -950
rect 8405 -1030 8435 -950
rect 8725 -1030 8755 -950
rect 9045 -1030 9075 -950
rect 9365 -1030 9395 -950
rect 9685 -1030 9715 -950
rect 10005 -1030 10035 -950
rect 10325 -1030 10355 -950
rect -75 -1730 -45 -1650
rect 245 -1730 275 -1650
rect 565 -1730 595 -1650
rect 10 -1795 190 -1765
rect 330 -1795 510 -1765
rect 885 -1730 915 -1650
rect 1205 -1730 1235 -1650
rect 650 -1795 830 -1765
rect 970 -1795 1150 -1765
rect 1525 -1730 1555 -1650
rect 1845 -1730 1875 -1650
rect 1290 -1795 1470 -1765
rect 1610 -1795 1790 -1765
rect 2165 -1730 2195 -1650
rect 2485 -1730 2515 -1650
rect 1930 -1795 2110 -1765
rect 2250 -1795 2430 -1765
rect 2805 -1730 2835 -1650
rect 3125 -1730 3155 -1650
rect 2570 -1795 2750 -1765
rect 2890 -1795 3070 -1765
rect 3445 -1730 3475 -1650
rect 3765 -1730 3795 -1650
rect 3210 -1795 3390 -1765
rect 3530 -1795 3710 -1765
rect 4085 -1730 4115 -1650
rect 4405 -1730 4435 -1650
rect 3850 -1795 4030 -1765
rect 4170 -1795 4350 -1765
rect 4725 -1730 4755 -1650
rect 5045 -1730 5075 -1650
rect 4490 -1795 4670 -1765
rect 4810 -1795 4990 -1765
rect 5205 -1730 5235 -1650
rect 5525 -1730 5555 -1650
rect 5845 -1730 5875 -1650
rect 6165 -1730 6195 -1650
rect 6485 -1730 6515 -1650
rect 6805 -1730 6835 -1650
rect 7125 -1730 7155 -1650
rect 7445 -1730 7475 -1650
rect 7765 -1730 7795 -1650
rect 8085 -1730 8115 -1650
rect 8405 -1730 8435 -1650
rect 8725 -1730 8755 -1650
rect 9045 -1730 9075 -1650
rect 9365 -1730 9395 -1650
rect 9685 -1730 9715 -1650
rect 10005 -1730 10035 -1650
rect 10325 -1730 10355 -1650
rect 5290 -1795 5470 -1765
rect 5610 -1795 5790 -1765
rect 5930 -1795 6110 -1765
rect 6250 -1795 6430 -1765
rect 6570 -1795 6750 -1765
rect 6890 -1795 7070 -1765
rect 7210 -1795 7390 -1765
rect 7530 -1795 7710 -1765
rect 7850 -1795 8030 -1765
rect 8170 -1795 8350 -1765
rect 8490 -1795 8670 -1765
rect 8810 -1795 8990 -1765
rect 9130 -1795 9310 -1765
rect 9450 -1795 9630 -1765
rect 9770 -1795 9950 -1765
rect 10090 -1795 10270 -1765
rect 10 -2275 190 -2245
rect 330 -2275 510 -2245
rect 650 -2275 830 -2245
rect 970 -2275 1150 -2245
rect 1290 -2275 1470 -2245
rect 1610 -2275 1790 -2245
rect 1930 -2275 2110 -2245
rect 2250 -2275 2430 -2245
rect -75 -2390 -45 -2310
rect 245 -2390 275 -2310
rect 565 -2390 595 -2310
rect 885 -2390 915 -2310
rect 1205 -2390 1235 -2310
rect 1525 -2390 1555 -2310
rect 1845 -2390 1875 -2310
rect 2165 -2390 2195 -2310
rect 2570 -2275 2750 -2245
rect 2890 -2275 3070 -2245
rect 3210 -2275 3390 -2245
rect 3530 -2275 3710 -2245
rect 3850 -2275 4030 -2245
rect 4170 -2275 4350 -2245
rect 4490 -2275 4670 -2245
rect 4810 -2275 4990 -2245
rect 2485 -2390 2515 -2310
rect 2805 -2390 2835 -2310
rect 3125 -2390 3155 -2310
rect 3445 -2390 3475 -2310
rect 3765 -2390 3795 -2310
rect 4085 -2390 4115 -2310
rect 4405 -2390 4435 -2310
rect 4725 -2390 4755 -2310
rect 5045 -2390 5075 -2310
rect 5290 -2275 5470 -2245
rect 5610 -2275 5790 -2245
rect 5930 -2275 6110 -2245
rect 6250 -2275 6430 -2245
rect 6570 -2275 6750 -2245
rect 6890 -2275 7070 -2245
rect 7210 -2275 7390 -2245
rect 7530 -2275 7710 -2245
rect 5205 -2390 5235 -2310
rect 5525 -2390 5555 -2310
rect 5845 -2390 5875 -2310
rect 6165 -2390 6195 -2310
rect 6485 -2390 6515 -2310
rect 6805 -2390 6835 -2310
rect 7125 -2390 7155 -2310
rect 7445 -2390 7475 -2310
rect 7850 -2275 8030 -2245
rect 8170 -2275 8350 -2245
rect 8490 -2275 8670 -2245
rect 8810 -2275 8990 -2245
rect 9130 -2275 9310 -2245
rect 9450 -2275 9630 -2245
rect 9770 -2275 9950 -2245
rect 10090 -2275 10270 -2245
rect 7765 -2390 7795 -2310
rect 8085 -2390 8115 -2310
rect 8405 -2390 8435 -2310
rect 8725 -2390 8755 -2310
rect 9045 -2390 9075 -2310
rect 9365 -2390 9395 -2310
rect 9685 -2390 9715 -2310
rect 10005 -2390 10035 -2310
rect 10325 -2390 10355 -2310
rect -75 -2770 -45 -2690
rect 245 -2770 275 -2690
rect 565 -2770 595 -2690
rect 885 -2770 915 -2690
rect 1205 -2770 1235 -2690
rect 1525 -2770 1555 -2690
rect 1845 -2770 1875 -2690
rect 2165 -2770 2195 -2690
rect 2485 -2770 2515 -2690
rect 10 -2835 190 -2805
rect 330 -2835 510 -2805
rect 650 -2835 830 -2805
rect 970 -2835 1150 -2805
rect 1290 -2835 1470 -2805
rect 1610 -2835 1790 -2805
rect 1930 -2835 2110 -2805
rect 2250 -2835 2430 -2805
rect 2805 -2770 2835 -2690
rect 3125 -2770 3155 -2690
rect 3445 -2770 3475 -2690
rect 3765 -2770 3795 -2690
rect 4085 -2770 4115 -2690
rect 4405 -2770 4435 -2690
rect 4725 -2770 4755 -2690
rect 5045 -2770 5075 -2690
rect 2570 -2835 2750 -2805
rect 2890 -2835 3070 -2805
rect 3210 -2835 3390 -2805
rect 3530 -2835 3710 -2805
rect 3850 -2835 4030 -2805
rect 4170 -2835 4350 -2805
rect 4490 -2835 4670 -2805
rect 4810 -2835 4990 -2805
rect 5205 -2770 5235 -2690
rect 5525 -2770 5555 -2690
rect 5845 -2770 5875 -2690
rect 6165 -2770 6195 -2690
rect 6485 -2770 6515 -2690
rect 6805 -2770 6835 -2690
rect 7125 -2770 7155 -2690
rect 7445 -2770 7475 -2690
rect 7765 -2770 7795 -2690
rect 5290 -2835 5470 -2805
rect 5610 -2835 5790 -2805
rect 5930 -2835 6110 -2805
rect 6250 -2835 6430 -2805
rect 6570 -2835 6750 -2805
rect 6890 -2835 7070 -2805
rect 7210 -2835 7390 -2805
rect 7530 -2835 7710 -2805
rect 8085 -2770 8115 -2690
rect 8405 -2770 8435 -2690
rect 8725 -2770 8755 -2690
rect 9045 -2770 9075 -2690
rect 9365 -2770 9395 -2690
rect 9685 -2770 9715 -2690
rect 10005 -2770 10035 -2690
rect 10325 -2770 10355 -2690
rect 7850 -2835 8030 -2805
rect 8170 -2835 8350 -2805
rect 8490 -2835 8670 -2805
rect 8810 -2835 8990 -2805
rect 9130 -2835 9310 -2805
rect 9450 -2835 9630 -2805
rect 9770 -2835 9950 -2805
rect 10090 -2835 10270 -2805
rect 10 -3315 190 -3285
rect 330 -3315 510 -3285
rect 650 -3315 830 -3285
rect 970 -3315 1150 -3285
rect 1290 -3315 1470 -3285
rect 1610 -3315 1790 -3285
rect 1930 -3315 2110 -3285
rect 2250 -3315 2430 -3285
rect 2570 -3315 2750 -3285
rect 2890 -3315 3070 -3285
rect 3210 -3315 3390 -3285
rect 3530 -3315 3710 -3285
rect 3850 -3315 4030 -3285
rect 4170 -3315 4350 -3285
rect 4490 -3315 4670 -3285
rect 4810 -3315 4990 -3285
rect -75 -3430 -45 -3350
rect 245 -3430 275 -3350
rect 565 -3430 595 -3350
rect 885 -3430 915 -3350
rect 1205 -3430 1235 -3350
rect 1525 -3430 1555 -3350
rect 1845 -3430 1875 -3350
rect 2165 -3430 2195 -3350
rect 2485 -3430 2515 -3350
rect 2805 -3430 2835 -3350
rect 3125 -3430 3155 -3350
rect 3445 -3430 3475 -3350
rect 3765 -3430 3795 -3350
rect 4085 -3430 4115 -3350
rect 4405 -3430 4435 -3350
rect 4725 -3430 4755 -3350
rect 5045 -3430 5075 -3350
rect 5290 -3315 5470 -3285
rect 5610 -3315 5790 -3285
rect 5205 -3430 5235 -3350
rect 5525 -3430 5555 -3350
rect 5930 -3315 6110 -3285
rect 6250 -3315 6430 -3285
rect 5845 -3430 5875 -3350
rect 6165 -3430 6195 -3350
rect 6570 -3315 6750 -3285
rect 6890 -3315 7070 -3285
rect 6485 -3430 6515 -3350
rect 6805 -3430 6835 -3350
rect 7210 -3315 7390 -3285
rect 7530 -3315 7710 -3285
rect 7125 -3430 7155 -3350
rect 7445 -3430 7475 -3350
rect 7850 -3315 8030 -3285
rect 8170 -3315 8350 -3285
rect 7765 -3430 7795 -3350
rect 8085 -3430 8115 -3350
rect 8490 -3315 8670 -3285
rect 8810 -3315 8990 -3285
rect 8405 -3430 8435 -3350
rect 8725 -3430 8755 -3350
rect 9130 -3315 9310 -3285
rect 9450 -3315 9630 -3285
rect 9045 -3430 9075 -3350
rect 9365 -3430 9395 -3350
rect 9770 -3315 9950 -3285
rect 10090 -3315 10270 -3285
rect 9685 -3430 9715 -3350
rect 10005 -3430 10035 -3350
rect 10325 -3430 10355 -3350
<< metal1 >>
rect -720 1035 -680 1040
rect -720 1005 -715 1035
rect -685 1005 -680 1035
rect -720 1000 -680 1005
rect -560 1035 -520 1040
rect -560 1005 -555 1035
rect -525 1005 -520 1035
rect -560 1000 -520 1005
rect -400 1035 -360 1040
rect -400 1005 -395 1035
rect -365 1005 -360 1035
rect -400 1000 -360 1005
rect 10640 1035 10680 1040
rect 10640 1005 10645 1035
rect 10675 1005 10680 1035
rect 10640 1000 10680 1005
rect 10800 1035 10840 1040
rect 10800 1005 10805 1035
rect 10835 1005 10840 1035
rect 10800 1000 10840 1005
rect 10960 1035 11000 1040
rect 10960 1005 10965 1035
rect 10995 1005 11000 1035
rect 10960 1000 11000 1005
rect -720 955 -680 960
rect -720 925 -715 955
rect -685 925 -680 955
rect -720 920 -680 925
rect -560 955 -520 960
rect -560 925 -555 955
rect -525 925 -520 955
rect -560 920 -520 925
rect -400 955 -360 960
rect -400 925 -395 955
rect -365 925 -360 955
rect -400 920 -360 925
rect 10640 955 10680 960
rect 10640 925 10645 955
rect 10675 925 10680 955
rect 10640 920 10680 925
rect 10800 955 10840 960
rect 10800 925 10805 955
rect 10835 925 10840 955
rect 10800 920 10840 925
rect 10960 955 11000 960
rect 10960 925 10965 955
rect 10995 925 11000 955
rect 10960 920 11000 925
rect -720 875 -680 880
rect -720 845 -715 875
rect -685 845 -680 875
rect -720 840 -680 845
rect -560 875 -520 880
rect -560 845 -555 875
rect -525 845 -520 875
rect -560 840 -520 845
rect -400 875 -360 880
rect -400 845 -395 875
rect -365 845 -360 875
rect -400 840 -360 845
rect 10640 875 10680 880
rect 10640 845 10645 875
rect 10675 845 10680 875
rect 10640 840 10680 845
rect 10800 875 10840 880
rect 10800 845 10805 875
rect 10835 845 10840 875
rect 10800 840 10840 845
rect 10960 875 11000 880
rect 10960 845 10965 875
rect 10995 845 11000 875
rect 10960 840 11000 845
rect -80 795 -40 800
rect -80 765 -75 795
rect -45 765 -40 795
rect -80 750 -40 765
rect 5200 795 5240 800
rect 5200 765 5205 795
rect 5235 765 5240 795
rect -80 670 -75 750
rect -45 670 -40 750
rect -80 660 -40 670
rect 240 750 280 760
rect 240 670 245 750
rect 275 670 280 750
rect 240 660 280 670
rect 560 750 600 760
rect 560 670 565 750
rect 595 670 600 750
rect 560 660 600 670
rect 880 750 920 760
rect 880 670 885 750
rect 915 670 920 750
rect 880 660 920 670
rect 1200 750 1240 760
rect 1200 670 1205 750
rect 1235 670 1240 750
rect 1200 660 1240 670
rect 1520 750 1560 760
rect 1520 670 1525 750
rect 1555 670 1560 750
rect 1520 660 1560 670
rect 1840 750 1880 760
rect 1840 670 1845 750
rect 1875 670 1880 750
rect 1840 660 1880 670
rect 2160 750 2200 760
rect 2160 670 2165 750
rect 2195 670 2200 750
rect 2160 660 2200 670
rect 2480 750 2520 760
rect 2480 670 2485 750
rect 2515 670 2520 750
rect 2480 660 2520 670
rect 2800 750 2840 760
rect 2800 670 2805 750
rect 2835 670 2840 750
rect 2800 660 2840 670
rect 3120 750 3160 760
rect 3120 670 3125 750
rect 3155 670 3160 750
rect 3120 660 3160 670
rect 3440 750 3480 760
rect 3440 670 3445 750
rect 3475 670 3480 750
rect 3440 660 3480 670
rect 3760 750 3800 760
rect 3760 670 3765 750
rect 3795 670 3800 750
rect 3760 660 3800 670
rect 4080 750 4120 760
rect 4080 670 4085 750
rect 4115 670 4120 750
rect 4080 660 4120 670
rect 4400 750 4440 760
rect 4400 670 4405 750
rect 4435 670 4440 750
rect 4400 660 4440 670
rect 4720 750 4760 760
rect 4720 670 4725 750
rect 4755 670 4760 750
rect 4720 660 4760 670
rect 5040 750 5080 760
rect 5040 670 5045 750
rect 5075 670 5080 750
rect -720 635 -680 640
rect -720 605 -715 635
rect -685 605 -680 635
rect -720 600 -680 605
rect -560 635 -520 640
rect -560 605 -555 635
rect -525 605 -520 635
rect -560 600 -520 605
rect -400 635 -360 640
rect -400 605 -395 635
rect -365 605 -360 635
rect -400 600 -360 605
rect 0 635 200 640
rect 0 605 10 635
rect 190 605 200 635
rect 0 600 200 605
rect 320 635 520 640
rect 320 605 330 635
rect 510 605 520 635
rect 320 600 520 605
rect 640 635 840 640
rect 640 605 650 635
rect 830 605 840 635
rect 640 600 840 605
rect 960 635 1160 640
rect 960 605 970 635
rect 1150 605 1160 635
rect 960 600 1160 605
rect 1280 635 1480 640
rect 1280 605 1290 635
rect 1470 605 1480 635
rect 1280 600 1480 605
rect 1600 635 1800 640
rect 1600 605 1610 635
rect 1790 605 1800 635
rect 1600 600 1800 605
rect 1920 635 2120 640
rect 1920 605 1930 635
rect 2110 605 2120 635
rect 1920 600 2120 605
rect 2240 635 2440 640
rect 2240 605 2250 635
rect 2430 605 2440 635
rect 2240 600 2440 605
rect 2560 635 2760 640
rect 2560 605 2570 635
rect 2750 605 2760 635
rect 2560 600 2760 605
rect 2880 635 3080 640
rect 2880 605 2890 635
rect 3070 605 3080 635
rect 2880 600 3080 605
rect 3200 635 3400 640
rect 3200 605 3210 635
rect 3390 605 3400 635
rect 3200 600 3400 605
rect 3520 635 3720 640
rect 3520 605 3530 635
rect 3710 605 3720 635
rect 3520 600 3720 605
rect 3840 635 4040 640
rect 3840 605 3850 635
rect 4030 605 4040 635
rect 3840 600 4040 605
rect 4160 635 4360 640
rect 4160 605 4170 635
rect 4350 605 4360 635
rect 4160 600 4360 605
rect 4480 635 4680 640
rect 4480 605 4490 635
rect 4670 605 4680 635
rect 4480 600 4680 605
rect 4800 635 5000 640
rect 4800 605 4810 635
rect 4990 605 5000 635
rect 4800 600 5000 605
rect -720 555 -680 560
rect -720 525 -715 555
rect -685 525 -680 555
rect -720 520 -680 525
rect -560 555 -520 560
rect -560 525 -555 555
rect -525 525 -520 555
rect -560 520 -520 525
rect -400 555 -360 560
rect -400 525 -395 555
rect -365 525 -360 555
rect -400 520 -360 525
rect -720 475 -680 480
rect -720 445 -715 475
rect -685 445 -680 475
rect -720 440 -680 445
rect -560 475 -520 480
rect -560 445 -555 475
rect -525 445 -520 475
rect -560 440 -520 445
rect 80 475 120 600
rect 80 445 85 475
rect 115 445 120 475
rect 80 440 120 445
rect 400 475 440 600
rect 400 445 405 475
rect 435 445 440 475
rect 400 440 440 445
rect 720 475 760 600
rect 720 445 725 475
rect 755 445 760 475
rect 720 440 760 445
rect 1040 475 1080 600
rect 1040 445 1045 475
rect 1075 445 1080 475
rect 1040 440 1080 445
rect 1360 475 1400 600
rect 1360 445 1365 475
rect 1395 445 1400 475
rect 1360 440 1400 445
rect 1680 475 1720 600
rect 1680 445 1685 475
rect 1715 445 1720 475
rect 1680 440 1720 445
rect 2000 475 2040 600
rect 2000 445 2005 475
rect 2035 445 2040 475
rect 2000 440 2040 445
rect 2320 475 2360 600
rect 2320 445 2325 475
rect 2355 445 2360 475
rect 2320 440 2360 445
rect 2640 475 2680 600
rect 2640 445 2645 475
rect 2675 445 2680 475
rect 2640 440 2680 445
rect 2960 475 3000 600
rect 2960 445 2965 475
rect 2995 445 3000 475
rect 2960 440 3000 445
rect 3280 475 3320 600
rect 3280 445 3285 475
rect 3315 445 3320 475
rect 3280 440 3320 445
rect 3600 475 3640 600
rect 3600 445 3605 475
rect 3635 445 3640 475
rect 3600 440 3640 445
rect 3920 475 3960 600
rect 3920 445 3925 475
rect 3955 445 3960 475
rect 3920 440 3960 445
rect 4240 475 4280 600
rect 4240 445 4245 475
rect 4275 445 4280 475
rect 4240 440 4280 445
rect 4560 475 4600 600
rect 4560 445 4565 475
rect 4595 445 4600 475
rect 4560 440 4600 445
rect 4880 475 4920 600
rect 4880 445 4885 475
rect 4915 445 4920 475
rect 4880 440 4920 445
rect -720 395 -680 400
rect -720 365 -715 395
rect -685 365 -680 395
rect -720 360 -680 365
rect -560 395 -520 400
rect -560 365 -555 395
rect -525 365 -520 395
rect -560 360 -520 365
rect -400 395 -360 400
rect -400 365 -395 395
rect -365 365 -360 395
rect -400 360 -360 365
rect -720 315 -680 320
rect -720 285 -715 315
rect -685 285 -680 315
rect -720 280 -680 285
rect -560 315 -520 320
rect -560 285 -555 315
rect -525 285 -520 315
rect -560 280 -520 285
rect -400 315 -360 320
rect -400 285 -395 315
rect -365 285 -360 315
rect -400 280 -360 285
rect -720 235 -680 240
rect -720 205 -715 235
rect -685 205 -680 235
rect -720 200 -680 205
rect -560 235 -520 240
rect -560 205 -555 235
rect -525 205 -520 235
rect -560 200 -520 205
rect -400 235 -360 240
rect -400 205 -395 235
rect -365 205 -360 235
rect -400 200 -360 205
rect -720 155 -680 160
rect -720 125 -715 155
rect -685 125 -680 155
rect -720 120 -680 125
rect -560 155 -520 160
rect -560 125 -555 155
rect -525 125 -520 155
rect -560 120 -520 125
rect -400 155 -360 160
rect -400 125 -395 155
rect -365 125 -360 155
rect -400 120 -360 125
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 120 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 120 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 120 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 120 1160 125
rect 1200 155 1240 160
rect 1200 125 1205 155
rect 1235 125 1240 155
rect -80 90 -40 100
rect -720 75 -680 80
rect -720 45 -715 75
rect -685 45 -680 75
rect -720 40 -680 45
rect -560 75 -520 80
rect -560 45 -555 75
rect -525 45 -520 75
rect -560 40 -520 45
rect -400 75 -360 80
rect -400 45 -395 75
rect -365 45 -360 75
rect -400 40 -360 45
rect -80 10 -75 90
rect -45 10 -40 90
rect -720 -5 -680 0
rect -720 -35 -715 -5
rect -685 -35 -680 -5
rect -720 -40 -680 -35
rect -560 -5 -520 0
rect -560 -35 -555 -5
rect -525 -35 -520 -5
rect -560 -40 -520 -35
rect -400 -5 -360 0
rect -400 -35 -395 -5
rect -365 -35 -360 -5
rect -400 -40 -360 -35
rect -80 -5 -40 10
rect 240 90 280 100
rect 240 10 245 90
rect 275 10 280 90
rect 240 0 280 10
rect 560 90 600 100
rect 560 10 565 90
rect 595 10 600 90
rect 560 0 600 10
rect 880 90 920 100
rect 880 10 885 90
rect 915 10 920 90
rect 880 0 920 10
rect 1200 90 1240 125
rect 1280 155 1480 160
rect 1280 125 1290 155
rect 1470 125 1480 155
rect 1280 120 1480 125
rect 1600 155 1800 160
rect 1600 125 1610 155
rect 1790 125 1800 155
rect 1600 120 1800 125
rect 1920 155 2120 160
rect 1920 125 1930 155
rect 2110 125 2120 155
rect 1920 120 2120 125
rect 2240 155 2440 160
rect 2240 125 2250 155
rect 2430 125 2440 155
rect 2240 120 2440 125
rect 2560 155 2760 160
rect 2560 125 2570 155
rect 2750 125 2760 155
rect 2560 120 2760 125
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 120 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 120 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 120 3720 125
rect 3760 155 3800 160
rect 3760 125 3765 155
rect 3795 125 3800 155
rect 1200 10 1205 90
rect 1235 10 1240 90
rect 1200 0 1240 10
rect 1520 90 1560 100
rect 1520 10 1525 90
rect 1555 10 1560 90
rect 1520 0 1560 10
rect 1840 90 1880 100
rect 1840 10 1845 90
rect 1875 10 1880 90
rect 1840 0 1880 10
rect 2160 90 2200 100
rect 2160 10 2165 90
rect 2195 10 2200 90
rect 2160 0 2200 10
rect 2480 90 2520 100
rect 2480 10 2485 90
rect 2515 10 2520 90
rect -80 -35 -75 -5
rect -45 -35 -40 -5
rect -80 -40 -40 -35
rect 2480 -5 2520 10
rect 2800 90 2840 100
rect 2800 10 2805 90
rect 2835 10 2840 90
rect 2800 0 2840 10
rect 3120 90 3160 100
rect 3120 10 3125 90
rect 3155 10 3160 90
rect 3120 0 3160 10
rect 3440 90 3480 100
rect 3440 10 3445 90
rect 3475 10 3480 90
rect 3440 0 3480 10
rect 3760 90 3800 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 120 4040 125
rect 4160 155 4360 160
rect 4160 125 4170 155
rect 4350 125 4360 155
rect 4160 120 4360 125
rect 4480 155 4680 160
rect 4480 125 4490 155
rect 4670 125 4680 155
rect 4480 120 4680 125
rect 4800 155 5000 160
rect 4800 125 4810 155
rect 4990 125 5000 155
rect 4800 120 5000 125
rect 5040 155 5080 670
rect 5200 750 5240 765
rect 5840 795 5880 800
rect 5840 765 5845 795
rect 5875 765 5880 795
rect 5200 670 5205 750
rect 5235 670 5240 750
rect 5200 660 5240 670
rect 5520 750 5560 760
rect 5520 670 5525 750
rect 5555 670 5560 750
rect 5280 635 5480 640
rect 5280 605 5290 635
rect 5470 605 5480 635
rect 5280 600 5480 605
rect 5360 315 5400 600
rect 5360 285 5365 315
rect 5395 285 5400 315
rect 5360 280 5400 285
rect 5520 315 5560 670
rect 5840 750 5880 765
rect 6480 795 6520 800
rect 6480 765 6485 795
rect 6515 765 6520 795
rect 5840 670 5845 750
rect 5875 670 5880 750
rect 5840 660 5880 670
rect 6160 750 6200 760
rect 6160 670 6165 750
rect 6195 670 6200 750
rect 6160 660 6200 670
rect 6480 750 6520 765
rect 7120 795 7160 800
rect 7120 765 7125 795
rect 7155 765 7160 795
rect 6480 670 6485 750
rect 6515 670 6520 750
rect 6480 660 6520 670
rect 6800 750 6840 760
rect 6800 670 6805 750
rect 6835 670 6840 750
rect 6800 660 6840 670
rect 7120 750 7160 765
rect 7760 795 7800 800
rect 7760 765 7765 795
rect 7795 765 7800 795
rect 7120 670 7125 750
rect 7155 670 7160 750
rect 7120 660 7160 670
rect 7440 750 7480 760
rect 7440 670 7445 750
rect 7475 670 7480 750
rect 7440 660 7480 670
rect 7760 750 7800 765
rect 8400 795 8440 800
rect 8400 765 8405 795
rect 8435 765 8440 795
rect 7760 670 7765 750
rect 7795 670 7800 750
rect 7760 660 7800 670
rect 8080 750 8120 760
rect 8080 670 8085 750
rect 8115 670 8120 750
rect 5600 635 5800 640
rect 5600 605 5610 635
rect 5790 605 5800 635
rect 5600 600 5800 605
rect 5920 635 6120 640
rect 5920 605 5930 635
rect 6110 605 6120 635
rect 5920 600 6120 605
rect 6240 635 6440 640
rect 6240 605 6250 635
rect 6430 605 6440 635
rect 6240 600 6440 605
rect 6560 635 6760 640
rect 6560 605 6570 635
rect 6750 605 6760 635
rect 6560 600 6760 605
rect 6880 635 7080 640
rect 6880 605 6890 635
rect 7070 605 7080 635
rect 6880 600 7080 605
rect 7200 635 7400 640
rect 7200 605 7210 635
rect 7390 605 7400 635
rect 7200 600 7400 605
rect 7520 635 7720 640
rect 7520 605 7530 635
rect 7710 605 7720 635
rect 7520 600 7720 605
rect 7840 635 8040 640
rect 7840 605 7850 635
rect 8030 605 8040 635
rect 7840 600 8040 605
rect 5520 285 5525 315
rect 5555 285 5560 315
rect 5520 280 5560 285
rect 5680 315 5720 600
rect 5680 285 5685 315
rect 5715 285 5720 315
rect 5680 280 5720 285
rect 6000 315 6040 600
rect 6000 285 6005 315
rect 6035 285 6040 315
rect 6000 280 6040 285
rect 6160 315 6200 600
rect 6160 285 6165 315
rect 6195 285 6200 315
rect 6160 280 6200 285
rect 6320 315 6360 600
rect 6320 285 6325 315
rect 6355 285 6360 315
rect 6320 280 6360 285
rect 6480 315 6520 320
rect 6480 285 6485 315
rect 6515 285 6520 315
rect 5040 125 5045 155
rect 5075 125 5080 155
rect 5040 120 5080 125
rect 5280 155 5480 160
rect 5280 125 5290 155
rect 5470 125 5480 155
rect 5280 120 5480 125
rect 5600 155 5800 160
rect 5600 125 5610 155
rect 5790 125 5800 155
rect 5600 120 5800 125
rect 5920 155 6120 160
rect 5920 125 5930 155
rect 6110 125 6120 155
rect 5920 120 6120 125
rect 6240 155 6440 160
rect 6240 125 6250 155
rect 6430 125 6440 155
rect 6240 120 6440 125
rect 3760 10 3765 90
rect 3795 10 3800 90
rect 3760 0 3800 10
rect 4080 90 4120 100
rect 4080 10 4085 90
rect 4115 10 4120 90
rect 4080 0 4120 10
rect 4400 90 4440 100
rect 4400 10 4405 90
rect 4435 10 4440 90
rect 4400 0 4440 10
rect 4720 90 4760 100
rect 4720 10 4725 90
rect 4755 10 4760 90
rect 4720 0 4760 10
rect 5040 90 5080 100
rect 5040 10 5045 90
rect 5075 10 5080 90
rect 2480 -35 2485 -5
rect 2515 -35 2520 -5
rect 2480 -40 2520 -35
rect 5040 -5 5080 10
rect 5040 -35 5045 -5
rect 5075 -35 5080 -5
rect 5040 -40 5080 -35
rect 5200 90 5240 100
rect 5200 10 5205 90
rect 5235 10 5240 90
rect 5200 -5 5240 10
rect 5520 90 5560 100
rect 5520 10 5525 90
rect 5555 10 5560 90
rect 5520 0 5560 10
rect 5840 90 5880 100
rect 5840 10 5845 90
rect 5875 10 5880 90
rect 5840 0 5880 10
rect 6160 90 6200 100
rect 6160 10 6165 90
rect 6195 10 6200 90
rect 6160 0 6200 10
rect 6480 90 6520 285
rect 6640 315 6680 600
rect 6640 285 6645 315
rect 6675 285 6680 315
rect 6640 280 6680 285
rect 6800 315 6840 600
rect 6800 285 6805 315
rect 6835 285 6840 315
rect 6800 280 6840 285
rect 6960 315 7000 600
rect 6960 285 6965 315
rect 6995 285 7000 315
rect 6960 280 7000 285
rect 7280 315 7320 600
rect 7280 285 7285 315
rect 7315 285 7320 315
rect 7280 280 7320 285
rect 7440 315 7480 600
rect 7440 285 7445 315
rect 7475 285 7480 315
rect 7440 280 7480 285
rect 7600 315 7640 600
rect 7600 285 7605 315
rect 7635 285 7640 315
rect 7600 280 7640 285
rect 7920 315 7960 600
rect 7920 285 7925 315
rect 7955 285 7960 315
rect 7920 280 7960 285
rect 8080 315 8120 670
rect 8400 750 8440 765
rect 9040 795 9080 800
rect 9040 765 9045 795
rect 9075 765 9080 795
rect 8400 670 8405 750
rect 8435 670 8440 750
rect 8400 660 8440 670
rect 8720 750 8760 760
rect 8720 670 8725 750
rect 8755 670 8760 750
rect 8160 635 8360 640
rect 8160 605 8170 635
rect 8350 605 8360 635
rect 8160 600 8360 605
rect 8480 635 8680 640
rect 8480 605 8490 635
rect 8670 605 8680 635
rect 8480 600 8680 605
rect 8080 285 8085 315
rect 8115 285 8120 315
rect 8080 280 8120 285
rect 8240 315 8280 600
rect 8240 285 8245 315
rect 8275 285 8280 315
rect 8240 280 8280 285
rect 8560 315 8600 600
rect 8560 285 8565 315
rect 8595 285 8600 315
rect 8560 280 8600 285
rect 8720 315 8760 670
rect 9040 750 9080 765
rect 9680 795 9720 800
rect 9680 765 9685 795
rect 9715 765 9720 795
rect 9040 670 9045 750
rect 9075 670 9080 750
rect 9040 660 9080 670
rect 9360 750 9400 760
rect 9360 670 9365 750
rect 9395 670 9400 750
rect 8800 635 9000 640
rect 8800 605 8810 635
rect 8990 605 9000 635
rect 8800 600 9000 605
rect 9120 635 9320 640
rect 9120 605 9130 635
rect 9310 605 9320 635
rect 9120 600 9320 605
rect 8720 285 8725 315
rect 8755 285 8760 315
rect 8720 280 8760 285
rect 8880 315 8920 600
rect 8880 285 8885 315
rect 8915 285 8920 315
rect 8880 280 8920 285
rect 9040 315 9080 320
rect 9040 285 9045 315
rect 9075 285 9080 315
rect 6560 155 6760 160
rect 6560 125 6570 155
rect 6750 125 6760 155
rect 6560 120 6760 125
rect 6880 155 7080 160
rect 6880 125 6890 155
rect 7070 125 7080 155
rect 6880 120 7080 125
rect 7200 155 7400 160
rect 7200 125 7210 155
rect 7390 125 7400 155
rect 7200 120 7400 125
rect 7520 155 7720 160
rect 7520 125 7530 155
rect 7710 125 7720 155
rect 7520 120 7720 125
rect 7840 155 8040 160
rect 7840 125 7850 155
rect 8030 125 8040 155
rect 7840 120 8040 125
rect 8160 155 8360 160
rect 8160 125 8170 155
rect 8350 125 8360 155
rect 8160 120 8360 125
rect 8480 155 8680 160
rect 8480 125 8490 155
rect 8670 125 8680 155
rect 8480 120 8680 125
rect 8800 155 9000 160
rect 8800 125 8810 155
rect 8990 125 9000 155
rect 8800 120 9000 125
rect 6480 10 6485 90
rect 6515 10 6520 90
rect 6480 0 6520 10
rect 6800 90 6840 100
rect 6800 10 6805 90
rect 6835 10 6840 90
rect 6800 0 6840 10
rect 7120 90 7160 100
rect 7120 10 7125 90
rect 7155 10 7160 90
rect 7120 0 7160 10
rect 7440 90 7480 100
rect 7440 10 7445 90
rect 7475 10 7480 90
rect 7440 0 7480 10
rect 7760 90 7800 100
rect 7760 10 7765 90
rect 7795 10 7800 90
rect 5200 -35 5205 -5
rect 5235 -35 5240 -5
rect 5200 -40 5240 -35
rect 7760 -5 7800 10
rect 8080 90 8120 100
rect 8080 10 8085 90
rect 8115 10 8120 90
rect 8080 0 8120 10
rect 8400 90 8440 100
rect 8400 10 8405 90
rect 8435 10 8440 90
rect 8400 0 8440 10
rect 8720 90 8760 100
rect 8720 10 8725 90
rect 8755 10 8760 90
rect 8720 0 8760 10
rect 9040 90 9080 285
rect 9200 315 9240 600
rect 9200 285 9205 315
rect 9235 285 9240 315
rect 9200 280 9240 285
rect 9360 315 9400 670
rect 9680 750 9720 765
rect 10320 795 10360 800
rect 10320 765 10325 795
rect 10355 765 10360 795
rect 9680 670 9685 750
rect 9715 670 9720 750
rect 9680 660 9720 670
rect 10000 750 10040 760
rect 10000 670 10005 750
rect 10035 670 10040 750
rect 9440 635 9640 640
rect 9440 605 9450 635
rect 9630 605 9640 635
rect 9440 600 9640 605
rect 9760 635 9960 640
rect 9760 605 9770 635
rect 9950 605 9960 635
rect 9760 600 9960 605
rect 9360 285 9365 315
rect 9395 285 9400 315
rect 9360 280 9400 285
rect 9520 315 9560 600
rect 9520 285 9525 315
rect 9555 285 9560 315
rect 9520 280 9560 285
rect 9840 315 9880 600
rect 9840 285 9845 315
rect 9875 285 9880 315
rect 9840 280 9880 285
rect 10000 315 10040 670
rect 10320 750 10360 765
rect 10640 795 10680 800
rect 10640 765 10645 795
rect 10675 765 10680 795
rect 10640 760 10680 765
rect 10800 795 10840 800
rect 10800 765 10805 795
rect 10835 765 10840 795
rect 10800 760 10840 765
rect 10960 795 11000 800
rect 10960 765 10965 795
rect 10995 765 11000 795
rect 10960 760 11000 765
rect 10320 670 10325 750
rect 10355 670 10360 750
rect 10640 715 10680 720
rect 10640 685 10645 715
rect 10675 685 10680 715
rect 10640 680 10680 685
rect 10800 715 10840 720
rect 10800 685 10805 715
rect 10835 685 10840 715
rect 10800 680 10840 685
rect 10960 715 11000 720
rect 10960 685 10965 715
rect 10995 685 11000 715
rect 10960 680 11000 685
rect 10320 660 10360 670
rect 10080 635 10280 640
rect 10080 605 10090 635
rect 10270 605 10280 635
rect 10080 600 10280 605
rect 10640 635 10680 640
rect 10640 605 10645 635
rect 10675 605 10680 635
rect 10640 600 10680 605
rect 10800 635 10840 640
rect 10800 605 10805 635
rect 10835 605 10840 635
rect 10800 600 10840 605
rect 10960 635 11000 640
rect 10960 605 10965 635
rect 10995 605 11000 635
rect 10960 600 11000 605
rect 10000 285 10005 315
rect 10035 285 10040 315
rect 10000 280 10040 285
rect 10160 315 10200 600
rect 10640 555 10680 560
rect 10640 525 10645 555
rect 10675 525 10680 555
rect 10640 520 10680 525
rect 10800 555 10840 560
rect 10800 525 10805 555
rect 10835 525 10840 555
rect 10800 520 10840 525
rect 10960 555 11000 560
rect 10960 525 10965 555
rect 10995 525 11000 555
rect 10960 520 11000 525
rect 10640 475 10680 480
rect 10640 445 10645 475
rect 10675 445 10680 475
rect 10640 440 10680 445
rect 10800 475 10840 480
rect 10800 445 10805 475
rect 10835 445 10840 475
rect 10800 440 10840 445
rect 10960 475 11000 480
rect 10960 445 10965 475
rect 10995 445 11000 475
rect 10960 440 11000 445
rect 10640 395 10680 400
rect 10640 365 10645 395
rect 10675 365 10680 395
rect 10640 360 10680 365
rect 10800 395 10840 400
rect 10800 365 10805 395
rect 10835 365 10840 395
rect 10800 360 10840 365
rect 10960 395 11000 400
rect 10960 365 10965 395
rect 10995 365 11000 395
rect 10960 360 11000 365
rect 10160 285 10165 315
rect 10195 285 10200 315
rect 10160 280 10200 285
rect 10640 235 10680 240
rect 10640 205 10645 235
rect 10675 205 10680 235
rect 10640 200 10680 205
rect 10800 235 10840 240
rect 10800 205 10805 235
rect 10835 205 10840 235
rect 10800 200 10840 205
rect 10960 235 11000 240
rect 10960 205 10965 235
rect 10995 205 11000 235
rect 10960 200 11000 205
rect 9120 155 9320 160
rect 9120 125 9130 155
rect 9310 125 9320 155
rect 9120 120 9320 125
rect 9440 155 9640 160
rect 9440 125 9450 155
rect 9630 125 9640 155
rect 9440 120 9640 125
rect 9760 155 9960 160
rect 9760 125 9770 155
rect 9950 125 9960 155
rect 9760 120 9960 125
rect 10080 155 10280 160
rect 10080 125 10090 155
rect 10270 125 10280 155
rect 10080 120 10280 125
rect 10800 155 10840 160
rect 10800 125 10805 155
rect 10835 125 10840 155
rect 10800 120 10840 125
rect 10960 155 11000 160
rect 10960 125 10965 155
rect 10995 125 11000 155
rect 10960 120 11000 125
rect 9040 10 9045 90
rect 9075 10 9080 90
rect 9040 0 9080 10
rect 9360 90 9400 100
rect 9360 10 9365 90
rect 9395 10 9400 90
rect 9360 0 9400 10
rect 9680 90 9720 100
rect 9680 10 9685 90
rect 9715 10 9720 90
rect 9680 0 9720 10
rect 10000 90 10040 100
rect 10000 10 10005 90
rect 10035 10 10040 90
rect 10000 0 10040 10
rect 10320 90 10360 100
rect 10320 10 10325 90
rect 10355 10 10360 90
rect 10640 75 10680 80
rect 10640 45 10645 75
rect 10675 45 10680 75
rect 10640 40 10680 45
rect 10800 75 10840 80
rect 10800 45 10805 75
rect 10835 45 10840 75
rect 10800 40 10840 45
rect 10960 75 11000 80
rect 10960 45 10965 75
rect 10995 45 11000 75
rect 10960 40 11000 45
rect 7760 -35 7765 -5
rect 7795 -35 7800 -5
rect 7760 -40 7800 -35
rect 10320 -5 10360 10
rect 10320 -35 10325 -5
rect 10355 -35 10360 -5
rect 10320 -40 10360 -35
rect 10640 -5 10680 0
rect 10640 -35 10645 -5
rect 10675 -35 10680 -5
rect 10640 -40 10680 -35
rect 10800 -5 10840 0
rect 10800 -35 10805 -5
rect 10835 -35 10840 -5
rect 10800 -40 10840 -35
rect 10960 -5 11000 0
rect 10960 -35 10965 -5
rect 10995 -35 11000 -5
rect 10960 -40 11000 -35
rect -720 -85 -680 -80
rect -720 -115 -715 -85
rect -685 -115 -680 -85
rect -720 -120 -680 -115
rect -560 -85 -520 -80
rect -560 -115 -555 -85
rect -525 -115 -520 -85
rect -560 -120 -520 -115
rect -400 -85 -360 -80
rect -400 -115 -395 -85
rect -365 -115 -360 -85
rect -400 -120 -360 -115
rect 10640 -85 10680 -80
rect 10640 -115 10645 -85
rect 10675 -115 10680 -85
rect 10640 -120 10680 -115
rect 10800 -85 10840 -80
rect 10800 -115 10805 -85
rect 10835 -115 10840 -85
rect 10800 -120 10840 -115
rect 10960 -85 11000 -80
rect 10960 -115 10965 -85
rect 10995 -115 11000 -85
rect 10960 -120 11000 -115
rect -720 -165 -680 -160
rect -720 -195 -715 -165
rect -685 -195 -680 -165
rect -720 -200 -680 -195
rect -560 -165 -520 -160
rect -560 -195 -555 -165
rect -525 -195 -520 -165
rect -560 -200 -520 -195
rect -400 -165 -360 -160
rect -400 -195 -395 -165
rect -365 -195 -360 -165
rect -400 -200 -360 -195
rect 10640 -165 10680 -160
rect 10640 -195 10645 -165
rect 10675 -195 10680 -165
rect 10640 -200 10680 -195
rect 10800 -165 10840 -160
rect 10800 -195 10805 -165
rect 10835 -195 10840 -165
rect 10800 -200 10840 -195
rect 10960 -165 11000 -160
rect 10960 -195 10965 -165
rect 10995 -195 11000 -165
rect 10960 -200 11000 -195
rect -720 -245 -680 -240
rect -720 -275 -715 -245
rect -685 -275 -680 -245
rect -720 -280 -680 -275
rect -560 -245 -520 -240
rect -560 -275 -555 -245
rect -525 -275 -520 -245
rect -560 -280 -520 -275
rect -400 -245 -360 -240
rect -400 -275 -395 -245
rect -365 -275 -360 -245
rect -400 -280 -360 -275
rect -80 -245 -40 -240
rect -80 -275 -75 -245
rect -45 -275 -40 -245
rect -80 -290 -40 -275
rect 2480 -245 2520 -240
rect 2480 -275 2485 -245
rect 2515 -275 2520 -245
rect -720 -325 -680 -320
rect -720 -355 -715 -325
rect -685 -355 -680 -325
rect -720 -360 -680 -355
rect -560 -325 -520 -320
rect -560 -355 -555 -325
rect -525 -355 -520 -325
rect -560 -360 -520 -355
rect -400 -325 -360 -320
rect -400 -355 -395 -325
rect -365 -355 -360 -325
rect -400 -360 -360 -355
rect -80 -370 -75 -290
rect -45 -370 -40 -290
rect -80 -380 -40 -370
rect 240 -290 280 -280
rect 240 -370 245 -290
rect 275 -370 280 -290
rect 240 -380 280 -370
rect 560 -290 600 -280
rect 560 -370 565 -290
rect 595 -370 600 -290
rect 560 -380 600 -370
rect 880 -290 920 -280
rect 880 -370 885 -290
rect 915 -370 920 -290
rect 880 -380 920 -370
rect 1200 -290 1240 -280
rect 1200 -370 1205 -290
rect 1235 -370 1240 -290
rect -720 -405 -680 -400
rect -720 -435 -715 -405
rect -685 -435 -680 -405
rect -720 -440 -680 -435
rect -560 -405 -520 -400
rect -560 -435 -555 -405
rect -525 -435 -520 -405
rect -560 -440 -520 -435
rect -400 -405 -360 -400
rect -400 -435 -395 -405
rect -365 -435 -360 -405
rect -400 -440 -360 -435
rect 0 -405 200 -400
rect 0 -435 10 -405
rect 190 -435 200 -405
rect 0 -440 200 -435
rect 320 -405 520 -400
rect 320 -435 330 -405
rect 510 -435 520 -405
rect 320 -440 520 -435
rect 640 -405 840 -400
rect 640 -435 650 -405
rect 830 -435 840 -405
rect 640 -440 840 -435
rect 960 -405 1160 -400
rect 960 -435 970 -405
rect 1150 -435 1160 -405
rect 960 -440 1160 -435
rect -720 -485 -680 -480
rect -720 -515 -715 -485
rect -685 -515 -680 -485
rect -720 -520 -680 -515
rect -560 -485 -520 -480
rect -560 -515 -555 -485
rect -525 -515 -520 -485
rect -560 -520 -520 -515
rect -400 -485 -360 -480
rect -400 -515 -395 -485
rect -365 -515 -360 -485
rect -400 -520 -360 -515
rect -720 -565 -680 -560
rect -720 -595 -715 -565
rect -685 -595 -680 -565
rect -720 -600 -680 -595
rect -560 -565 -520 -560
rect -560 -595 -555 -565
rect -525 -595 -520 -565
rect -560 -600 -520 -595
rect -400 -565 -360 -560
rect -400 -595 -395 -565
rect -365 -595 -360 -565
rect -400 -600 -360 -595
rect 80 -565 120 -560
rect 80 -595 85 -565
rect 115 -595 120 -565
rect -720 -645 -680 -640
rect -720 -675 -715 -645
rect -685 -675 -680 -645
rect -720 -680 -680 -675
rect -560 -645 -520 -640
rect -560 -675 -555 -645
rect -525 -675 -520 -645
rect -560 -680 -520 -675
rect -400 -645 -360 -640
rect -400 -675 -395 -645
rect -365 -675 -360 -645
rect -400 -680 -360 -675
rect -720 -725 -680 -720
rect -720 -755 -715 -725
rect -685 -755 -680 -725
rect -720 -760 -680 -755
rect -560 -725 -520 -720
rect -560 -755 -555 -725
rect -525 -755 -520 -725
rect -560 -760 -520 -755
rect -720 -805 -680 -800
rect -720 -835 -715 -805
rect -685 -835 -680 -805
rect -720 -840 -680 -835
rect -560 -805 -520 -800
rect -560 -835 -555 -805
rect -525 -835 -520 -805
rect -560 -840 -520 -835
rect -400 -805 -360 -800
rect -400 -835 -395 -805
rect -365 -835 -360 -805
rect -400 -840 -360 -835
rect 80 -880 120 -595
rect 240 -565 280 -560
rect 240 -595 245 -565
rect 275 -595 280 -565
rect -720 -885 -680 -880
rect -720 -915 -715 -885
rect -685 -915 -680 -885
rect -720 -920 -680 -915
rect -560 -885 -520 -880
rect -560 -915 -555 -885
rect -525 -915 -520 -885
rect -560 -920 -520 -915
rect -400 -885 -360 -880
rect -400 -915 -395 -885
rect -365 -915 -360 -885
rect -400 -920 -360 -915
rect 0 -885 200 -880
rect 0 -915 10 -885
rect 190 -915 200 -885
rect 0 -920 200 -915
rect -80 -950 -40 -940
rect -80 -1030 -75 -950
rect -45 -1030 -40 -950
rect -80 -1045 -40 -1030
rect 240 -950 280 -595
rect 400 -565 440 -560
rect 400 -595 405 -565
rect 435 -595 440 -565
rect 400 -880 440 -595
rect 720 -565 760 -560
rect 720 -595 725 -565
rect 755 -595 760 -565
rect 720 -880 760 -595
rect 880 -565 920 -560
rect 880 -595 885 -565
rect 915 -595 920 -565
rect 320 -885 520 -880
rect 320 -915 330 -885
rect 510 -915 520 -885
rect 320 -920 520 -915
rect 640 -885 840 -880
rect 640 -915 650 -885
rect 830 -915 840 -885
rect 640 -920 840 -915
rect 240 -1030 245 -950
rect 275 -1030 280 -950
rect 240 -1040 280 -1030
rect 560 -950 600 -940
rect 560 -1030 565 -950
rect 595 -1030 600 -950
rect -80 -1075 -75 -1045
rect -45 -1075 -40 -1045
rect -80 -1080 -40 -1075
rect 560 -1045 600 -1030
rect 880 -950 920 -595
rect 1040 -565 1080 -560
rect 1040 -595 1045 -565
rect 1075 -595 1080 -565
rect 1040 -880 1080 -595
rect 1200 -565 1240 -370
rect 1520 -290 1560 -280
rect 1520 -370 1525 -290
rect 1555 -370 1560 -290
rect 1520 -380 1560 -370
rect 1840 -290 1880 -280
rect 1840 -370 1845 -290
rect 1875 -370 1880 -290
rect 1840 -380 1880 -370
rect 2160 -290 2200 -280
rect 2160 -370 2165 -290
rect 2195 -370 2200 -290
rect 2160 -380 2200 -370
rect 2480 -290 2520 -275
rect 5040 -245 5080 -240
rect 5040 -275 5045 -245
rect 5075 -275 5080 -245
rect 2480 -370 2485 -290
rect 2515 -370 2520 -290
rect 2480 -380 2520 -370
rect 2800 -290 2840 -280
rect 2800 -370 2805 -290
rect 2835 -370 2840 -290
rect 2800 -380 2840 -370
rect 3120 -290 3160 -280
rect 3120 -370 3125 -290
rect 3155 -370 3160 -290
rect 3120 -380 3160 -370
rect 3440 -290 3480 -280
rect 3440 -370 3445 -290
rect 3475 -370 3480 -290
rect 3440 -380 3480 -370
rect 3760 -290 3800 -280
rect 3760 -370 3765 -290
rect 3795 -370 3800 -290
rect 1280 -405 1480 -400
rect 1280 -435 1290 -405
rect 1470 -435 1480 -405
rect 1280 -440 1480 -435
rect 1600 -405 1800 -400
rect 1600 -435 1610 -405
rect 1790 -435 1800 -405
rect 1600 -440 1800 -435
rect 1920 -405 2120 -400
rect 1920 -435 1930 -405
rect 2110 -435 2120 -405
rect 1920 -440 2120 -435
rect 2240 -405 2440 -400
rect 2240 -435 2250 -405
rect 2430 -435 2440 -405
rect 2240 -440 2440 -435
rect 2560 -405 2760 -400
rect 2560 -435 2570 -405
rect 2750 -435 2760 -405
rect 2560 -440 2760 -435
rect 2880 -405 3080 -400
rect 2880 -435 2890 -405
rect 3070 -435 3080 -405
rect 2880 -440 3080 -435
rect 3200 -405 3400 -400
rect 3200 -435 3210 -405
rect 3390 -435 3400 -405
rect 3200 -440 3400 -435
rect 3520 -405 3720 -400
rect 3520 -435 3530 -405
rect 3710 -435 3720 -405
rect 3520 -440 3720 -435
rect 1200 -595 1205 -565
rect 1235 -595 1240 -565
rect 1200 -600 1240 -595
rect 1360 -565 1400 -560
rect 1360 -595 1365 -565
rect 1395 -595 1400 -565
rect 1360 -880 1400 -595
rect 1520 -565 1560 -560
rect 1520 -595 1525 -565
rect 1555 -595 1560 -565
rect 960 -885 1160 -880
rect 960 -915 970 -885
rect 1150 -915 1160 -885
rect 960 -920 1160 -915
rect 1280 -885 1480 -880
rect 1280 -915 1290 -885
rect 1470 -915 1480 -885
rect 1280 -920 1480 -915
rect 880 -1030 885 -950
rect 915 -1030 920 -950
rect 880 -1040 920 -1030
rect 1200 -950 1240 -940
rect 1200 -1030 1205 -950
rect 1235 -1030 1240 -950
rect 560 -1075 565 -1045
rect 595 -1075 600 -1045
rect 560 -1080 600 -1075
rect 1200 -1045 1240 -1030
rect 1520 -950 1560 -595
rect 1680 -565 1720 -560
rect 1680 -595 1685 -565
rect 1715 -595 1720 -565
rect 1680 -880 1720 -595
rect 2000 -565 2040 -560
rect 2000 -595 2005 -565
rect 2035 -595 2040 -565
rect 2000 -880 2040 -595
rect 2160 -565 2200 -560
rect 2160 -595 2165 -565
rect 2195 -595 2200 -565
rect 1600 -885 1800 -880
rect 1600 -915 1610 -885
rect 1790 -915 1800 -885
rect 1600 -920 1800 -915
rect 1920 -885 2120 -880
rect 1920 -915 1930 -885
rect 2110 -915 2120 -885
rect 1920 -920 2120 -915
rect 1520 -1030 1525 -950
rect 1555 -1030 1560 -950
rect 1520 -1040 1560 -1030
rect 1840 -950 1880 -940
rect 1840 -1030 1845 -950
rect 1875 -1030 1880 -950
rect 1200 -1075 1205 -1045
rect 1235 -1075 1240 -1045
rect 1200 -1080 1240 -1075
rect 1840 -1045 1880 -1030
rect 2160 -950 2200 -595
rect 2320 -565 2360 -560
rect 2320 -595 2325 -565
rect 2355 -595 2360 -565
rect 2320 -880 2360 -595
rect 2640 -565 2680 -560
rect 2640 -595 2645 -565
rect 2675 -595 2680 -565
rect 2640 -880 2680 -595
rect 2800 -565 2840 -560
rect 2800 -595 2805 -565
rect 2835 -595 2840 -565
rect 2240 -885 2440 -880
rect 2240 -915 2250 -885
rect 2430 -915 2440 -885
rect 2240 -920 2440 -915
rect 2560 -885 2760 -880
rect 2560 -915 2570 -885
rect 2750 -915 2760 -885
rect 2560 -920 2760 -915
rect 2160 -1030 2165 -950
rect 2195 -1030 2200 -950
rect 2160 -1040 2200 -1030
rect 2480 -950 2520 -940
rect 2480 -1030 2485 -950
rect 2515 -1030 2520 -950
rect 1840 -1075 1845 -1045
rect 1875 -1075 1880 -1045
rect 1840 -1080 1880 -1075
rect 2480 -1045 2520 -1030
rect 2800 -950 2840 -595
rect 2960 -565 3000 -560
rect 2960 -595 2965 -565
rect 2995 -595 3000 -565
rect 2960 -880 3000 -595
rect 3280 -565 3320 -560
rect 3280 -595 3285 -565
rect 3315 -595 3320 -565
rect 3280 -880 3320 -595
rect 3440 -565 3480 -560
rect 3440 -595 3445 -565
rect 3475 -595 3480 -565
rect 2880 -885 3080 -880
rect 2880 -915 2890 -885
rect 3070 -915 3080 -885
rect 2880 -920 3080 -915
rect 3200 -885 3400 -880
rect 3200 -915 3210 -885
rect 3390 -915 3400 -885
rect 3200 -920 3400 -915
rect 2800 -1030 2805 -950
rect 2835 -1030 2840 -950
rect 2800 -1040 2840 -1030
rect 3120 -950 3160 -940
rect 3120 -1030 3125 -950
rect 3155 -1030 3160 -950
rect 2480 -1075 2485 -1045
rect 2515 -1075 2520 -1045
rect 2480 -1080 2520 -1075
rect 3120 -1045 3160 -1030
rect 3440 -950 3480 -595
rect 3600 -565 3640 -560
rect 3600 -595 3605 -565
rect 3635 -595 3640 -565
rect 3600 -880 3640 -595
rect 3760 -565 3800 -370
rect 4080 -290 4120 -280
rect 4080 -370 4085 -290
rect 4115 -370 4120 -290
rect 4080 -380 4120 -370
rect 4400 -290 4440 -280
rect 4400 -370 4405 -290
rect 4435 -370 4440 -290
rect 4400 -380 4440 -370
rect 4720 -290 4760 -280
rect 4720 -370 4725 -290
rect 4755 -370 4760 -290
rect 4720 -380 4760 -370
rect 5040 -290 5080 -275
rect 5040 -370 5045 -290
rect 5075 -370 5080 -290
rect 5040 -380 5080 -370
rect 5200 -245 5240 -240
rect 5200 -275 5205 -245
rect 5235 -275 5240 -245
rect 5200 -290 5240 -275
rect 7760 -245 7800 -240
rect 7760 -275 7765 -245
rect 7795 -275 7800 -245
rect 5200 -370 5205 -290
rect 5235 -370 5240 -290
rect 5200 -380 5240 -370
rect 5520 -290 5560 -280
rect 5520 -370 5525 -290
rect 5555 -370 5560 -290
rect 5520 -380 5560 -370
rect 5840 -290 5880 -280
rect 5840 -370 5845 -290
rect 5875 -370 5880 -290
rect 5840 -380 5880 -370
rect 6160 -290 6200 -280
rect 6160 -370 6165 -290
rect 6195 -370 6200 -290
rect 6160 -380 6200 -370
rect 6480 -290 6520 -280
rect 6480 -370 6485 -290
rect 6515 -370 6520 -290
rect 3840 -405 4040 -400
rect 3840 -435 3850 -405
rect 4030 -435 4040 -405
rect 3840 -440 4040 -435
rect 4160 -405 4360 -400
rect 4160 -435 4170 -405
rect 4350 -435 4360 -405
rect 4160 -440 4360 -435
rect 4480 -405 4680 -400
rect 4480 -435 4490 -405
rect 4670 -435 4680 -405
rect 4480 -440 4680 -435
rect 4800 -405 5000 -400
rect 4800 -435 4810 -405
rect 4990 -435 5000 -405
rect 4800 -440 5000 -435
rect 5200 -405 5240 -400
rect 5200 -435 5205 -405
rect 5235 -435 5240 -405
rect 3760 -595 3765 -565
rect 3795 -595 3800 -565
rect 3760 -600 3800 -595
rect 3920 -565 3960 -560
rect 3920 -595 3925 -565
rect 3955 -595 3960 -565
rect 3920 -880 3960 -595
rect 4080 -565 4120 -560
rect 4080 -595 4085 -565
rect 4115 -595 4120 -565
rect 3520 -885 3720 -880
rect 3520 -915 3530 -885
rect 3710 -915 3720 -885
rect 3520 -920 3720 -915
rect 3840 -885 4040 -880
rect 3840 -915 3850 -885
rect 4030 -915 4040 -885
rect 3840 -920 4040 -915
rect 3440 -1030 3445 -950
rect 3475 -1030 3480 -950
rect 3440 -1040 3480 -1030
rect 3760 -950 3800 -940
rect 3760 -1030 3765 -950
rect 3795 -1030 3800 -950
rect 3120 -1075 3125 -1045
rect 3155 -1075 3160 -1045
rect 3120 -1080 3160 -1075
rect 3760 -1045 3800 -1030
rect 4080 -950 4120 -595
rect 4240 -565 4280 -560
rect 4240 -595 4245 -565
rect 4275 -595 4280 -565
rect 4240 -880 4280 -595
rect 4560 -565 4600 -560
rect 4560 -595 4565 -565
rect 4595 -595 4600 -565
rect 4560 -880 4600 -595
rect 4720 -565 4760 -560
rect 4720 -595 4725 -565
rect 4755 -595 4760 -565
rect 4160 -885 4360 -880
rect 4160 -915 4170 -885
rect 4350 -915 4360 -885
rect 4160 -920 4360 -915
rect 4480 -885 4680 -880
rect 4480 -915 4490 -885
rect 4670 -915 4680 -885
rect 4480 -920 4680 -915
rect 4080 -1030 4085 -950
rect 4115 -1030 4120 -950
rect 4080 -1040 4120 -1030
rect 4400 -950 4440 -940
rect 4400 -1030 4405 -950
rect 4435 -1030 4440 -950
rect 3760 -1075 3765 -1045
rect 3795 -1075 3800 -1045
rect 3760 -1080 3800 -1075
rect 4400 -1045 4440 -1030
rect 4720 -950 4760 -595
rect 4880 -565 4920 -560
rect 4880 -595 4885 -565
rect 4915 -595 4920 -565
rect 4880 -880 4920 -595
rect 4800 -885 5000 -880
rect 4800 -915 4810 -885
rect 4990 -915 5000 -885
rect 4800 -920 5000 -915
rect 4720 -1030 4725 -950
rect 4755 -1030 4760 -950
rect 4720 -1040 4760 -1030
rect 5040 -950 5080 -940
rect 5040 -1030 5045 -950
rect 5075 -1030 5080 -950
rect 4400 -1075 4405 -1045
rect 4435 -1075 4440 -1045
rect 4400 -1080 4440 -1075
rect 5040 -1045 5080 -1030
rect 5200 -950 5240 -435
rect 5280 -405 5480 -400
rect 5280 -435 5290 -405
rect 5470 -435 5480 -405
rect 5280 -440 5480 -435
rect 5600 -405 5800 -400
rect 5600 -435 5610 -405
rect 5790 -435 5800 -405
rect 5600 -440 5800 -435
rect 5920 -405 6120 -400
rect 5920 -435 5930 -405
rect 6110 -435 6120 -405
rect 5920 -440 6120 -435
rect 6240 -405 6440 -400
rect 6240 -435 6250 -405
rect 6430 -435 6440 -405
rect 6240 -440 6440 -435
rect 6480 -405 6520 -370
rect 6800 -290 6840 -280
rect 6800 -370 6805 -290
rect 6835 -370 6840 -290
rect 6800 -380 6840 -370
rect 7120 -290 7160 -280
rect 7120 -370 7125 -290
rect 7155 -370 7160 -290
rect 7120 -380 7160 -370
rect 7440 -290 7480 -280
rect 7440 -370 7445 -290
rect 7475 -370 7480 -290
rect 7440 -380 7480 -370
rect 7760 -290 7800 -275
rect 10320 -245 10360 -240
rect 10320 -275 10325 -245
rect 10355 -275 10360 -245
rect 7760 -370 7765 -290
rect 7795 -370 7800 -290
rect 7760 -380 7800 -370
rect 8080 -290 8120 -280
rect 8080 -370 8085 -290
rect 8115 -370 8120 -290
rect 8080 -380 8120 -370
rect 8400 -290 8440 -280
rect 8400 -370 8405 -290
rect 8435 -370 8440 -290
rect 8400 -380 8440 -370
rect 8720 -290 8760 -280
rect 8720 -370 8725 -290
rect 8755 -370 8760 -290
rect 8720 -380 8760 -370
rect 9040 -290 9080 -280
rect 9040 -370 9045 -290
rect 9075 -370 9080 -290
rect 6480 -435 6485 -405
rect 6515 -435 6520 -405
rect 6480 -440 6520 -435
rect 6560 -405 6760 -400
rect 6560 -435 6570 -405
rect 6750 -435 6760 -405
rect 6560 -440 6760 -435
rect 6880 -405 7080 -400
rect 6880 -435 6890 -405
rect 7070 -435 7080 -405
rect 6880 -440 7080 -435
rect 7200 -405 7400 -400
rect 7200 -435 7210 -405
rect 7390 -435 7400 -405
rect 7200 -440 7400 -435
rect 7520 -405 7720 -400
rect 7520 -435 7530 -405
rect 7710 -435 7720 -405
rect 7520 -440 7720 -435
rect 7840 -405 8040 -400
rect 7840 -435 7850 -405
rect 8030 -435 8040 -405
rect 7840 -440 8040 -435
rect 8160 -405 8360 -400
rect 8160 -435 8170 -405
rect 8350 -435 8360 -405
rect 8160 -440 8360 -435
rect 8480 -405 8680 -400
rect 8480 -435 8490 -405
rect 8670 -435 8680 -405
rect 8480 -440 8680 -435
rect 8800 -405 9000 -400
rect 8800 -435 8810 -405
rect 8990 -435 9000 -405
rect 8800 -440 9000 -435
rect 9040 -405 9080 -370
rect 9360 -290 9400 -280
rect 9360 -370 9365 -290
rect 9395 -370 9400 -290
rect 9360 -380 9400 -370
rect 9680 -290 9720 -280
rect 9680 -370 9685 -290
rect 9715 -370 9720 -290
rect 9680 -380 9720 -370
rect 10000 -290 10040 -280
rect 10000 -370 10005 -290
rect 10035 -370 10040 -290
rect 10000 -380 10040 -370
rect 10320 -290 10360 -275
rect 10640 -245 10680 -240
rect 10640 -275 10645 -245
rect 10675 -275 10680 -245
rect 10640 -280 10680 -275
rect 10800 -245 10840 -240
rect 10800 -275 10805 -245
rect 10835 -275 10840 -245
rect 10800 -280 10840 -275
rect 10960 -245 11000 -240
rect 10960 -275 10965 -245
rect 10995 -275 11000 -245
rect 10960 -280 11000 -275
rect 10320 -370 10325 -290
rect 10355 -370 10360 -290
rect 10640 -325 10680 -320
rect 10640 -355 10645 -325
rect 10675 -355 10680 -325
rect 10640 -360 10680 -355
rect 10800 -325 10840 -320
rect 10800 -355 10805 -325
rect 10835 -355 10840 -325
rect 10800 -360 10840 -355
rect 10960 -325 11000 -320
rect 10960 -355 10965 -325
rect 10995 -355 11000 -325
rect 10960 -360 11000 -355
rect 10320 -380 10360 -370
rect 9040 -435 9045 -405
rect 9075 -435 9080 -405
rect 9040 -440 9080 -435
rect 9120 -405 9320 -400
rect 9120 -435 9130 -405
rect 9310 -435 9320 -405
rect 9120 -440 9320 -435
rect 9440 -405 9640 -400
rect 9440 -435 9450 -405
rect 9630 -435 9640 -405
rect 9440 -440 9640 -435
rect 9760 -405 9960 -400
rect 9760 -435 9770 -405
rect 9950 -435 9960 -405
rect 9760 -440 9960 -435
rect 10080 -405 10280 -400
rect 10080 -435 10090 -405
rect 10270 -435 10280 -405
rect 10080 -440 10280 -435
rect 10800 -405 10840 -400
rect 10800 -435 10805 -405
rect 10835 -435 10840 -405
rect 10800 -440 10840 -435
rect 10960 -405 11000 -400
rect 10960 -435 10965 -405
rect 10995 -435 11000 -405
rect 10960 -440 11000 -435
rect 10640 -485 10680 -480
rect 10640 -515 10645 -485
rect 10675 -515 10680 -485
rect 10640 -520 10680 -515
rect 10800 -485 10840 -480
rect 10800 -515 10805 -485
rect 10835 -515 10840 -485
rect 10800 -520 10840 -515
rect 10960 -485 11000 -480
rect 10960 -515 10965 -485
rect 10995 -515 11000 -485
rect 10960 -520 11000 -515
rect 10640 -645 10680 -640
rect 10640 -675 10645 -645
rect 10675 -675 10680 -645
rect 10640 -680 10680 -675
rect 10800 -645 10840 -640
rect 10800 -675 10805 -645
rect 10835 -675 10840 -645
rect 10800 -680 10840 -675
rect 10960 -645 11000 -640
rect 10960 -675 10965 -645
rect 10995 -675 11000 -645
rect 10960 -680 11000 -675
rect 5360 -725 5400 -720
rect 5360 -755 5365 -725
rect 5395 -755 5400 -725
rect 5360 -880 5400 -755
rect 5680 -725 5720 -720
rect 5680 -755 5685 -725
rect 5715 -755 5720 -725
rect 5680 -880 5720 -755
rect 6000 -725 6040 -720
rect 6000 -755 6005 -725
rect 6035 -755 6040 -725
rect 6000 -880 6040 -755
rect 6320 -725 6360 -720
rect 6320 -755 6325 -725
rect 6355 -755 6360 -725
rect 6320 -880 6360 -755
rect 6640 -725 6680 -720
rect 6640 -755 6645 -725
rect 6675 -755 6680 -725
rect 6640 -880 6680 -755
rect 6960 -725 7000 -720
rect 6960 -755 6965 -725
rect 6995 -755 7000 -725
rect 6960 -880 7000 -755
rect 7280 -725 7320 -720
rect 7280 -755 7285 -725
rect 7315 -755 7320 -725
rect 7280 -880 7320 -755
rect 7600 -725 7640 -720
rect 7600 -755 7605 -725
rect 7635 -755 7640 -725
rect 7600 -880 7640 -755
rect 7920 -725 7960 -720
rect 7920 -755 7925 -725
rect 7955 -755 7960 -725
rect 7920 -880 7960 -755
rect 8240 -725 8280 -720
rect 8240 -755 8245 -725
rect 8275 -755 8280 -725
rect 8240 -880 8280 -755
rect 8560 -725 8600 -720
rect 8560 -755 8565 -725
rect 8595 -755 8600 -725
rect 8560 -880 8600 -755
rect 8880 -725 8920 -720
rect 8880 -755 8885 -725
rect 8915 -755 8920 -725
rect 8880 -880 8920 -755
rect 9200 -725 9240 -720
rect 9200 -755 9205 -725
rect 9235 -755 9240 -725
rect 9200 -880 9240 -755
rect 9520 -725 9560 -720
rect 9520 -755 9525 -725
rect 9555 -755 9560 -725
rect 9520 -880 9560 -755
rect 9840 -725 9880 -720
rect 9840 -755 9845 -725
rect 9875 -755 9880 -725
rect 9840 -880 9880 -755
rect 10160 -725 10200 -720
rect 10160 -755 10165 -725
rect 10195 -755 10200 -725
rect 10160 -880 10200 -755
rect 10640 -725 10680 -720
rect 10640 -755 10645 -725
rect 10675 -755 10680 -725
rect 10640 -760 10680 -755
rect 10800 -725 10840 -720
rect 10800 -755 10805 -725
rect 10835 -755 10840 -725
rect 10800 -760 10840 -755
rect 10960 -725 11000 -720
rect 10960 -755 10965 -725
rect 10995 -755 11000 -725
rect 10960 -760 11000 -755
rect 10640 -805 10680 -800
rect 10640 -835 10645 -805
rect 10675 -835 10680 -805
rect 10640 -840 10680 -835
rect 10800 -805 10840 -800
rect 10800 -835 10805 -805
rect 10835 -835 10840 -805
rect 10800 -840 10840 -835
rect 10960 -805 11000 -800
rect 10960 -835 10965 -805
rect 10995 -835 11000 -805
rect 10960 -840 11000 -835
rect 5280 -885 5480 -880
rect 5280 -915 5290 -885
rect 5470 -915 5480 -885
rect 5280 -920 5480 -915
rect 5600 -885 5800 -880
rect 5600 -915 5610 -885
rect 5790 -915 5800 -885
rect 5600 -920 5800 -915
rect 5920 -885 6120 -880
rect 5920 -915 5930 -885
rect 6110 -915 6120 -885
rect 5920 -920 6120 -915
rect 6240 -885 6440 -880
rect 6240 -915 6250 -885
rect 6430 -915 6440 -885
rect 6240 -920 6440 -915
rect 6560 -885 6760 -880
rect 6560 -915 6570 -885
rect 6750 -915 6760 -885
rect 6560 -920 6760 -915
rect 6880 -885 7080 -880
rect 6880 -915 6890 -885
rect 7070 -915 7080 -885
rect 6880 -920 7080 -915
rect 7200 -885 7400 -880
rect 7200 -915 7210 -885
rect 7390 -915 7400 -885
rect 7200 -920 7400 -915
rect 7520 -885 7720 -880
rect 7520 -915 7530 -885
rect 7710 -915 7720 -885
rect 7520 -920 7720 -915
rect 7840 -885 8040 -880
rect 7840 -915 7850 -885
rect 8030 -915 8040 -885
rect 7840 -920 8040 -915
rect 8160 -885 8360 -880
rect 8160 -915 8170 -885
rect 8350 -915 8360 -885
rect 8160 -920 8360 -915
rect 8480 -885 8680 -880
rect 8480 -915 8490 -885
rect 8670 -915 8680 -885
rect 8480 -920 8680 -915
rect 8800 -885 9000 -880
rect 8800 -915 8810 -885
rect 8990 -915 9000 -885
rect 8800 -920 9000 -915
rect 9120 -885 9320 -880
rect 9120 -915 9130 -885
rect 9310 -915 9320 -885
rect 9120 -920 9320 -915
rect 9440 -885 9640 -880
rect 9440 -915 9450 -885
rect 9630 -915 9640 -885
rect 9440 -920 9640 -915
rect 9760 -885 9960 -880
rect 9760 -915 9770 -885
rect 9950 -915 9960 -885
rect 9760 -920 9960 -915
rect 10080 -885 10280 -880
rect 10080 -915 10090 -885
rect 10270 -915 10280 -885
rect 10080 -920 10280 -915
rect 10640 -885 10680 -880
rect 10640 -915 10645 -885
rect 10675 -915 10680 -885
rect 10640 -920 10680 -915
rect 10800 -885 10840 -880
rect 10800 -915 10805 -885
rect 10835 -915 10840 -885
rect 10800 -920 10840 -915
rect 10960 -885 11000 -880
rect 10960 -915 10965 -885
rect 10995 -915 11000 -885
rect 10960 -920 11000 -915
rect 5200 -1030 5205 -950
rect 5235 -1030 5240 -950
rect 5200 -1040 5240 -1030
rect 5520 -950 5560 -940
rect 5520 -1030 5525 -950
rect 5555 -1030 5560 -950
rect 5520 -1040 5560 -1030
rect 5840 -950 5880 -940
rect 5840 -1030 5845 -950
rect 5875 -1030 5880 -950
rect 5840 -1040 5880 -1030
rect 6160 -950 6200 -940
rect 6160 -1030 6165 -950
rect 6195 -1030 6200 -950
rect 6160 -1040 6200 -1030
rect 6480 -950 6520 -940
rect 6480 -1030 6485 -950
rect 6515 -1030 6520 -950
rect 6480 -1040 6520 -1030
rect 6800 -950 6840 -940
rect 6800 -1030 6805 -950
rect 6835 -1030 6840 -950
rect 6800 -1040 6840 -1030
rect 7120 -950 7160 -940
rect 7120 -1030 7125 -950
rect 7155 -1030 7160 -950
rect 7120 -1040 7160 -1030
rect 7440 -950 7480 -940
rect 7440 -1030 7445 -950
rect 7475 -1030 7480 -950
rect 7440 -1040 7480 -1030
rect 7760 -950 7800 -940
rect 7760 -1030 7765 -950
rect 7795 -1030 7800 -950
rect 7760 -1040 7800 -1030
rect 8080 -950 8120 -940
rect 8080 -1030 8085 -950
rect 8115 -1030 8120 -950
rect 8080 -1040 8120 -1030
rect 8400 -950 8440 -940
rect 8400 -1030 8405 -950
rect 8435 -1030 8440 -950
rect 8400 -1040 8440 -1030
rect 8720 -950 8760 -940
rect 8720 -1030 8725 -950
rect 8755 -1030 8760 -950
rect 8720 -1040 8760 -1030
rect 9040 -950 9080 -940
rect 9040 -1030 9045 -950
rect 9075 -1030 9080 -950
rect 9040 -1040 9080 -1030
rect 9360 -950 9400 -940
rect 9360 -1030 9365 -950
rect 9395 -1030 9400 -950
rect 9360 -1040 9400 -1030
rect 9680 -950 9720 -940
rect 9680 -1030 9685 -950
rect 9715 -1030 9720 -950
rect 9680 -1040 9720 -1030
rect 10000 -950 10040 -940
rect 10000 -1030 10005 -950
rect 10035 -1030 10040 -950
rect 10000 -1040 10040 -1030
rect 10320 -950 10360 -940
rect 10320 -1030 10325 -950
rect 10355 -1030 10360 -950
rect 10640 -965 10680 -960
rect 10640 -995 10645 -965
rect 10675 -995 10680 -965
rect 10640 -1000 10680 -995
rect 10800 -965 10840 -960
rect 10800 -995 10805 -965
rect 10835 -995 10840 -965
rect 10800 -1000 10840 -995
rect 10960 -965 11000 -960
rect 10960 -995 10965 -965
rect 10995 -995 11000 -965
rect 10960 -1000 11000 -995
rect 5040 -1075 5045 -1045
rect 5075 -1075 5080 -1045
rect 5040 -1080 5080 -1075
rect 10320 -1045 10360 -1030
rect 10320 -1075 10325 -1045
rect 10355 -1075 10360 -1045
rect 10320 -1080 10360 -1075
rect 10640 -1045 10680 -1040
rect 10640 -1075 10645 -1045
rect 10675 -1075 10680 -1045
rect 10640 -1080 10680 -1075
rect 10800 -1045 10840 -1040
rect 10800 -1075 10805 -1045
rect 10835 -1075 10840 -1045
rect 10800 -1080 10840 -1075
rect 10960 -1045 11000 -1040
rect 10960 -1075 10965 -1045
rect 10995 -1075 11000 -1045
rect 10960 -1080 11000 -1075
rect -720 -1125 -680 -1120
rect -720 -1155 -715 -1125
rect -685 -1155 -680 -1125
rect -720 -1160 -680 -1155
rect -560 -1125 -520 -1120
rect -560 -1155 -555 -1125
rect -525 -1155 -520 -1125
rect -560 -1160 -520 -1155
rect -400 -1125 -360 -1120
rect -400 -1155 -395 -1125
rect -365 -1155 -360 -1125
rect -400 -1160 -360 -1155
rect 10640 -1125 10680 -1120
rect 10640 -1155 10645 -1125
rect 10675 -1155 10680 -1125
rect 10640 -1160 10680 -1155
rect 10800 -1125 10840 -1120
rect 10800 -1155 10805 -1125
rect 10835 -1155 10840 -1125
rect 10800 -1160 10840 -1155
rect 10960 -1125 11000 -1120
rect 10960 -1155 10965 -1125
rect 10995 -1155 11000 -1125
rect 10960 -1160 11000 -1155
rect -720 -1205 -680 -1200
rect -720 -1235 -715 -1205
rect -685 -1235 -680 -1205
rect -720 -1240 -680 -1235
rect -560 -1205 -520 -1200
rect -560 -1235 -555 -1205
rect -525 -1235 -520 -1205
rect -560 -1240 -520 -1235
rect -400 -1205 -360 -1200
rect -400 -1235 -395 -1205
rect -365 -1235 -360 -1205
rect -400 -1240 -360 -1235
rect 10640 -1205 10680 -1200
rect 10640 -1235 10645 -1205
rect 10675 -1235 10680 -1205
rect 10640 -1240 10680 -1235
rect 10800 -1205 10840 -1200
rect 10800 -1235 10805 -1205
rect 10835 -1235 10840 -1205
rect 10800 -1240 10840 -1235
rect 10960 -1205 11000 -1200
rect 10960 -1235 10965 -1205
rect 10995 -1235 11000 -1205
rect 10960 -1240 11000 -1235
rect -720 -1285 -680 -1280
rect -720 -1315 -715 -1285
rect -685 -1315 -680 -1285
rect -720 -1320 -680 -1315
rect -560 -1285 -520 -1280
rect -560 -1315 -555 -1285
rect -525 -1315 -520 -1285
rect -560 -1320 -520 -1315
rect -400 -1285 -360 -1280
rect -400 -1315 -395 -1285
rect -365 -1315 -360 -1285
rect -400 -1320 -360 -1315
rect 10640 -1285 10680 -1280
rect 10640 -1315 10645 -1285
rect 10675 -1315 10680 -1285
rect 10640 -1320 10680 -1315
rect 10800 -1285 10840 -1280
rect 10800 -1315 10805 -1285
rect 10835 -1315 10840 -1285
rect 10800 -1320 10840 -1315
rect 10960 -1285 11000 -1280
rect 10960 -1315 10965 -1285
rect 10995 -1315 11000 -1285
rect 10960 -1320 11000 -1315
rect -720 -1365 -680 -1360
rect -720 -1395 -715 -1365
rect -685 -1395 -680 -1365
rect -720 -1400 -680 -1395
rect -560 -1365 -520 -1360
rect -560 -1395 -555 -1365
rect -525 -1395 -520 -1365
rect -560 -1400 -520 -1395
rect -400 -1365 -360 -1360
rect -400 -1395 -395 -1365
rect -365 -1395 -360 -1365
rect -400 -1400 -360 -1395
rect 10640 -1365 10680 -1360
rect 10640 -1395 10645 -1365
rect 10675 -1395 10680 -1365
rect 10640 -1400 10680 -1395
rect 10800 -1365 10840 -1360
rect 10800 -1395 10805 -1365
rect 10835 -1395 10840 -1365
rect 10800 -1400 10840 -1395
rect 10960 -1365 11000 -1360
rect 10960 -1395 10965 -1365
rect 10995 -1395 11000 -1365
rect 10960 -1400 11000 -1395
rect -720 -1445 -680 -1440
rect -720 -1475 -715 -1445
rect -685 -1475 -680 -1445
rect -720 -1480 -680 -1475
rect -560 -1445 -520 -1440
rect -560 -1475 -555 -1445
rect -525 -1475 -520 -1445
rect -560 -1480 -520 -1475
rect -400 -1445 -360 -1440
rect -400 -1475 -395 -1445
rect -365 -1475 -360 -1445
rect -400 -1480 -360 -1475
rect 10640 -1445 10680 -1440
rect 10640 -1475 10645 -1445
rect 10675 -1475 10680 -1445
rect 10640 -1480 10680 -1475
rect 10800 -1445 10840 -1440
rect 10800 -1475 10805 -1445
rect 10835 -1475 10840 -1445
rect 10800 -1480 10840 -1475
rect 10960 -1445 11000 -1440
rect 10960 -1475 10965 -1445
rect 10995 -1475 11000 -1445
rect 10960 -1480 11000 -1475
rect -720 -1525 -680 -1520
rect -720 -1555 -715 -1525
rect -685 -1555 -680 -1525
rect -720 -1560 -680 -1555
rect -560 -1525 -520 -1520
rect -560 -1555 -555 -1525
rect -525 -1555 -520 -1525
rect -560 -1560 -520 -1555
rect -400 -1525 -360 -1520
rect -400 -1555 -395 -1525
rect -365 -1555 -360 -1525
rect -400 -1560 -360 -1555
rect 10640 -1525 10680 -1520
rect 10640 -1555 10645 -1525
rect 10675 -1555 10680 -1525
rect 10640 -1560 10680 -1555
rect 10800 -1525 10840 -1520
rect 10800 -1555 10805 -1525
rect 10835 -1555 10840 -1525
rect 10800 -1560 10840 -1555
rect 10960 -1525 11000 -1520
rect 10960 -1555 10965 -1525
rect 10995 -1555 11000 -1525
rect 10960 -1560 11000 -1555
rect -80 -1605 -40 -1600
rect -80 -1635 -75 -1605
rect -45 -1635 -40 -1605
rect -80 -1650 -40 -1635
rect 560 -1605 600 -1600
rect 560 -1635 565 -1605
rect 595 -1635 600 -1605
rect -80 -1730 -75 -1650
rect -45 -1730 -40 -1650
rect -80 -1740 -40 -1730
rect 240 -1650 280 -1640
rect 240 -1730 245 -1650
rect 275 -1730 280 -1650
rect -720 -1765 -680 -1760
rect -720 -1795 -715 -1765
rect -685 -1795 -680 -1765
rect -720 -1800 -680 -1795
rect -560 -1765 -520 -1760
rect -560 -1795 -555 -1765
rect -525 -1795 -520 -1765
rect -560 -1800 -520 -1795
rect -400 -1765 -360 -1760
rect -400 -1795 -395 -1765
rect -365 -1795 -360 -1765
rect -400 -1800 -360 -1795
rect 0 -1765 200 -1760
rect 0 -1795 10 -1765
rect 190 -1795 200 -1765
rect 0 -1800 200 -1795
rect -720 -1845 -680 -1840
rect -720 -1875 -715 -1845
rect -685 -1875 -680 -1845
rect -720 -1880 -680 -1875
rect -560 -1845 -520 -1840
rect -560 -1875 -555 -1845
rect -525 -1875 -520 -1845
rect -560 -1880 -520 -1875
rect -400 -1845 -360 -1840
rect -400 -1875 -395 -1845
rect -365 -1875 -360 -1845
rect -400 -1880 -360 -1875
rect -720 -1925 -680 -1920
rect -720 -1955 -715 -1925
rect -685 -1955 -680 -1925
rect -720 -1960 -680 -1955
rect -560 -1925 -520 -1920
rect -560 -1955 -555 -1925
rect -525 -1955 -520 -1925
rect -560 -1960 -520 -1955
rect -720 -2005 -680 -2000
rect -720 -2035 -715 -2005
rect -685 -2035 -680 -2005
rect -720 -2040 -680 -2035
rect -560 -2005 -520 -2000
rect -560 -2035 -555 -2005
rect -525 -2035 -520 -2005
rect -560 -2040 -520 -2035
rect -400 -2005 -360 -2000
rect -400 -2035 -395 -2005
rect -365 -2035 -360 -2005
rect -400 -2040 -360 -2035
rect -720 -2085 -680 -2080
rect -720 -2115 -715 -2085
rect -685 -2115 -680 -2085
rect -720 -2120 -680 -2115
rect -560 -2085 -520 -2080
rect -560 -2115 -555 -2085
rect -525 -2115 -520 -2085
rect -560 -2120 -520 -2115
rect -400 -2085 -360 -2080
rect -400 -2115 -395 -2085
rect -365 -2115 -360 -2085
rect -400 -2120 -360 -2115
rect 80 -2085 120 -1800
rect 80 -2115 85 -2085
rect 115 -2115 120 -2085
rect 80 -2120 120 -2115
rect 240 -2085 280 -1730
rect 560 -1650 600 -1635
rect 1200 -1605 1240 -1600
rect 1200 -1635 1205 -1605
rect 1235 -1635 1240 -1605
rect 560 -1730 565 -1650
rect 595 -1730 600 -1650
rect 560 -1740 600 -1730
rect 880 -1650 920 -1640
rect 880 -1730 885 -1650
rect 915 -1730 920 -1650
rect 320 -1765 520 -1760
rect 320 -1795 330 -1765
rect 510 -1795 520 -1765
rect 320 -1800 520 -1795
rect 640 -1765 840 -1760
rect 640 -1795 650 -1765
rect 830 -1795 840 -1765
rect 640 -1800 840 -1795
rect 240 -2115 245 -2085
rect 275 -2115 280 -2085
rect 240 -2120 280 -2115
rect 400 -2085 440 -1800
rect 400 -2115 405 -2085
rect 435 -2115 440 -2085
rect 400 -2120 440 -2115
rect 720 -2085 760 -1800
rect 720 -2115 725 -2085
rect 755 -2115 760 -2085
rect 720 -2120 760 -2115
rect 880 -2085 920 -1730
rect 1200 -1650 1240 -1635
rect 1840 -1605 1880 -1600
rect 1840 -1635 1845 -1605
rect 1875 -1635 1880 -1605
rect 1200 -1730 1205 -1650
rect 1235 -1730 1240 -1650
rect 1200 -1740 1240 -1730
rect 1520 -1650 1560 -1640
rect 1520 -1730 1525 -1650
rect 1555 -1730 1560 -1650
rect 960 -1765 1160 -1760
rect 960 -1795 970 -1765
rect 1150 -1795 1160 -1765
rect 960 -1800 1160 -1795
rect 1280 -1765 1480 -1760
rect 1280 -1795 1290 -1765
rect 1470 -1795 1480 -1765
rect 1280 -1800 1480 -1795
rect 880 -2115 885 -2085
rect 915 -2115 920 -2085
rect 880 -2120 920 -2115
rect 1040 -2085 1080 -1800
rect 1040 -2115 1045 -2085
rect 1075 -2115 1080 -2085
rect 1040 -2120 1080 -2115
rect 1200 -2085 1240 -2080
rect 1200 -2115 1205 -2085
rect 1235 -2115 1240 -2085
rect -720 -2165 -680 -2160
rect -720 -2195 -715 -2165
rect -685 -2195 -680 -2165
rect -720 -2200 -680 -2195
rect -560 -2165 -520 -2160
rect -560 -2195 -555 -2165
rect -525 -2195 -520 -2165
rect -560 -2200 -520 -2195
rect -400 -2165 -360 -2160
rect -400 -2195 -395 -2165
rect -365 -2195 -360 -2165
rect -400 -2200 -360 -2195
rect -720 -2245 -680 -2240
rect -720 -2275 -715 -2245
rect -685 -2275 -680 -2245
rect -720 -2280 -680 -2275
rect -560 -2245 -520 -2240
rect -560 -2275 -555 -2245
rect -525 -2275 -520 -2245
rect -560 -2280 -520 -2275
rect -400 -2245 -360 -2240
rect -400 -2275 -395 -2245
rect -365 -2275 -360 -2245
rect -400 -2280 -360 -2275
rect 0 -2245 200 -2240
rect 0 -2275 10 -2245
rect 190 -2275 200 -2245
rect 0 -2280 200 -2275
rect 320 -2245 520 -2240
rect 320 -2275 330 -2245
rect 510 -2275 520 -2245
rect 320 -2280 520 -2275
rect 640 -2245 840 -2240
rect 640 -2275 650 -2245
rect 830 -2275 840 -2245
rect 640 -2280 840 -2275
rect 960 -2245 1160 -2240
rect 960 -2275 970 -2245
rect 1150 -2275 1160 -2245
rect 960 -2280 1160 -2275
rect -80 -2310 -40 -2300
rect -720 -2325 -680 -2320
rect -720 -2355 -715 -2325
rect -685 -2355 -680 -2325
rect -720 -2360 -680 -2355
rect -560 -2325 -520 -2320
rect -560 -2355 -555 -2325
rect -525 -2355 -520 -2325
rect -560 -2360 -520 -2355
rect -400 -2325 -360 -2320
rect -400 -2355 -395 -2325
rect -365 -2355 -360 -2325
rect -400 -2360 -360 -2355
rect -80 -2390 -75 -2310
rect -45 -2390 -40 -2310
rect -720 -2405 -680 -2400
rect -720 -2435 -715 -2405
rect -685 -2435 -680 -2405
rect -720 -2440 -680 -2435
rect -560 -2405 -520 -2400
rect -560 -2435 -555 -2405
rect -525 -2435 -520 -2405
rect -560 -2440 -520 -2435
rect -400 -2405 -360 -2400
rect -400 -2435 -395 -2405
rect -365 -2435 -360 -2405
rect -400 -2440 -360 -2435
rect -80 -2405 -40 -2390
rect 240 -2310 280 -2300
rect 240 -2390 245 -2310
rect 275 -2390 280 -2310
rect 240 -2400 280 -2390
rect 560 -2310 600 -2300
rect 560 -2390 565 -2310
rect 595 -2390 600 -2310
rect 560 -2400 600 -2390
rect 880 -2310 920 -2300
rect 880 -2390 885 -2310
rect 915 -2390 920 -2310
rect 880 -2400 920 -2390
rect 1200 -2310 1240 -2115
rect 1360 -2085 1400 -1800
rect 1360 -2115 1365 -2085
rect 1395 -2115 1400 -2085
rect 1360 -2120 1400 -2115
rect 1520 -2085 1560 -1730
rect 1840 -1650 1880 -1635
rect 2480 -1605 2520 -1600
rect 2480 -1635 2485 -1605
rect 2515 -1635 2520 -1605
rect 1840 -1730 1845 -1650
rect 1875 -1730 1880 -1650
rect 1840 -1740 1880 -1730
rect 2160 -1650 2200 -1640
rect 2160 -1730 2165 -1650
rect 2195 -1730 2200 -1650
rect 1600 -1765 1800 -1760
rect 1600 -1795 1610 -1765
rect 1790 -1795 1800 -1765
rect 1600 -1800 1800 -1795
rect 1920 -1765 2120 -1760
rect 1920 -1795 1930 -1765
rect 2110 -1795 2120 -1765
rect 1920 -1800 2120 -1795
rect 1520 -2115 1525 -2085
rect 1555 -2115 1560 -2085
rect 1520 -2120 1560 -2115
rect 1680 -2085 1720 -1800
rect 1680 -2115 1685 -2085
rect 1715 -2115 1720 -2085
rect 1680 -2120 1720 -2115
rect 2000 -2085 2040 -1800
rect 2000 -2115 2005 -2085
rect 2035 -2115 2040 -2085
rect 2000 -2120 2040 -2115
rect 2160 -2085 2200 -1730
rect 2480 -1650 2520 -1635
rect 3120 -1605 3160 -1600
rect 3120 -1635 3125 -1605
rect 3155 -1635 3160 -1605
rect 2480 -1730 2485 -1650
rect 2515 -1730 2520 -1650
rect 2480 -1740 2520 -1730
rect 2800 -1650 2840 -1640
rect 2800 -1730 2805 -1650
rect 2835 -1730 2840 -1650
rect 2240 -1765 2440 -1760
rect 2240 -1795 2250 -1765
rect 2430 -1795 2440 -1765
rect 2240 -1800 2440 -1795
rect 2560 -1765 2760 -1760
rect 2560 -1795 2570 -1765
rect 2750 -1795 2760 -1765
rect 2560 -1800 2760 -1795
rect 2160 -2115 2165 -2085
rect 2195 -2115 2200 -2085
rect 2160 -2120 2200 -2115
rect 2320 -2085 2360 -1800
rect 2320 -2115 2325 -2085
rect 2355 -2115 2360 -2085
rect 2320 -2120 2360 -2115
rect 2640 -2085 2680 -1800
rect 2640 -2115 2645 -2085
rect 2675 -2115 2680 -2085
rect 2640 -2120 2680 -2115
rect 2800 -2085 2840 -1730
rect 3120 -1650 3160 -1635
rect 3760 -1605 3800 -1600
rect 3760 -1635 3765 -1605
rect 3795 -1635 3800 -1605
rect 3120 -1730 3125 -1650
rect 3155 -1730 3160 -1650
rect 3120 -1740 3160 -1730
rect 3440 -1650 3480 -1640
rect 3440 -1730 3445 -1650
rect 3475 -1730 3480 -1650
rect 2880 -1765 3080 -1760
rect 2880 -1795 2890 -1765
rect 3070 -1795 3080 -1765
rect 2880 -1800 3080 -1795
rect 3200 -1765 3400 -1760
rect 3200 -1795 3210 -1765
rect 3390 -1795 3400 -1765
rect 3200 -1800 3400 -1795
rect 2800 -2115 2805 -2085
rect 2835 -2115 2840 -2085
rect 2800 -2120 2840 -2115
rect 2960 -2085 3000 -1800
rect 2960 -2115 2965 -2085
rect 2995 -2115 3000 -2085
rect 2960 -2120 3000 -2115
rect 3280 -2085 3320 -1800
rect 3280 -2115 3285 -2085
rect 3315 -2115 3320 -2085
rect 3280 -2120 3320 -2115
rect 3440 -2085 3480 -1730
rect 3760 -1650 3800 -1635
rect 4400 -1605 4440 -1600
rect 4400 -1635 4405 -1605
rect 4435 -1635 4440 -1605
rect 3760 -1730 3765 -1650
rect 3795 -1730 3800 -1650
rect 3760 -1740 3800 -1730
rect 4080 -1650 4120 -1640
rect 4080 -1730 4085 -1650
rect 4115 -1730 4120 -1650
rect 3520 -1765 3720 -1760
rect 3520 -1795 3530 -1765
rect 3710 -1795 3720 -1765
rect 3520 -1800 3720 -1795
rect 3840 -1765 4040 -1760
rect 3840 -1795 3850 -1765
rect 4030 -1795 4040 -1765
rect 3840 -1800 4040 -1795
rect 3440 -2115 3445 -2085
rect 3475 -2115 3480 -2085
rect 3440 -2120 3480 -2115
rect 3600 -2085 3640 -1800
rect 3600 -2115 3605 -2085
rect 3635 -2115 3640 -2085
rect 3600 -2120 3640 -2115
rect 3760 -2085 3800 -2080
rect 3760 -2115 3765 -2085
rect 3795 -2115 3800 -2085
rect 1280 -2245 1480 -2240
rect 1280 -2275 1290 -2245
rect 1470 -2275 1480 -2245
rect 1280 -2280 1480 -2275
rect 1600 -2245 1800 -2240
rect 1600 -2275 1610 -2245
rect 1790 -2275 1800 -2245
rect 1600 -2280 1800 -2275
rect 1920 -2245 2120 -2240
rect 1920 -2275 1930 -2245
rect 2110 -2275 2120 -2245
rect 1920 -2280 2120 -2275
rect 2240 -2245 2440 -2240
rect 2240 -2275 2250 -2245
rect 2430 -2275 2440 -2245
rect 2240 -2280 2440 -2275
rect 2560 -2245 2760 -2240
rect 2560 -2275 2570 -2245
rect 2750 -2275 2760 -2245
rect 2560 -2280 2760 -2275
rect 2880 -2245 3080 -2240
rect 2880 -2275 2890 -2245
rect 3070 -2275 3080 -2245
rect 2880 -2280 3080 -2275
rect 3200 -2245 3400 -2240
rect 3200 -2275 3210 -2245
rect 3390 -2275 3400 -2245
rect 3200 -2280 3400 -2275
rect 3520 -2245 3720 -2240
rect 3520 -2275 3530 -2245
rect 3710 -2275 3720 -2245
rect 3520 -2280 3720 -2275
rect 1200 -2390 1205 -2310
rect 1235 -2390 1240 -2310
rect 1200 -2400 1240 -2390
rect 1520 -2310 1560 -2300
rect 1520 -2390 1525 -2310
rect 1555 -2390 1560 -2310
rect 1520 -2400 1560 -2390
rect 1840 -2310 1880 -2300
rect 1840 -2390 1845 -2310
rect 1875 -2390 1880 -2310
rect 1840 -2400 1880 -2390
rect 2160 -2310 2200 -2300
rect 2160 -2390 2165 -2310
rect 2195 -2390 2200 -2310
rect 2160 -2400 2200 -2390
rect 2480 -2310 2520 -2300
rect 2480 -2390 2485 -2310
rect 2515 -2390 2520 -2310
rect -80 -2435 -75 -2405
rect -45 -2435 -40 -2405
rect -80 -2440 -40 -2435
rect 2480 -2405 2520 -2390
rect 2800 -2310 2840 -2300
rect 2800 -2390 2805 -2310
rect 2835 -2390 2840 -2310
rect 2800 -2400 2840 -2390
rect 3120 -2310 3160 -2300
rect 3120 -2390 3125 -2310
rect 3155 -2390 3160 -2310
rect 3120 -2400 3160 -2390
rect 3440 -2310 3480 -2300
rect 3440 -2390 3445 -2310
rect 3475 -2390 3480 -2310
rect 3440 -2400 3480 -2390
rect 3760 -2310 3800 -2115
rect 3920 -2085 3960 -1800
rect 3920 -2115 3925 -2085
rect 3955 -2115 3960 -2085
rect 3920 -2120 3960 -2115
rect 4080 -2085 4120 -1730
rect 4400 -1650 4440 -1635
rect 5040 -1605 5080 -1600
rect 5040 -1635 5045 -1605
rect 5075 -1635 5080 -1605
rect 4400 -1730 4405 -1650
rect 4435 -1730 4440 -1650
rect 4400 -1740 4440 -1730
rect 4720 -1650 4760 -1640
rect 4720 -1730 4725 -1650
rect 4755 -1730 4760 -1650
rect 4160 -1765 4360 -1760
rect 4160 -1795 4170 -1765
rect 4350 -1795 4360 -1765
rect 4160 -1800 4360 -1795
rect 4480 -1765 4680 -1760
rect 4480 -1795 4490 -1765
rect 4670 -1795 4680 -1765
rect 4480 -1800 4680 -1795
rect 4080 -2115 4085 -2085
rect 4115 -2115 4120 -2085
rect 4080 -2120 4120 -2115
rect 4240 -2085 4280 -1800
rect 4240 -2115 4245 -2085
rect 4275 -2115 4280 -2085
rect 4240 -2120 4280 -2115
rect 4560 -2085 4600 -1800
rect 4560 -2115 4565 -2085
rect 4595 -2115 4600 -2085
rect 4560 -2120 4600 -2115
rect 4720 -2085 4760 -1730
rect 5040 -1650 5080 -1635
rect 10320 -1605 10360 -1600
rect 10320 -1635 10325 -1605
rect 10355 -1635 10360 -1605
rect 5040 -1730 5045 -1650
rect 5075 -1730 5080 -1650
rect 5040 -1740 5080 -1730
rect 5200 -1650 5240 -1640
rect 5200 -1730 5205 -1650
rect 5235 -1730 5240 -1650
rect 4800 -1765 5000 -1760
rect 4800 -1795 4810 -1765
rect 4990 -1795 5000 -1765
rect 4800 -1800 5000 -1795
rect 4720 -2115 4725 -2085
rect 4755 -2115 4760 -2085
rect 4720 -2120 4760 -2115
rect 4880 -2085 4920 -1800
rect 4880 -2115 4885 -2085
rect 4915 -2115 4920 -2085
rect 4880 -2120 4920 -2115
rect 3840 -2245 4040 -2240
rect 3840 -2275 3850 -2245
rect 4030 -2275 4040 -2245
rect 3840 -2280 4040 -2275
rect 4160 -2245 4360 -2240
rect 4160 -2275 4170 -2245
rect 4350 -2275 4360 -2245
rect 4160 -2280 4360 -2275
rect 4480 -2245 4680 -2240
rect 4480 -2275 4490 -2245
rect 4670 -2275 4680 -2245
rect 4480 -2280 4680 -2275
rect 4800 -2245 5000 -2240
rect 4800 -2275 4810 -2245
rect 4990 -2275 5000 -2245
rect 4800 -2280 5000 -2275
rect 5200 -2245 5240 -1730
rect 5520 -1650 5560 -1640
rect 5520 -1730 5525 -1650
rect 5555 -1730 5560 -1650
rect 5520 -1740 5560 -1730
rect 5840 -1650 5880 -1640
rect 5840 -1730 5845 -1650
rect 5875 -1730 5880 -1650
rect 5840 -1740 5880 -1730
rect 6160 -1650 6200 -1640
rect 6160 -1730 6165 -1650
rect 6195 -1730 6200 -1650
rect 6160 -1740 6200 -1730
rect 6480 -1650 6520 -1640
rect 6480 -1730 6485 -1650
rect 6515 -1730 6520 -1650
rect 6480 -1740 6520 -1730
rect 6800 -1650 6840 -1640
rect 6800 -1730 6805 -1650
rect 6835 -1730 6840 -1650
rect 6800 -1740 6840 -1730
rect 7120 -1650 7160 -1640
rect 7120 -1730 7125 -1650
rect 7155 -1730 7160 -1650
rect 7120 -1740 7160 -1730
rect 7440 -1650 7480 -1640
rect 7440 -1730 7445 -1650
rect 7475 -1730 7480 -1650
rect 7440 -1740 7480 -1730
rect 7760 -1650 7800 -1640
rect 7760 -1730 7765 -1650
rect 7795 -1730 7800 -1650
rect 7760 -1740 7800 -1730
rect 8080 -1650 8120 -1640
rect 8080 -1730 8085 -1650
rect 8115 -1730 8120 -1650
rect 8080 -1740 8120 -1730
rect 8400 -1650 8440 -1640
rect 8400 -1730 8405 -1650
rect 8435 -1730 8440 -1650
rect 8400 -1740 8440 -1730
rect 8720 -1650 8760 -1640
rect 8720 -1730 8725 -1650
rect 8755 -1730 8760 -1650
rect 8720 -1740 8760 -1730
rect 9040 -1650 9080 -1640
rect 9040 -1730 9045 -1650
rect 9075 -1730 9080 -1650
rect 9040 -1740 9080 -1730
rect 9360 -1650 9400 -1640
rect 9360 -1730 9365 -1650
rect 9395 -1730 9400 -1650
rect 9360 -1740 9400 -1730
rect 9680 -1650 9720 -1640
rect 9680 -1730 9685 -1650
rect 9715 -1730 9720 -1650
rect 9680 -1740 9720 -1730
rect 10000 -1650 10040 -1640
rect 10000 -1730 10005 -1650
rect 10035 -1730 10040 -1650
rect 10000 -1740 10040 -1730
rect 10320 -1650 10360 -1635
rect 10640 -1605 10680 -1600
rect 10640 -1635 10645 -1605
rect 10675 -1635 10680 -1605
rect 10640 -1640 10680 -1635
rect 10800 -1605 10840 -1600
rect 10800 -1635 10805 -1605
rect 10835 -1635 10840 -1605
rect 10800 -1640 10840 -1635
rect 10960 -1605 11000 -1600
rect 10960 -1635 10965 -1605
rect 10995 -1635 11000 -1605
rect 10960 -1640 11000 -1635
rect 10320 -1730 10325 -1650
rect 10355 -1730 10360 -1650
rect 10640 -1685 10680 -1680
rect 10640 -1715 10645 -1685
rect 10675 -1715 10680 -1685
rect 10640 -1720 10680 -1715
rect 10800 -1685 10840 -1680
rect 10800 -1715 10805 -1685
rect 10835 -1715 10840 -1685
rect 10800 -1720 10840 -1715
rect 10960 -1685 11000 -1680
rect 10960 -1715 10965 -1685
rect 10995 -1715 11000 -1685
rect 10960 -1720 11000 -1715
rect 10320 -1740 10360 -1730
rect 5280 -1765 5480 -1760
rect 5280 -1795 5290 -1765
rect 5470 -1795 5480 -1765
rect 5280 -1800 5480 -1795
rect 5600 -1765 5800 -1760
rect 5600 -1795 5610 -1765
rect 5790 -1795 5800 -1765
rect 5600 -1800 5800 -1795
rect 5920 -1765 6120 -1760
rect 5920 -1795 5930 -1765
rect 6110 -1795 6120 -1765
rect 5920 -1800 6120 -1795
rect 6240 -1765 6440 -1760
rect 6240 -1795 6250 -1765
rect 6430 -1795 6440 -1765
rect 6240 -1800 6440 -1795
rect 6560 -1765 6760 -1760
rect 6560 -1795 6570 -1765
rect 6750 -1795 6760 -1765
rect 6560 -1800 6760 -1795
rect 6880 -1765 7080 -1760
rect 6880 -1795 6890 -1765
rect 7070 -1795 7080 -1765
rect 6880 -1800 7080 -1795
rect 7200 -1765 7400 -1760
rect 7200 -1795 7210 -1765
rect 7390 -1795 7400 -1765
rect 7200 -1800 7400 -1795
rect 7520 -1765 7720 -1760
rect 7520 -1795 7530 -1765
rect 7710 -1795 7720 -1765
rect 7520 -1800 7720 -1795
rect 7840 -1765 8040 -1760
rect 7840 -1795 7850 -1765
rect 8030 -1795 8040 -1765
rect 7840 -1800 8040 -1795
rect 8160 -1765 8360 -1760
rect 8160 -1795 8170 -1765
rect 8350 -1795 8360 -1765
rect 8160 -1800 8360 -1795
rect 8480 -1765 8680 -1760
rect 8480 -1795 8490 -1765
rect 8670 -1795 8680 -1765
rect 8480 -1800 8680 -1795
rect 8800 -1765 9000 -1760
rect 8800 -1795 8810 -1765
rect 8990 -1795 9000 -1765
rect 8800 -1800 9000 -1795
rect 9120 -1765 9320 -1760
rect 9120 -1795 9130 -1765
rect 9310 -1795 9320 -1765
rect 9120 -1800 9320 -1795
rect 9440 -1765 9640 -1760
rect 9440 -1795 9450 -1765
rect 9630 -1795 9640 -1765
rect 9440 -1800 9640 -1795
rect 9760 -1765 9960 -1760
rect 9760 -1795 9770 -1765
rect 9950 -1795 9960 -1765
rect 9760 -1800 9960 -1795
rect 10080 -1765 10280 -1760
rect 10080 -1795 10090 -1765
rect 10270 -1795 10280 -1765
rect 10080 -1800 10280 -1795
rect 10640 -1765 10680 -1760
rect 10640 -1795 10645 -1765
rect 10675 -1795 10680 -1765
rect 10640 -1800 10680 -1795
rect 10800 -1765 10840 -1760
rect 10800 -1795 10805 -1765
rect 10835 -1795 10840 -1765
rect 10800 -1800 10840 -1795
rect 10960 -1765 11000 -1760
rect 10960 -1795 10965 -1765
rect 10995 -1795 11000 -1765
rect 10960 -1800 11000 -1795
rect 5360 -1925 5400 -1800
rect 5360 -1955 5365 -1925
rect 5395 -1955 5400 -1925
rect 5360 -1960 5400 -1955
rect 5680 -1925 5720 -1800
rect 5680 -1955 5685 -1925
rect 5715 -1955 5720 -1925
rect 5680 -1960 5720 -1955
rect 6000 -1925 6040 -1800
rect 6000 -1955 6005 -1925
rect 6035 -1955 6040 -1925
rect 6000 -1960 6040 -1955
rect 6320 -1925 6360 -1800
rect 6320 -1955 6325 -1925
rect 6355 -1955 6360 -1925
rect 6320 -1960 6360 -1955
rect 6640 -1925 6680 -1800
rect 6640 -1955 6645 -1925
rect 6675 -1955 6680 -1925
rect 6640 -1960 6680 -1955
rect 6960 -1925 7000 -1800
rect 6960 -1955 6965 -1925
rect 6995 -1955 7000 -1925
rect 6960 -1960 7000 -1955
rect 7280 -1925 7320 -1800
rect 7280 -1955 7285 -1925
rect 7315 -1955 7320 -1925
rect 7280 -1960 7320 -1955
rect 7600 -1925 7640 -1800
rect 7600 -1955 7605 -1925
rect 7635 -1955 7640 -1925
rect 7600 -1960 7640 -1955
rect 7920 -1925 7960 -1800
rect 7920 -1955 7925 -1925
rect 7955 -1955 7960 -1925
rect 7920 -1960 7960 -1955
rect 8240 -1925 8280 -1800
rect 8240 -1955 8245 -1925
rect 8275 -1955 8280 -1925
rect 8240 -1960 8280 -1955
rect 8560 -1925 8600 -1800
rect 8560 -1955 8565 -1925
rect 8595 -1955 8600 -1925
rect 8560 -1960 8600 -1955
rect 8880 -1925 8920 -1800
rect 8880 -1955 8885 -1925
rect 8915 -1955 8920 -1925
rect 8880 -1960 8920 -1955
rect 9200 -1925 9240 -1800
rect 9200 -1955 9205 -1925
rect 9235 -1955 9240 -1925
rect 9200 -1960 9240 -1955
rect 9520 -1925 9560 -1800
rect 9520 -1955 9525 -1925
rect 9555 -1955 9560 -1925
rect 9520 -1960 9560 -1955
rect 9840 -1925 9880 -1800
rect 9840 -1955 9845 -1925
rect 9875 -1955 9880 -1925
rect 9840 -1960 9880 -1955
rect 10160 -1925 10200 -1800
rect 10640 -1845 10680 -1840
rect 10640 -1875 10645 -1845
rect 10675 -1875 10680 -1845
rect 10640 -1880 10680 -1875
rect 10800 -1845 10840 -1840
rect 10800 -1875 10805 -1845
rect 10835 -1875 10840 -1845
rect 10800 -1880 10840 -1875
rect 10960 -1845 11000 -1840
rect 10960 -1875 10965 -1845
rect 10995 -1875 11000 -1845
rect 10960 -1880 11000 -1875
rect 10160 -1955 10165 -1925
rect 10195 -1955 10200 -1925
rect 10160 -1960 10200 -1955
rect 10640 -1925 10680 -1920
rect 10640 -1955 10645 -1925
rect 10675 -1955 10680 -1925
rect 10640 -1960 10680 -1955
rect 10800 -1925 10840 -1920
rect 10800 -1955 10805 -1925
rect 10835 -1955 10840 -1925
rect 10800 -1960 10840 -1955
rect 10960 -1925 11000 -1920
rect 10960 -1955 10965 -1925
rect 10995 -1955 11000 -1925
rect 10960 -1960 11000 -1955
rect 10640 -2005 10680 -2000
rect 10640 -2035 10645 -2005
rect 10675 -2035 10680 -2005
rect 10640 -2040 10680 -2035
rect 10800 -2005 10840 -2000
rect 10800 -2035 10805 -2005
rect 10835 -2035 10840 -2005
rect 10800 -2040 10840 -2035
rect 10960 -2005 11000 -2000
rect 10960 -2035 10965 -2005
rect 10995 -2035 11000 -2005
rect 10960 -2040 11000 -2035
rect 10640 -2165 10680 -2160
rect 10640 -2195 10645 -2165
rect 10675 -2195 10680 -2165
rect 10640 -2200 10680 -2195
rect 10800 -2165 10840 -2160
rect 10800 -2195 10805 -2165
rect 10835 -2195 10840 -2165
rect 10800 -2200 10840 -2195
rect 10960 -2165 11000 -2160
rect 10960 -2195 10965 -2165
rect 10995 -2195 11000 -2165
rect 10960 -2200 11000 -2195
rect 5200 -2275 5205 -2245
rect 5235 -2275 5240 -2245
rect 5200 -2280 5240 -2275
rect 5280 -2245 5480 -2240
rect 5280 -2275 5290 -2245
rect 5470 -2275 5480 -2245
rect 5280 -2280 5480 -2275
rect 5600 -2245 5800 -2240
rect 5600 -2275 5610 -2245
rect 5790 -2275 5800 -2245
rect 5600 -2280 5800 -2275
rect 5920 -2245 6120 -2240
rect 5920 -2275 5930 -2245
rect 6110 -2275 6120 -2245
rect 5920 -2280 6120 -2275
rect 6240 -2245 6440 -2240
rect 6240 -2275 6250 -2245
rect 6430 -2275 6440 -2245
rect 6240 -2280 6440 -2275
rect 6480 -2245 6520 -2240
rect 6480 -2275 6485 -2245
rect 6515 -2275 6520 -2245
rect 3760 -2390 3765 -2310
rect 3795 -2390 3800 -2310
rect 3760 -2400 3800 -2390
rect 4080 -2310 4120 -2300
rect 4080 -2390 4085 -2310
rect 4115 -2390 4120 -2310
rect 4080 -2400 4120 -2390
rect 4400 -2310 4440 -2300
rect 4400 -2390 4405 -2310
rect 4435 -2390 4440 -2310
rect 4400 -2400 4440 -2390
rect 4720 -2310 4760 -2300
rect 4720 -2390 4725 -2310
rect 4755 -2390 4760 -2310
rect 4720 -2400 4760 -2390
rect 5040 -2310 5080 -2300
rect 5040 -2390 5045 -2310
rect 5075 -2390 5080 -2310
rect 2480 -2435 2485 -2405
rect 2515 -2435 2520 -2405
rect 2480 -2440 2520 -2435
rect 5040 -2405 5080 -2390
rect 5040 -2435 5045 -2405
rect 5075 -2435 5080 -2405
rect 5040 -2440 5080 -2435
rect 5200 -2310 5240 -2300
rect 5200 -2390 5205 -2310
rect 5235 -2390 5240 -2310
rect 5200 -2405 5240 -2390
rect 5520 -2310 5560 -2300
rect 5520 -2390 5525 -2310
rect 5555 -2390 5560 -2310
rect 5520 -2400 5560 -2390
rect 5840 -2310 5880 -2300
rect 5840 -2390 5845 -2310
rect 5875 -2390 5880 -2310
rect 5840 -2400 5880 -2390
rect 6160 -2310 6200 -2300
rect 6160 -2390 6165 -2310
rect 6195 -2390 6200 -2310
rect 6160 -2400 6200 -2390
rect 6480 -2310 6520 -2275
rect 6560 -2245 6760 -2240
rect 6560 -2275 6570 -2245
rect 6750 -2275 6760 -2245
rect 6560 -2280 6760 -2275
rect 6880 -2245 7080 -2240
rect 6880 -2275 6890 -2245
rect 7070 -2275 7080 -2245
rect 6880 -2280 7080 -2275
rect 7200 -2245 7400 -2240
rect 7200 -2275 7210 -2245
rect 7390 -2275 7400 -2245
rect 7200 -2280 7400 -2275
rect 7520 -2245 7720 -2240
rect 7520 -2275 7530 -2245
rect 7710 -2275 7720 -2245
rect 7520 -2280 7720 -2275
rect 7840 -2245 8040 -2240
rect 7840 -2275 7850 -2245
rect 8030 -2275 8040 -2245
rect 7840 -2280 8040 -2275
rect 8160 -2245 8360 -2240
rect 8160 -2275 8170 -2245
rect 8350 -2275 8360 -2245
rect 8160 -2280 8360 -2275
rect 8480 -2245 8680 -2240
rect 8480 -2275 8490 -2245
rect 8670 -2275 8680 -2245
rect 8480 -2280 8680 -2275
rect 8800 -2245 9000 -2240
rect 8800 -2275 8810 -2245
rect 8990 -2275 9000 -2245
rect 8800 -2280 9000 -2275
rect 9040 -2245 9080 -2240
rect 9040 -2275 9045 -2245
rect 9075 -2275 9080 -2245
rect 6480 -2390 6485 -2310
rect 6515 -2390 6520 -2310
rect 6480 -2400 6520 -2390
rect 6800 -2310 6840 -2300
rect 6800 -2390 6805 -2310
rect 6835 -2390 6840 -2310
rect 6800 -2400 6840 -2390
rect 7120 -2310 7160 -2300
rect 7120 -2390 7125 -2310
rect 7155 -2390 7160 -2310
rect 7120 -2400 7160 -2390
rect 7440 -2310 7480 -2300
rect 7440 -2390 7445 -2310
rect 7475 -2390 7480 -2310
rect 7440 -2400 7480 -2390
rect 7760 -2310 7800 -2300
rect 7760 -2390 7765 -2310
rect 7795 -2390 7800 -2310
rect 5200 -2435 5205 -2405
rect 5235 -2435 5240 -2405
rect 5200 -2440 5240 -2435
rect 7760 -2405 7800 -2390
rect 8080 -2310 8120 -2300
rect 8080 -2390 8085 -2310
rect 8115 -2390 8120 -2310
rect 8080 -2400 8120 -2390
rect 8400 -2310 8440 -2300
rect 8400 -2390 8405 -2310
rect 8435 -2390 8440 -2310
rect 8400 -2400 8440 -2390
rect 8720 -2310 8760 -2300
rect 8720 -2390 8725 -2310
rect 8755 -2390 8760 -2310
rect 8720 -2400 8760 -2390
rect 9040 -2310 9080 -2275
rect 9120 -2245 9320 -2240
rect 9120 -2275 9130 -2245
rect 9310 -2275 9320 -2245
rect 9120 -2280 9320 -2275
rect 9440 -2245 9640 -2240
rect 9440 -2275 9450 -2245
rect 9630 -2275 9640 -2245
rect 9440 -2280 9640 -2275
rect 9760 -2245 9960 -2240
rect 9760 -2275 9770 -2245
rect 9950 -2275 9960 -2245
rect 9760 -2280 9960 -2275
rect 10080 -2245 10280 -2240
rect 10080 -2275 10090 -2245
rect 10270 -2275 10280 -2245
rect 10080 -2280 10280 -2275
rect 10800 -2245 10840 -2240
rect 10800 -2275 10805 -2245
rect 10835 -2275 10840 -2245
rect 10800 -2280 10840 -2275
rect 10960 -2245 11000 -2240
rect 10960 -2275 10965 -2245
rect 10995 -2275 11000 -2245
rect 10960 -2280 11000 -2275
rect 9040 -2390 9045 -2310
rect 9075 -2390 9080 -2310
rect 9040 -2400 9080 -2390
rect 9360 -2310 9400 -2300
rect 9360 -2390 9365 -2310
rect 9395 -2390 9400 -2310
rect 9360 -2400 9400 -2390
rect 9680 -2310 9720 -2300
rect 9680 -2390 9685 -2310
rect 9715 -2390 9720 -2310
rect 9680 -2400 9720 -2390
rect 10000 -2310 10040 -2300
rect 10000 -2390 10005 -2310
rect 10035 -2390 10040 -2310
rect 10000 -2400 10040 -2390
rect 10320 -2310 10360 -2300
rect 10320 -2390 10325 -2310
rect 10355 -2390 10360 -2310
rect 10640 -2325 10680 -2320
rect 10640 -2355 10645 -2325
rect 10675 -2355 10680 -2325
rect 10640 -2360 10680 -2355
rect 10800 -2325 10840 -2320
rect 10800 -2355 10805 -2325
rect 10835 -2355 10840 -2325
rect 10800 -2360 10840 -2355
rect 10960 -2325 11000 -2320
rect 10960 -2355 10965 -2325
rect 10995 -2355 11000 -2325
rect 10960 -2360 11000 -2355
rect 7760 -2435 7765 -2405
rect 7795 -2435 7800 -2405
rect 7760 -2440 7800 -2435
rect 10320 -2405 10360 -2390
rect 10320 -2435 10325 -2405
rect 10355 -2435 10360 -2405
rect 10320 -2440 10360 -2435
rect 10640 -2405 10680 -2400
rect 10640 -2435 10645 -2405
rect 10675 -2435 10680 -2405
rect 10640 -2440 10680 -2435
rect 10800 -2405 10840 -2400
rect 10800 -2435 10805 -2405
rect 10835 -2435 10840 -2405
rect 10800 -2440 10840 -2435
rect 10960 -2405 11000 -2400
rect 10960 -2435 10965 -2405
rect 10995 -2435 11000 -2405
rect 10960 -2440 11000 -2435
rect -720 -2485 -680 -2480
rect -720 -2515 -715 -2485
rect -685 -2515 -680 -2485
rect -720 -2520 -680 -2515
rect -560 -2485 -520 -2480
rect -560 -2515 -555 -2485
rect -525 -2515 -520 -2485
rect -560 -2520 -520 -2515
rect -400 -2485 -360 -2480
rect -400 -2515 -395 -2485
rect -365 -2515 -360 -2485
rect -400 -2520 -360 -2515
rect 10640 -2485 10680 -2480
rect 10640 -2515 10645 -2485
rect 10675 -2515 10680 -2485
rect 10640 -2520 10680 -2515
rect 10800 -2485 10840 -2480
rect 10800 -2515 10805 -2485
rect 10835 -2515 10840 -2485
rect 10800 -2520 10840 -2515
rect 10960 -2485 11000 -2480
rect 10960 -2515 10965 -2485
rect 10995 -2515 11000 -2485
rect 10960 -2520 11000 -2515
rect -720 -2565 -680 -2560
rect -720 -2595 -715 -2565
rect -685 -2595 -680 -2565
rect -720 -2600 -680 -2595
rect -560 -2565 -520 -2560
rect -560 -2595 -555 -2565
rect -525 -2595 -520 -2565
rect -560 -2600 -520 -2595
rect -400 -2565 -360 -2560
rect -400 -2595 -395 -2565
rect -365 -2595 -360 -2565
rect -400 -2600 -360 -2595
rect 10640 -2565 10680 -2560
rect 10640 -2595 10645 -2565
rect 10675 -2595 10680 -2565
rect 10640 -2600 10680 -2595
rect 10800 -2565 10840 -2560
rect 10800 -2595 10805 -2565
rect 10835 -2595 10840 -2565
rect 10800 -2600 10840 -2595
rect 10960 -2565 11000 -2560
rect 10960 -2595 10965 -2565
rect 10995 -2595 11000 -2565
rect 10960 -2600 11000 -2595
rect -720 -2645 -680 -2640
rect -720 -2675 -715 -2645
rect -685 -2675 -680 -2645
rect -720 -2680 -680 -2675
rect -560 -2645 -520 -2640
rect -560 -2675 -555 -2645
rect -525 -2675 -520 -2645
rect -560 -2680 -520 -2675
rect -400 -2645 -360 -2640
rect -400 -2675 -395 -2645
rect -365 -2675 -360 -2645
rect -400 -2680 -360 -2675
rect -80 -2645 -40 -2640
rect -80 -2675 -75 -2645
rect -45 -2675 -40 -2645
rect -80 -2690 -40 -2675
rect 2480 -2645 2520 -2640
rect 2480 -2675 2485 -2645
rect 2515 -2675 2520 -2645
rect -720 -2725 -680 -2720
rect -720 -2755 -715 -2725
rect -685 -2755 -680 -2725
rect -720 -2760 -680 -2755
rect -560 -2725 -520 -2720
rect -560 -2755 -555 -2725
rect -525 -2755 -520 -2725
rect -560 -2760 -520 -2755
rect -400 -2725 -360 -2720
rect -400 -2755 -395 -2725
rect -365 -2755 -360 -2725
rect -400 -2760 -360 -2755
rect -80 -2770 -75 -2690
rect -45 -2770 -40 -2690
rect -80 -2780 -40 -2770
rect 240 -2690 280 -2680
rect 240 -2770 245 -2690
rect 275 -2770 280 -2690
rect 240 -2780 280 -2770
rect 560 -2690 600 -2680
rect 560 -2770 565 -2690
rect 595 -2770 600 -2690
rect 560 -2780 600 -2770
rect 880 -2690 920 -2680
rect 880 -2770 885 -2690
rect 915 -2770 920 -2690
rect 880 -2780 920 -2770
rect 1200 -2690 1240 -2680
rect 1200 -2770 1205 -2690
rect 1235 -2770 1240 -2690
rect -720 -2805 -680 -2800
rect -720 -2835 -715 -2805
rect -685 -2835 -680 -2805
rect -720 -2840 -680 -2835
rect -560 -2805 -520 -2800
rect -560 -2835 -555 -2805
rect -525 -2835 -520 -2805
rect -560 -2840 -520 -2835
rect -400 -2805 -360 -2800
rect -400 -2835 -395 -2805
rect -365 -2835 -360 -2805
rect -400 -2840 -360 -2835
rect 0 -2805 200 -2800
rect 0 -2835 10 -2805
rect 190 -2835 200 -2805
rect 0 -2840 200 -2835
rect 320 -2805 520 -2800
rect 320 -2835 330 -2805
rect 510 -2835 520 -2805
rect 320 -2840 520 -2835
rect 640 -2805 840 -2800
rect 640 -2835 650 -2805
rect 830 -2835 840 -2805
rect 640 -2840 840 -2835
rect 960 -2805 1160 -2800
rect 960 -2835 970 -2805
rect 1150 -2835 1160 -2805
rect 960 -2840 1160 -2835
rect 1200 -2805 1240 -2770
rect 1520 -2690 1560 -2680
rect 1520 -2770 1525 -2690
rect 1555 -2770 1560 -2690
rect 1520 -2780 1560 -2770
rect 1840 -2690 1880 -2680
rect 1840 -2770 1845 -2690
rect 1875 -2770 1880 -2690
rect 1840 -2780 1880 -2770
rect 2160 -2690 2200 -2680
rect 2160 -2770 2165 -2690
rect 2195 -2770 2200 -2690
rect 2160 -2780 2200 -2770
rect 2480 -2690 2520 -2675
rect 5040 -2645 5080 -2640
rect 5040 -2675 5045 -2645
rect 5075 -2675 5080 -2645
rect 2480 -2770 2485 -2690
rect 2515 -2770 2520 -2690
rect 2480 -2780 2520 -2770
rect 2800 -2690 2840 -2680
rect 2800 -2770 2805 -2690
rect 2835 -2770 2840 -2690
rect 2800 -2780 2840 -2770
rect 3120 -2690 3160 -2680
rect 3120 -2770 3125 -2690
rect 3155 -2770 3160 -2690
rect 3120 -2780 3160 -2770
rect 3440 -2690 3480 -2680
rect 3440 -2770 3445 -2690
rect 3475 -2770 3480 -2690
rect 3440 -2780 3480 -2770
rect 3760 -2690 3800 -2680
rect 3760 -2770 3765 -2690
rect 3795 -2770 3800 -2690
rect 1200 -2835 1205 -2805
rect 1235 -2835 1240 -2805
rect 1200 -2840 1240 -2835
rect 1280 -2805 1480 -2800
rect 1280 -2835 1290 -2805
rect 1470 -2835 1480 -2805
rect 1280 -2840 1480 -2835
rect 1600 -2805 1800 -2800
rect 1600 -2835 1610 -2805
rect 1790 -2835 1800 -2805
rect 1600 -2840 1800 -2835
rect 1920 -2805 2120 -2800
rect 1920 -2835 1930 -2805
rect 2110 -2835 2120 -2805
rect 1920 -2840 2120 -2835
rect 2240 -2805 2440 -2800
rect 2240 -2835 2250 -2805
rect 2430 -2835 2440 -2805
rect 2240 -2840 2440 -2835
rect 2560 -2805 2760 -2800
rect 2560 -2835 2570 -2805
rect 2750 -2835 2760 -2805
rect 2560 -2840 2760 -2835
rect 2880 -2805 3080 -2800
rect 2880 -2835 2890 -2805
rect 3070 -2835 3080 -2805
rect 2880 -2840 3080 -2835
rect 3200 -2805 3400 -2800
rect 3200 -2835 3210 -2805
rect 3390 -2835 3400 -2805
rect 3200 -2840 3400 -2835
rect 3520 -2805 3720 -2800
rect 3520 -2835 3530 -2805
rect 3710 -2835 3720 -2805
rect 3520 -2840 3720 -2835
rect 3760 -2805 3800 -2770
rect 4080 -2690 4120 -2680
rect 4080 -2770 4085 -2690
rect 4115 -2770 4120 -2690
rect 4080 -2780 4120 -2770
rect 4400 -2690 4440 -2680
rect 4400 -2770 4405 -2690
rect 4435 -2770 4440 -2690
rect 4400 -2780 4440 -2770
rect 4720 -2690 4760 -2680
rect 4720 -2770 4725 -2690
rect 4755 -2770 4760 -2690
rect 4720 -2780 4760 -2770
rect 5040 -2690 5080 -2675
rect 5040 -2770 5045 -2690
rect 5075 -2770 5080 -2690
rect 5040 -2780 5080 -2770
rect 5200 -2645 5240 -2640
rect 5200 -2675 5205 -2645
rect 5235 -2675 5240 -2645
rect 5200 -2690 5240 -2675
rect 7760 -2645 7800 -2640
rect 7760 -2675 7765 -2645
rect 7795 -2675 7800 -2645
rect 5200 -2770 5205 -2690
rect 5235 -2770 5240 -2690
rect 5200 -2780 5240 -2770
rect 5520 -2690 5560 -2680
rect 5520 -2770 5525 -2690
rect 5555 -2770 5560 -2690
rect 5520 -2780 5560 -2770
rect 5840 -2690 5880 -2680
rect 5840 -2770 5845 -2690
rect 5875 -2770 5880 -2690
rect 5840 -2780 5880 -2770
rect 6160 -2690 6200 -2680
rect 6160 -2770 6165 -2690
rect 6195 -2770 6200 -2690
rect 6160 -2780 6200 -2770
rect 6480 -2690 6520 -2680
rect 6480 -2770 6485 -2690
rect 6515 -2770 6520 -2690
rect 3760 -2835 3765 -2805
rect 3795 -2835 3800 -2805
rect 3760 -2840 3800 -2835
rect 3840 -2805 4040 -2800
rect 3840 -2835 3850 -2805
rect 4030 -2835 4040 -2805
rect 3840 -2840 4040 -2835
rect 4160 -2805 4360 -2800
rect 4160 -2835 4170 -2805
rect 4350 -2835 4360 -2805
rect 4160 -2840 4360 -2835
rect 4480 -2805 4680 -2800
rect 4480 -2835 4490 -2805
rect 4670 -2835 4680 -2805
rect 4480 -2840 4680 -2835
rect 4800 -2805 5000 -2800
rect 4800 -2835 4810 -2805
rect 4990 -2835 5000 -2805
rect 4800 -2840 5000 -2835
rect 5040 -2805 5080 -2800
rect 5040 -2835 5045 -2805
rect 5075 -2835 5080 -2805
rect -720 -2885 -680 -2880
rect -720 -2915 -715 -2885
rect -685 -2915 -680 -2885
rect -720 -2920 -680 -2915
rect -560 -2885 -520 -2880
rect -560 -2915 -555 -2885
rect -525 -2915 -520 -2885
rect -560 -2920 -520 -2915
rect -400 -2885 -360 -2880
rect -400 -2915 -395 -2885
rect -365 -2915 -360 -2885
rect -400 -2920 -360 -2915
rect -720 -2965 -680 -2960
rect -720 -2995 -715 -2965
rect -685 -2995 -680 -2965
rect -720 -3000 -680 -2995
rect -560 -2965 -520 -2960
rect -560 -2995 -555 -2965
rect -525 -2995 -520 -2965
rect -560 -3000 -520 -2995
rect -400 -2965 -360 -2960
rect -400 -2995 -395 -2965
rect -365 -2995 -360 -2965
rect -400 -3000 -360 -2995
rect -720 -3045 -680 -3040
rect -720 -3075 -715 -3045
rect -685 -3075 -680 -3045
rect -720 -3080 -680 -3075
rect -560 -3045 -520 -3040
rect -560 -3075 -555 -3045
rect -525 -3075 -520 -3045
rect -560 -3080 -520 -3075
rect -400 -3045 -360 -3040
rect -400 -3075 -395 -3045
rect -365 -3075 -360 -3045
rect -400 -3080 -360 -3075
rect -720 -3125 -680 -3120
rect -720 -3155 -715 -3125
rect -685 -3155 -680 -3125
rect -720 -3160 -680 -3155
rect -560 -3125 -520 -3120
rect -560 -3155 -555 -3125
rect -525 -3155 -520 -3125
rect -560 -3160 -520 -3155
rect 80 -3125 120 -3120
rect 80 -3155 85 -3125
rect 115 -3155 120 -3125
rect -720 -3205 -680 -3200
rect -720 -3235 -715 -3205
rect -685 -3235 -680 -3205
rect -720 -3240 -680 -3235
rect -560 -3205 -520 -3200
rect -560 -3235 -555 -3205
rect -525 -3235 -520 -3205
rect -560 -3240 -520 -3235
rect -400 -3205 -360 -3200
rect -400 -3235 -395 -3205
rect -365 -3235 -360 -3205
rect -400 -3240 -360 -3235
rect 80 -3280 120 -3155
rect 400 -3125 440 -3120
rect 400 -3155 405 -3125
rect 435 -3155 440 -3125
rect 400 -3280 440 -3155
rect 720 -3125 760 -3120
rect 720 -3155 725 -3125
rect 755 -3155 760 -3125
rect 720 -3280 760 -3155
rect 1040 -3125 1080 -3120
rect 1040 -3155 1045 -3125
rect 1075 -3155 1080 -3125
rect 1040 -3280 1080 -3155
rect 1360 -3125 1400 -3120
rect 1360 -3155 1365 -3125
rect 1395 -3155 1400 -3125
rect 1360 -3280 1400 -3155
rect 1680 -3125 1720 -3120
rect 1680 -3155 1685 -3125
rect 1715 -3155 1720 -3125
rect 1680 -3280 1720 -3155
rect 2000 -3125 2040 -3120
rect 2000 -3155 2005 -3125
rect 2035 -3155 2040 -3125
rect 2000 -3280 2040 -3155
rect 2320 -3125 2360 -3120
rect 2320 -3155 2325 -3125
rect 2355 -3155 2360 -3125
rect 2320 -3280 2360 -3155
rect 2640 -3125 2680 -3120
rect 2640 -3155 2645 -3125
rect 2675 -3155 2680 -3125
rect 2640 -3280 2680 -3155
rect 2960 -3125 3000 -3120
rect 2960 -3155 2965 -3125
rect 2995 -3155 3000 -3125
rect 2960 -3280 3000 -3155
rect 3280 -3125 3320 -3120
rect 3280 -3155 3285 -3125
rect 3315 -3155 3320 -3125
rect 3280 -3280 3320 -3155
rect 3600 -3125 3640 -3120
rect 3600 -3155 3605 -3125
rect 3635 -3155 3640 -3125
rect 3600 -3280 3640 -3155
rect 3920 -3125 3960 -3120
rect 3920 -3155 3925 -3125
rect 3955 -3155 3960 -3125
rect 3920 -3280 3960 -3155
rect 4240 -3125 4280 -3120
rect 4240 -3155 4245 -3125
rect 4275 -3155 4280 -3125
rect 4240 -3280 4280 -3155
rect 4560 -3125 4600 -3120
rect 4560 -3155 4565 -3125
rect 4595 -3155 4600 -3125
rect 4560 -3280 4600 -3155
rect 4880 -3125 4920 -3120
rect 4880 -3155 4885 -3125
rect 4915 -3155 4920 -3125
rect 4880 -3280 4920 -3155
rect -720 -3285 -680 -3280
rect -720 -3315 -715 -3285
rect -685 -3315 -680 -3285
rect -720 -3320 -680 -3315
rect -560 -3285 -520 -3280
rect -560 -3315 -555 -3285
rect -525 -3315 -520 -3285
rect -560 -3320 -520 -3315
rect -400 -3285 -360 -3280
rect -400 -3315 -395 -3285
rect -365 -3315 -360 -3285
rect -400 -3320 -360 -3315
rect 0 -3285 200 -3280
rect 0 -3315 10 -3285
rect 190 -3315 200 -3285
rect 0 -3320 200 -3315
rect 320 -3285 520 -3280
rect 320 -3315 330 -3285
rect 510 -3315 520 -3285
rect 320 -3320 520 -3315
rect 640 -3285 840 -3280
rect 640 -3315 650 -3285
rect 830 -3315 840 -3285
rect 640 -3320 840 -3315
rect 960 -3285 1160 -3280
rect 960 -3315 970 -3285
rect 1150 -3315 1160 -3285
rect 960 -3320 1160 -3315
rect 1280 -3285 1480 -3280
rect 1280 -3315 1290 -3285
rect 1470 -3315 1480 -3285
rect 1280 -3320 1480 -3315
rect 1600 -3285 1800 -3280
rect 1600 -3315 1610 -3285
rect 1790 -3315 1800 -3285
rect 1600 -3320 1800 -3315
rect 1920 -3285 2120 -3280
rect 1920 -3315 1930 -3285
rect 2110 -3315 2120 -3285
rect 1920 -3320 2120 -3315
rect 2240 -3285 2440 -3280
rect 2240 -3315 2250 -3285
rect 2430 -3315 2440 -3285
rect 2240 -3320 2440 -3315
rect 2560 -3285 2760 -3280
rect 2560 -3315 2570 -3285
rect 2750 -3315 2760 -3285
rect 2560 -3320 2760 -3315
rect 2880 -3285 3080 -3280
rect 2880 -3315 2890 -3285
rect 3070 -3315 3080 -3285
rect 2880 -3320 3080 -3315
rect 3200 -3285 3400 -3280
rect 3200 -3315 3210 -3285
rect 3390 -3315 3400 -3285
rect 3200 -3320 3400 -3315
rect 3520 -3285 3720 -3280
rect 3520 -3315 3530 -3285
rect 3710 -3315 3720 -3285
rect 3520 -3320 3720 -3315
rect 3840 -3285 4040 -3280
rect 3840 -3315 3850 -3285
rect 4030 -3315 4040 -3285
rect 3840 -3320 4040 -3315
rect 4160 -3285 4360 -3280
rect 4160 -3315 4170 -3285
rect 4350 -3315 4360 -3285
rect 4160 -3320 4360 -3315
rect 4480 -3285 4680 -3280
rect 4480 -3315 4490 -3285
rect 4670 -3315 4680 -3285
rect 4480 -3320 4680 -3315
rect 4800 -3285 5000 -3280
rect 4800 -3315 4810 -3285
rect 4990 -3315 5000 -3285
rect 4800 -3320 5000 -3315
rect -80 -3350 -40 -3340
rect -80 -3430 -75 -3350
rect -45 -3430 -40 -3350
rect -80 -3445 -40 -3430
rect 240 -3350 280 -3340
rect 240 -3430 245 -3350
rect 275 -3430 280 -3350
rect 240 -3440 280 -3430
rect 560 -3350 600 -3340
rect 560 -3430 565 -3350
rect 595 -3430 600 -3350
rect 560 -3440 600 -3430
rect 880 -3350 920 -3340
rect 880 -3430 885 -3350
rect 915 -3430 920 -3350
rect 880 -3440 920 -3430
rect 1200 -3350 1240 -3340
rect 1200 -3430 1205 -3350
rect 1235 -3430 1240 -3350
rect 1200 -3440 1240 -3430
rect 1520 -3350 1560 -3340
rect 1520 -3430 1525 -3350
rect 1555 -3430 1560 -3350
rect 1520 -3440 1560 -3430
rect 1840 -3350 1880 -3340
rect 1840 -3430 1845 -3350
rect 1875 -3430 1880 -3350
rect 1840 -3440 1880 -3430
rect 2160 -3350 2200 -3340
rect 2160 -3430 2165 -3350
rect 2195 -3430 2200 -3350
rect 2160 -3440 2200 -3430
rect 2480 -3350 2520 -3340
rect 2480 -3430 2485 -3350
rect 2515 -3430 2520 -3350
rect 2480 -3440 2520 -3430
rect 2800 -3350 2840 -3340
rect 2800 -3430 2805 -3350
rect 2835 -3430 2840 -3350
rect 2800 -3440 2840 -3430
rect 3120 -3350 3160 -3340
rect 3120 -3430 3125 -3350
rect 3155 -3430 3160 -3350
rect 3120 -3440 3160 -3430
rect 3440 -3350 3480 -3340
rect 3440 -3430 3445 -3350
rect 3475 -3430 3480 -3350
rect 3440 -3440 3480 -3430
rect 3760 -3350 3800 -3340
rect 3760 -3430 3765 -3350
rect 3795 -3430 3800 -3350
rect 3760 -3440 3800 -3430
rect 4080 -3350 4120 -3340
rect 4080 -3430 4085 -3350
rect 4115 -3430 4120 -3350
rect 4080 -3440 4120 -3430
rect 4400 -3350 4440 -3340
rect 4400 -3430 4405 -3350
rect 4435 -3430 4440 -3350
rect 4400 -3440 4440 -3430
rect 4720 -3350 4760 -3340
rect 4720 -3430 4725 -3350
rect 4755 -3430 4760 -3350
rect 4720 -3440 4760 -3430
rect 5040 -3350 5080 -2835
rect 5280 -2805 5480 -2800
rect 5280 -2835 5290 -2805
rect 5470 -2835 5480 -2805
rect 5280 -2840 5480 -2835
rect 5600 -2805 5800 -2800
rect 5600 -2835 5610 -2805
rect 5790 -2835 5800 -2805
rect 5600 -2840 5800 -2835
rect 5920 -2805 6120 -2800
rect 5920 -2835 5930 -2805
rect 6110 -2835 6120 -2805
rect 5920 -2840 6120 -2835
rect 6240 -2805 6440 -2800
rect 6240 -2835 6250 -2805
rect 6430 -2835 6440 -2805
rect 6240 -2840 6440 -2835
rect 5360 -2965 5400 -2960
rect 5360 -2995 5365 -2965
rect 5395 -2995 5400 -2965
rect 5360 -3280 5400 -2995
rect 5520 -2965 5560 -2960
rect 5520 -2995 5525 -2965
rect 5555 -2995 5560 -2965
rect 5280 -3285 5480 -3280
rect 5280 -3315 5290 -3285
rect 5470 -3315 5480 -3285
rect 5280 -3320 5480 -3315
rect 5040 -3430 5045 -3350
rect 5075 -3430 5080 -3350
rect 5040 -3440 5080 -3430
rect 5200 -3350 5240 -3340
rect 5200 -3430 5205 -3350
rect 5235 -3430 5240 -3350
rect -80 -3475 -75 -3445
rect -45 -3475 -40 -3445
rect -80 -3480 -40 -3475
rect 5200 -3445 5240 -3430
rect 5520 -3350 5560 -2995
rect 5680 -2965 5720 -2960
rect 5680 -2995 5685 -2965
rect 5715 -2995 5720 -2965
rect 5680 -3280 5720 -2995
rect 6000 -2965 6040 -2960
rect 6000 -2995 6005 -2965
rect 6035 -2995 6040 -2965
rect 6000 -3280 6040 -2995
rect 6160 -2965 6200 -2960
rect 6160 -2995 6165 -2965
rect 6195 -2995 6200 -2965
rect 6160 -3280 6200 -2995
rect 6320 -2965 6360 -2960
rect 6320 -2995 6325 -2965
rect 6355 -2995 6360 -2965
rect 6320 -3280 6360 -2995
rect 6480 -2965 6520 -2770
rect 6800 -2690 6840 -2680
rect 6800 -2770 6805 -2690
rect 6835 -2770 6840 -2690
rect 6800 -2780 6840 -2770
rect 7120 -2690 7160 -2680
rect 7120 -2770 7125 -2690
rect 7155 -2770 7160 -2690
rect 7120 -2780 7160 -2770
rect 7440 -2690 7480 -2680
rect 7440 -2770 7445 -2690
rect 7475 -2770 7480 -2690
rect 7440 -2780 7480 -2770
rect 7760 -2690 7800 -2675
rect 10320 -2645 10360 -2640
rect 10320 -2675 10325 -2645
rect 10355 -2675 10360 -2645
rect 7760 -2770 7765 -2690
rect 7795 -2770 7800 -2690
rect 7760 -2780 7800 -2770
rect 8080 -2690 8120 -2680
rect 8080 -2770 8085 -2690
rect 8115 -2770 8120 -2690
rect 8080 -2780 8120 -2770
rect 8400 -2690 8440 -2680
rect 8400 -2770 8405 -2690
rect 8435 -2770 8440 -2690
rect 8400 -2780 8440 -2770
rect 8720 -2690 8760 -2680
rect 8720 -2770 8725 -2690
rect 8755 -2770 8760 -2690
rect 8720 -2780 8760 -2770
rect 9040 -2690 9080 -2680
rect 9040 -2770 9045 -2690
rect 9075 -2770 9080 -2690
rect 6560 -2805 6760 -2800
rect 6560 -2835 6570 -2805
rect 6750 -2835 6760 -2805
rect 6560 -2840 6760 -2835
rect 6880 -2805 7080 -2800
rect 6880 -2835 6890 -2805
rect 7070 -2835 7080 -2805
rect 6880 -2840 7080 -2835
rect 7200 -2805 7400 -2800
rect 7200 -2835 7210 -2805
rect 7390 -2835 7400 -2805
rect 7200 -2840 7400 -2835
rect 7520 -2805 7720 -2800
rect 7520 -2835 7530 -2805
rect 7710 -2835 7720 -2805
rect 7520 -2840 7720 -2835
rect 7840 -2805 8040 -2800
rect 7840 -2835 7850 -2805
rect 8030 -2835 8040 -2805
rect 7840 -2840 8040 -2835
rect 8160 -2805 8360 -2800
rect 8160 -2835 8170 -2805
rect 8350 -2835 8360 -2805
rect 8160 -2840 8360 -2835
rect 8480 -2805 8680 -2800
rect 8480 -2835 8490 -2805
rect 8670 -2835 8680 -2805
rect 8480 -2840 8680 -2835
rect 8800 -2805 9000 -2800
rect 8800 -2835 8810 -2805
rect 8990 -2835 9000 -2805
rect 8800 -2840 9000 -2835
rect 6480 -2995 6485 -2965
rect 6515 -2995 6520 -2965
rect 6480 -3000 6520 -2995
rect 6640 -2965 6680 -2960
rect 6640 -2995 6645 -2965
rect 6675 -2995 6680 -2965
rect 6640 -3280 6680 -2995
rect 6800 -2965 6840 -2960
rect 6800 -2995 6805 -2965
rect 6835 -2995 6840 -2965
rect 6800 -3280 6840 -2995
rect 6960 -2965 7000 -2960
rect 6960 -2995 6965 -2965
rect 6995 -2995 7000 -2965
rect 6960 -3280 7000 -2995
rect 7280 -2965 7320 -2960
rect 7280 -2995 7285 -2965
rect 7315 -2995 7320 -2965
rect 7280 -3280 7320 -2995
rect 7440 -2965 7480 -2960
rect 7440 -2995 7445 -2965
rect 7475 -2995 7480 -2965
rect 7440 -3280 7480 -2995
rect 7600 -2965 7640 -2960
rect 7600 -2995 7605 -2965
rect 7635 -2995 7640 -2965
rect 7600 -3280 7640 -2995
rect 7920 -2965 7960 -2960
rect 7920 -2995 7925 -2965
rect 7955 -2995 7960 -2965
rect 7920 -3280 7960 -2995
rect 8080 -2965 8120 -2960
rect 8080 -2995 8085 -2965
rect 8115 -2995 8120 -2965
rect 5600 -3285 5800 -3280
rect 5600 -3315 5610 -3285
rect 5790 -3315 5800 -3285
rect 5600 -3320 5800 -3315
rect 5920 -3285 6120 -3280
rect 5920 -3315 5930 -3285
rect 6110 -3315 6120 -3285
rect 5920 -3320 6120 -3315
rect 6240 -3285 6440 -3280
rect 6240 -3315 6250 -3285
rect 6430 -3315 6440 -3285
rect 6240 -3320 6440 -3315
rect 6560 -3285 6760 -3280
rect 6560 -3315 6570 -3285
rect 6750 -3315 6760 -3285
rect 6560 -3320 6760 -3315
rect 6880 -3285 7080 -3280
rect 6880 -3315 6890 -3285
rect 7070 -3315 7080 -3285
rect 6880 -3320 7080 -3315
rect 7200 -3285 7400 -3280
rect 7200 -3315 7210 -3285
rect 7390 -3315 7400 -3285
rect 7200 -3320 7400 -3315
rect 7520 -3285 7720 -3280
rect 7520 -3315 7530 -3285
rect 7710 -3315 7720 -3285
rect 7520 -3320 7720 -3315
rect 7840 -3285 8040 -3280
rect 7840 -3315 7850 -3285
rect 8030 -3315 8040 -3285
rect 7840 -3320 8040 -3315
rect 5520 -3430 5525 -3350
rect 5555 -3430 5560 -3350
rect 5520 -3440 5560 -3430
rect 5840 -3350 5880 -3340
rect 5840 -3430 5845 -3350
rect 5875 -3430 5880 -3350
rect 5200 -3475 5205 -3445
rect 5235 -3475 5240 -3445
rect 5200 -3480 5240 -3475
rect 5840 -3445 5880 -3430
rect 6160 -3350 6200 -3340
rect 6160 -3430 6165 -3350
rect 6195 -3430 6200 -3350
rect 6160 -3440 6200 -3430
rect 6480 -3350 6520 -3340
rect 6480 -3430 6485 -3350
rect 6515 -3430 6520 -3350
rect 5840 -3475 5845 -3445
rect 5875 -3475 5880 -3445
rect 5840 -3480 5880 -3475
rect 6480 -3445 6520 -3430
rect 6800 -3350 6840 -3340
rect 6800 -3430 6805 -3350
rect 6835 -3430 6840 -3350
rect 6800 -3440 6840 -3430
rect 7120 -3350 7160 -3340
rect 7120 -3430 7125 -3350
rect 7155 -3430 7160 -3350
rect 6480 -3475 6485 -3445
rect 6515 -3475 6520 -3445
rect 6480 -3480 6520 -3475
rect 7120 -3445 7160 -3430
rect 7440 -3350 7480 -3340
rect 7440 -3430 7445 -3350
rect 7475 -3430 7480 -3350
rect 7440 -3440 7480 -3430
rect 7760 -3350 7800 -3340
rect 7760 -3430 7765 -3350
rect 7795 -3430 7800 -3350
rect 7120 -3475 7125 -3445
rect 7155 -3475 7160 -3445
rect 7120 -3480 7160 -3475
rect 7760 -3445 7800 -3430
rect 8080 -3350 8120 -2995
rect 8240 -2965 8280 -2960
rect 8240 -2995 8245 -2965
rect 8275 -2995 8280 -2965
rect 8240 -3280 8280 -2995
rect 8560 -2965 8600 -2960
rect 8560 -2995 8565 -2965
rect 8595 -2995 8600 -2965
rect 8560 -3280 8600 -2995
rect 8720 -2965 8760 -2960
rect 8720 -2995 8725 -2965
rect 8755 -2995 8760 -2965
rect 8160 -3285 8360 -3280
rect 8160 -3315 8170 -3285
rect 8350 -3315 8360 -3285
rect 8160 -3320 8360 -3315
rect 8480 -3285 8680 -3280
rect 8480 -3315 8490 -3285
rect 8670 -3315 8680 -3285
rect 8480 -3320 8680 -3315
rect 8080 -3430 8085 -3350
rect 8115 -3430 8120 -3350
rect 8080 -3440 8120 -3430
rect 8400 -3350 8440 -3340
rect 8400 -3430 8405 -3350
rect 8435 -3430 8440 -3350
rect 7760 -3475 7765 -3445
rect 7795 -3475 7800 -3445
rect 7760 -3480 7800 -3475
rect 8400 -3445 8440 -3430
rect 8720 -3350 8760 -2995
rect 8880 -2965 8920 -2960
rect 8880 -2995 8885 -2965
rect 8915 -2995 8920 -2965
rect 8880 -3280 8920 -2995
rect 9040 -2965 9080 -2770
rect 9360 -2690 9400 -2680
rect 9360 -2770 9365 -2690
rect 9395 -2770 9400 -2690
rect 9360 -2780 9400 -2770
rect 9680 -2690 9720 -2680
rect 9680 -2770 9685 -2690
rect 9715 -2770 9720 -2690
rect 9680 -2780 9720 -2770
rect 10000 -2690 10040 -2680
rect 10000 -2770 10005 -2690
rect 10035 -2770 10040 -2690
rect 10000 -2780 10040 -2770
rect 10320 -2690 10360 -2675
rect 10640 -2645 10680 -2640
rect 10640 -2675 10645 -2645
rect 10675 -2675 10680 -2645
rect 10640 -2680 10680 -2675
rect 10800 -2645 10840 -2640
rect 10800 -2675 10805 -2645
rect 10835 -2675 10840 -2645
rect 10800 -2680 10840 -2675
rect 10960 -2645 11000 -2640
rect 10960 -2675 10965 -2645
rect 10995 -2675 11000 -2645
rect 10960 -2680 11000 -2675
rect 10320 -2770 10325 -2690
rect 10355 -2770 10360 -2690
rect 10640 -2725 10680 -2720
rect 10640 -2755 10645 -2725
rect 10675 -2755 10680 -2725
rect 10640 -2760 10680 -2755
rect 10800 -2725 10840 -2720
rect 10800 -2755 10805 -2725
rect 10835 -2755 10840 -2725
rect 10800 -2760 10840 -2755
rect 10960 -2725 11000 -2720
rect 10960 -2755 10965 -2725
rect 10995 -2755 11000 -2725
rect 10960 -2760 11000 -2755
rect 10320 -2780 10360 -2770
rect 9120 -2805 9320 -2800
rect 9120 -2835 9130 -2805
rect 9310 -2835 9320 -2805
rect 9120 -2840 9320 -2835
rect 9440 -2805 9640 -2800
rect 9440 -2835 9450 -2805
rect 9630 -2835 9640 -2805
rect 9440 -2840 9640 -2835
rect 9760 -2805 9960 -2800
rect 9760 -2835 9770 -2805
rect 9950 -2835 9960 -2805
rect 9760 -2840 9960 -2835
rect 10080 -2805 10280 -2800
rect 10080 -2835 10090 -2805
rect 10270 -2835 10280 -2805
rect 10080 -2840 10280 -2835
rect 10800 -2805 10840 -2800
rect 10800 -2835 10805 -2805
rect 10835 -2835 10840 -2805
rect 10800 -2840 10840 -2835
rect 10960 -2805 11000 -2800
rect 10960 -2835 10965 -2805
rect 10995 -2835 11000 -2805
rect 10960 -2840 11000 -2835
rect 10640 -2885 10680 -2880
rect 10640 -2915 10645 -2885
rect 10675 -2915 10680 -2885
rect 10640 -2920 10680 -2915
rect 10800 -2885 10840 -2880
rect 10800 -2915 10805 -2885
rect 10835 -2915 10840 -2885
rect 10800 -2920 10840 -2915
rect 10960 -2885 11000 -2880
rect 10960 -2915 10965 -2885
rect 10995 -2915 11000 -2885
rect 10960 -2920 11000 -2915
rect 9040 -2995 9045 -2965
rect 9075 -2995 9080 -2965
rect 9040 -3000 9080 -2995
rect 9200 -2965 9240 -2960
rect 9200 -2995 9205 -2965
rect 9235 -2995 9240 -2965
rect 9200 -3280 9240 -2995
rect 9360 -2965 9400 -2960
rect 9360 -2995 9365 -2965
rect 9395 -2995 9400 -2965
rect 8800 -3285 9000 -3280
rect 8800 -3315 8810 -3285
rect 8990 -3315 9000 -3285
rect 8800 -3320 9000 -3315
rect 9120 -3285 9320 -3280
rect 9120 -3315 9130 -3285
rect 9310 -3315 9320 -3285
rect 9120 -3320 9320 -3315
rect 8720 -3430 8725 -3350
rect 8755 -3430 8760 -3350
rect 8720 -3440 8760 -3430
rect 9040 -3350 9080 -3340
rect 9040 -3430 9045 -3350
rect 9075 -3430 9080 -3350
rect 8400 -3475 8405 -3445
rect 8435 -3475 8440 -3445
rect 8400 -3480 8440 -3475
rect 9040 -3445 9080 -3430
rect 9360 -3350 9400 -2995
rect 9520 -2965 9560 -2960
rect 9520 -2995 9525 -2965
rect 9555 -2995 9560 -2965
rect 9520 -3280 9560 -2995
rect 9840 -2965 9880 -2960
rect 9840 -2995 9845 -2965
rect 9875 -2995 9880 -2965
rect 9840 -3280 9880 -2995
rect 10000 -2965 10040 -2960
rect 10000 -2995 10005 -2965
rect 10035 -2995 10040 -2965
rect 9440 -3285 9640 -3280
rect 9440 -3315 9450 -3285
rect 9630 -3315 9640 -3285
rect 9440 -3320 9640 -3315
rect 9760 -3285 9960 -3280
rect 9760 -3315 9770 -3285
rect 9950 -3315 9960 -3285
rect 9760 -3320 9960 -3315
rect 9360 -3430 9365 -3350
rect 9395 -3430 9400 -3350
rect 9360 -3440 9400 -3430
rect 9680 -3350 9720 -3340
rect 9680 -3430 9685 -3350
rect 9715 -3430 9720 -3350
rect 9040 -3475 9045 -3445
rect 9075 -3475 9080 -3445
rect 9040 -3480 9080 -3475
rect 9680 -3445 9720 -3430
rect 10000 -3350 10040 -2995
rect 10160 -2965 10200 -2960
rect 10160 -2995 10165 -2965
rect 10195 -2995 10200 -2965
rect 10160 -3280 10200 -2995
rect 10640 -3045 10680 -3040
rect 10640 -3075 10645 -3045
rect 10675 -3075 10680 -3045
rect 10640 -3080 10680 -3075
rect 10800 -3045 10840 -3040
rect 10800 -3075 10805 -3045
rect 10835 -3075 10840 -3045
rect 10800 -3080 10840 -3075
rect 10960 -3045 11000 -3040
rect 10960 -3075 10965 -3045
rect 10995 -3075 11000 -3045
rect 10960 -3080 11000 -3075
rect 10640 -3125 10680 -3120
rect 10640 -3155 10645 -3125
rect 10675 -3155 10680 -3125
rect 10640 -3160 10680 -3155
rect 10800 -3125 10840 -3120
rect 10800 -3155 10805 -3125
rect 10835 -3155 10840 -3125
rect 10800 -3160 10840 -3155
rect 10960 -3125 11000 -3120
rect 10960 -3155 10965 -3125
rect 10995 -3155 11000 -3125
rect 10960 -3160 11000 -3155
rect 10640 -3205 10680 -3200
rect 10640 -3235 10645 -3205
rect 10675 -3235 10680 -3205
rect 10640 -3240 10680 -3235
rect 10800 -3205 10840 -3200
rect 10800 -3235 10805 -3205
rect 10835 -3235 10840 -3205
rect 10800 -3240 10840 -3235
rect 10960 -3205 11000 -3200
rect 10960 -3235 10965 -3205
rect 10995 -3235 11000 -3205
rect 10960 -3240 11000 -3235
rect 10080 -3285 10280 -3280
rect 10080 -3315 10090 -3285
rect 10270 -3315 10280 -3285
rect 10080 -3320 10280 -3315
rect 10640 -3285 10680 -3280
rect 10640 -3315 10645 -3285
rect 10675 -3315 10680 -3285
rect 10640 -3320 10680 -3315
rect 10800 -3285 10840 -3280
rect 10800 -3315 10805 -3285
rect 10835 -3315 10840 -3285
rect 10800 -3320 10840 -3315
rect 10960 -3285 11000 -3280
rect 10960 -3315 10965 -3285
rect 10995 -3315 11000 -3285
rect 10960 -3320 11000 -3315
rect 10000 -3430 10005 -3350
rect 10035 -3430 10040 -3350
rect 10000 -3440 10040 -3430
rect 10320 -3350 10360 -3340
rect 10320 -3430 10325 -3350
rect 10355 -3430 10360 -3350
rect 10640 -3365 10680 -3360
rect 10640 -3395 10645 -3365
rect 10675 -3395 10680 -3365
rect 10640 -3400 10680 -3395
rect 10800 -3365 10840 -3360
rect 10800 -3395 10805 -3365
rect 10835 -3395 10840 -3365
rect 10800 -3400 10840 -3395
rect 10960 -3365 11000 -3360
rect 10960 -3395 10965 -3365
rect 10995 -3395 11000 -3365
rect 10960 -3400 11000 -3395
rect 9680 -3475 9685 -3445
rect 9715 -3475 9720 -3445
rect 9680 -3480 9720 -3475
rect 10320 -3445 10360 -3430
rect 10320 -3475 10325 -3445
rect 10355 -3475 10360 -3445
rect 10320 -3480 10360 -3475
rect 10640 -3445 10680 -3440
rect 10640 -3475 10645 -3445
rect 10675 -3475 10680 -3445
rect 10640 -3480 10680 -3475
rect 10800 -3445 10840 -3440
rect 10800 -3475 10805 -3445
rect 10835 -3475 10840 -3445
rect 10800 -3480 10840 -3475
rect 10960 -3445 11000 -3440
rect 10960 -3475 10965 -3445
rect 10995 -3475 11000 -3445
rect 10960 -3480 11000 -3475
rect -720 -3525 -680 -3520
rect -720 -3555 -715 -3525
rect -685 -3555 -680 -3525
rect -720 -3560 -680 -3555
rect -560 -3525 -520 -3520
rect -560 -3555 -555 -3525
rect -525 -3555 -520 -3525
rect -560 -3560 -520 -3555
rect -400 -3525 -360 -3520
rect -400 -3555 -395 -3525
rect -365 -3555 -360 -3525
rect -400 -3560 -360 -3555
rect 10640 -3525 10680 -3520
rect 10640 -3555 10645 -3525
rect 10675 -3555 10680 -3525
rect 10640 -3560 10680 -3555
rect 10800 -3525 10840 -3520
rect 10800 -3555 10805 -3525
rect 10835 -3555 10840 -3525
rect 10800 -3560 10840 -3555
rect 10960 -3525 11000 -3520
rect 10960 -3555 10965 -3525
rect 10995 -3555 11000 -3525
rect 10960 -3560 11000 -3555
rect -720 -3605 -680 -3600
rect -720 -3635 -715 -3605
rect -685 -3635 -680 -3605
rect -720 -3640 -680 -3635
rect -560 -3605 -520 -3600
rect -560 -3635 -555 -3605
rect -525 -3635 -520 -3605
rect -560 -3640 -520 -3635
rect -400 -3605 -360 -3600
rect -400 -3635 -395 -3605
rect -365 -3635 -360 -3605
rect -400 -3640 -360 -3635
rect 10640 -3605 10680 -3600
rect 10640 -3635 10645 -3605
rect 10675 -3635 10680 -3605
rect 10640 -3640 10680 -3635
rect 10800 -3605 10840 -3600
rect 10800 -3635 10805 -3605
rect 10835 -3635 10840 -3605
rect 10800 -3640 10840 -3635
rect 10960 -3605 11000 -3600
rect 10960 -3635 10965 -3605
rect 10995 -3635 11000 -3605
rect 10960 -3640 11000 -3635
rect -720 -3685 -680 -3680
rect -720 -3715 -715 -3685
rect -685 -3715 -680 -3685
rect -720 -3720 -680 -3715
rect -560 -3685 -520 -3680
rect -560 -3715 -555 -3685
rect -525 -3715 -520 -3685
rect -560 -3720 -520 -3715
rect -400 -3685 -360 -3680
rect -400 -3715 -395 -3685
rect -365 -3715 -360 -3685
rect -400 -3720 -360 -3715
rect 10640 -3685 10680 -3680
rect 10640 -3715 10645 -3685
rect 10675 -3715 10680 -3685
rect 10640 -3720 10680 -3715
rect 10800 -3685 10840 -3680
rect 10800 -3715 10805 -3685
rect 10835 -3715 10840 -3685
rect 10800 -3720 10840 -3715
rect 10960 -3685 11000 -3680
rect 10960 -3715 10965 -3685
rect 10995 -3715 11000 -3685
rect 10960 -3720 11000 -3715
<< via1 >>
rect -715 1005 -685 1035
rect -555 1005 -525 1035
rect -395 1005 -365 1035
rect 10645 1005 10675 1035
rect 10805 1005 10835 1035
rect 10965 1005 10995 1035
rect -715 925 -685 955
rect -555 925 -525 955
rect -395 925 -365 955
rect 10645 925 10675 955
rect 10805 925 10835 955
rect 10965 925 10995 955
rect -715 845 -685 875
rect -555 845 -525 875
rect -395 845 -365 875
rect 10645 845 10675 875
rect 10805 845 10835 875
rect 10965 845 10995 875
rect -75 765 -45 795
rect 5205 765 5235 795
rect -75 685 -45 715
rect -715 605 -685 635
rect -555 605 -525 635
rect -395 605 -365 635
rect -715 525 -685 555
rect -555 525 -525 555
rect -395 525 -365 555
rect -715 445 -685 475
rect -555 445 -525 475
rect 85 445 115 475
rect 405 445 435 475
rect 725 445 755 475
rect 1045 445 1075 475
rect 1365 445 1395 475
rect 1685 445 1715 475
rect 2005 445 2035 475
rect 2325 445 2355 475
rect 2645 445 2675 475
rect 2965 445 2995 475
rect 3285 445 3315 475
rect 3605 445 3635 475
rect 3925 445 3955 475
rect 4245 445 4275 475
rect 4565 445 4595 475
rect 4885 445 4915 475
rect -715 365 -685 395
rect -555 365 -525 395
rect -395 365 -365 395
rect -715 285 -685 315
rect -555 285 -525 315
rect -395 285 -365 315
rect -715 205 -685 235
rect -555 205 -525 235
rect -395 205 -365 235
rect -715 125 -685 155
rect -555 125 -525 155
rect -395 125 -365 155
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect 1205 125 1235 155
rect -715 45 -685 75
rect -555 45 -525 75
rect -395 45 -365 75
rect -75 45 -45 75
rect -715 -35 -685 -5
rect -555 -35 -525 -5
rect -395 -35 -365 -5
rect 1290 125 1470 155
rect 1610 125 1790 155
rect 1930 125 2110 155
rect 2250 125 2430 155
rect 2570 125 2750 155
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3765 125 3795 155
rect 2485 45 2515 75
rect -75 -35 -45 -5
rect 3850 125 4030 155
rect 4170 125 4350 155
rect 4490 125 4670 155
rect 4810 125 4990 155
rect 5845 765 5875 795
rect 5205 685 5235 715
rect 5365 285 5395 315
rect 6485 765 6515 795
rect 5845 685 5875 715
rect 7125 765 7155 795
rect 6485 685 6515 715
rect 7765 765 7795 795
rect 7125 685 7155 715
rect 8405 765 8435 795
rect 7765 685 7795 715
rect 5525 285 5555 315
rect 5685 285 5715 315
rect 6005 285 6035 315
rect 6165 285 6195 315
rect 6325 285 6355 315
rect 6485 285 6515 315
rect 5045 125 5075 155
rect 5290 125 5470 155
rect 5610 125 5790 155
rect 5930 125 6110 155
rect 6250 125 6430 155
rect 5045 45 5075 75
rect 2485 -35 2515 -5
rect 5045 -35 5075 -5
rect 5205 45 5235 75
rect 6645 285 6675 315
rect 6805 285 6835 315
rect 6965 285 6995 315
rect 7285 285 7315 315
rect 7445 285 7475 315
rect 7605 285 7635 315
rect 7925 285 7955 315
rect 9045 765 9075 795
rect 8405 685 8435 715
rect 8085 285 8115 315
rect 8245 285 8275 315
rect 8565 285 8595 315
rect 9685 765 9715 795
rect 9045 685 9075 715
rect 8725 285 8755 315
rect 8885 285 8915 315
rect 9045 285 9075 315
rect 6570 125 6750 155
rect 6890 125 7070 155
rect 7210 125 7390 155
rect 7530 125 7710 155
rect 7850 125 8030 155
rect 8170 125 8350 155
rect 8490 125 8670 155
rect 8810 125 8990 155
rect 7765 45 7795 75
rect 5205 -35 5235 -5
rect 9205 285 9235 315
rect 10325 765 10355 795
rect 9685 685 9715 715
rect 9365 285 9395 315
rect 9525 285 9555 315
rect 9845 285 9875 315
rect 10645 765 10675 795
rect 10805 765 10835 795
rect 10965 765 10995 795
rect 10325 685 10355 715
rect 10645 685 10675 715
rect 10805 685 10835 715
rect 10965 685 10995 715
rect 10645 605 10675 635
rect 10805 605 10835 635
rect 10965 605 10995 635
rect 10005 285 10035 315
rect 10645 525 10675 555
rect 10805 525 10835 555
rect 10965 525 10995 555
rect 10645 445 10675 475
rect 10805 445 10835 475
rect 10965 445 10995 475
rect 10645 365 10675 395
rect 10805 365 10835 395
rect 10965 365 10995 395
rect 10165 285 10195 315
rect 10645 205 10675 235
rect 10805 205 10835 235
rect 10965 205 10995 235
rect 9130 125 9310 155
rect 9450 125 9630 155
rect 9770 125 9950 155
rect 10090 125 10270 155
rect 10805 125 10835 155
rect 10965 125 10995 155
rect 10325 45 10355 75
rect 10645 45 10675 75
rect 10805 45 10835 75
rect 10965 45 10995 75
rect 7765 -35 7795 -5
rect 10325 -35 10355 -5
rect 10645 -35 10675 -5
rect 10805 -35 10835 -5
rect 10965 -35 10995 -5
rect -715 -115 -685 -85
rect -555 -115 -525 -85
rect -395 -115 -365 -85
rect 10645 -115 10675 -85
rect 10805 -115 10835 -85
rect 10965 -115 10995 -85
rect -715 -195 -685 -165
rect -555 -195 -525 -165
rect -395 -195 -365 -165
rect 10645 -195 10675 -165
rect 10805 -195 10835 -165
rect 10965 -195 10995 -165
rect -715 -275 -685 -245
rect -555 -275 -525 -245
rect -395 -275 -365 -245
rect -75 -275 -45 -245
rect 2485 -275 2515 -245
rect -715 -355 -685 -325
rect -555 -355 -525 -325
rect -395 -355 -365 -325
rect -75 -355 -45 -325
rect -715 -435 -685 -405
rect -555 -435 -525 -405
rect -395 -435 -365 -405
rect 10 -435 190 -405
rect 330 -435 510 -405
rect 650 -435 830 -405
rect 970 -435 1150 -405
rect -715 -515 -685 -485
rect -555 -515 -525 -485
rect -395 -515 -365 -485
rect -715 -595 -685 -565
rect -555 -595 -525 -565
rect -395 -595 -365 -565
rect 85 -595 115 -565
rect -715 -675 -685 -645
rect -555 -675 -525 -645
rect -395 -675 -365 -645
rect -715 -755 -685 -725
rect -555 -755 -525 -725
rect -715 -835 -685 -805
rect -555 -835 -525 -805
rect -395 -835 -365 -805
rect 245 -595 275 -565
rect -715 -915 -685 -885
rect -555 -915 -525 -885
rect -395 -915 -365 -885
rect -75 -995 -45 -965
rect 405 -595 435 -565
rect 725 -595 755 -565
rect 885 -595 915 -565
rect 565 -995 595 -965
rect -75 -1075 -45 -1045
rect 1045 -595 1075 -565
rect 5045 -275 5075 -245
rect 2485 -355 2515 -325
rect 1290 -435 1470 -405
rect 1610 -435 1790 -405
rect 1930 -435 2110 -405
rect 2250 -435 2430 -405
rect 2570 -435 2750 -405
rect 2890 -435 3070 -405
rect 3210 -435 3390 -405
rect 3530 -435 3710 -405
rect 1205 -595 1235 -565
rect 1365 -595 1395 -565
rect 1525 -595 1555 -565
rect 1205 -995 1235 -965
rect 565 -1075 595 -1045
rect 1685 -595 1715 -565
rect 2005 -595 2035 -565
rect 2165 -595 2195 -565
rect 1845 -995 1875 -965
rect 1205 -1075 1235 -1045
rect 2325 -595 2355 -565
rect 2645 -595 2675 -565
rect 2805 -595 2835 -565
rect 2485 -995 2515 -965
rect 1845 -1075 1875 -1045
rect 2965 -595 2995 -565
rect 3285 -595 3315 -565
rect 3445 -595 3475 -565
rect 3125 -995 3155 -965
rect 2485 -1075 2515 -1045
rect 3605 -595 3635 -565
rect 5045 -355 5075 -325
rect 5205 -275 5235 -245
rect 7765 -275 7795 -245
rect 5205 -355 5235 -325
rect 3850 -435 4030 -405
rect 4170 -435 4350 -405
rect 4490 -435 4670 -405
rect 4810 -435 4990 -405
rect 5205 -435 5235 -405
rect 3765 -595 3795 -565
rect 3925 -595 3955 -565
rect 4085 -595 4115 -565
rect 3765 -995 3795 -965
rect 3125 -1075 3155 -1045
rect 4245 -595 4275 -565
rect 4565 -595 4595 -565
rect 4725 -595 4755 -565
rect 4405 -995 4435 -965
rect 3765 -1075 3795 -1045
rect 4885 -595 4915 -565
rect 5045 -995 5075 -965
rect 4405 -1075 4435 -1045
rect 5290 -435 5470 -405
rect 5610 -435 5790 -405
rect 5930 -435 6110 -405
rect 6250 -435 6430 -405
rect 10325 -275 10355 -245
rect 7765 -355 7795 -325
rect 6485 -435 6515 -405
rect 6570 -435 6750 -405
rect 6890 -435 7070 -405
rect 7210 -435 7390 -405
rect 7530 -435 7710 -405
rect 7850 -435 8030 -405
rect 8170 -435 8350 -405
rect 8490 -435 8670 -405
rect 8810 -435 8990 -405
rect 10645 -275 10675 -245
rect 10805 -275 10835 -245
rect 10965 -275 10995 -245
rect 10325 -355 10355 -325
rect 10645 -355 10675 -325
rect 10805 -355 10835 -325
rect 10965 -355 10995 -325
rect 9045 -435 9075 -405
rect 9130 -435 9310 -405
rect 9450 -435 9630 -405
rect 9770 -435 9950 -405
rect 10090 -435 10270 -405
rect 10805 -435 10835 -405
rect 10965 -435 10995 -405
rect 10645 -515 10675 -485
rect 10805 -515 10835 -485
rect 10965 -515 10995 -485
rect 10645 -675 10675 -645
rect 10805 -675 10835 -645
rect 10965 -675 10995 -645
rect 5365 -755 5395 -725
rect 5685 -755 5715 -725
rect 6005 -755 6035 -725
rect 6325 -755 6355 -725
rect 6645 -755 6675 -725
rect 6965 -755 6995 -725
rect 7285 -755 7315 -725
rect 7605 -755 7635 -725
rect 7925 -755 7955 -725
rect 8245 -755 8275 -725
rect 8565 -755 8595 -725
rect 8885 -755 8915 -725
rect 9205 -755 9235 -725
rect 9525 -755 9555 -725
rect 9845 -755 9875 -725
rect 10165 -755 10195 -725
rect 10645 -755 10675 -725
rect 10805 -755 10835 -725
rect 10965 -755 10995 -725
rect 10645 -835 10675 -805
rect 10805 -835 10835 -805
rect 10965 -835 10995 -805
rect 10645 -915 10675 -885
rect 10805 -915 10835 -885
rect 10965 -915 10995 -885
rect 10325 -995 10355 -965
rect 10645 -995 10675 -965
rect 10805 -995 10835 -965
rect 10965 -995 10995 -965
rect 5045 -1075 5075 -1045
rect 10325 -1075 10355 -1045
rect 10645 -1075 10675 -1045
rect 10805 -1075 10835 -1045
rect 10965 -1075 10995 -1045
rect -715 -1155 -685 -1125
rect -555 -1155 -525 -1125
rect -395 -1155 -365 -1125
rect 10645 -1155 10675 -1125
rect 10805 -1155 10835 -1125
rect 10965 -1155 10995 -1125
rect -715 -1235 -685 -1205
rect -555 -1235 -525 -1205
rect -395 -1235 -365 -1205
rect 10645 -1235 10675 -1205
rect 10805 -1235 10835 -1205
rect 10965 -1235 10995 -1205
rect -715 -1315 -685 -1285
rect -555 -1315 -525 -1285
rect -395 -1315 -365 -1285
rect 10645 -1315 10675 -1285
rect 10805 -1315 10835 -1285
rect 10965 -1315 10995 -1285
rect -715 -1395 -685 -1365
rect -555 -1395 -525 -1365
rect -395 -1395 -365 -1365
rect 10645 -1395 10675 -1365
rect 10805 -1395 10835 -1365
rect 10965 -1395 10995 -1365
rect -715 -1475 -685 -1445
rect -555 -1475 -525 -1445
rect -395 -1475 -365 -1445
rect 10645 -1475 10675 -1445
rect 10805 -1475 10835 -1445
rect 10965 -1475 10995 -1445
rect -715 -1555 -685 -1525
rect -555 -1555 -525 -1525
rect -395 -1555 -365 -1525
rect 10645 -1555 10675 -1525
rect 10805 -1555 10835 -1525
rect 10965 -1555 10995 -1525
rect -75 -1635 -45 -1605
rect 565 -1635 595 -1605
rect -75 -1715 -45 -1685
rect -715 -1795 -685 -1765
rect -555 -1795 -525 -1765
rect -395 -1795 -365 -1765
rect -715 -1875 -685 -1845
rect -555 -1875 -525 -1845
rect -395 -1875 -365 -1845
rect -715 -1955 -685 -1925
rect -555 -1955 -525 -1925
rect -715 -2035 -685 -2005
rect -555 -2035 -525 -2005
rect -395 -2035 -365 -2005
rect -715 -2115 -685 -2085
rect -555 -2115 -525 -2085
rect -395 -2115 -365 -2085
rect 85 -2115 115 -2085
rect 1205 -1635 1235 -1605
rect 565 -1715 595 -1685
rect 245 -2115 275 -2085
rect 405 -2115 435 -2085
rect 725 -2115 755 -2085
rect 1845 -1635 1875 -1605
rect 1205 -1715 1235 -1685
rect 885 -2115 915 -2085
rect 1045 -2115 1075 -2085
rect 1205 -2115 1235 -2085
rect -715 -2195 -685 -2165
rect -555 -2195 -525 -2165
rect -395 -2195 -365 -2165
rect -715 -2275 -685 -2245
rect -555 -2275 -525 -2245
rect -395 -2275 -365 -2245
rect 10 -2275 190 -2245
rect 330 -2275 510 -2245
rect 650 -2275 830 -2245
rect 970 -2275 1150 -2245
rect -715 -2355 -685 -2325
rect -555 -2355 -525 -2325
rect -395 -2355 -365 -2325
rect -75 -2355 -45 -2325
rect -715 -2435 -685 -2405
rect -555 -2435 -525 -2405
rect -395 -2435 -365 -2405
rect 1365 -2115 1395 -2085
rect 2485 -1635 2515 -1605
rect 1845 -1715 1875 -1685
rect 1525 -2115 1555 -2085
rect 1685 -2115 1715 -2085
rect 2005 -2115 2035 -2085
rect 3125 -1635 3155 -1605
rect 2485 -1715 2515 -1685
rect 2165 -2115 2195 -2085
rect 2325 -2115 2355 -2085
rect 2645 -2115 2675 -2085
rect 3765 -1635 3795 -1605
rect 3125 -1715 3155 -1685
rect 2805 -2115 2835 -2085
rect 2965 -2115 2995 -2085
rect 3285 -2115 3315 -2085
rect 4405 -1635 4435 -1605
rect 3765 -1715 3795 -1685
rect 3445 -2115 3475 -2085
rect 3605 -2115 3635 -2085
rect 3765 -2115 3795 -2085
rect 1290 -2275 1470 -2245
rect 1610 -2275 1790 -2245
rect 1930 -2275 2110 -2245
rect 2250 -2275 2430 -2245
rect 2570 -2275 2750 -2245
rect 2890 -2275 3070 -2245
rect 3210 -2275 3390 -2245
rect 3530 -2275 3710 -2245
rect 2485 -2355 2515 -2325
rect -75 -2435 -45 -2405
rect 3925 -2115 3955 -2085
rect 5045 -1635 5075 -1605
rect 4405 -1715 4435 -1685
rect 4085 -2115 4115 -2085
rect 4245 -2115 4275 -2085
rect 4565 -2115 4595 -2085
rect 10325 -1635 10355 -1605
rect 5045 -1715 5075 -1685
rect 4725 -2115 4755 -2085
rect 4885 -2115 4915 -2085
rect 3850 -2275 4030 -2245
rect 4170 -2275 4350 -2245
rect 4490 -2275 4670 -2245
rect 4810 -2275 4990 -2245
rect 10645 -1635 10675 -1605
rect 10805 -1635 10835 -1605
rect 10965 -1635 10995 -1605
rect 10325 -1715 10355 -1685
rect 10645 -1715 10675 -1685
rect 10805 -1715 10835 -1685
rect 10965 -1715 10995 -1685
rect 10645 -1795 10675 -1765
rect 10805 -1795 10835 -1765
rect 10965 -1795 10995 -1765
rect 5365 -1955 5395 -1925
rect 5685 -1955 5715 -1925
rect 6005 -1955 6035 -1925
rect 6325 -1955 6355 -1925
rect 6645 -1955 6675 -1925
rect 6965 -1955 6995 -1925
rect 7285 -1955 7315 -1925
rect 7605 -1955 7635 -1925
rect 7925 -1955 7955 -1925
rect 8245 -1955 8275 -1925
rect 8565 -1955 8595 -1925
rect 8885 -1955 8915 -1925
rect 9205 -1955 9235 -1925
rect 9525 -1955 9555 -1925
rect 9845 -1955 9875 -1925
rect 10645 -1875 10675 -1845
rect 10805 -1875 10835 -1845
rect 10965 -1875 10995 -1845
rect 10165 -1955 10195 -1925
rect 10645 -1955 10675 -1925
rect 10805 -1955 10835 -1925
rect 10965 -1955 10995 -1925
rect 10645 -2035 10675 -2005
rect 10805 -2035 10835 -2005
rect 10965 -2035 10995 -2005
rect 10645 -2195 10675 -2165
rect 10805 -2195 10835 -2165
rect 10965 -2195 10995 -2165
rect 5205 -2275 5235 -2245
rect 5290 -2275 5470 -2245
rect 5610 -2275 5790 -2245
rect 5930 -2275 6110 -2245
rect 6250 -2275 6430 -2245
rect 6485 -2275 6515 -2245
rect 5045 -2355 5075 -2325
rect 2485 -2435 2515 -2405
rect 5045 -2435 5075 -2405
rect 5205 -2355 5235 -2325
rect 6570 -2275 6750 -2245
rect 6890 -2275 7070 -2245
rect 7210 -2275 7390 -2245
rect 7530 -2275 7710 -2245
rect 7850 -2275 8030 -2245
rect 8170 -2275 8350 -2245
rect 8490 -2275 8670 -2245
rect 8810 -2275 8990 -2245
rect 9045 -2275 9075 -2245
rect 7765 -2355 7795 -2325
rect 5205 -2435 5235 -2405
rect 9130 -2275 9310 -2245
rect 9450 -2275 9630 -2245
rect 9770 -2275 9950 -2245
rect 10090 -2275 10270 -2245
rect 10805 -2275 10835 -2245
rect 10965 -2275 10995 -2245
rect 10325 -2355 10355 -2325
rect 10645 -2355 10675 -2325
rect 10805 -2355 10835 -2325
rect 10965 -2355 10995 -2325
rect 7765 -2435 7795 -2405
rect 10325 -2435 10355 -2405
rect 10645 -2435 10675 -2405
rect 10805 -2435 10835 -2405
rect 10965 -2435 10995 -2405
rect -715 -2515 -685 -2485
rect -555 -2515 -525 -2485
rect -395 -2515 -365 -2485
rect 10645 -2515 10675 -2485
rect 10805 -2515 10835 -2485
rect 10965 -2515 10995 -2485
rect -715 -2595 -685 -2565
rect -555 -2595 -525 -2565
rect -395 -2595 -365 -2565
rect 10645 -2595 10675 -2565
rect 10805 -2595 10835 -2565
rect 10965 -2595 10995 -2565
rect -715 -2675 -685 -2645
rect -555 -2675 -525 -2645
rect -395 -2675 -365 -2645
rect -75 -2675 -45 -2645
rect 2485 -2675 2515 -2645
rect -715 -2755 -685 -2725
rect -555 -2755 -525 -2725
rect -395 -2755 -365 -2725
rect -75 -2755 -45 -2725
rect -715 -2835 -685 -2805
rect -555 -2835 -525 -2805
rect -395 -2835 -365 -2805
rect 10 -2835 190 -2805
rect 330 -2835 510 -2805
rect 650 -2835 830 -2805
rect 970 -2835 1150 -2805
rect 5045 -2675 5075 -2645
rect 2485 -2755 2515 -2725
rect 1205 -2835 1235 -2805
rect 1290 -2835 1470 -2805
rect 1610 -2835 1790 -2805
rect 1930 -2835 2110 -2805
rect 2250 -2835 2430 -2805
rect 2570 -2835 2750 -2805
rect 2890 -2835 3070 -2805
rect 3210 -2835 3390 -2805
rect 3530 -2835 3710 -2805
rect 5045 -2755 5075 -2725
rect 5205 -2675 5235 -2645
rect 7765 -2675 7795 -2645
rect 5205 -2755 5235 -2725
rect 3765 -2835 3795 -2805
rect 3850 -2835 4030 -2805
rect 4170 -2835 4350 -2805
rect 4490 -2835 4670 -2805
rect 4810 -2835 4990 -2805
rect 5045 -2835 5075 -2805
rect -715 -2915 -685 -2885
rect -555 -2915 -525 -2885
rect -395 -2915 -365 -2885
rect -715 -2995 -685 -2965
rect -555 -2995 -525 -2965
rect -395 -2995 -365 -2965
rect -715 -3075 -685 -3045
rect -555 -3075 -525 -3045
rect -395 -3075 -365 -3045
rect -715 -3155 -685 -3125
rect -555 -3155 -525 -3125
rect 85 -3155 115 -3125
rect -715 -3235 -685 -3205
rect -555 -3235 -525 -3205
rect -395 -3235 -365 -3205
rect 405 -3155 435 -3125
rect 725 -3155 755 -3125
rect 1045 -3155 1075 -3125
rect 1365 -3155 1395 -3125
rect 1685 -3155 1715 -3125
rect 2005 -3155 2035 -3125
rect 2325 -3155 2355 -3125
rect 2645 -3155 2675 -3125
rect 2965 -3155 2995 -3125
rect 3285 -3155 3315 -3125
rect 3605 -3155 3635 -3125
rect 3925 -3155 3955 -3125
rect 4245 -3155 4275 -3125
rect 4565 -3155 4595 -3125
rect 4885 -3155 4915 -3125
rect -715 -3315 -685 -3285
rect -555 -3315 -525 -3285
rect -395 -3315 -365 -3285
rect -75 -3395 -45 -3365
rect 5290 -2835 5470 -2805
rect 5610 -2835 5790 -2805
rect 5930 -2835 6110 -2805
rect 6250 -2835 6430 -2805
rect 5365 -2995 5395 -2965
rect 5525 -2995 5555 -2965
rect 5205 -3395 5235 -3365
rect -75 -3475 -45 -3445
rect 5685 -2995 5715 -2965
rect 6005 -2995 6035 -2965
rect 6165 -2995 6195 -2965
rect 6325 -2995 6355 -2965
rect 10325 -2675 10355 -2645
rect 7765 -2755 7795 -2725
rect 6570 -2835 6750 -2805
rect 6890 -2835 7070 -2805
rect 7210 -2835 7390 -2805
rect 7530 -2835 7710 -2805
rect 7850 -2835 8030 -2805
rect 8170 -2835 8350 -2805
rect 8490 -2835 8670 -2805
rect 8810 -2835 8990 -2805
rect 6485 -2995 6515 -2965
rect 6645 -2995 6675 -2965
rect 6805 -2995 6835 -2965
rect 6965 -2995 6995 -2965
rect 7285 -2995 7315 -2965
rect 7445 -2995 7475 -2965
rect 7605 -2995 7635 -2965
rect 7925 -2995 7955 -2965
rect 8085 -2995 8115 -2965
rect 5845 -3395 5875 -3365
rect 5205 -3475 5235 -3445
rect 6485 -3395 6515 -3365
rect 5845 -3475 5875 -3445
rect 7125 -3395 7155 -3365
rect 6485 -3475 6515 -3445
rect 7765 -3395 7795 -3365
rect 7125 -3475 7155 -3445
rect 8245 -2995 8275 -2965
rect 8565 -2995 8595 -2965
rect 8725 -2995 8755 -2965
rect 8405 -3395 8435 -3365
rect 7765 -3475 7795 -3445
rect 8885 -2995 8915 -2965
rect 10645 -2675 10675 -2645
rect 10805 -2675 10835 -2645
rect 10965 -2675 10995 -2645
rect 10325 -2755 10355 -2725
rect 10645 -2755 10675 -2725
rect 10805 -2755 10835 -2725
rect 10965 -2755 10995 -2725
rect 9130 -2835 9310 -2805
rect 9450 -2835 9630 -2805
rect 9770 -2835 9950 -2805
rect 10090 -2835 10270 -2805
rect 10805 -2835 10835 -2805
rect 10965 -2835 10995 -2805
rect 10645 -2915 10675 -2885
rect 10805 -2915 10835 -2885
rect 10965 -2915 10995 -2885
rect 9045 -2995 9075 -2965
rect 9205 -2995 9235 -2965
rect 9365 -2995 9395 -2965
rect 9045 -3395 9075 -3365
rect 8405 -3475 8435 -3445
rect 9525 -2995 9555 -2965
rect 9845 -2995 9875 -2965
rect 10005 -2995 10035 -2965
rect 9685 -3395 9715 -3365
rect 9045 -3475 9075 -3445
rect 10165 -2995 10195 -2965
rect 10645 -3075 10675 -3045
rect 10805 -3075 10835 -3045
rect 10965 -3075 10995 -3045
rect 10645 -3155 10675 -3125
rect 10805 -3155 10835 -3125
rect 10965 -3155 10995 -3125
rect 10645 -3235 10675 -3205
rect 10805 -3235 10835 -3205
rect 10965 -3235 10995 -3205
rect 10645 -3315 10675 -3285
rect 10805 -3315 10835 -3285
rect 10965 -3315 10995 -3285
rect 10325 -3395 10355 -3365
rect 10645 -3395 10675 -3365
rect 10805 -3395 10835 -3365
rect 10965 -3395 10995 -3365
rect 9685 -3475 9715 -3445
rect 10325 -3475 10355 -3445
rect 10645 -3475 10675 -3445
rect 10805 -3475 10835 -3445
rect 10965 -3475 10995 -3445
rect -715 -3555 -685 -3525
rect -555 -3555 -525 -3525
rect -395 -3555 -365 -3525
rect 10645 -3555 10675 -3525
rect 10805 -3555 10835 -3525
rect 10965 -3555 10995 -3525
rect -715 -3635 -685 -3605
rect -555 -3635 -525 -3605
rect -395 -3635 -365 -3605
rect 10645 -3635 10675 -3605
rect 10805 -3635 10835 -3605
rect 10965 -3635 10995 -3605
rect -715 -3715 -685 -3685
rect -555 -3715 -525 -3685
rect -395 -3715 -365 -3685
rect 10645 -3715 10675 -3685
rect 10805 -3715 10835 -3685
rect 10965 -3715 10995 -3685
<< metal2 >>
rect -720 1035 11000 1040
rect -720 1005 -715 1035
rect -685 1005 -555 1035
rect -525 1005 -395 1035
rect -365 1005 -315 1035
rect -285 1005 -235 1035
rect -205 1005 -155 1035
rect -125 1005 -75 1035
rect -45 1005 5 1035
rect 35 1005 85 1035
rect 115 1005 165 1035
rect 195 1005 245 1035
rect 275 1005 325 1035
rect 355 1005 405 1035
rect 435 1005 485 1035
rect 515 1005 565 1035
rect 595 1005 645 1035
rect 675 1005 725 1035
rect 755 1005 805 1035
rect 835 1005 885 1035
rect 915 1005 965 1035
rect 995 1005 1045 1035
rect 1075 1005 1125 1035
rect 1155 1005 1205 1035
rect 1235 1005 1285 1035
rect 1315 1005 1365 1035
rect 1395 1005 1445 1035
rect 1475 1005 1525 1035
rect 1555 1005 1605 1035
rect 1635 1005 1685 1035
rect 1715 1005 1765 1035
rect 1795 1005 1845 1035
rect 1875 1005 1925 1035
rect 1955 1005 2005 1035
rect 2035 1005 2085 1035
rect 2115 1005 2165 1035
rect 2195 1005 2245 1035
rect 2275 1005 2325 1035
rect 2355 1005 2405 1035
rect 2435 1005 2485 1035
rect 2515 1005 2565 1035
rect 2595 1005 2645 1035
rect 2675 1005 2725 1035
rect 2755 1005 2805 1035
rect 2835 1005 2885 1035
rect 2915 1005 2965 1035
rect 2995 1005 3045 1035
rect 3075 1005 3125 1035
rect 3155 1005 3205 1035
rect 3235 1005 3285 1035
rect 3315 1005 3365 1035
rect 3395 1005 3445 1035
rect 3475 1005 3525 1035
rect 3555 1005 3605 1035
rect 3635 1005 3685 1035
rect 3715 1005 3765 1035
rect 3795 1005 3845 1035
rect 3875 1005 3925 1035
rect 3955 1005 4005 1035
rect 4035 1005 4085 1035
rect 4115 1005 4165 1035
rect 4195 1005 4245 1035
rect 4275 1005 4325 1035
rect 4355 1005 4405 1035
rect 4435 1005 4485 1035
rect 4515 1005 4565 1035
rect 4595 1005 4645 1035
rect 4675 1005 4725 1035
rect 4755 1005 4805 1035
rect 4835 1005 4885 1035
rect 4915 1005 4965 1035
rect 4995 1005 5045 1035
rect 5075 1005 5125 1035
rect 5155 1005 5205 1035
rect 5235 1005 5285 1035
rect 5315 1005 5365 1035
rect 5395 1005 5445 1035
rect 5475 1005 5525 1035
rect 5555 1005 5605 1035
rect 5635 1005 5685 1035
rect 5715 1005 5765 1035
rect 5795 1005 5845 1035
rect 5875 1005 5925 1035
rect 5955 1005 6005 1035
rect 6035 1005 6085 1035
rect 6115 1005 6165 1035
rect 6195 1005 6245 1035
rect 6275 1005 6325 1035
rect 6355 1005 6405 1035
rect 6435 1005 6485 1035
rect 6515 1005 6565 1035
rect 6595 1005 6645 1035
rect 6675 1005 6725 1035
rect 6755 1005 6805 1035
rect 6835 1005 6885 1035
rect 6915 1005 6965 1035
rect 6995 1005 7045 1035
rect 7075 1005 7125 1035
rect 7155 1005 7205 1035
rect 7235 1005 7285 1035
rect 7315 1005 7365 1035
rect 7395 1005 7445 1035
rect 7475 1005 7525 1035
rect 7555 1005 7605 1035
rect 7635 1005 7685 1035
rect 7715 1005 7765 1035
rect 7795 1005 7845 1035
rect 7875 1005 7925 1035
rect 7955 1005 8005 1035
rect 8035 1005 8085 1035
rect 8115 1005 8165 1035
rect 8195 1005 8245 1035
rect 8275 1005 8325 1035
rect 8355 1005 8405 1035
rect 8435 1005 8485 1035
rect 8515 1005 8565 1035
rect 8595 1005 8645 1035
rect 8675 1005 8725 1035
rect 8755 1005 8805 1035
rect 8835 1005 8885 1035
rect 8915 1005 8965 1035
rect 8995 1005 9045 1035
rect 9075 1005 9125 1035
rect 9155 1005 9205 1035
rect 9235 1005 9285 1035
rect 9315 1005 9365 1035
rect 9395 1005 9445 1035
rect 9475 1005 9525 1035
rect 9555 1005 9605 1035
rect 9635 1005 9685 1035
rect 9715 1005 9765 1035
rect 9795 1005 9845 1035
rect 9875 1005 9925 1035
rect 9955 1005 10005 1035
rect 10035 1005 10085 1035
rect 10115 1005 10165 1035
rect 10195 1005 10245 1035
rect 10275 1005 10325 1035
rect 10355 1005 10405 1035
rect 10435 1005 10485 1035
rect 10515 1005 10645 1035
rect 10675 1005 10805 1035
rect 10835 1005 10965 1035
rect 10995 1005 11000 1035
rect -720 1000 11000 1005
rect -720 955 11000 960
rect -720 925 -715 955
rect -685 925 -555 955
rect -525 925 -395 955
rect -365 925 -315 955
rect -285 925 -235 955
rect -205 925 -155 955
rect -125 925 -75 955
rect -45 925 5 955
rect 35 925 85 955
rect 115 925 165 955
rect 195 925 245 955
rect 275 925 325 955
rect 355 925 405 955
rect 435 925 485 955
rect 515 925 565 955
rect 595 925 645 955
rect 675 925 725 955
rect 755 925 805 955
rect 835 925 885 955
rect 915 925 965 955
rect 995 925 1045 955
rect 1075 925 1125 955
rect 1155 925 1205 955
rect 1235 925 1285 955
rect 1315 925 1365 955
rect 1395 925 1445 955
rect 1475 925 1525 955
rect 1555 925 1605 955
rect 1635 925 1685 955
rect 1715 925 1765 955
rect 1795 925 1845 955
rect 1875 925 1925 955
rect 1955 925 2005 955
rect 2035 925 2085 955
rect 2115 925 2165 955
rect 2195 925 2245 955
rect 2275 925 2325 955
rect 2355 925 2405 955
rect 2435 925 2485 955
rect 2515 925 2565 955
rect 2595 925 2645 955
rect 2675 925 2725 955
rect 2755 925 2805 955
rect 2835 925 2885 955
rect 2915 925 2965 955
rect 2995 925 3045 955
rect 3075 925 3125 955
rect 3155 925 3205 955
rect 3235 925 3285 955
rect 3315 925 3365 955
rect 3395 925 3445 955
rect 3475 925 3525 955
rect 3555 925 3605 955
rect 3635 925 3685 955
rect 3715 925 3765 955
rect 3795 925 3845 955
rect 3875 925 3925 955
rect 3955 925 4005 955
rect 4035 925 4085 955
rect 4115 925 4165 955
rect 4195 925 4245 955
rect 4275 925 4325 955
rect 4355 925 4405 955
rect 4435 925 4485 955
rect 4515 925 4565 955
rect 4595 925 4645 955
rect 4675 925 4725 955
rect 4755 925 4805 955
rect 4835 925 4885 955
rect 4915 925 4965 955
rect 4995 925 5045 955
rect 5075 925 5125 955
rect 5155 925 5205 955
rect 5235 925 5285 955
rect 5315 925 5365 955
rect 5395 925 5445 955
rect 5475 925 5525 955
rect 5555 925 5605 955
rect 5635 925 5685 955
rect 5715 925 5765 955
rect 5795 925 5845 955
rect 5875 925 5925 955
rect 5955 925 6005 955
rect 6035 925 6085 955
rect 6115 925 6165 955
rect 6195 925 6245 955
rect 6275 925 6325 955
rect 6355 925 6405 955
rect 6435 925 6485 955
rect 6515 925 6565 955
rect 6595 925 6645 955
rect 6675 925 6725 955
rect 6755 925 6805 955
rect 6835 925 6885 955
rect 6915 925 6965 955
rect 6995 925 7045 955
rect 7075 925 7125 955
rect 7155 925 7205 955
rect 7235 925 7285 955
rect 7315 925 7365 955
rect 7395 925 7445 955
rect 7475 925 7525 955
rect 7555 925 7605 955
rect 7635 925 7685 955
rect 7715 925 7765 955
rect 7795 925 7845 955
rect 7875 925 7925 955
rect 7955 925 8005 955
rect 8035 925 8085 955
rect 8115 925 8165 955
rect 8195 925 8245 955
rect 8275 925 8325 955
rect 8355 925 8405 955
rect 8435 925 8485 955
rect 8515 925 8565 955
rect 8595 925 8645 955
rect 8675 925 8725 955
rect 8755 925 8805 955
rect 8835 925 8885 955
rect 8915 925 8965 955
rect 8995 925 9045 955
rect 9075 925 9125 955
rect 9155 925 9205 955
rect 9235 925 9285 955
rect 9315 925 9365 955
rect 9395 925 9445 955
rect 9475 925 9525 955
rect 9555 925 9605 955
rect 9635 925 9685 955
rect 9715 925 9765 955
rect 9795 925 9845 955
rect 9875 925 9925 955
rect 9955 925 10005 955
rect 10035 925 10085 955
rect 10115 925 10165 955
rect 10195 925 10245 955
rect 10275 925 10325 955
rect 10355 925 10405 955
rect 10435 925 10485 955
rect 10515 925 10645 955
rect 10675 925 10805 955
rect 10835 925 10965 955
rect 10995 925 11000 955
rect -720 920 11000 925
rect -720 875 11000 880
rect -720 845 -715 875
rect -685 845 -555 875
rect -525 845 -395 875
rect -365 845 -315 875
rect -285 845 -235 875
rect -205 845 -155 875
rect -125 845 -75 875
rect -45 845 5 875
rect 35 845 85 875
rect 115 845 165 875
rect 195 845 245 875
rect 275 845 325 875
rect 355 845 405 875
rect 435 845 485 875
rect 515 845 565 875
rect 595 845 645 875
rect 675 845 725 875
rect 755 845 805 875
rect 835 845 885 875
rect 915 845 965 875
rect 995 845 1045 875
rect 1075 845 1125 875
rect 1155 845 1205 875
rect 1235 845 1285 875
rect 1315 845 1365 875
rect 1395 845 1445 875
rect 1475 845 1525 875
rect 1555 845 1605 875
rect 1635 845 1685 875
rect 1715 845 1765 875
rect 1795 845 1845 875
rect 1875 845 1925 875
rect 1955 845 2005 875
rect 2035 845 2085 875
rect 2115 845 2165 875
rect 2195 845 2245 875
rect 2275 845 2325 875
rect 2355 845 2405 875
rect 2435 845 2485 875
rect 2515 845 2565 875
rect 2595 845 2645 875
rect 2675 845 2725 875
rect 2755 845 2805 875
rect 2835 845 2885 875
rect 2915 845 2965 875
rect 2995 845 3045 875
rect 3075 845 3125 875
rect 3155 845 3205 875
rect 3235 845 3285 875
rect 3315 845 3365 875
rect 3395 845 3445 875
rect 3475 845 3525 875
rect 3555 845 3605 875
rect 3635 845 3685 875
rect 3715 845 3765 875
rect 3795 845 3845 875
rect 3875 845 3925 875
rect 3955 845 4005 875
rect 4035 845 4085 875
rect 4115 845 4165 875
rect 4195 845 4245 875
rect 4275 845 4325 875
rect 4355 845 4405 875
rect 4435 845 4485 875
rect 4515 845 4565 875
rect 4595 845 4645 875
rect 4675 845 4725 875
rect 4755 845 4805 875
rect 4835 845 4885 875
rect 4915 845 4965 875
rect 4995 845 5045 875
rect 5075 845 5125 875
rect 5155 845 5205 875
rect 5235 845 5285 875
rect 5315 845 5365 875
rect 5395 845 5445 875
rect 5475 845 5525 875
rect 5555 845 5605 875
rect 5635 845 5685 875
rect 5715 845 5765 875
rect 5795 845 5845 875
rect 5875 845 5925 875
rect 5955 845 6005 875
rect 6035 845 6085 875
rect 6115 845 6165 875
rect 6195 845 6245 875
rect 6275 845 6325 875
rect 6355 845 6405 875
rect 6435 845 6485 875
rect 6515 845 6565 875
rect 6595 845 6645 875
rect 6675 845 6725 875
rect 6755 845 6805 875
rect 6835 845 6885 875
rect 6915 845 6965 875
rect 6995 845 7045 875
rect 7075 845 7125 875
rect 7155 845 7205 875
rect 7235 845 7285 875
rect 7315 845 7365 875
rect 7395 845 7445 875
rect 7475 845 7525 875
rect 7555 845 7605 875
rect 7635 845 7685 875
rect 7715 845 7765 875
rect 7795 845 7845 875
rect 7875 845 7925 875
rect 7955 845 8005 875
rect 8035 845 8085 875
rect 8115 845 8165 875
rect 8195 845 8245 875
rect 8275 845 8325 875
rect 8355 845 8405 875
rect 8435 845 8485 875
rect 8515 845 8565 875
rect 8595 845 8645 875
rect 8675 845 8725 875
rect 8755 845 8805 875
rect 8835 845 8885 875
rect 8915 845 8965 875
rect 8995 845 9045 875
rect 9075 845 9125 875
rect 9155 845 9205 875
rect 9235 845 9285 875
rect 9315 845 9365 875
rect 9395 845 9445 875
rect 9475 845 9525 875
rect 9555 845 9605 875
rect 9635 845 9685 875
rect 9715 845 9765 875
rect 9795 845 9845 875
rect 9875 845 9925 875
rect 9955 845 10005 875
rect 10035 845 10085 875
rect 10115 845 10165 875
rect 10195 845 10245 875
rect 10275 845 10325 875
rect 10355 845 10405 875
rect 10435 845 10485 875
rect 10515 845 10645 875
rect 10675 845 10805 875
rect 10835 845 10965 875
rect 10995 845 11000 875
rect -720 840 11000 845
rect -640 795 10600 800
rect -640 765 -635 795
rect -605 765 -75 795
rect -45 765 5205 795
rect 5235 765 5845 795
rect 5875 765 6485 795
rect 6515 765 7125 795
rect 7155 765 7765 795
rect 7795 765 8405 795
rect 8435 765 9045 795
rect 9075 765 9685 795
rect 9715 765 10325 795
rect 10355 765 10600 795
rect -640 760 10600 765
rect 10640 795 11000 800
rect 10640 765 10645 795
rect 10675 765 10805 795
rect 10835 765 10965 795
rect 10995 765 11000 795
rect 10640 760 11000 765
rect -640 715 10600 720
rect -640 685 -635 715
rect -605 685 -75 715
rect -45 685 5205 715
rect 5235 685 5845 715
rect 5875 685 6485 715
rect 6515 685 7125 715
rect 7155 685 7765 715
rect 7795 685 8405 715
rect 8435 685 9045 715
rect 9075 685 9685 715
rect 9715 685 10325 715
rect 10355 685 10600 715
rect -640 680 10600 685
rect 10640 715 11000 720
rect 10640 685 10645 715
rect 10675 685 10805 715
rect 10835 685 10965 715
rect 10995 685 11000 715
rect 10640 680 11000 685
rect -720 635 11000 640
rect -720 605 -715 635
rect -685 605 -555 635
rect -525 605 -395 635
rect -365 605 -315 635
rect -285 605 -235 635
rect -205 605 -155 635
rect -125 605 -75 635
rect -45 605 5 635
rect 35 605 85 635
rect 115 605 165 635
rect 195 605 245 635
rect 275 605 325 635
rect 355 605 405 635
rect 435 605 485 635
rect 515 605 565 635
rect 595 605 645 635
rect 675 605 725 635
rect 755 605 805 635
rect 835 605 885 635
rect 915 605 965 635
rect 995 605 1045 635
rect 1075 605 1125 635
rect 1155 605 1205 635
rect 1235 605 1285 635
rect 1315 605 1365 635
rect 1395 605 1445 635
rect 1475 605 1525 635
rect 1555 605 1605 635
rect 1635 605 1685 635
rect 1715 605 1765 635
rect 1795 605 1845 635
rect 1875 605 1925 635
rect 1955 605 2005 635
rect 2035 605 2085 635
rect 2115 605 2165 635
rect 2195 605 2245 635
rect 2275 605 2325 635
rect 2355 605 2405 635
rect 2435 605 2485 635
rect 2515 605 2565 635
rect 2595 605 2645 635
rect 2675 605 2725 635
rect 2755 605 2805 635
rect 2835 605 2885 635
rect 2915 605 2965 635
rect 2995 605 3045 635
rect 3075 605 3125 635
rect 3155 605 3205 635
rect 3235 605 3285 635
rect 3315 605 3365 635
rect 3395 605 3445 635
rect 3475 605 3525 635
rect 3555 605 3605 635
rect 3635 605 3685 635
rect 3715 605 3765 635
rect 3795 605 3845 635
rect 3875 605 3925 635
rect 3955 605 4005 635
rect 4035 605 4085 635
rect 4115 605 4165 635
rect 4195 605 4245 635
rect 4275 605 4325 635
rect 4355 605 4405 635
rect 4435 605 4485 635
rect 4515 605 4565 635
rect 4595 605 4645 635
rect 4675 605 4725 635
rect 4755 605 4805 635
rect 4835 605 4885 635
rect 4915 605 4965 635
rect 4995 605 5045 635
rect 5075 605 5125 635
rect 5155 605 5205 635
rect 5235 605 5285 635
rect 5315 605 5365 635
rect 5395 605 5445 635
rect 5475 605 5525 635
rect 5555 605 5605 635
rect 5635 605 5685 635
rect 5715 605 5765 635
rect 5795 605 5845 635
rect 5875 605 5925 635
rect 5955 605 6005 635
rect 6035 605 6085 635
rect 6115 605 6165 635
rect 6195 605 6245 635
rect 6275 605 6325 635
rect 6355 605 6405 635
rect 6435 605 6485 635
rect 6515 605 6565 635
rect 6595 605 6645 635
rect 6675 605 6725 635
rect 6755 605 6805 635
rect 6835 605 6885 635
rect 6915 605 6965 635
rect 6995 605 7045 635
rect 7075 605 7125 635
rect 7155 605 7205 635
rect 7235 605 7285 635
rect 7315 605 7365 635
rect 7395 605 7445 635
rect 7475 605 7525 635
rect 7555 605 7605 635
rect 7635 605 7685 635
rect 7715 605 7765 635
rect 7795 605 7845 635
rect 7875 605 7925 635
rect 7955 605 8005 635
rect 8035 605 8085 635
rect 8115 605 8165 635
rect 8195 605 8245 635
rect 8275 605 8325 635
rect 8355 605 8405 635
rect 8435 605 8485 635
rect 8515 605 8565 635
rect 8595 605 8645 635
rect 8675 605 8725 635
rect 8755 605 8805 635
rect 8835 605 8885 635
rect 8915 605 8965 635
rect 8995 605 9045 635
rect 9075 605 9125 635
rect 9155 605 9205 635
rect 9235 605 9285 635
rect 9315 605 9365 635
rect 9395 605 9445 635
rect 9475 605 9525 635
rect 9555 605 9605 635
rect 9635 605 9685 635
rect 9715 605 9765 635
rect 9795 605 9845 635
rect 9875 605 9925 635
rect 9955 605 10005 635
rect 10035 605 10085 635
rect 10115 605 10165 635
rect 10195 605 10245 635
rect 10275 605 10325 635
rect 10355 605 10405 635
rect 10435 605 10485 635
rect 10515 605 10645 635
rect 10675 605 10805 635
rect 10835 605 10965 635
rect 10995 605 11000 635
rect -720 600 11000 605
rect -720 555 11000 560
rect -720 525 -715 555
rect -685 525 -555 555
rect -525 525 -395 555
rect -365 525 -315 555
rect -285 525 -235 555
rect -205 525 -155 555
rect -125 525 -75 555
rect -45 525 5 555
rect 35 525 85 555
rect 115 525 165 555
rect 195 525 245 555
rect 275 525 325 555
rect 355 525 405 555
rect 435 525 485 555
rect 515 525 565 555
rect 595 525 645 555
rect 675 525 725 555
rect 755 525 805 555
rect 835 525 885 555
rect 915 525 965 555
rect 995 525 1045 555
rect 1075 525 1125 555
rect 1155 525 1205 555
rect 1235 525 1285 555
rect 1315 525 1365 555
rect 1395 525 1445 555
rect 1475 525 1525 555
rect 1555 525 1605 555
rect 1635 525 1685 555
rect 1715 525 1765 555
rect 1795 525 1845 555
rect 1875 525 1925 555
rect 1955 525 2005 555
rect 2035 525 2085 555
rect 2115 525 2165 555
rect 2195 525 2245 555
rect 2275 525 2325 555
rect 2355 525 2405 555
rect 2435 525 2485 555
rect 2515 525 2565 555
rect 2595 525 2645 555
rect 2675 525 2725 555
rect 2755 525 2805 555
rect 2835 525 2885 555
rect 2915 525 2965 555
rect 2995 525 3045 555
rect 3075 525 3125 555
rect 3155 525 3205 555
rect 3235 525 3285 555
rect 3315 525 3365 555
rect 3395 525 3445 555
rect 3475 525 3525 555
rect 3555 525 3605 555
rect 3635 525 3685 555
rect 3715 525 3765 555
rect 3795 525 3845 555
rect 3875 525 3925 555
rect 3955 525 4005 555
rect 4035 525 4085 555
rect 4115 525 4165 555
rect 4195 525 4245 555
rect 4275 525 4325 555
rect 4355 525 4405 555
rect 4435 525 4485 555
rect 4515 525 4565 555
rect 4595 525 4645 555
rect 4675 525 4725 555
rect 4755 525 4805 555
rect 4835 525 4885 555
rect 4915 525 4965 555
rect 4995 525 5045 555
rect 5075 525 5125 555
rect 5155 525 5205 555
rect 5235 525 5285 555
rect 5315 525 5365 555
rect 5395 525 5445 555
rect 5475 525 5525 555
rect 5555 525 5605 555
rect 5635 525 5685 555
rect 5715 525 5765 555
rect 5795 525 5845 555
rect 5875 525 5925 555
rect 5955 525 6005 555
rect 6035 525 6085 555
rect 6115 525 6165 555
rect 6195 525 6245 555
rect 6275 525 6325 555
rect 6355 525 6405 555
rect 6435 525 6485 555
rect 6515 525 6565 555
rect 6595 525 6645 555
rect 6675 525 6725 555
rect 6755 525 6805 555
rect 6835 525 6885 555
rect 6915 525 6965 555
rect 6995 525 7045 555
rect 7075 525 7125 555
rect 7155 525 7205 555
rect 7235 525 7285 555
rect 7315 525 7365 555
rect 7395 525 7445 555
rect 7475 525 7525 555
rect 7555 525 7605 555
rect 7635 525 7685 555
rect 7715 525 7765 555
rect 7795 525 7845 555
rect 7875 525 7925 555
rect 7955 525 8005 555
rect 8035 525 8085 555
rect 8115 525 8165 555
rect 8195 525 8245 555
rect 8275 525 8325 555
rect 8355 525 8405 555
rect 8435 525 8485 555
rect 8515 525 8565 555
rect 8595 525 8645 555
rect 8675 525 8725 555
rect 8755 525 8805 555
rect 8835 525 8885 555
rect 8915 525 8965 555
rect 8995 525 9045 555
rect 9075 525 9125 555
rect 9155 525 9205 555
rect 9235 525 9285 555
rect 9315 525 9365 555
rect 9395 525 9445 555
rect 9475 525 9525 555
rect 9555 525 9605 555
rect 9635 525 9685 555
rect 9715 525 9765 555
rect 9795 525 9845 555
rect 9875 525 9925 555
rect 9955 525 10005 555
rect 10035 525 10085 555
rect 10115 525 10165 555
rect 10195 525 10245 555
rect 10275 525 10325 555
rect 10355 525 10405 555
rect 10435 525 10485 555
rect 10515 525 10645 555
rect 10675 525 10805 555
rect 10835 525 10965 555
rect 10995 525 11000 555
rect -720 520 11000 525
rect -720 475 -520 480
rect -720 445 -715 475
rect -685 445 -555 475
rect -525 445 -520 475
rect -720 440 -520 445
rect -480 475 10600 480
rect -480 445 -475 475
rect -445 445 85 475
rect 115 445 405 475
rect 435 445 725 475
rect 755 445 1045 475
rect 1075 445 1365 475
rect 1395 445 1685 475
rect 1715 445 2005 475
rect 2035 445 2325 475
rect 2355 445 2645 475
rect 2675 445 2965 475
rect 2995 445 3285 475
rect 3315 445 3605 475
rect 3635 445 3925 475
rect 3955 445 4245 475
rect 4275 445 4565 475
rect 4595 445 4885 475
rect 4915 445 10600 475
rect -480 440 10600 445
rect 10640 475 11000 480
rect 10640 445 10645 475
rect 10675 445 10805 475
rect 10835 445 10965 475
rect 10995 445 11000 475
rect 10640 440 11000 445
rect -720 395 11000 400
rect -720 365 -715 395
rect -685 365 -555 395
rect -525 365 -395 395
rect -365 365 -315 395
rect -285 365 -235 395
rect -205 365 -155 395
rect -125 365 -75 395
rect -45 365 5 395
rect 35 365 85 395
rect 115 365 165 395
rect 195 365 245 395
rect 275 365 325 395
rect 355 365 405 395
rect 435 365 485 395
rect 515 365 565 395
rect 595 365 645 395
rect 675 365 725 395
rect 755 365 805 395
rect 835 365 885 395
rect 915 365 965 395
rect 995 365 1045 395
rect 1075 365 1125 395
rect 1155 365 1205 395
rect 1235 365 1285 395
rect 1315 365 1365 395
rect 1395 365 1445 395
rect 1475 365 1525 395
rect 1555 365 1605 395
rect 1635 365 1685 395
rect 1715 365 1765 395
rect 1795 365 1845 395
rect 1875 365 1925 395
rect 1955 365 2005 395
rect 2035 365 2085 395
rect 2115 365 2165 395
rect 2195 365 2245 395
rect 2275 365 2325 395
rect 2355 365 2405 395
rect 2435 365 2485 395
rect 2515 365 2565 395
rect 2595 365 2645 395
rect 2675 365 2725 395
rect 2755 365 2805 395
rect 2835 365 2885 395
rect 2915 365 2965 395
rect 2995 365 3045 395
rect 3075 365 3125 395
rect 3155 365 3205 395
rect 3235 365 3285 395
rect 3315 365 3365 395
rect 3395 365 3445 395
rect 3475 365 3525 395
rect 3555 365 3605 395
rect 3635 365 3685 395
rect 3715 365 3765 395
rect 3795 365 3845 395
rect 3875 365 3925 395
rect 3955 365 4005 395
rect 4035 365 4085 395
rect 4115 365 4165 395
rect 4195 365 4245 395
rect 4275 365 4325 395
rect 4355 365 4405 395
rect 4435 365 4485 395
rect 4515 365 4565 395
rect 4595 365 4645 395
rect 4675 365 4725 395
rect 4755 365 4805 395
rect 4835 365 4885 395
rect 4915 365 4965 395
rect 4995 365 5045 395
rect 5075 365 5125 395
rect 5155 365 5205 395
rect 5235 365 5285 395
rect 5315 365 5365 395
rect 5395 365 5445 395
rect 5475 365 5525 395
rect 5555 365 5605 395
rect 5635 365 5685 395
rect 5715 365 5765 395
rect 5795 365 5845 395
rect 5875 365 5925 395
rect 5955 365 6005 395
rect 6035 365 6085 395
rect 6115 365 6165 395
rect 6195 365 6245 395
rect 6275 365 6325 395
rect 6355 365 6405 395
rect 6435 365 6485 395
rect 6515 365 6565 395
rect 6595 365 6645 395
rect 6675 365 6725 395
rect 6755 365 6805 395
rect 6835 365 6885 395
rect 6915 365 6965 395
rect 6995 365 7045 395
rect 7075 365 7125 395
rect 7155 365 7205 395
rect 7235 365 7285 395
rect 7315 365 7365 395
rect 7395 365 7445 395
rect 7475 365 7525 395
rect 7555 365 7605 395
rect 7635 365 7685 395
rect 7715 365 7765 395
rect 7795 365 7845 395
rect 7875 365 7925 395
rect 7955 365 8005 395
rect 8035 365 8085 395
rect 8115 365 8165 395
rect 8195 365 8245 395
rect 8275 365 8325 395
rect 8355 365 8405 395
rect 8435 365 8485 395
rect 8515 365 8565 395
rect 8595 365 8645 395
rect 8675 365 8725 395
rect 8755 365 8805 395
rect 8835 365 8885 395
rect 8915 365 8965 395
rect 8995 365 9045 395
rect 9075 365 9125 395
rect 9155 365 9205 395
rect 9235 365 9285 395
rect 9315 365 9365 395
rect 9395 365 9445 395
rect 9475 365 9525 395
rect 9555 365 9605 395
rect 9635 365 9685 395
rect 9715 365 9765 395
rect 9795 365 9845 395
rect 9875 365 9925 395
rect 9955 365 10005 395
rect 10035 365 10085 395
rect 10115 365 10165 395
rect 10195 365 10245 395
rect 10275 365 10325 395
rect 10355 365 10405 395
rect 10435 365 10485 395
rect 10515 365 10645 395
rect 10675 365 10805 395
rect 10835 365 10965 395
rect 10995 365 11000 395
rect -720 360 11000 365
rect -720 315 -360 320
rect -720 285 -715 315
rect -685 285 -555 315
rect -525 285 -395 315
rect -365 285 -360 315
rect -720 280 -360 285
rect -320 315 10920 320
rect -320 285 5365 315
rect 5395 285 5525 315
rect 5555 285 5685 315
rect 5715 285 6005 315
rect 6035 285 6165 315
rect 6195 285 6325 315
rect 6355 285 6485 315
rect 6515 285 6645 315
rect 6675 285 6805 315
rect 6835 285 6965 315
rect 6995 285 7285 315
rect 7315 285 7445 315
rect 7475 285 7605 315
rect 7635 285 7925 315
rect 7955 285 8085 315
rect 8115 285 8245 315
rect 8275 285 8565 315
rect 8595 285 8725 315
rect 8755 285 8885 315
rect 8915 285 9045 315
rect 9075 285 9205 315
rect 9235 285 9365 315
rect 9395 285 9525 315
rect 9555 285 9845 315
rect 9875 285 10005 315
rect 10035 285 10165 315
rect 10195 285 10885 315
rect 10915 285 10920 315
rect -320 280 10920 285
rect 10960 280 11000 320
rect -720 235 11000 240
rect -720 205 -715 235
rect -685 205 -555 235
rect -525 205 -395 235
rect -365 205 -315 235
rect -285 205 -235 235
rect -205 205 -155 235
rect -125 205 -75 235
rect -45 205 5 235
rect 35 205 85 235
rect 115 205 165 235
rect 195 205 245 235
rect 275 205 325 235
rect 355 205 405 235
rect 435 205 485 235
rect 515 205 565 235
rect 595 205 645 235
rect 675 205 725 235
rect 755 205 805 235
rect 835 205 885 235
rect 915 205 965 235
rect 995 205 1045 235
rect 1075 205 1125 235
rect 1155 205 1205 235
rect 1235 205 1285 235
rect 1315 205 1365 235
rect 1395 205 1445 235
rect 1475 205 1525 235
rect 1555 205 1605 235
rect 1635 205 1685 235
rect 1715 205 1765 235
rect 1795 205 1845 235
rect 1875 205 1925 235
rect 1955 205 2005 235
rect 2035 205 2085 235
rect 2115 205 2165 235
rect 2195 205 2245 235
rect 2275 205 2325 235
rect 2355 205 2405 235
rect 2435 205 2485 235
rect 2515 205 2565 235
rect 2595 205 2645 235
rect 2675 205 2725 235
rect 2755 205 2805 235
rect 2835 205 2885 235
rect 2915 205 2965 235
rect 2995 205 3045 235
rect 3075 205 3125 235
rect 3155 205 3205 235
rect 3235 205 3285 235
rect 3315 205 3365 235
rect 3395 205 3445 235
rect 3475 205 3525 235
rect 3555 205 3605 235
rect 3635 205 3685 235
rect 3715 205 3765 235
rect 3795 205 3845 235
rect 3875 205 3925 235
rect 3955 205 4005 235
rect 4035 205 4085 235
rect 4115 205 4165 235
rect 4195 205 4245 235
rect 4275 205 4325 235
rect 4355 205 4405 235
rect 4435 205 4485 235
rect 4515 205 4565 235
rect 4595 205 4645 235
rect 4675 205 4725 235
rect 4755 205 4805 235
rect 4835 205 4885 235
rect 4915 205 4965 235
rect 4995 205 5045 235
rect 5075 205 5125 235
rect 5155 205 5205 235
rect 5235 205 5285 235
rect 5315 205 5365 235
rect 5395 205 5445 235
rect 5475 205 5525 235
rect 5555 205 5605 235
rect 5635 205 5685 235
rect 5715 205 5765 235
rect 5795 205 5845 235
rect 5875 205 5925 235
rect 5955 205 6005 235
rect 6035 205 6085 235
rect 6115 205 6165 235
rect 6195 205 6245 235
rect 6275 205 6325 235
rect 6355 205 6405 235
rect 6435 205 6485 235
rect 6515 205 6565 235
rect 6595 205 6645 235
rect 6675 205 6725 235
rect 6755 205 6805 235
rect 6835 205 6885 235
rect 6915 205 6965 235
rect 6995 205 7045 235
rect 7075 205 7125 235
rect 7155 205 7205 235
rect 7235 205 7285 235
rect 7315 205 7365 235
rect 7395 205 7445 235
rect 7475 205 7525 235
rect 7555 205 7605 235
rect 7635 205 7685 235
rect 7715 205 7765 235
rect 7795 205 7845 235
rect 7875 205 7925 235
rect 7955 205 8005 235
rect 8035 205 8085 235
rect 8115 205 8165 235
rect 8195 205 8245 235
rect 8275 205 8325 235
rect 8355 205 8405 235
rect 8435 205 8485 235
rect 8515 205 8565 235
rect 8595 205 8645 235
rect 8675 205 8725 235
rect 8755 205 8805 235
rect 8835 205 8885 235
rect 8915 205 8965 235
rect 8995 205 9045 235
rect 9075 205 9125 235
rect 9155 205 9205 235
rect 9235 205 9285 235
rect 9315 205 9365 235
rect 9395 205 9445 235
rect 9475 205 9525 235
rect 9555 205 9605 235
rect 9635 205 9685 235
rect 9715 205 9765 235
rect 9795 205 9845 235
rect 9875 205 9925 235
rect 9955 205 10005 235
rect 10035 205 10085 235
rect 10115 205 10165 235
rect 10195 205 10245 235
rect 10275 205 10325 235
rect 10355 205 10405 235
rect 10435 205 10485 235
rect 10515 205 10645 235
rect 10675 205 10805 235
rect 10835 205 10965 235
rect 10995 205 11000 235
rect -720 200 11000 205
rect -720 155 -360 160
rect -720 125 -715 155
rect -685 125 -555 155
rect -525 125 -395 155
rect -365 125 -360 155
rect -720 120 -360 125
rect -320 155 10760 160
rect -320 125 10 155
rect 190 125 330 155
rect 510 125 650 155
rect 830 125 970 155
rect 1150 125 1205 155
rect 1235 125 1290 155
rect 1470 125 1610 155
rect 1790 125 1930 155
rect 2110 125 2250 155
rect 2430 125 2570 155
rect 2750 125 2890 155
rect 3070 125 3210 155
rect 3390 125 3530 155
rect 3710 125 3765 155
rect 3795 125 3850 155
rect 4030 125 4170 155
rect 4350 125 4490 155
rect 4670 125 4810 155
rect 4990 125 5045 155
rect 5075 125 5290 155
rect 5470 125 5610 155
rect 5790 125 5930 155
rect 6110 125 6250 155
rect 6430 125 6570 155
rect 6750 125 6890 155
rect 7070 125 7210 155
rect 7390 125 7530 155
rect 7710 125 7850 155
rect 8030 125 8170 155
rect 8350 125 8490 155
rect 8670 125 8810 155
rect 8990 125 9130 155
rect 9310 125 9450 155
rect 9630 125 9770 155
rect 9950 125 10090 155
rect 10270 125 10725 155
rect 10755 125 10760 155
rect -320 120 10760 125
rect 10800 155 11000 160
rect 10800 125 10805 155
rect 10835 125 10965 155
rect 10995 125 11000 155
rect 10800 120 11000 125
rect -720 75 11000 80
rect -720 45 -715 75
rect -685 45 -555 75
rect -525 45 -395 75
rect -365 45 -315 75
rect -285 45 -235 75
rect -205 45 -155 75
rect -125 45 -75 75
rect -45 45 5 75
rect 35 45 85 75
rect 115 45 165 75
rect 195 45 245 75
rect 275 45 325 75
rect 355 45 405 75
rect 435 45 485 75
rect 515 45 565 75
rect 595 45 645 75
rect 675 45 725 75
rect 755 45 805 75
rect 835 45 885 75
rect 915 45 965 75
rect 995 45 1045 75
rect 1075 45 1125 75
rect 1155 45 1205 75
rect 1235 45 1285 75
rect 1315 45 1365 75
rect 1395 45 1445 75
rect 1475 45 1525 75
rect 1555 45 1605 75
rect 1635 45 1685 75
rect 1715 45 1765 75
rect 1795 45 1845 75
rect 1875 45 1925 75
rect 1955 45 2005 75
rect 2035 45 2085 75
rect 2115 45 2165 75
rect 2195 45 2245 75
rect 2275 45 2325 75
rect 2355 45 2405 75
rect 2435 45 2485 75
rect 2515 45 2565 75
rect 2595 45 2645 75
rect 2675 45 2725 75
rect 2755 45 2805 75
rect 2835 45 2885 75
rect 2915 45 2965 75
rect 2995 45 3045 75
rect 3075 45 3125 75
rect 3155 45 3205 75
rect 3235 45 3285 75
rect 3315 45 3365 75
rect 3395 45 3445 75
rect 3475 45 3525 75
rect 3555 45 3605 75
rect 3635 45 3685 75
rect 3715 45 3765 75
rect 3795 45 3845 75
rect 3875 45 3925 75
rect 3955 45 4005 75
rect 4035 45 4085 75
rect 4115 45 4165 75
rect 4195 45 4245 75
rect 4275 45 4325 75
rect 4355 45 4405 75
rect 4435 45 4485 75
rect 4515 45 4565 75
rect 4595 45 4645 75
rect 4675 45 4725 75
rect 4755 45 4805 75
rect 4835 45 4885 75
rect 4915 45 4965 75
rect 4995 45 5045 75
rect 5075 45 5125 75
rect 5155 45 5205 75
rect 5235 45 5285 75
rect 5315 45 5365 75
rect 5395 45 5445 75
rect 5475 45 5525 75
rect 5555 45 5605 75
rect 5635 45 5685 75
rect 5715 45 5765 75
rect 5795 45 5845 75
rect 5875 45 5925 75
rect 5955 45 6005 75
rect 6035 45 6085 75
rect 6115 45 6165 75
rect 6195 45 6245 75
rect 6275 45 6325 75
rect 6355 45 6405 75
rect 6435 45 6485 75
rect 6515 45 6565 75
rect 6595 45 6645 75
rect 6675 45 6725 75
rect 6755 45 6805 75
rect 6835 45 6885 75
rect 6915 45 6965 75
rect 6995 45 7045 75
rect 7075 45 7125 75
rect 7155 45 7205 75
rect 7235 45 7285 75
rect 7315 45 7365 75
rect 7395 45 7445 75
rect 7475 45 7525 75
rect 7555 45 7605 75
rect 7635 45 7685 75
rect 7715 45 7765 75
rect 7795 45 7845 75
rect 7875 45 7925 75
rect 7955 45 8005 75
rect 8035 45 8085 75
rect 8115 45 8165 75
rect 8195 45 8245 75
rect 8275 45 8325 75
rect 8355 45 8405 75
rect 8435 45 8485 75
rect 8515 45 8565 75
rect 8595 45 8645 75
rect 8675 45 8725 75
rect 8755 45 8805 75
rect 8835 45 8885 75
rect 8915 45 8965 75
rect 8995 45 9045 75
rect 9075 45 9125 75
rect 9155 45 9205 75
rect 9235 45 9285 75
rect 9315 45 9365 75
rect 9395 45 9445 75
rect 9475 45 9525 75
rect 9555 45 9605 75
rect 9635 45 9685 75
rect 9715 45 9765 75
rect 9795 45 9845 75
rect 9875 45 9925 75
rect 9955 45 10005 75
rect 10035 45 10085 75
rect 10115 45 10165 75
rect 10195 45 10245 75
rect 10275 45 10325 75
rect 10355 45 10405 75
rect 10435 45 10485 75
rect 10515 45 10645 75
rect 10675 45 10805 75
rect 10835 45 10965 75
rect 10995 45 11000 75
rect -720 40 11000 45
rect -720 -5 11000 0
rect -720 -35 -715 -5
rect -685 -35 -555 -5
rect -525 -35 -395 -5
rect -365 -35 -315 -5
rect -285 -35 -235 -5
rect -205 -35 -155 -5
rect -125 -35 -75 -5
rect -45 -35 5 -5
rect 35 -35 85 -5
rect 115 -35 165 -5
rect 195 -35 245 -5
rect 275 -35 325 -5
rect 355 -35 405 -5
rect 435 -35 485 -5
rect 515 -35 565 -5
rect 595 -35 645 -5
rect 675 -35 725 -5
rect 755 -35 805 -5
rect 835 -35 885 -5
rect 915 -35 965 -5
rect 995 -35 1045 -5
rect 1075 -35 1125 -5
rect 1155 -35 1205 -5
rect 1235 -35 1285 -5
rect 1315 -35 1365 -5
rect 1395 -35 1445 -5
rect 1475 -35 1525 -5
rect 1555 -35 1605 -5
rect 1635 -35 1685 -5
rect 1715 -35 1765 -5
rect 1795 -35 1845 -5
rect 1875 -35 1925 -5
rect 1955 -35 2005 -5
rect 2035 -35 2085 -5
rect 2115 -35 2165 -5
rect 2195 -35 2245 -5
rect 2275 -35 2325 -5
rect 2355 -35 2405 -5
rect 2435 -35 2485 -5
rect 2515 -35 2565 -5
rect 2595 -35 2645 -5
rect 2675 -35 2725 -5
rect 2755 -35 2805 -5
rect 2835 -35 2885 -5
rect 2915 -35 2965 -5
rect 2995 -35 3045 -5
rect 3075 -35 3125 -5
rect 3155 -35 3205 -5
rect 3235 -35 3285 -5
rect 3315 -35 3365 -5
rect 3395 -35 3445 -5
rect 3475 -35 3525 -5
rect 3555 -35 3605 -5
rect 3635 -35 3685 -5
rect 3715 -35 3765 -5
rect 3795 -35 3845 -5
rect 3875 -35 3925 -5
rect 3955 -35 4005 -5
rect 4035 -35 4085 -5
rect 4115 -35 4165 -5
rect 4195 -35 4245 -5
rect 4275 -35 4325 -5
rect 4355 -35 4405 -5
rect 4435 -35 4485 -5
rect 4515 -35 4565 -5
rect 4595 -35 4645 -5
rect 4675 -35 4725 -5
rect 4755 -35 4805 -5
rect 4835 -35 4885 -5
rect 4915 -35 4965 -5
rect 4995 -35 5045 -5
rect 5075 -35 5125 -5
rect 5155 -35 5205 -5
rect 5235 -35 5285 -5
rect 5315 -35 5365 -5
rect 5395 -35 5445 -5
rect 5475 -35 5525 -5
rect 5555 -35 5605 -5
rect 5635 -35 5685 -5
rect 5715 -35 5765 -5
rect 5795 -35 5845 -5
rect 5875 -35 5925 -5
rect 5955 -35 6005 -5
rect 6035 -35 6085 -5
rect 6115 -35 6165 -5
rect 6195 -35 6245 -5
rect 6275 -35 6325 -5
rect 6355 -35 6405 -5
rect 6435 -35 6485 -5
rect 6515 -35 6565 -5
rect 6595 -35 6645 -5
rect 6675 -35 6725 -5
rect 6755 -35 6805 -5
rect 6835 -35 6885 -5
rect 6915 -35 6965 -5
rect 6995 -35 7045 -5
rect 7075 -35 7125 -5
rect 7155 -35 7205 -5
rect 7235 -35 7285 -5
rect 7315 -35 7365 -5
rect 7395 -35 7445 -5
rect 7475 -35 7525 -5
rect 7555 -35 7605 -5
rect 7635 -35 7685 -5
rect 7715 -35 7765 -5
rect 7795 -35 7845 -5
rect 7875 -35 7925 -5
rect 7955 -35 8005 -5
rect 8035 -35 8085 -5
rect 8115 -35 8165 -5
rect 8195 -35 8245 -5
rect 8275 -35 8325 -5
rect 8355 -35 8405 -5
rect 8435 -35 8485 -5
rect 8515 -35 8565 -5
rect 8595 -35 8645 -5
rect 8675 -35 8725 -5
rect 8755 -35 8805 -5
rect 8835 -35 8885 -5
rect 8915 -35 8965 -5
rect 8995 -35 9045 -5
rect 9075 -35 9125 -5
rect 9155 -35 9205 -5
rect 9235 -35 9285 -5
rect 9315 -35 9365 -5
rect 9395 -35 9445 -5
rect 9475 -35 9525 -5
rect 9555 -35 9605 -5
rect 9635 -35 9685 -5
rect 9715 -35 9765 -5
rect 9795 -35 9845 -5
rect 9875 -35 9925 -5
rect 9955 -35 10005 -5
rect 10035 -35 10085 -5
rect 10115 -35 10165 -5
rect 10195 -35 10245 -5
rect 10275 -35 10325 -5
rect 10355 -35 10405 -5
rect 10435 -35 10485 -5
rect 10515 -35 10645 -5
rect 10675 -35 10805 -5
rect 10835 -35 10965 -5
rect 10995 -35 11000 -5
rect -720 -40 11000 -35
rect -720 -85 11000 -80
rect -720 -115 -715 -85
rect -685 -115 -555 -85
rect -525 -115 -395 -85
rect -365 -115 -315 -85
rect -285 -115 -235 -85
rect -205 -115 -155 -85
rect -125 -115 -75 -85
rect -45 -115 5 -85
rect 35 -115 85 -85
rect 115 -115 165 -85
rect 195 -115 245 -85
rect 275 -115 325 -85
rect 355 -115 405 -85
rect 435 -115 485 -85
rect 515 -115 565 -85
rect 595 -115 645 -85
rect 675 -115 725 -85
rect 755 -115 805 -85
rect 835 -115 885 -85
rect 915 -115 965 -85
rect 995 -115 1045 -85
rect 1075 -115 1125 -85
rect 1155 -115 1205 -85
rect 1235 -115 1285 -85
rect 1315 -115 1365 -85
rect 1395 -115 1445 -85
rect 1475 -115 1525 -85
rect 1555 -115 1605 -85
rect 1635 -115 1685 -85
rect 1715 -115 1765 -85
rect 1795 -115 1845 -85
rect 1875 -115 1925 -85
rect 1955 -115 2005 -85
rect 2035 -115 2085 -85
rect 2115 -115 2165 -85
rect 2195 -115 2245 -85
rect 2275 -115 2325 -85
rect 2355 -115 2405 -85
rect 2435 -115 2485 -85
rect 2515 -115 2565 -85
rect 2595 -115 2645 -85
rect 2675 -115 2725 -85
rect 2755 -115 2805 -85
rect 2835 -115 2885 -85
rect 2915 -115 2965 -85
rect 2995 -115 3045 -85
rect 3075 -115 3125 -85
rect 3155 -115 3205 -85
rect 3235 -115 3285 -85
rect 3315 -115 3365 -85
rect 3395 -115 3445 -85
rect 3475 -115 3525 -85
rect 3555 -115 3605 -85
rect 3635 -115 3685 -85
rect 3715 -115 3765 -85
rect 3795 -115 3845 -85
rect 3875 -115 3925 -85
rect 3955 -115 4005 -85
rect 4035 -115 4085 -85
rect 4115 -115 4165 -85
rect 4195 -115 4245 -85
rect 4275 -115 4325 -85
rect 4355 -115 4405 -85
rect 4435 -115 4485 -85
rect 4515 -115 4565 -85
rect 4595 -115 4645 -85
rect 4675 -115 4725 -85
rect 4755 -115 4805 -85
rect 4835 -115 4885 -85
rect 4915 -115 4965 -85
rect 4995 -115 5045 -85
rect 5075 -115 5125 -85
rect 5155 -115 5205 -85
rect 5235 -115 5285 -85
rect 5315 -115 5365 -85
rect 5395 -115 5445 -85
rect 5475 -115 5525 -85
rect 5555 -115 5605 -85
rect 5635 -115 5685 -85
rect 5715 -115 5765 -85
rect 5795 -115 5845 -85
rect 5875 -115 5925 -85
rect 5955 -115 6005 -85
rect 6035 -115 6085 -85
rect 6115 -115 6165 -85
rect 6195 -115 6245 -85
rect 6275 -115 6325 -85
rect 6355 -115 6405 -85
rect 6435 -115 6485 -85
rect 6515 -115 6565 -85
rect 6595 -115 6645 -85
rect 6675 -115 6725 -85
rect 6755 -115 6805 -85
rect 6835 -115 6885 -85
rect 6915 -115 6965 -85
rect 6995 -115 7045 -85
rect 7075 -115 7125 -85
rect 7155 -115 7205 -85
rect 7235 -115 7285 -85
rect 7315 -115 7365 -85
rect 7395 -115 7445 -85
rect 7475 -115 7525 -85
rect 7555 -115 7605 -85
rect 7635 -115 7685 -85
rect 7715 -115 7765 -85
rect 7795 -115 7845 -85
rect 7875 -115 7925 -85
rect 7955 -115 8005 -85
rect 8035 -115 8085 -85
rect 8115 -115 8165 -85
rect 8195 -115 8245 -85
rect 8275 -115 8325 -85
rect 8355 -115 8405 -85
rect 8435 -115 8485 -85
rect 8515 -115 8565 -85
rect 8595 -115 8645 -85
rect 8675 -115 8725 -85
rect 8755 -115 8805 -85
rect 8835 -115 8885 -85
rect 8915 -115 8965 -85
rect 8995 -115 9045 -85
rect 9075 -115 9125 -85
rect 9155 -115 9205 -85
rect 9235 -115 9285 -85
rect 9315 -115 9365 -85
rect 9395 -115 9445 -85
rect 9475 -115 9525 -85
rect 9555 -115 9605 -85
rect 9635 -115 9685 -85
rect 9715 -115 9765 -85
rect 9795 -115 9845 -85
rect 9875 -115 9925 -85
rect 9955 -115 10005 -85
rect 10035 -115 10085 -85
rect 10115 -115 10165 -85
rect 10195 -115 10245 -85
rect 10275 -115 10325 -85
rect 10355 -115 10405 -85
rect 10435 -115 10485 -85
rect 10515 -115 10645 -85
rect 10675 -115 10805 -85
rect 10835 -115 10965 -85
rect 10995 -115 11000 -85
rect -720 -120 11000 -115
rect -720 -165 11000 -160
rect -720 -195 -715 -165
rect -685 -195 -555 -165
rect -525 -195 -395 -165
rect -365 -195 -235 -165
rect -205 -195 -155 -165
rect -125 -195 -75 -165
rect -45 -195 5 -165
rect 35 -195 85 -165
rect 115 -195 165 -165
rect 195 -195 245 -165
rect 275 -195 325 -165
rect 355 -195 405 -165
rect 435 -195 485 -165
rect 515 -195 565 -165
rect 595 -195 645 -165
rect 675 -195 725 -165
rect 755 -195 805 -165
rect 835 -195 885 -165
rect 915 -195 965 -165
rect 995 -195 1045 -165
rect 1075 -195 1125 -165
rect 1155 -195 1205 -165
rect 1235 -195 1285 -165
rect 1315 -195 1365 -165
rect 1395 -195 1445 -165
rect 1475 -195 1525 -165
rect 1555 -195 1605 -165
rect 1635 -195 1685 -165
rect 1715 -195 1765 -165
rect 1795 -195 1845 -165
rect 1875 -195 1925 -165
rect 1955 -195 2005 -165
rect 2035 -195 2085 -165
rect 2115 -195 2165 -165
rect 2195 -195 2245 -165
rect 2275 -195 2325 -165
rect 2355 -195 2405 -165
rect 2435 -195 2485 -165
rect 2515 -195 2565 -165
rect 2595 -195 2645 -165
rect 2675 -195 2725 -165
rect 2755 -195 2805 -165
rect 2835 -195 2885 -165
rect 2915 -195 2965 -165
rect 2995 -195 3045 -165
rect 3075 -195 3125 -165
rect 3155 -195 3205 -165
rect 3235 -195 3285 -165
rect 3315 -195 3365 -165
rect 3395 -195 3445 -165
rect 3475 -195 3525 -165
rect 3555 -195 3605 -165
rect 3635 -195 3685 -165
rect 3715 -195 3765 -165
rect 3795 -195 3845 -165
rect 3875 -195 3925 -165
rect 3955 -195 4005 -165
rect 4035 -195 4085 -165
rect 4115 -195 4165 -165
rect 4195 -195 4245 -165
rect 4275 -195 4325 -165
rect 4355 -195 4405 -165
rect 4435 -195 4485 -165
rect 4515 -195 4565 -165
rect 4595 -195 4645 -165
rect 4675 -195 4725 -165
rect 4755 -195 4805 -165
rect 4835 -195 4885 -165
rect 4915 -195 4965 -165
rect 4995 -195 5045 -165
rect 5075 -195 5125 -165
rect 5155 -195 5205 -165
rect 5235 -195 5285 -165
rect 5315 -195 5365 -165
rect 5395 -195 5445 -165
rect 5475 -195 5525 -165
rect 5555 -195 5605 -165
rect 5635 -195 5685 -165
rect 5715 -195 5765 -165
rect 5795 -195 5845 -165
rect 5875 -195 5925 -165
rect 5955 -195 6005 -165
rect 6035 -195 6085 -165
rect 6115 -195 6165 -165
rect 6195 -195 6245 -165
rect 6275 -195 6325 -165
rect 6355 -195 6405 -165
rect 6435 -195 6485 -165
rect 6515 -195 6565 -165
rect 6595 -195 6645 -165
rect 6675 -195 6725 -165
rect 6755 -195 6805 -165
rect 6835 -195 6885 -165
rect 6915 -195 6965 -165
rect 6995 -195 7045 -165
rect 7075 -195 7125 -165
rect 7155 -195 7205 -165
rect 7235 -195 7285 -165
rect 7315 -195 7365 -165
rect 7395 -195 7445 -165
rect 7475 -195 7525 -165
rect 7555 -195 7605 -165
rect 7635 -195 7685 -165
rect 7715 -195 7765 -165
rect 7795 -195 7845 -165
rect 7875 -195 7925 -165
rect 7955 -195 8005 -165
rect 8035 -195 8085 -165
rect 8115 -195 8165 -165
rect 8195 -195 8245 -165
rect 8275 -195 8325 -165
rect 8355 -195 8405 -165
rect 8435 -195 8485 -165
rect 8515 -195 8565 -165
rect 8595 -195 8645 -165
rect 8675 -195 8725 -165
rect 8755 -195 8805 -165
rect 8835 -195 8885 -165
rect 8915 -195 8965 -165
rect 8995 -195 9045 -165
rect 9075 -195 9125 -165
rect 9155 -195 9205 -165
rect 9235 -195 9285 -165
rect 9315 -195 9365 -165
rect 9395 -195 9445 -165
rect 9475 -195 9525 -165
rect 9555 -195 9605 -165
rect 9635 -195 9685 -165
rect 9715 -195 9765 -165
rect 9795 -195 9845 -165
rect 9875 -195 9925 -165
rect 9955 -195 10005 -165
rect 10035 -195 10085 -165
rect 10115 -195 10165 -165
rect 10195 -195 10245 -165
rect 10275 -195 10325 -165
rect 10355 -195 10405 -165
rect 10435 -195 10485 -165
rect 10515 -195 10565 -165
rect 10595 -195 10645 -165
rect 10675 -195 10805 -165
rect 10835 -195 10965 -165
rect 10995 -195 11000 -165
rect -720 -200 11000 -195
rect -720 -245 11000 -240
rect -720 -275 -715 -245
rect -685 -275 -555 -245
rect -525 -275 -395 -245
rect -365 -275 -235 -245
rect -205 -275 -155 -245
rect -125 -275 -75 -245
rect -45 -275 5 -245
rect 35 -275 85 -245
rect 115 -275 165 -245
rect 195 -275 245 -245
rect 275 -275 325 -245
rect 355 -275 405 -245
rect 435 -275 485 -245
rect 515 -275 565 -245
rect 595 -275 645 -245
rect 675 -275 725 -245
rect 755 -275 805 -245
rect 835 -275 885 -245
rect 915 -275 965 -245
rect 995 -275 1045 -245
rect 1075 -275 1125 -245
rect 1155 -275 1205 -245
rect 1235 -275 1285 -245
rect 1315 -275 1365 -245
rect 1395 -275 1445 -245
rect 1475 -275 1525 -245
rect 1555 -275 1605 -245
rect 1635 -275 1685 -245
rect 1715 -275 1765 -245
rect 1795 -275 1845 -245
rect 1875 -275 1925 -245
rect 1955 -275 2005 -245
rect 2035 -275 2085 -245
rect 2115 -275 2165 -245
rect 2195 -275 2245 -245
rect 2275 -275 2325 -245
rect 2355 -275 2405 -245
rect 2435 -275 2485 -245
rect 2515 -275 2565 -245
rect 2595 -275 2645 -245
rect 2675 -275 2725 -245
rect 2755 -275 2805 -245
rect 2835 -275 2885 -245
rect 2915 -275 2965 -245
rect 2995 -275 3045 -245
rect 3075 -275 3125 -245
rect 3155 -275 3205 -245
rect 3235 -275 3285 -245
rect 3315 -275 3365 -245
rect 3395 -275 3445 -245
rect 3475 -275 3525 -245
rect 3555 -275 3605 -245
rect 3635 -275 3685 -245
rect 3715 -275 3765 -245
rect 3795 -275 3845 -245
rect 3875 -275 3925 -245
rect 3955 -275 4005 -245
rect 4035 -275 4085 -245
rect 4115 -275 4165 -245
rect 4195 -275 4245 -245
rect 4275 -275 4325 -245
rect 4355 -275 4405 -245
rect 4435 -275 4485 -245
rect 4515 -275 4565 -245
rect 4595 -275 4645 -245
rect 4675 -275 4725 -245
rect 4755 -275 4805 -245
rect 4835 -275 4885 -245
rect 4915 -275 4965 -245
rect 4995 -275 5045 -245
rect 5075 -275 5125 -245
rect 5155 -275 5205 -245
rect 5235 -275 5285 -245
rect 5315 -275 5365 -245
rect 5395 -275 5445 -245
rect 5475 -275 5525 -245
rect 5555 -275 5605 -245
rect 5635 -275 5685 -245
rect 5715 -275 5765 -245
rect 5795 -275 5845 -245
rect 5875 -275 5925 -245
rect 5955 -275 6005 -245
rect 6035 -275 6085 -245
rect 6115 -275 6165 -245
rect 6195 -275 6245 -245
rect 6275 -275 6325 -245
rect 6355 -275 6405 -245
rect 6435 -275 6485 -245
rect 6515 -275 6565 -245
rect 6595 -275 6645 -245
rect 6675 -275 6725 -245
rect 6755 -275 6805 -245
rect 6835 -275 6885 -245
rect 6915 -275 6965 -245
rect 6995 -275 7045 -245
rect 7075 -275 7125 -245
rect 7155 -275 7205 -245
rect 7235 -275 7285 -245
rect 7315 -275 7365 -245
rect 7395 -275 7445 -245
rect 7475 -275 7525 -245
rect 7555 -275 7605 -245
rect 7635 -275 7685 -245
rect 7715 -275 7765 -245
rect 7795 -275 7845 -245
rect 7875 -275 7925 -245
rect 7955 -275 8005 -245
rect 8035 -275 8085 -245
rect 8115 -275 8165 -245
rect 8195 -275 8245 -245
rect 8275 -275 8325 -245
rect 8355 -275 8405 -245
rect 8435 -275 8485 -245
rect 8515 -275 8565 -245
rect 8595 -275 8645 -245
rect 8675 -275 8725 -245
rect 8755 -275 8805 -245
rect 8835 -275 8885 -245
rect 8915 -275 8965 -245
rect 8995 -275 9045 -245
rect 9075 -275 9125 -245
rect 9155 -275 9205 -245
rect 9235 -275 9285 -245
rect 9315 -275 9365 -245
rect 9395 -275 9445 -245
rect 9475 -275 9525 -245
rect 9555 -275 9605 -245
rect 9635 -275 9685 -245
rect 9715 -275 9765 -245
rect 9795 -275 9845 -245
rect 9875 -275 9925 -245
rect 9955 -275 10005 -245
rect 10035 -275 10085 -245
rect 10115 -275 10165 -245
rect 10195 -275 10245 -245
rect 10275 -275 10325 -245
rect 10355 -275 10405 -245
rect 10435 -275 10485 -245
rect 10515 -275 10565 -245
rect 10595 -275 10645 -245
rect 10675 -275 10805 -245
rect 10835 -275 10965 -245
rect 10995 -275 11000 -245
rect -720 -280 11000 -275
rect -720 -325 11000 -320
rect -720 -355 -715 -325
rect -685 -355 -555 -325
rect -525 -355 -395 -325
rect -365 -355 -235 -325
rect -205 -355 -155 -325
rect -125 -355 -75 -325
rect -45 -355 5 -325
rect 35 -355 85 -325
rect 115 -355 165 -325
rect 195 -355 245 -325
rect 275 -355 325 -325
rect 355 -355 405 -325
rect 435 -355 485 -325
rect 515 -355 565 -325
rect 595 -355 645 -325
rect 675 -355 725 -325
rect 755 -355 805 -325
rect 835 -355 885 -325
rect 915 -355 965 -325
rect 995 -355 1045 -325
rect 1075 -355 1125 -325
rect 1155 -355 1205 -325
rect 1235 -355 1285 -325
rect 1315 -355 1365 -325
rect 1395 -355 1445 -325
rect 1475 -355 1525 -325
rect 1555 -355 1605 -325
rect 1635 -355 1685 -325
rect 1715 -355 1765 -325
rect 1795 -355 1845 -325
rect 1875 -355 1925 -325
rect 1955 -355 2005 -325
rect 2035 -355 2085 -325
rect 2115 -355 2165 -325
rect 2195 -355 2245 -325
rect 2275 -355 2325 -325
rect 2355 -355 2405 -325
rect 2435 -355 2485 -325
rect 2515 -355 2565 -325
rect 2595 -355 2645 -325
rect 2675 -355 2725 -325
rect 2755 -355 2805 -325
rect 2835 -355 2885 -325
rect 2915 -355 2965 -325
rect 2995 -355 3045 -325
rect 3075 -355 3125 -325
rect 3155 -355 3205 -325
rect 3235 -355 3285 -325
rect 3315 -355 3365 -325
rect 3395 -355 3445 -325
rect 3475 -355 3525 -325
rect 3555 -355 3605 -325
rect 3635 -355 3685 -325
rect 3715 -355 3765 -325
rect 3795 -355 3845 -325
rect 3875 -355 3925 -325
rect 3955 -355 4005 -325
rect 4035 -355 4085 -325
rect 4115 -355 4165 -325
rect 4195 -355 4245 -325
rect 4275 -355 4325 -325
rect 4355 -355 4405 -325
rect 4435 -355 4485 -325
rect 4515 -355 4565 -325
rect 4595 -355 4645 -325
rect 4675 -355 4725 -325
rect 4755 -355 4805 -325
rect 4835 -355 4885 -325
rect 4915 -355 4965 -325
rect 4995 -355 5045 -325
rect 5075 -355 5125 -325
rect 5155 -355 5205 -325
rect 5235 -355 5285 -325
rect 5315 -355 5365 -325
rect 5395 -355 5445 -325
rect 5475 -355 5525 -325
rect 5555 -355 5605 -325
rect 5635 -355 5685 -325
rect 5715 -355 5765 -325
rect 5795 -355 5845 -325
rect 5875 -355 5925 -325
rect 5955 -355 6005 -325
rect 6035 -355 6085 -325
rect 6115 -355 6165 -325
rect 6195 -355 6245 -325
rect 6275 -355 6325 -325
rect 6355 -355 6405 -325
rect 6435 -355 6485 -325
rect 6515 -355 6565 -325
rect 6595 -355 6645 -325
rect 6675 -355 6725 -325
rect 6755 -355 6805 -325
rect 6835 -355 6885 -325
rect 6915 -355 6965 -325
rect 6995 -355 7045 -325
rect 7075 -355 7125 -325
rect 7155 -355 7205 -325
rect 7235 -355 7285 -325
rect 7315 -355 7365 -325
rect 7395 -355 7445 -325
rect 7475 -355 7525 -325
rect 7555 -355 7605 -325
rect 7635 -355 7685 -325
rect 7715 -355 7765 -325
rect 7795 -355 7845 -325
rect 7875 -355 7925 -325
rect 7955 -355 8005 -325
rect 8035 -355 8085 -325
rect 8115 -355 8165 -325
rect 8195 -355 8245 -325
rect 8275 -355 8325 -325
rect 8355 -355 8405 -325
rect 8435 -355 8485 -325
rect 8515 -355 8565 -325
rect 8595 -355 8645 -325
rect 8675 -355 8725 -325
rect 8755 -355 8805 -325
rect 8835 -355 8885 -325
rect 8915 -355 8965 -325
rect 8995 -355 9045 -325
rect 9075 -355 9125 -325
rect 9155 -355 9205 -325
rect 9235 -355 9285 -325
rect 9315 -355 9365 -325
rect 9395 -355 9445 -325
rect 9475 -355 9525 -325
rect 9555 -355 9605 -325
rect 9635 -355 9685 -325
rect 9715 -355 9765 -325
rect 9795 -355 9845 -325
rect 9875 -355 9925 -325
rect 9955 -355 10005 -325
rect 10035 -355 10085 -325
rect 10115 -355 10165 -325
rect 10195 -355 10245 -325
rect 10275 -355 10325 -325
rect 10355 -355 10405 -325
rect 10435 -355 10485 -325
rect 10515 -355 10565 -325
rect 10595 -355 10645 -325
rect 10675 -355 10805 -325
rect 10835 -355 10965 -325
rect 10995 -355 11000 -325
rect -720 -360 11000 -355
rect -720 -405 -360 -400
rect -720 -435 -715 -405
rect -685 -435 -555 -405
rect -525 -435 -395 -405
rect -365 -435 -360 -405
rect -720 -440 -360 -435
rect -320 -405 10760 -400
rect -320 -435 10 -405
rect 190 -435 330 -405
rect 510 -435 650 -405
rect 830 -435 970 -405
rect 1150 -435 1290 -405
rect 1470 -435 1610 -405
rect 1790 -435 1930 -405
rect 2110 -435 2250 -405
rect 2430 -435 2570 -405
rect 2750 -435 2890 -405
rect 3070 -435 3210 -405
rect 3390 -435 3530 -405
rect 3710 -435 3850 -405
rect 4030 -435 4170 -405
rect 4350 -435 4490 -405
rect 4670 -435 4810 -405
rect 4990 -435 5205 -405
rect 5235 -435 5290 -405
rect 5470 -435 5610 -405
rect 5790 -435 5930 -405
rect 6110 -435 6250 -405
rect 6430 -435 6485 -405
rect 6515 -435 6570 -405
rect 6750 -435 6890 -405
rect 7070 -435 7210 -405
rect 7390 -435 7530 -405
rect 7710 -435 7850 -405
rect 8030 -435 8170 -405
rect 8350 -435 8490 -405
rect 8670 -435 8810 -405
rect 8990 -435 9045 -405
rect 9075 -435 9130 -405
rect 9310 -435 9450 -405
rect 9630 -435 9770 -405
rect 9950 -435 10090 -405
rect 10270 -435 10725 -405
rect 10755 -435 10760 -405
rect -320 -440 10760 -435
rect 10800 -405 11000 -400
rect 10800 -435 10805 -405
rect 10835 -435 10965 -405
rect 10995 -435 11000 -405
rect 10800 -440 11000 -435
rect -720 -485 11000 -480
rect -720 -515 -715 -485
rect -685 -515 -555 -485
rect -525 -515 -395 -485
rect -365 -515 -235 -485
rect -205 -515 -155 -485
rect -125 -515 -75 -485
rect -45 -515 5 -485
rect 35 -515 85 -485
rect 115 -515 165 -485
rect 195 -515 245 -485
rect 275 -515 325 -485
rect 355 -515 405 -485
rect 435 -515 485 -485
rect 515 -515 565 -485
rect 595 -515 645 -485
rect 675 -515 725 -485
rect 755 -515 805 -485
rect 835 -515 885 -485
rect 915 -515 965 -485
rect 995 -515 1045 -485
rect 1075 -515 1125 -485
rect 1155 -515 1205 -485
rect 1235 -515 1285 -485
rect 1315 -515 1365 -485
rect 1395 -515 1445 -485
rect 1475 -515 1525 -485
rect 1555 -515 1605 -485
rect 1635 -515 1685 -485
rect 1715 -515 1765 -485
rect 1795 -515 1845 -485
rect 1875 -515 1925 -485
rect 1955 -515 2005 -485
rect 2035 -515 2085 -485
rect 2115 -515 2165 -485
rect 2195 -515 2245 -485
rect 2275 -515 2325 -485
rect 2355 -515 2405 -485
rect 2435 -515 2485 -485
rect 2515 -515 2565 -485
rect 2595 -515 2645 -485
rect 2675 -515 2725 -485
rect 2755 -515 2805 -485
rect 2835 -515 2885 -485
rect 2915 -515 2965 -485
rect 2995 -515 3045 -485
rect 3075 -515 3125 -485
rect 3155 -515 3205 -485
rect 3235 -515 3285 -485
rect 3315 -515 3365 -485
rect 3395 -515 3445 -485
rect 3475 -515 3525 -485
rect 3555 -515 3605 -485
rect 3635 -515 3685 -485
rect 3715 -515 3765 -485
rect 3795 -515 3845 -485
rect 3875 -515 3925 -485
rect 3955 -515 4005 -485
rect 4035 -515 4085 -485
rect 4115 -515 4165 -485
rect 4195 -515 4245 -485
rect 4275 -515 4325 -485
rect 4355 -515 4405 -485
rect 4435 -515 4485 -485
rect 4515 -515 4565 -485
rect 4595 -515 4645 -485
rect 4675 -515 4725 -485
rect 4755 -515 4805 -485
rect 4835 -515 4885 -485
rect 4915 -515 4965 -485
rect 4995 -515 5045 -485
rect 5075 -515 5125 -485
rect 5155 -515 5205 -485
rect 5235 -515 5285 -485
rect 5315 -515 5365 -485
rect 5395 -515 5445 -485
rect 5475 -515 5525 -485
rect 5555 -515 5605 -485
rect 5635 -515 5685 -485
rect 5715 -515 5765 -485
rect 5795 -515 5845 -485
rect 5875 -515 5925 -485
rect 5955 -515 6005 -485
rect 6035 -515 6085 -485
rect 6115 -515 6165 -485
rect 6195 -515 6245 -485
rect 6275 -515 6325 -485
rect 6355 -515 6405 -485
rect 6435 -515 6485 -485
rect 6515 -515 6565 -485
rect 6595 -515 6645 -485
rect 6675 -515 6725 -485
rect 6755 -515 6805 -485
rect 6835 -515 6885 -485
rect 6915 -515 6965 -485
rect 6995 -515 7045 -485
rect 7075 -515 7125 -485
rect 7155 -515 7205 -485
rect 7235 -515 7285 -485
rect 7315 -515 7365 -485
rect 7395 -515 7445 -485
rect 7475 -515 7525 -485
rect 7555 -515 7605 -485
rect 7635 -515 7685 -485
rect 7715 -515 7765 -485
rect 7795 -515 7845 -485
rect 7875 -515 7925 -485
rect 7955 -515 8005 -485
rect 8035 -515 8085 -485
rect 8115 -515 8165 -485
rect 8195 -515 8245 -485
rect 8275 -515 8325 -485
rect 8355 -515 8405 -485
rect 8435 -515 8485 -485
rect 8515 -515 8565 -485
rect 8595 -515 8645 -485
rect 8675 -515 8725 -485
rect 8755 -515 8805 -485
rect 8835 -515 8885 -485
rect 8915 -515 8965 -485
rect 8995 -515 9045 -485
rect 9075 -515 9125 -485
rect 9155 -515 9205 -485
rect 9235 -515 9285 -485
rect 9315 -515 9365 -485
rect 9395 -515 9445 -485
rect 9475 -515 9525 -485
rect 9555 -515 9605 -485
rect 9635 -515 9685 -485
rect 9715 -515 9765 -485
rect 9795 -515 9845 -485
rect 9875 -515 9925 -485
rect 9955 -515 10005 -485
rect 10035 -515 10085 -485
rect 10115 -515 10165 -485
rect 10195 -515 10245 -485
rect 10275 -515 10325 -485
rect 10355 -515 10405 -485
rect 10435 -515 10485 -485
rect 10515 -515 10565 -485
rect 10595 -515 10645 -485
rect 10675 -515 10805 -485
rect 10835 -515 10965 -485
rect 10995 -515 11000 -485
rect -720 -520 11000 -515
rect -720 -565 -360 -560
rect -720 -595 -715 -565
rect -685 -595 -555 -565
rect -525 -595 -395 -565
rect -365 -595 -360 -565
rect -720 -600 -360 -595
rect -320 -565 10920 -560
rect -320 -595 85 -565
rect 115 -595 245 -565
rect 275 -595 405 -565
rect 435 -595 725 -565
rect 755 -595 885 -565
rect 915 -595 1045 -565
rect 1075 -595 1205 -565
rect 1235 -595 1365 -565
rect 1395 -595 1525 -565
rect 1555 -595 1685 -565
rect 1715 -595 2005 -565
rect 2035 -595 2165 -565
rect 2195 -595 2325 -565
rect 2355 -595 2645 -565
rect 2675 -595 2805 -565
rect 2835 -595 2965 -565
rect 2995 -595 3285 -565
rect 3315 -595 3445 -565
rect 3475 -595 3605 -565
rect 3635 -595 3765 -565
rect 3795 -595 3925 -565
rect 3955 -595 4085 -565
rect 4115 -595 4245 -565
rect 4275 -595 4565 -565
rect 4595 -595 4725 -565
rect 4755 -595 4885 -565
rect 4915 -595 10885 -565
rect 10915 -595 10920 -565
rect -320 -600 10920 -595
rect 10960 -600 11000 -560
rect -720 -645 11000 -640
rect -720 -675 -715 -645
rect -685 -675 -555 -645
rect -525 -675 -395 -645
rect -365 -675 -235 -645
rect -205 -675 -155 -645
rect -125 -675 -75 -645
rect -45 -675 5 -645
rect 35 -675 85 -645
rect 115 -675 165 -645
rect 195 -675 245 -645
rect 275 -675 325 -645
rect 355 -675 405 -645
rect 435 -675 485 -645
rect 515 -675 565 -645
rect 595 -675 645 -645
rect 675 -675 725 -645
rect 755 -675 805 -645
rect 835 -675 885 -645
rect 915 -675 965 -645
rect 995 -675 1045 -645
rect 1075 -675 1125 -645
rect 1155 -675 1205 -645
rect 1235 -675 1285 -645
rect 1315 -675 1365 -645
rect 1395 -675 1445 -645
rect 1475 -675 1525 -645
rect 1555 -675 1605 -645
rect 1635 -675 1685 -645
rect 1715 -675 1765 -645
rect 1795 -675 1845 -645
rect 1875 -675 1925 -645
rect 1955 -675 2005 -645
rect 2035 -675 2085 -645
rect 2115 -675 2165 -645
rect 2195 -675 2245 -645
rect 2275 -675 2325 -645
rect 2355 -675 2405 -645
rect 2435 -675 2485 -645
rect 2515 -675 2565 -645
rect 2595 -675 2645 -645
rect 2675 -675 2725 -645
rect 2755 -675 2805 -645
rect 2835 -675 2885 -645
rect 2915 -675 2965 -645
rect 2995 -675 3045 -645
rect 3075 -675 3125 -645
rect 3155 -675 3205 -645
rect 3235 -675 3285 -645
rect 3315 -675 3365 -645
rect 3395 -675 3445 -645
rect 3475 -675 3525 -645
rect 3555 -675 3605 -645
rect 3635 -675 3685 -645
rect 3715 -675 3765 -645
rect 3795 -675 3845 -645
rect 3875 -675 3925 -645
rect 3955 -675 4005 -645
rect 4035 -675 4085 -645
rect 4115 -675 4165 -645
rect 4195 -675 4245 -645
rect 4275 -675 4325 -645
rect 4355 -675 4405 -645
rect 4435 -675 4485 -645
rect 4515 -675 4565 -645
rect 4595 -675 4645 -645
rect 4675 -675 4725 -645
rect 4755 -675 4805 -645
rect 4835 -675 4885 -645
rect 4915 -675 4965 -645
rect 4995 -675 5045 -645
rect 5075 -675 5125 -645
rect 5155 -675 5205 -645
rect 5235 -675 5285 -645
rect 5315 -675 5365 -645
rect 5395 -675 5445 -645
rect 5475 -675 5525 -645
rect 5555 -675 5605 -645
rect 5635 -675 5685 -645
rect 5715 -675 5765 -645
rect 5795 -675 5845 -645
rect 5875 -675 5925 -645
rect 5955 -675 6005 -645
rect 6035 -675 6085 -645
rect 6115 -675 6165 -645
rect 6195 -675 6245 -645
rect 6275 -675 6325 -645
rect 6355 -675 6405 -645
rect 6435 -675 6485 -645
rect 6515 -675 6565 -645
rect 6595 -675 6645 -645
rect 6675 -675 6725 -645
rect 6755 -675 6805 -645
rect 6835 -675 6885 -645
rect 6915 -675 6965 -645
rect 6995 -675 7045 -645
rect 7075 -675 7125 -645
rect 7155 -675 7205 -645
rect 7235 -675 7285 -645
rect 7315 -675 7365 -645
rect 7395 -675 7445 -645
rect 7475 -675 7525 -645
rect 7555 -675 7605 -645
rect 7635 -675 7685 -645
rect 7715 -675 7765 -645
rect 7795 -675 7845 -645
rect 7875 -675 7925 -645
rect 7955 -675 8005 -645
rect 8035 -675 8085 -645
rect 8115 -675 8165 -645
rect 8195 -675 8245 -645
rect 8275 -675 8325 -645
rect 8355 -675 8405 -645
rect 8435 -675 8485 -645
rect 8515 -675 8565 -645
rect 8595 -675 8645 -645
rect 8675 -675 8725 -645
rect 8755 -675 8805 -645
rect 8835 -675 8885 -645
rect 8915 -675 8965 -645
rect 8995 -675 9045 -645
rect 9075 -675 9125 -645
rect 9155 -675 9205 -645
rect 9235 -675 9285 -645
rect 9315 -675 9365 -645
rect 9395 -675 9445 -645
rect 9475 -675 9525 -645
rect 9555 -675 9605 -645
rect 9635 -675 9685 -645
rect 9715 -675 9765 -645
rect 9795 -675 9845 -645
rect 9875 -675 9925 -645
rect 9955 -675 10005 -645
rect 10035 -675 10085 -645
rect 10115 -675 10165 -645
rect 10195 -675 10245 -645
rect 10275 -675 10325 -645
rect 10355 -675 10405 -645
rect 10435 -675 10485 -645
rect 10515 -675 10565 -645
rect 10595 -675 10645 -645
rect 10675 -675 10805 -645
rect 10835 -675 10965 -645
rect 10995 -675 11000 -645
rect -720 -680 11000 -675
rect -720 -725 -520 -720
rect -720 -755 -715 -725
rect -685 -755 -555 -725
rect -525 -755 -520 -725
rect -720 -760 -520 -755
rect -480 -725 10600 -720
rect -480 -755 -475 -725
rect -445 -755 5365 -725
rect 5395 -755 5685 -725
rect 5715 -755 6005 -725
rect 6035 -755 6325 -725
rect 6355 -755 6645 -725
rect 6675 -755 6965 -725
rect 6995 -755 7285 -725
rect 7315 -755 7605 -725
rect 7635 -755 7925 -725
rect 7955 -755 8245 -725
rect 8275 -755 8565 -725
rect 8595 -755 8885 -725
rect 8915 -755 9205 -725
rect 9235 -755 9525 -725
rect 9555 -755 9845 -725
rect 9875 -755 10165 -725
rect 10195 -755 10600 -725
rect -480 -760 10600 -755
rect 10640 -725 11000 -720
rect 10640 -755 10645 -725
rect 10675 -755 10805 -725
rect 10835 -755 10965 -725
rect 10995 -755 11000 -725
rect 10640 -760 11000 -755
rect -720 -805 11000 -800
rect -720 -835 -715 -805
rect -685 -835 -555 -805
rect -525 -835 -395 -805
rect -365 -835 -235 -805
rect -205 -835 -155 -805
rect -125 -835 -75 -805
rect -45 -835 5 -805
rect 35 -835 85 -805
rect 115 -835 165 -805
rect 195 -835 245 -805
rect 275 -835 325 -805
rect 355 -835 405 -805
rect 435 -835 485 -805
rect 515 -835 565 -805
rect 595 -835 645 -805
rect 675 -835 725 -805
rect 755 -835 805 -805
rect 835 -835 885 -805
rect 915 -835 965 -805
rect 995 -835 1045 -805
rect 1075 -835 1125 -805
rect 1155 -835 1205 -805
rect 1235 -835 1285 -805
rect 1315 -835 1365 -805
rect 1395 -835 1445 -805
rect 1475 -835 1525 -805
rect 1555 -835 1605 -805
rect 1635 -835 1685 -805
rect 1715 -835 1765 -805
rect 1795 -835 1845 -805
rect 1875 -835 1925 -805
rect 1955 -835 2005 -805
rect 2035 -835 2085 -805
rect 2115 -835 2165 -805
rect 2195 -835 2245 -805
rect 2275 -835 2325 -805
rect 2355 -835 2405 -805
rect 2435 -835 2485 -805
rect 2515 -835 2565 -805
rect 2595 -835 2645 -805
rect 2675 -835 2725 -805
rect 2755 -835 2805 -805
rect 2835 -835 2885 -805
rect 2915 -835 2965 -805
rect 2995 -835 3045 -805
rect 3075 -835 3125 -805
rect 3155 -835 3205 -805
rect 3235 -835 3285 -805
rect 3315 -835 3365 -805
rect 3395 -835 3445 -805
rect 3475 -835 3525 -805
rect 3555 -835 3605 -805
rect 3635 -835 3685 -805
rect 3715 -835 3765 -805
rect 3795 -835 3845 -805
rect 3875 -835 3925 -805
rect 3955 -835 4005 -805
rect 4035 -835 4085 -805
rect 4115 -835 4165 -805
rect 4195 -835 4245 -805
rect 4275 -835 4325 -805
rect 4355 -835 4405 -805
rect 4435 -835 4485 -805
rect 4515 -835 4565 -805
rect 4595 -835 4645 -805
rect 4675 -835 4725 -805
rect 4755 -835 4805 -805
rect 4835 -835 4885 -805
rect 4915 -835 4965 -805
rect 4995 -835 5045 -805
rect 5075 -835 5125 -805
rect 5155 -835 5205 -805
rect 5235 -835 5285 -805
rect 5315 -835 5365 -805
rect 5395 -835 5445 -805
rect 5475 -835 5525 -805
rect 5555 -835 5605 -805
rect 5635 -835 5685 -805
rect 5715 -835 5765 -805
rect 5795 -835 5845 -805
rect 5875 -835 5925 -805
rect 5955 -835 6005 -805
rect 6035 -835 6085 -805
rect 6115 -835 6165 -805
rect 6195 -835 6245 -805
rect 6275 -835 6325 -805
rect 6355 -835 6405 -805
rect 6435 -835 6485 -805
rect 6515 -835 6565 -805
rect 6595 -835 6645 -805
rect 6675 -835 6725 -805
rect 6755 -835 6805 -805
rect 6835 -835 6885 -805
rect 6915 -835 6965 -805
rect 6995 -835 7045 -805
rect 7075 -835 7125 -805
rect 7155 -835 7205 -805
rect 7235 -835 7285 -805
rect 7315 -835 7365 -805
rect 7395 -835 7445 -805
rect 7475 -835 7525 -805
rect 7555 -835 7605 -805
rect 7635 -835 7685 -805
rect 7715 -835 7765 -805
rect 7795 -835 7845 -805
rect 7875 -835 7925 -805
rect 7955 -835 8005 -805
rect 8035 -835 8085 -805
rect 8115 -835 8165 -805
rect 8195 -835 8245 -805
rect 8275 -835 8325 -805
rect 8355 -835 8405 -805
rect 8435 -835 8485 -805
rect 8515 -835 8565 -805
rect 8595 -835 8645 -805
rect 8675 -835 8725 -805
rect 8755 -835 8805 -805
rect 8835 -835 8885 -805
rect 8915 -835 8965 -805
rect 8995 -835 9045 -805
rect 9075 -835 9125 -805
rect 9155 -835 9205 -805
rect 9235 -835 9285 -805
rect 9315 -835 9365 -805
rect 9395 -835 9445 -805
rect 9475 -835 9525 -805
rect 9555 -835 9605 -805
rect 9635 -835 9685 -805
rect 9715 -835 9765 -805
rect 9795 -835 9845 -805
rect 9875 -835 9925 -805
rect 9955 -835 10005 -805
rect 10035 -835 10085 -805
rect 10115 -835 10165 -805
rect 10195 -835 10245 -805
rect 10275 -835 10325 -805
rect 10355 -835 10405 -805
rect 10435 -835 10485 -805
rect 10515 -835 10565 -805
rect 10595 -835 10645 -805
rect 10675 -835 10805 -805
rect 10835 -835 10965 -805
rect 10995 -835 11000 -805
rect -720 -840 11000 -835
rect -720 -885 11000 -880
rect -720 -915 -715 -885
rect -685 -915 -555 -885
rect -525 -915 -395 -885
rect -365 -915 -235 -885
rect -205 -915 -155 -885
rect -125 -915 -75 -885
rect -45 -915 5 -885
rect 35 -915 85 -885
rect 115 -915 165 -885
rect 195 -915 245 -885
rect 275 -915 325 -885
rect 355 -915 405 -885
rect 435 -915 485 -885
rect 515 -915 565 -885
rect 595 -915 645 -885
rect 675 -915 725 -885
rect 755 -915 805 -885
rect 835 -915 885 -885
rect 915 -915 965 -885
rect 995 -915 1045 -885
rect 1075 -915 1125 -885
rect 1155 -915 1205 -885
rect 1235 -915 1285 -885
rect 1315 -915 1365 -885
rect 1395 -915 1445 -885
rect 1475 -915 1525 -885
rect 1555 -915 1605 -885
rect 1635 -915 1685 -885
rect 1715 -915 1765 -885
rect 1795 -915 1845 -885
rect 1875 -915 1925 -885
rect 1955 -915 2005 -885
rect 2035 -915 2085 -885
rect 2115 -915 2165 -885
rect 2195 -915 2245 -885
rect 2275 -915 2325 -885
rect 2355 -915 2405 -885
rect 2435 -915 2485 -885
rect 2515 -915 2565 -885
rect 2595 -915 2645 -885
rect 2675 -915 2725 -885
rect 2755 -915 2805 -885
rect 2835 -915 2885 -885
rect 2915 -915 2965 -885
rect 2995 -915 3045 -885
rect 3075 -915 3125 -885
rect 3155 -915 3205 -885
rect 3235 -915 3285 -885
rect 3315 -915 3365 -885
rect 3395 -915 3445 -885
rect 3475 -915 3525 -885
rect 3555 -915 3605 -885
rect 3635 -915 3685 -885
rect 3715 -915 3765 -885
rect 3795 -915 3845 -885
rect 3875 -915 3925 -885
rect 3955 -915 4005 -885
rect 4035 -915 4085 -885
rect 4115 -915 4165 -885
rect 4195 -915 4245 -885
rect 4275 -915 4325 -885
rect 4355 -915 4405 -885
rect 4435 -915 4485 -885
rect 4515 -915 4565 -885
rect 4595 -915 4645 -885
rect 4675 -915 4725 -885
rect 4755 -915 4805 -885
rect 4835 -915 4885 -885
rect 4915 -915 4965 -885
rect 4995 -915 5045 -885
rect 5075 -915 5125 -885
rect 5155 -915 5205 -885
rect 5235 -915 5285 -885
rect 5315 -915 5365 -885
rect 5395 -915 5445 -885
rect 5475 -915 5525 -885
rect 5555 -915 5605 -885
rect 5635 -915 5685 -885
rect 5715 -915 5765 -885
rect 5795 -915 5845 -885
rect 5875 -915 5925 -885
rect 5955 -915 6005 -885
rect 6035 -915 6085 -885
rect 6115 -915 6165 -885
rect 6195 -915 6245 -885
rect 6275 -915 6325 -885
rect 6355 -915 6405 -885
rect 6435 -915 6485 -885
rect 6515 -915 6565 -885
rect 6595 -915 6645 -885
rect 6675 -915 6725 -885
rect 6755 -915 6805 -885
rect 6835 -915 6885 -885
rect 6915 -915 6965 -885
rect 6995 -915 7045 -885
rect 7075 -915 7125 -885
rect 7155 -915 7205 -885
rect 7235 -915 7285 -885
rect 7315 -915 7365 -885
rect 7395 -915 7445 -885
rect 7475 -915 7525 -885
rect 7555 -915 7605 -885
rect 7635 -915 7685 -885
rect 7715 -915 7765 -885
rect 7795 -915 7845 -885
rect 7875 -915 7925 -885
rect 7955 -915 8005 -885
rect 8035 -915 8085 -885
rect 8115 -915 8165 -885
rect 8195 -915 8245 -885
rect 8275 -915 8325 -885
rect 8355 -915 8405 -885
rect 8435 -915 8485 -885
rect 8515 -915 8565 -885
rect 8595 -915 8645 -885
rect 8675 -915 8725 -885
rect 8755 -915 8805 -885
rect 8835 -915 8885 -885
rect 8915 -915 8965 -885
rect 8995 -915 9045 -885
rect 9075 -915 9125 -885
rect 9155 -915 9205 -885
rect 9235 -915 9285 -885
rect 9315 -915 9365 -885
rect 9395 -915 9445 -885
rect 9475 -915 9525 -885
rect 9555 -915 9605 -885
rect 9635 -915 9685 -885
rect 9715 -915 9765 -885
rect 9795 -915 9845 -885
rect 9875 -915 9925 -885
rect 9955 -915 10005 -885
rect 10035 -915 10085 -885
rect 10115 -915 10165 -885
rect 10195 -915 10245 -885
rect 10275 -915 10325 -885
rect 10355 -915 10405 -885
rect 10435 -915 10485 -885
rect 10515 -915 10565 -885
rect 10595 -915 10645 -885
rect 10675 -915 10805 -885
rect 10835 -915 10965 -885
rect 10995 -915 11000 -885
rect -720 -920 11000 -915
rect -640 -965 10600 -960
rect -640 -995 -635 -965
rect -605 -995 -75 -965
rect -45 -995 565 -965
rect 595 -995 1205 -965
rect 1235 -995 1845 -965
rect 1875 -995 2485 -965
rect 2515 -995 3125 -965
rect 3155 -995 3765 -965
rect 3795 -995 4405 -965
rect 4435 -995 5045 -965
rect 5075 -995 10325 -965
rect 10355 -995 10600 -965
rect -640 -1000 10600 -995
rect 10640 -965 11000 -960
rect 10640 -995 10645 -965
rect 10675 -995 10805 -965
rect 10835 -995 10965 -965
rect 10995 -995 11000 -965
rect 10640 -1000 11000 -995
rect -640 -1045 10600 -1040
rect -640 -1075 -635 -1045
rect -605 -1075 -75 -1045
rect -45 -1075 565 -1045
rect 595 -1075 1205 -1045
rect 1235 -1075 1845 -1045
rect 1875 -1075 2485 -1045
rect 2515 -1075 3125 -1045
rect 3155 -1075 3765 -1045
rect 3795 -1075 4405 -1045
rect 4435 -1075 5045 -1045
rect 5075 -1075 10325 -1045
rect 10355 -1075 10600 -1045
rect -640 -1080 10600 -1075
rect 10640 -1045 11000 -1040
rect 10640 -1075 10645 -1045
rect 10675 -1075 10805 -1045
rect 10835 -1075 10965 -1045
rect 10995 -1075 11000 -1045
rect 10640 -1080 11000 -1075
rect -720 -1125 11000 -1120
rect -720 -1155 -715 -1125
rect -685 -1155 -555 -1125
rect -525 -1155 -395 -1125
rect -365 -1155 -235 -1125
rect -205 -1155 -155 -1125
rect -125 -1155 -75 -1125
rect -45 -1155 5 -1125
rect 35 -1155 85 -1125
rect 115 -1155 165 -1125
rect 195 -1155 245 -1125
rect 275 -1155 325 -1125
rect 355 -1155 405 -1125
rect 435 -1155 485 -1125
rect 515 -1155 565 -1125
rect 595 -1155 645 -1125
rect 675 -1155 725 -1125
rect 755 -1155 805 -1125
rect 835 -1155 885 -1125
rect 915 -1155 965 -1125
rect 995 -1155 1045 -1125
rect 1075 -1155 1125 -1125
rect 1155 -1155 1205 -1125
rect 1235 -1155 1285 -1125
rect 1315 -1155 1365 -1125
rect 1395 -1155 1445 -1125
rect 1475 -1155 1525 -1125
rect 1555 -1155 1605 -1125
rect 1635 -1155 1685 -1125
rect 1715 -1155 1765 -1125
rect 1795 -1155 1845 -1125
rect 1875 -1155 1925 -1125
rect 1955 -1155 2005 -1125
rect 2035 -1155 2085 -1125
rect 2115 -1155 2165 -1125
rect 2195 -1155 2245 -1125
rect 2275 -1155 2325 -1125
rect 2355 -1155 2405 -1125
rect 2435 -1155 2485 -1125
rect 2515 -1155 2565 -1125
rect 2595 -1155 2645 -1125
rect 2675 -1155 2725 -1125
rect 2755 -1155 2805 -1125
rect 2835 -1155 2885 -1125
rect 2915 -1155 2965 -1125
rect 2995 -1155 3045 -1125
rect 3075 -1155 3125 -1125
rect 3155 -1155 3205 -1125
rect 3235 -1155 3285 -1125
rect 3315 -1155 3365 -1125
rect 3395 -1155 3445 -1125
rect 3475 -1155 3525 -1125
rect 3555 -1155 3605 -1125
rect 3635 -1155 3685 -1125
rect 3715 -1155 3765 -1125
rect 3795 -1155 3845 -1125
rect 3875 -1155 3925 -1125
rect 3955 -1155 4005 -1125
rect 4035 -1155 4085 -1125
rect 4115 -1155 4165 -1125
rect 4195 -1155 4245 -1125
rect 4275 -1155 4325 -1125
rect 4355 -1155 4405 -1125
rect 4435 -1155 4485 -1125
rect 4515 -1155 4565 -1125
rect 4595 -1155 4645 -1125
rect 4675 -1155 4725 -1125
rect 4755 -1155 4805 -1125
rect 4835 -1155 4885 -1125
rect 4915 -1155 4965 -1125
rect 4995 -1155 5045 -1125
rect 5075 -1155 5125 -1125
rect 5155 -1155 5205 -1125
rect 5235 -1155 5285 -1125
rect 5315 -1155 5365 -1125
rect 5395 -1155 5445 -1125
rect 5475 -1155 5525 -1125
rect 5555 -1155 5605 -1125
rect 5635 -1155 5685 -1125
rect 5715 -1155 5765 -1125
rect 5795 -1155 5845 -1125
rect 5875 -1155 5925 -1125
rect 5955 -1155 6005 -1125
rect 6035 -1155 6085 -1125
rect 6115 -1155 6165 -1125
rect 6195 -1155 6245 -1125
rect 6275 -1155 6325 -1125
rect 6355 -1155 6405 -1125
rect 6435 -1155 6485 -1125
rect 6515 -1155 6565 -1125
rect 6595 -1155 6645 -1125
rect 6675 -1155 6725 -1125
rect 6755 -1155 6805 -1125
rect 6835 -1155 6885 -1125
rect 6915 -1155 6965 -1125
rect 6995 -1155 7045 -1125
rect 7075 -1155 7125 -1125
rect 7155 -1155 7205 -1125
rect 7235 -1155 7285 -1125
rect 7315 -1155 7365 -1125
rect 7395 -1155 7445 -1125
rect 7475 -1155 7525 -1125
rect 7555 -1155 7605 -1125
rect 7635 -1155 7685 -1125
rect 7715 -1155 7765 -1125
rect 7795 -1155 7845 -1125
rect 7875 -1155 7925 -1125
rect 7955 -1155 8005 -1125
rect 8035 -1155 8085 -1125
rect 8115 -1155 8165 -1125
rect 8195 -1155 8245 -1125
rect 8275 -1155 8325 -1125
rect 8355 -1155 8405 -1125
rect 8435 -1155 8485 -1125
rect 8515 -1155 8565 -1125
rect 8595 -1155 8645 -1125
rect 8675 -1155 8725 -1125
rect 8755 -1155 8805 -1125
rect 8835 -1155 8885 -1125
rect 8915 -1155 8965 -1125
rect 8995 -1155 9045 -1125
rect 9075 -1155 9125 -1125
rect 9155 -1155 9205 -1125
rect 9235 -1155 9285 -1125
rect 9315 -1155 9365 -1125
rect 9395 -1155 9445 -1125
rect 9475 -1155 9525 -1125
rect 9555 -1155 9605 -1125
rect 9635 -1155 9685 -1125
rect 9715 -1155 9765 -1125
rect 9795 -1155 9845 -1125
rect 9875 -1155 9925 -1125
rect 9955 -1155 10005 -1125
rect 10035 -1155 10085 -1125
rect 10115 -1155 10165 -1125
rect 10195 -1155 10245 -1125
rect 10275 -1155 10325 -1125
rect 10355 -1155 10405 -1125
rect 10435 -1155 10485 -1125
rect 10515 -1155 10565 -1125
rect 10595 -1155 10645 -1125
rect 10675 -1155 10805 -1125
rect 10835 -1155 10965 -1125
rect 10995 -1155 11000 -1125
rect -720 -1160 11000 -1155
rect -720 -1205 11000 -1200
rect -720 -1235 -715 -1205
rect -685 -1235 -555 -1205
rect -525 -1235 -395 -1205
rect -365 -1235 -235 -1205
rect -205 -1235 -155 -1205
rect -125 -1235 -75 -1205
rect -45 -1235 5 -1205
rect 35 -1235 85 -1205
rect 115 -1235 165 -1205
rect 195 -1235 245 -1205
rect 275 -1235 325 -1205
rect 355 -1235 405 -1205
rect 435 -1235 485 -1205
rect 515 -1235 565 -1205
rect 595 -1235 645 -1205
rect 675 -1235 725 -1205
rect 755 -1235 805 -1205
rect 835 -1235 885 -1205
rect 915 -1235 965 -1205
rect 995 -1235 1045 -1205
rect 1075 -1235 1125 -1205
rect 1155 -1235 1205 -1205
rect 1235 -1235 1285 -1205
rect 1315 -1235 1365 -1205
rect 1395 -1235 1445 -1205
rect 1475 -1235 1525 -1205
rect 1555 -1235 1605 -1205
rect 1635 -1235 1685 -1205
rect 1715 -1235 1765 -1205
rect 1795 -1235 1845 -1205
rect 1875 -1235 1925 -1205
rect 1955 -1235 2005 -1205
rect 2035 -1235 2085 -1205
rect 2115 -1235 2165 -1205
rect 2195 -1235 2245 -1205
rect 2275 -1235 2325 -1205
rect 2355 -1235 2405 -1205
rect 2435 -1235 2485 -1205
rect 2515 -1235 2565 -1205
rect 2595 -1235 2645 -1205
rect 2675 -1235 2725 -1205
rect 2755 -1235 2805 -1205
rect 2835 -1235 2885 -1205
rect 2915 -1235 2965 -1205
rect 2995 -1235 3045 -1205
rect 3075 -1235 3125 -1205
rect 3155 -1235 3205 -1205
rect 3235 -1235 3285 -1205
rect 3315 -1235 3365 -1205
rect 3395 -1235 3445 -1205
rect 3475 -1235 3525 -1205
rect 3555 -1235 3605 -1205
rect 3635 -1235 3685 -1205
rect 3715 -1235 3765 -1205
rect 3795 -1235 3845 -1205
rect 3875 -1235 3925 -1205
rect 3955 -1235 4005 -1205
rect 4035 -1235 4085 -1205
rect 4115 -1235 4165 -1205
rect 4195 -1235 4245 -1205
rect 4275 -1235 4325 -1205
rect 4355 -1235 4405 -1205
rect 4435 -1235 4485 -1205
rect 4515 -1235 4565 -1205
rect 4595 -1235 4645 -1205
rect 4675 -1235 4725 -1205
rect 4755 -1235 4805 -1205
rect 4835 -1235 4885 -1205
rect 4915 -1235 4965 -1205
rect 4995 -1235 5045 -1205
rect 5075 -1235 5125 -1205
rect 5155 -1235 5205 -1205
rect 5235 -1235 5285 -1205
rect 5315 -1235 5365 -1205
rect 5395 -1235 5445 -1205
rect 5475 -1235 5525 -1205
rect 5555 -1235 5605 -1205
rect 5635 -1235 5685 -1205
rect 5715 -1235 5765 -1205
rect 5795 -1235 5845 -1205
rect 5875 -1235 5925 -1205
rect 5955 -1235 6005 -1205
rect 6035 -1235 6085 -1205
rect 6115 -1235 6165 -1205
rect 6195 -1235 6245 -1205
rect 6275 -1235 6325 -1205
rect 6355 -1235 6405 -1205
rect 6435 -1235 6485 -1205
rect 6515 -1235 6565 -1205
rect 6595 -1235 6645 -1205
rect 6675 -1235 6725 -1205
rect 6755 -1235 6805 -1205
rect 6835 -1235 6885 -1205
rect 6915 -1235 6965 -1205
rect 6995 -1235 7045 -1205
rect 7075 -1235 7125 -1205
rect 7155 -1235 7205 -1205
rect 7235 -1235 7285 -1205
rect 7315 -1235 7365 -1205
rect 7395 -1235 7445 -1205
rect 7475 -1235 7525 -1205
rect 7555 -1235 7605 -1205
rect 7635 -1235 7685 -1205
rect 7715 -1235 7765 -1205
rect 7795 -1235 7845 -1205
rect 7875 -1235 7925 -1205
rect 7955 -1235 8005 -1205
rect 8035 -1235 8085 -1205
rect 8115 -1235 8165 -1205
rect 8195 -1235 8245 -1205
rect 8275 -1235 8325 -1205
rect 8355 -1235 8405 -1205
rect 8435 -1235 8485 -1205
rect 8515 -1235 8565 -1205
rect 8595 -1235 8645 -1205
rect 8675 -1235 8725 -1205
rect 8755 -1235 8805 -1205
rect 8835 -1235 8885 -1205
rect 8915 -1235 8965 -1205
rect 8995 -1235 9045 -1205
rect 9075 -1235 9125 -1205
rect 9155 -1235 9205 -1205
rect 9235 -1235 9285 -1205
rect 9315 -1235 9365 -1205
rect 9395 -1235 9445 -1205
rect 9475 -1235 9525 -1205
rect 9555 -1235 9605 -1205
rect 9635 -1235 9685 -1205
rect 9715 -1235 9765 -1205
rect 9795 -1235 9845 -1205
rect 9875 -1235 9925 -1205
rect 9955 -1235 10005 -1205
rect 10035 -1235 10085 -1205
rect 10115 -1235 10165 -1205
rect 10195 -1235 10245 -1205
rect 10275 -1235 10325 -1205
rect 10355 -1235 10405 -1205
rect 10435 -1235 10485 -1205
rect 10515 -1235 10565 -1205
rect 10595 -1235 10645 -1205
rect 10675 -1235 10805 -1205
rect 10835 -1235 10965 -1205
rect 10995 -1235 11000 -1205
rect -720 -1240 11000 -1235
rect -720 -1285 11000 -1280
rect -720 -1315 -715 -1285
rect -685 -1315 -555 -1285
rect -525 -1315 -395 -1285
rect -365 -1315 -235 -1285
rect -205 -1315 -155 -1285
rect -125 -1315 -75 -1285
rect -45 -1315 5 -1285
rect 35 -1315 85 -1285
rect 115 -1315 165 -1285
rect 195 -1315 245 -1285
rect 275 -1315 325 -1285
rect 355 -1315 405 -1285
rect 435 -1315 485 -1285
rect 515 -1315 565 -1285
rect 595 -1315 645 -1285
rect 675 -1315 725 -1285
rect 755 -1315 805 -1285
rect 835 -1315 885 -1285
rect 915 -1315 965 -1285
rect 995 -1315 1045 -1285
rect 1075 -1315 1125 -1285
rect 1155 -1315 1205 -1285
rect 1235 -1315 1285 -1285
rect 1315 -1315 1365 -1285
rect 1395 -1315 1445 -1285
rect 1475 -1315 1525 -1285
rect 1555 -1315 1605 -1285
rect 1635 -1315 1685 -1285
rect 1715 -1315 1765 -1285
rect 1795 -1315 1845 -1285
rect 1875 -1315 1925 -1285
rect 1955 -1315 2005 -1285
rect 2035 -1315 2085 -1285
rect 2115 -1315 2165 -1285
rect 2195 -1315 2245 -1285
rect 2275 -1315 2325 -1285
rect 2355 -1315 2405 -1285
rect 2435 -1315 2485 -1285
rect 2515 -1315 2565 -1285
rect 2595 -1315 2645 -1285
rect 2675 -1315 2725 -1285
rect 2755 -1315 2805 -1285
rect 2835 -1315 2885 -1285
rect 2915 -1315 2965 -1285
rect 2995 -1315 3045 -1285
rect 3075 -1315 3125 -1285
rect 3155 -1315 3205 -1285
rect 3235 -1315 3285 -1285
rect 3315 -1315 3365 -1285
rect 3395 -1315 3445 -1285
rect 3475 -1315 3525 -1285
rect 3555 -1315 3605 -1285
rect 3635 -1315 3685 -1285
rect 3715 -1315 3765 -1285
rect 3795 -1315 3845 -1285
rect 3875 -1315 3925 -1285
rect 3955 -1315 4005 -1285
rect 4035 -1315 4085 -1285
rect 4115 -1315 4165 -1285
rect 4195 -1315 4245 -1285
rect 4275 -1315 4325 -1285
rect 4355 -1315 4405 -1285
rect 4435 -1315 4485 -1285
rect 4515 -1315 4565 -1285
rect 4595 -1315 4645 -1285
rect 4675 -1315 4725 -1285
rect 4755 -1315 4805 -1285
rect 4835 -1315 4885 -1285
rect 4915 -1315 4965 -1285
rect 4995 -1315 5045 -1285
rect 5075 -1315 5125 -1285
rect 5155 -1315 5205 -1285
rect 5235 -1315 5285 -1285
rect 5315 -1315 5365 -1285
rect 5395 -1315 5445 -1285
rect 5475 -1315 5525 -1285
rect 5555 -1315 5605 -1285
rect 5635 -1315 5685 -1285
rect 5715 -1315 5765 -1285
rect 5795 -1315 5845 -1285
rect 5875 -1315 5925 -1285
rect 5955 -1315 6005 -1285
rect 6035 -1315 6085 -1285
rect 6115 -1315 6165 -1285
rect 6195 -1315 6245 -1285
rect 6275 -1315 6325 -1285
rect 6355 -1315 6405 -1285
rect 6435 -1315 6485 -1285
rect 6515 -1315 6565 -1285
rect 6595 -1315 6645 -1285
rect 6675 -1315 6725 -1285
rect 6755 -1315 6805 -1285
rect 6835 -1315 6885 -1285
rect 6915 -1315 6965 -1285
rect 6995 -1315 7045 -1285
rect 7075 -1315 7125 -1285
rect 7155 -1315 7205 -1285
rect 7235 -1315 7285 -1285
rect 7315 -1315 7365 -1285
rect 7395 -1315 7445 -1285
rect 7475 -1315 7525 -1285
rect 7555 -1315 7605 -1285
rect 7635 -1315 7685 -1285
rect 7715 -1315 7765 -1285
rect 7795 -1315 7845 -1285
rect 7875 -1315 7925 -1285
rect 7955 -1315 8005 -1285
rect 8035 -1315 8085 -1285
rect 8115 -1315 8165 -1285
rect 8195 -1315 8245 -1285
rect 8275 -1315 8325 -1285
rect 8355 -1315 8405 -1285
rect 8435 -1315 8485 -1285
rect 8515 -1315 8565 -1285
rect 8595 -1315 8645 -1285
rect 8675 -1315 8725 -1285
rect 8755 -1315 8805 -1285
rect 8835 -1315 8885 -1285
rect 8915 -1315 8965 -1285
rect 8995 -1315 9045 -1285
rect 9075 -1315 9125 -1285
rect 9155 -1315 9205 -1285
rect 9235 -1315 9285 -1285
rect 9315 -1315 9365 -1285
rect 9395 -1315 9445 -1285
rect 9475 -1315 9525 -1285
rect 9555 -1315 9605 -1285
rect 9635 -1315 9685 -1285
rect 9715 -1315 9765 -1285
rect 9795 -1315 9845 -1285
rect 9875 -1315 9925 -1285
rect 9955 -1315 10005 -1285
rect 10035 -1315 10085 -1285
rect 10115 -1315 10165 -1285
rect 10195 -1315 10245 -1285
rect 10275 -1315 10325 -1285
rect 10355 -1315 10405 -1285
rect 10435 -1315 10485 -1285
rect 10515 -1315 10565 -1285
rect 10595 -1315 10645 -1285
rect 10675 -1315 10805 -1285
rect 10835 -1315 10965 -1285
rect 10995 -1315 11000 -1285
rect -720 -1320 11000 -1315
rect -720 -1365 11000 -1360
rect -720 -1395 -715 -1365
rect -685 -1395 -555 -1365
rect -525 -1395 -395 -1365
rect -365 -1395 -235 -1365
rect -205 -1395 -155 -1365
rect -125 -1395 -75 -1365
rect -45 -1395 5 -1365
rect 35 -1395 85 -1365
rect 115 -1395 165 -1365
rect 195 -1395 245 -1365
rect 275 -1395 325 -1365
rect 355 -1395 405 -1365
rect 435 -1395 485 -1365
rect 515 -1395 565 -1365
rect 595 -1395 645 -1365
rect 675 -1395 725 -1365
rect 755 -1395 805 -1365
rect 835 -1395 885 -1365
rect 915 -1395 965 -1365
rect 995 -1395 1045 -1365
rect 1075 -1395 1125 -1365
rect 1155 -1395 1205 -1365
rect 1235 -1395 1285 -1365
rect 1315 -1395 1365 -1365
rect 1395 -1395 1445 -1365
rect 1475 -1395 1525 -1365
rect 1555 -1395 1605 -1365
rect 1635 -1395 1685 -1365
rect 1715 -1395 1765 -1365
rect 1795 -1395 1845 -1365
rect 1875 -1395 1925 -1365
rect 1955 -1395 2005 -1365
rect 2035 -1395 2085 -1365
rect 2115 -1395 2165 -1365
rect 2195 -1395 2245 -1365
rect 2275 -1395 2325 -1365
rect 2355 -1395 2405 -1365
rect 2435 -1395 2485 -1365
rect 2515 -1395 2565 -1365
rect 2595 -1395 2645 -1365
rect 2675 -1395 2725 -1365
rect 2755 -1395 2805 -1365
rect 2835 -1395 2885 -1365
rect 2915 -1395 2965 -1365
rect 2995 -1395 3045 -1365
rect 3075 -1395 3125 -1365
rect 3155 -1395 3205 -1365
rect 3235 -1395 3285 -1365
rect 3315 -1395 3365 -1365
rect 3395 -1395 3445 -1365
rect 3475 -1395 3525 -1365
rect 3555 -1395 3605 -1365
rect 3635 -1395 3685 -1365
rect 3715 -1395 3765 -1365
rect 3795 -1395 3845 -1365
rect 3875 -1395 3925 -1365
rect 3955 -1395 4005 -1365
rect 4035 -1395 4085 -1365
rect 4115 -1395 4165 -1365
rect 4195 -1395 4245 -1365
rect 4275 -1395 4325 -1365
rect 4355 -1395 4405 -1365
rect 4435 -1395 4485 -1365
rect 4515 -1395 4565 -1365
rect 4595 -1395 4645 -1365
rect 4675 -1395 4725 -1365
rect 4755 -1395 4805 -1365
rect 4835 -1395 4885 -1365
rect 4915 -1395 4965 -1365
rect 4995 -1395 5045 -1365
rect 5075 -1395 5125 -1365
rect 5155 -1395 5205 -1365
rect 5235 -1395 5285 -1365
rect 5315 -1395 5365 -1365
rect 5395 -1395 5445 -1365
rect 5475 -1395 5525 -1365
rect 5555 -1395 5605 -1365
rect 5635 -1395 5685 -1365
rect 5715 -1395 5765 -1365
rect 5795 -1395 5845 -1365
rect 5875 -1395 5925 -1365
rect 5955 -1395 6005 -1365
rect 6035 -1395 6085 -1365
rect 6115 -1395 6165 -1365
rect 6195 -1395 6245 -1365
rect 6275 -1395 6325 -1365
rect 6355 -1395 6405 -1365
rect 6435 -1395 6485 -1365
rect 6515 -1395 6565 -1365
rect 6595 -1395 6645 -1365
rect 6675 -1395 6725 -1365
rect 6755 -1395 6805 -1365
rect 6835 -1395 6885 -1365
rect 6915 -1395 6965 -1365
rect 6995 -1395 7045 -1365
rect 7075 -1395 7125 -1365
rect 7155 -1395 7205 -1365
rect 7235 -1395 7285 -1365
rect 7315 -1395 7365 -1365
rect 7395 -1395 7445 -1365
rect 7475 -1395 7525 -1365
rect 7555 -1395 7605 -1365
rect 7635 -1395 7685 -1365
rect 7715 -1395 7765 -1365
rect 7795 -1395 7845 -1365
rect 7875 -1395 7925 -1365
rect 7955 -1395 8005 -1365
rect 8035 -1395 8085 -1365
rect 8115 -1395 8165 -1365
rect 8195 -1395 8245 -1365
rect 8275 -1395 8325 -1365
rect 8355 -1395 8405 -1365
rect 8435 -1395 8485 -1365
rect 8515 -1395 8565 -1365
rect 8595 -1395 8645 -1365
rect 8675 -1395 8725 -1365
rect 8755 -1395 8805 -1365
rect 8835 -1395 8885 -1365
rect 8915 -1395 8965 -1365
rect 8995 -1395 9045 -1365
rect 9075 -1395 9125 -1365
rect 9155 -1395 9205 -1365
rect 9235 -1395 9285 -1365
rect 9315 -1395 9365 -1365
rect 9395 -1395 9445 -1365
rect 9475 -1395 9525 -1365
rect 9555 -1395 9605 -1365
rect 9635 -1395 9685 -1365
rect 9715 -1395 9765 -1365
rect 9795 -1395 9845 -1365
rect 9875 -1395 9925 -1365
rect 9955 -1395 10005 -1365
rect 10035 -1395 10085 -1365
rect 10115 -1395 10165 -1365
rect 10195 -1395 10245 -1365
rect 10275 -1395 10325 -1365
rect 10355 -1395 10405 -1365
rect 10435 -1395 10485 -1365
rect 10515 -1395 10565 -1365
rect 10595 -1395 10645 -1365
rect 10675 -1395 10805 -1365
rect 10835 -1395 10965 -1365
rect 10995 -1395 11000 -1365
rect -720 -1400 11000 -1395
rect -720 -1445 11000 -1440
rect -720 -1475 -715 -1445
rect -685 -1475 -555 -1445
rect -525 -1475 -395 -1445
rect -365 -1475 -235 -1445
rect -205 -1475 -155 -1445
rect -125 -1475 -75 -1445
rect -45 -1475 5 -1445
rect 35 -1475 85 -1445
rect 115 -1475 165 -1445
rect 195 -1475 245 -1445
rect 275 -1475 325 -1445
rect 355 -1475 405 -1445
rect 435 -1475 485 -1445
rect 515 -1475 565 -1445
rect 595 -1475 645 -1445
rect 675 -1475 725 -1445
rect 755 -1475 805 -1445
rect 835 -1475 885 -1445
rect 915 -1475 965 -1445
rect 995 -1475 1045 -1445
rect 1075 -1475 1125 -1445
rect 1155 -1475 1205 -1445
rect 1235 -1475 1285 -1445
rect 1315 -1475 1365 -1445
rect 1395 -1475 1445 -1445
rect 1475 -1475 1525 -1445
rect 1555 -1475 1605 -1445
rect 1635 -1475 1685 -1445
rect 1715 -1475 1765 -1445
rect 1795 -1475 1845 -1445
rect 1875 -1475 1925 -1445
rect 1955 -1475 2005 -1445
rect 2035 -1475 2085 -1445
rect 2115 -1475 2165 -1445
rect 2195 -1475 2245 -1445
rect 2275 -1475 2325 -1445
rect 2355 -1475 2405 -1445
rect 2435 -1475 2485 -1445
rect 2515 -1475 2565 -1445
rect 2595 -1475 2645 -1445
rect 2675 -1475 2725 -1445
rect 2755 -1475 2805 -1445
rect 2835 -1475 2885 -1445
rect 2915 -1475 2965 -1445
rect 2995 -1475 3045 -1445
rect 3075 -1475 3125 -1445
rect 3155 -1475 3205 -1445
rect 3235 -1475 3285 -1445
rect 3315 -1475 3365 -1445
rect 3395 -1475 3445 -1445
rect 3475 -1475 3525 -1445
rect 3555 -1475 3605 -1445
rect 3635 -1475 3685 -1445
rect 3715 -1475 3765 -1445
rect 3795 -1475 3845 -1445
rect 3875 -1475 3925 -1445
rect 3955 -1475 4005 -1445
rect 4035 -1475 4085 -1445
rect 4115 -1475 4165 -1445
rect 4195 -1475 4245 -1445
rect 4275 -1475 4325 -1445
rect 4355 -1475 4405 -1445
rect 4435 -1475 4485 -1445
rect 4515 -1475 4565 -1445
rect 4595 -1475 4645 -1445
rect 4675 -1475 4725 -1445
rect 4755 -1475 4805 -1445
rect 4835 -1475 4885 -1445
rect 4915 -1475 4965 -1445
rect 4995 -1475 5045 -1445
rect 5075 -1475 5125 -1445
rect 5155 -1475 5205 -1445
rect 5235 -1475 5285 -1445
rect 5315 -1475 5365 -1445
rect 5395 -1475 5445 -1445
rect 5475 -1475 5525 -1445
rect 5555 -1475 5605 -1445
rect 5635 -1475 5685 -1445
rect 5715 -1475 5765 -1445
rect 5795 -1475 5845 -1445
rect 5875 -1475 5925 -1445
rect 5955 -1475 6005 -1445
rect 6035 -1475 6085 -1445
rect 6115 -1475 6165 -1445
rect 6195 -1475 6245 -1445
rect 6275 -1475 6325 -1445
rect 6355 -1475 6405 -1445
rect 6435 -1475 6485 -1445
rect 6515 -1475 6565 -1445
rect 6595 -1475 6645 -1445
rect 6675 -1475 6725 -1445
rect 6755 -1475 6805 -1445
rect 6835 -1475 6885 -1445
rect 6915 -1475 6965 -1445
rect 6995 -1475 7045 -1445
rect 7075 -1475 7125 -1445
rect 7155 -1475 7205 -1445
rect 7235 -1475 7285 -1445
rect 7315 -1475 7365 -1445
rect 7395 -1475 7445 -1445
rect 7475 -1475 7525 -1445
rect 7555 -1475 7605 -1445
rect 7635 -1475 7685 -1445
rect 7715 -1475 7765 -1445
rect 7795 -1475 7845 -1445
rect 7875 -1475 7925 -1445
rect 7955 -1475 8005 -1445
rect 8035 -1475 8085 -1445
rect 8115 -1475 8165 -1445
rect 8195 -1475 8245 -1445
rect 8275 -1475 8325 -1445
rect 8355 -1475 8405 -1445
rect 8435 -1475 8485 -1445
rect 8515 -1475 8565 -1445
rect 8595 -1475 8645 -1445
rect 8675 -1475 8725 -1445
rect 8755 -1475 8805 -1445
rect 8835 -1475 8885 -1445
rect 8915 -1475 8965 -1445
rect 8995 -1475 9045 -1445
rect 9075 -1475 9125 -1445
rect 9155 -1475 9205 -1445
rect 9235 -1475 9285 -1445
rect 9315 -1475 9365 -1445
rect 9395 -1475 9445 -1445
rect 9475 -1475 9525 -1445
rect 9555 -1475 9605 -1445
rect 9635 -1475 9685 -1445
rect 9715 -1475 9765 -1445
rect 9795 -1475 9845 -1445
rect 9875 -1475 9925 -1445
rect 9955 -1475 10005 -1445
rect 10035 -1475 10085 -1445
rect 10115 -1475 10165 -1445
rect 10195 -1475 10245 -1445
rect 10275 -1475 10325 -1445
rect 10355 -1475 10405 -1445
rect 10435 -1475 10485 -1445
rect 10515 -1475 10565 -1445
rect 10595 -1475 10645 -1445
rect 10675 -1475 10805 -1445
rect 10835 -1475 10965 -1445
rect 10995 -1475 11000 -1445
rect -720 -1480 11000 -1475
rect -720 -1525 11000 -1520
rect -720 -1555 -715 -1525
rect -685 -1555 -555 -1525
rect -525 -1555 -395 -1525
rect -365 -1555 -235 -1525
rect -205 -1555 -155 -1525
rect -125 -1555 -75 -1525
rect -45 -1555 5 -1525
rect 35 -1555 85 -1525
rect 115 -1555 165 -1525
rect 195 -1555 245 -1525
rect 275 -1555 325 -1525
rect 355 -1555 405 -1525
rect 435 -1555 485 -1525
rect 515 -1555 565 -1525
rect 595 -1555 645 -1525
rect 675 -1555 725 -1525
rect 755 -1555 805 -1525
rect 835 -1555 885 -1525
rect 915 -1555 965 -1525
rect 995 -1555 1045 -1525
rect 1075 -1555 1125 -1525
rect 1155 -1555 1205 -1525
rect 1235 -1555 1285 -1525
rect 1315 -1555 1365 -1525
rect 1395 -1555 1445 -1525
rect 1475 -1555 1525 -1525
rect 1555 -1555 1605 -1525
rect 1635 -1555 1685 -1525
rect 1715 -1555 1765 -1525
rect 1795 -1555 1845 -1525
rect 1875 -1555 1925 -1525
rect 1955 -1555 2005 -1525
rect 2035 -1555 2085 -1525
rect 2115 -1555 2165 -1525
rect 2195 -1555 2245 -1525
rect 2275 -1555 2325 -1525
rect 2355 -1555 2405 -1525
rect 2435 -1555 2485 -1525
rect 2515 -1555 2565 -1525
rect 2595 -1555 2645 -1525
rect 2675 -1555 2725 -1525
rect 2755 -1555 2805 -1525
rect 2835 -1555 2885 -1525
rect 2915 -1555 2965 -1525
rect 2995 -1555 3045 -1525
rect 3075 -1555 3125 -1525
rect 3155 -1555 3205 -1525
rect 3235 -1555 3285 -1525
rect 3315 -1555 3365 -1525
rect 3395 -1555 3445 -1525
rect 3475 -1555 3525 -1525
rect 3555 -1555 3605 -1525
rect 3635 -1555 3685 -1525
rect 3715 -1555 3765 -1525
rect 3795 -1555 3845 -1525
rect 3875 -1555 3925 -1525
rect 3955 -1555 4005 -1525
rect 4035 -1555 4085 -1525
rect 4115 -1555 4165 -1525
rect 4195 -1555 4245 -1525
rect 4275 -1555 4325 -1525
rect 4355 -1555 4405 -1525
rect 4435 -1555 4485 -1525
rect 4515 -1555 4565 -1525
rect 4595 -1555 4645 -1525
rect 4675 -1555 4725 -1525
rect 4755 -1555 4805 -1525
rect 4835 -1555 4885 -1525
rect 4915 -1555 4965 -1525
rect 4995 -1555 5045 -1525
rect 5075 -1555 5125 -1525
rect 5155 -1555 5205 -1525
rect 5235 -1555 5285 -1525
rect 5315 -1555 5365 -1525
rect 5395 -1555 5445 -1525
rect 5475 -1555 5525 -1525
rect 5555 -1555 5605 -1525
rect 5635 -1555 5685 -1525
rect 5715 -1555 5765 -1525
rect 5795 -1555 5845 -1525
rect 5875 -1555 5925 -1525
rect 5955 -1555 6005 -1525
rect 6035 -1555 6085 -1525
rect 6115 -1555 6165 -1525
rect 6195 -1555 6245 -1525
rect 6275 -1555 6325 -1525
rect 6355 -1555 6405 -1525
rect 6435 -1555 6485 -1525
rect 6515 -1555 6565 -1525
rect 6595 -1555 6645 -1525
rect 6675 -1555 6725 -1525
rect 6755 -1555 6805 -1525
rect 6835 -1555 6885 -1525
rect 6915 -1555 6965 -1525
rect 6995 -1555 7045 -1525
rect 7075 -1555 7125 -1525
rect 7155 -1555 7205 -1525
rect 7235 -1555 7285 -1525
rect 7315 -1555 7365 -1525
rect 7395 -1555 7445 -1525
rect 7475 -1555 7525 -1525
rect 7555 -1555 7605 -1525
rect 7635 -1555 7685 -1525
rect 7715 -1555 7765 -1525
rect 7795 -1555 7845 -1525
rect 7875 -1555 7925 -1525
rect 7955 -1555 8005 -1525
rect 8035 -1555 8085 -1525
rect 8115 -1555 8165 -1525
rect 8195 -1555 8245 -1525
rect 8275 -1555 8325 -1525
rect 8355 -1555 8405 -1525
rect 8435 -1555 8485 -1525
rect 8515 -1555 8565 -1525
rect 8595 -1555 8645 -1525
rect 8675 -1555 8725 -1525
rect 8755 -1555 8805 -1525
rect 8835 -1555 8885 -1525
rect 8915 -1555 8965 -1525
rect 8995 -1555 9045 -1525
rect 9075 -1555 9125 -1525
rect 9155 -1555 9205 -1525
rect 9235 -1555 9285 -1525
rect 9315 -1555 9365 -1525
rect 9395 -1555 9445 -1525
rect 9475 -1555 9525 -1525
rect 9555 -1555 9605 -1525
rect 9635 -1555 9685 -1525
rect 9715 -1555 9765 -1525
rect 9795 -1555 9845 -1525
rect 9875 -1555 9925 -1525
rect 9955 -1555 10005 -1525
rect 10035 -1555 10085 -1525
rect 10115 -1555 10165 -1525
rect 10195 -1555 10245 -1525
rect 10275 -1555 10325 -1525
rect 10355 -1555 10405 -1525
rect 10435 -1555 10485 -1525
rect 10515 -1555 10565 -1525
rect 10595 -1555 10645 -1525
rect 10675 -1555 10805 -1525
rect 10835 -1555 10965 -1525
rect 10995 -1555 11000 -1525
rect -720 -1560 11000 -1555
rect -640 -1605 10600 -1600
rect -640 -1635 -635 -1605
rect -605 -1635 -75 -1605
rect -45 -1635 565 -1605
rect 595 -1635 1205 -1605
rect 1235 -1635 1845 -1605
rect 1875 -1635 2485 -1605
rect 2515 -1635 3125 -1605
rect 3155 -1635 3765 -1605
rect 3795 -1635 4405 -1605
rect 4435 -1635 5045 -1605
rect 5075 -1635 10325 -1605
rect 10355 -1635 10600 -1605
rect -640 -1640 10600 -1635
rect 10640 -1605 11000 -1600
rect 10640 -1635 10645 -1605
rect 10675 -1635 10805 -1605
rect 10835 -1635 10965 -1605
rect 10995 -1635 11000 -1605
rect 10640 -1640 11000 -1635
rect -640 -1685 10600 -1680
rect -640 -1715 -635 -1685
rect -605 -1715 -75 -1685
rect -45 -1715 565 -1685
rect 595 -1715 1205 -1685
rect 1235 -1715 1845 -1685
rect 1875 -1715 2485 -1685
rect 2515 -1715 3125 -1685
rect 3155 -1715 3765 -1685
rect 3795 -1715 4405 -1685
rect 4435 -1715 5045 -1685
rect 5075 -1715 10325 -1685
rect 10355 -1715 10600 -1685
rect -640 -1720 10600 -1715
rect 10640 -1685 11000 -1680
rect 10640 -1715 10645 -1685
rect 10675 -1715 10805 -1685
rect 10835 -1715 10965 -1685
rect 10995 -1715 11000 -1685
rect 10640 -1720 11000 -1715
rect -720 -1765 11000 -1760
rect -720 -1795 -715 -1765
rect -685 -1795 -555 -1765
rect -525 -1795 -395 -1765
rect -365 -1795 -235 -1765
rect -205 -1795 -155 -1765
rect -125 -1795 -75 -1765
rect -45 -1795 5 -1765
rect 35 -1795 85 -1765
rect 115 -1795 165 -1765
rect 195 -1795 245 -1765
rect 275 -1795 325 -1765
rect 355 -1795 405 -1765
rect 435 -1795 485 -1765
rect 515 -1795 565 -1765
rect 595 -1795 645 -1765
rect 675 -1795 725 -1765
rect 755 -1795 805 -1765
rect 835 -1795 885 -1765
rect 915 -1795 965 -1765
rect 995 -1795 1045 -1765
rect 1075 -1795 1125 -1765
rect 1155 -1795 1205 -1765
rect 1235 -1795 1285 -1765
rect 1315 -1795 1365 -1765
rect 1395 -1795 1445 -1765
rect 1475 -1795 1525 -1765
rect 1555 -1795 1605 -1765
rect 1635 -1795 1685 -1765
rect 1715 -1795 1765 -1765
rect 1795 -1795 1845 -1765
rect 1875 -1795 1925 -1765
rect 1955 -1795 2005 -1765
rect 2035 -1795 2085 -1765
rect 2115 -1795 2165 -1765
rect 2195 -1795 2245 -1765
rect 2275 -1795 2325 -1765
rect 2355 -1795 2405 -1765
rect 2435 -1795 2485 -1765
rect 2515 -1795 2565 -1765
rect 2595 -1795 2645 -1765
rect 2675 -1795 2725 -1765
rect 2755 -1795 2805 -1765
rect 2835 -1795 2885 -1765
rect 2915 -1795 2965 -1765
rect 2995 -1795 3045 -1765
rect 3075 -1795 3125 -1765
rect 3155 -1795 3205 -1765
rect 3235 -1795 3285 -1765
rect 3315 -1795 3365 -1765
rect 3395 -1795 3445 -1765
rect 3475 -1795 3525 -1765
rect 3555 -1795 3605 -1765
rect 3635 -1795 3685 -1765
rect 3715 -1795 3765 -1765
rect 3795 -1795 3845 -1765
rect 3875 -1795 3925 -1765
rect 3955 -1795 4005 -1765
rect 4035 -1795 4085 -1765
rect 4115 -1795 4165 -1765
rect 4195 -1795 4245 -1765
rect 4275 -1795 4325 -1765
rect 4355 -1795 4405 -1765
rect 4435 -1795 4485 -1765
rect 4515 -1795 4565 -1765
rect 4595 -1795 4645 -1765
rect 4675 -1795 4725 -1765
rect 4755 -1795 4805 -1765
rect 4835 -1795 4885 -1765
rect 4915 -1795 4965 -1765
rect 4995 -1795 5045 -1765
rect 5075 -1795 5125 -1765
rect 5155 -1795 5205 -1765
rect 5235 -1795 5285 -1765
rect 5315 -1795 5365 -1765
rect 5395 -1795 5445 -1765
rect 5475 -1795 5525 -1765
rect 5555 -1795 5605 -1765
rect 5635 -1795 5685 -1765
rect 5715 -1795 5765 -1765
rect 5795 -1795 5845 -1765
rect 5875 -1795 5925 -1765
rect 5955 -1795 6005 -1765
rect 6035 -1795 6085 -1765
rect 6115 -1795 6165 -1765
rect 6195 -1795 6245 -1765
rect 6275 -1795 6325 -1765
rect 6355 -1795 6405 -1765
rect 6435 -1795 6485 -1765
rect 6515 -1795 6565 -1765
rect 6595 -1795 6645 -1765
rect 6675 -1795 6725 -1765
rect 6755 -1795 6805 -1765
rect 6835 -1795 6885 -1765
rect 6915 -1795 6965 -1765
rect 6995 -1795 7045 -1765
rect 7075 -1795 7125 -1765
rect 7155 -1795 7205 -1765
rect 7235 -1795 7285 -1765
rect 7315 -1795 7365 -1765
rect 7395 -1795 7445 -1765
rect 7475 -1795 7525 -1765
rect 7555 -1795 7605 -1765
rect 7635 -1795 7685 -1765
rect 7715 -1795 7765 -1765
rect 7795 -1795 7845 -1765
rect 7875 -1795 7925 -1765
rect 7955 -1795 8005 -1765
rect 8035 -1795 8085 -1765
rect 8115 -1795 8165 -1765
rect 8195 -1795 8245 -1765
rect 8275 -1795 8325 -1765
rect 8355 -1795 8405 -1765
rect 8435 -1795 8485 -1765
rect 8515 -1795 8565 -1765
rect 8595 -1795 8645 -1765
rect 8675 -1795 8725 -1765
rect 8755 -1795 8805 -1765
rect 8835 -1795 8885 -1765
rect 8915 -1795 8965 -1765
rect 8995 -1795 9045 -1765
rect 9075 -1795 9125 -1765
rect 9155 -1795 9205 -1765
rect 9235 -1795 9285 -1765
rect 9315 -1795 9365 -1765
rect 9395 -1795 9445 -1765
rect 9475 -1795 9525 -1765
rect 9555 -1795 9605 -1765
rect 9635 -1795 9685 -1765
rect 9715 -1795 9765 -1765
rect 9795 -1795 9845 -1765
rect 9875 -1795 9925 -1765
rect 9955 -1795 10005 -1765
rect 10035 -1795 10085 -1765
rect 10115 -1795 10165 -1765
rect 10195 -1795 10245 -1765
rect 10275 -1795 10325 -1765
rect 10355 -1795 10405 -1765
rect 10435 -1795 10485 -1765
rect 10515 -1795 10565 -1765
rect 10595 -1795 10645 -1765
rect 10675 -1795 10805 -1765
rect 10835 -1795 10965 -1765
rect 10995 -1795 11000 -1765
rect -720 -1800 11000 -1795
rect -720 -1845 11000 -1840
rect -720 -1875 -715 -1845
rect -685 -1875 -555 -1845
rect -525 -1875 -395 -1845
rect -365 -1875 -235 -1845
rect -205 -1875 -155 -1845
rect -125 -1875 -75 -1845
rect -45 -1875 5 -1845
rect 35 -1875 85 -1845
rect 115 -1875 165 -1845
rect 195 -1875 245 -1845
rect 275 -1875 325 -1845
rect 355 -1875 405 -1845
rect 435 -1875 485 -1845
rect 515 -1875 565 -1845
rect 595 -1875 645 -1845
rect 675 -1875 725 -1845
rect 755 -1875 805 -1845
rect 835 -1875 885 -1845
rect 915 -1875 965 -1845
rect 995 -1875 1045 -1845
rect 1075 -1875 1125 -1845
rect 1155 -1875 1205 -1845
rect 1235 -1875 1285 -1845
rect 1315 -1875 1365 -1845
rect 1395 -1875 1445 -1845
rect 1475 -1875 1525 -1845
rect 1555 -1875 1605 -1845
rect 1635 -1875 1685 -1845
rect 1715 -1875 1765 -1845
rect 1795 -1875 1845 -1845
rect 1875 -1875 1925 -1845
rect 1955 -1875 2005 -1845
rect 2035 -1875 2085 -1845
rect 2115 -1875 2165 -1845
rect 2195 -1875 2245 -1845
rect 2275 -1875 2325 -1845
rect 2355 -1875 2405 -1845
rect 2435 -1875 2485 -1845
rect 2515 -1875 2565 -1845
rect 2595 -1875 2645 -1845
rect 2675 -1875 2725 -1845
rect 2755 -1875 2805 -1845
rect 2835 -1875 2885 -1845
rect 2915 -1875 2965 -1845
rect 2995 -1875 3045 -1845
rect 3075 -1875 3125 -1845
rect 3155 -1875 3205 -1845
rect 3235 -1875 3285 -1845
rect 3315 -1875 3365 -1845
rect 3395 -1875 3445 -1845
rect 3475 -1875 3525 -1845
rect 3555 -1875 3605 -1845
rect 3635 -1875 3685 -1845
rect 3715 -1875 3765 -1845
rect 3795 -1875 3845 -1845
rect 3875 -1875 3925 -1845
rect 3955 -1875 4005 -1845
rect 4035 -1875 4085 -1845
rect 4115 -1875 4165 -1845
rect 4195 -1875 4245 -1845
rect 4275 -1875 4325 -1845
rect 4355 -1875 4405 -1845
rect 4435 -1875 4485 -1845
rect 4515 -1875 4565 -1845
rect 4595 -1875 4645 -1845
rect 4675 -1875 4725 -1845
rect 4755 -1875 4805 -1845
rect 4835 -1875 4885 -1845
rect 4915 -1875 4965 -1845
rect 4995 -1875 5045 -1845
rect 5075 -1875 5125 -1845
rect 5155 -1875 5205 -1845
rect 5235 -1875 5285 -1845
rect 5315 -1875 5365 -1845
rect 5395 -1875 5445 -1845
rect 5475 -1875 5525 -1845
rect 5555 -1875 5605 -1845
rect 5635 -1875 5685 -1845
rect 5715 -1875 5765 -1845
rect 5795 -1875 5845 -1845
rect 5875 -1875 5925 -1845
rect 5955 -1875 6005 -1845
rect 6035 -1875 6085 -1845
rect 6115 -1875 6165 -1845
rect 6195 -1875 6245 -1845
rect 6275 -1875 6325 -1845
rect 6355 -1875 6405 -1845
rect 6435 -1875 6485 -1845
rect 6515 -1875 6565 -1845
rect 6595 -1875 6645 -1845
rect 6675 -1875 6725 -1845
rect 6755 -1875 6805 -1845
rect 6835 -1875 6885 -1845
rect 6915 -1875 6965 -1845
rect 6995 -1875 7045 -1845
rect 7075 -1875 7125 -1845
rect 7155 -1875 7205 -1845
rect 7235 -1875 7285 -1845
rect 7315 -1875 7365 -1845
rect 7395 -1875 7445 -1845
rect 7475 -1875 7525 -1845
rect 7555 -1875 7605 -1845
rect 7635 -1875 7685 -1845
rect 7715 -1875 7765 -1845
rect 7795 -1875 7845 -1845
rect 7875 -1875 7925 -1845
rect 7955 -1875 8005 -1845
rect 8035 -1875 8085 -1845
rect 8115 -1875 8165 -1845
rect 8195 -1875 8245 -1845
rect 8275 -1875 8325 -1845
rect 8355 -1875 8405 -1845
rect 8435 -1875 8485 -1845
rect 8515 -1875 8565 -1845
rect 8595 -1875 8645 -1845
rect 8675 -1875 8725 -1845
rect 8755 -1875 8805 -1845
rect 8835 -1875 8885 -1845
rect 8915 -1875 8965 -1845
rect 8995 -1875 9045 -1845
rect 9075 -1875 9125 -1845
rect 9155 -1875 9205 -1845
rect 9235 -1875 9285 -1845
rect 9315 -1875 9365 -1845
rect 9395 -1875 9445 -1845
rect 9475 -1875 9525 -1845
rect 9555 -1875 9605 -1845
rect 9635 -1875 9685 -1845
rect 9715 -1875 9765 -1845
rect 9795 -1875 9845 -1845
rect 9875 -1875 9925 -1845
rect 9955 -1875 10005 -1845
rect 10035 -1875 10085 -1845
rect 10115 -1875 10165 -1845
rect 10195 -1875 10245 -1845
rect 10275 -1875 10325 -1845
rect 10355 -1875 10405 -1845
rect 10435 -1875 10485 -1845
rect 10515 -1875 10565 -1845
rect 10595 -1875 10645 -1845
rect 10675 -1875 10805 -1845
rect 10835 -1875 10965 -1845
rect 10995 -1875 11000 -1845
rect -720 -1880 11000 -1875
rect -720 -1925 -520 -1920
rect -720 -1955 -715 -1925
rect -685 -1955 -555 -1925
rect -525 -1955 -520 -1925
rect -720 -1960 -520 -1955
rect -480 -1925 10600 -1920
rect -480 -1955 -475 -1925
rect -445 -1955 5365 -1925
rect 5395 -1955 5685 -1925
rect 5715 -1955 6005 -1925
rect 6035 -1955 6325 -1925
rect 6355 -1955 6645 -1925
rect 6675 -1955 6965 -1925
rect 6995 -1955 7285 -1925
rect 7315 -1955 7605 -1925
rect 7635 -1955 7925 -1925
rect 7955 -1955 8245 -1925
rect 8275 -1955 8565 -1925
rect 8595 -1955 8885 -1925
rect 8915 -1955 9205 -1925
rect 9235 -1955 9525 -1925
rect 9555 -1955 9845 -1925
rect 9875 -1955 10165 -1925
rect 10195 -1955 10600 -1925
rect -480 -1960 10600 -1955
rect 10640 -1925 11000 -1920
rect 10640 -1955 10645 -1925
rect 10675 -1955 10805 -1925
rect 10835 -1955 10965 -1925
rect 10995 -1955 11000 -1925
rect 10640 -1960 11000 -1955
rect -720 -2005 11000 -2000
rect -720 -2035 -715 -2005
rect -685 -2035 -555 -2005
rect -525 -2035 -395 -2005
rect -365 -2035 -235 -2005
rect -205 -2035 -155 -2005
rect -125 -2035 -75 -2005
rect -45 -2035 5 -2005
rect 35 -2035 85 -2005
rect 115 -2035 165 -2005
rect 195 -2035 245 -2005
rect 275 -2035 325 -2005
rect 355 -2035 405 -2005
rect 435 -2035 485 -2005
rect 515 -2035 565 -2005
rect 595 -2035 645 -2005
rect 675 -2035 725 -2005
rect 755 -2035 805 -2005
rect 835 -2035 885 -2005
rect 915 -2035 965 -2005
rect 995 -2035 1045 -2005
rect 1075 -2035 1125 -2005
rect 1155 -2035 1205 -2005
rect 1235 -2035 1285 -2005
rect 1315 -2035 1365 -2005
rect 1395 -2035 1445 -2005
rect 1475 -2035 1525 -2005
rect 1555 -2035 1605 -2005
rect 1635 -2035 1685 -2005
rect 1715 -2035 1765 -2005
rect 1795 -2035 1845 -2005
rect 1875 -2035 1925 -2005
rect 1955 -2035 2005 -2005
rect 2035 -2035 2085 -2005
rect 2115 -2035 2165 -2005
rect 2195 -2035 2245 -2005
rect 2275 -2035 2325 -2005
rect 2355 -2035 2405 -2005
rect 2435 -2035 2485 -2005
rect 2515 -2035 2565 -2005
rect 2595 -2035 2645 -2005
rect 2675 -2035 2725 -2005
rect 2755 -2035 2805 -2005
rect 2835 -2035 2885 -2005
rect 2915 -2035 2965 -2005
rect 2995 -2035 3045 -2005
rect 3075 -2035 3125 -2005
rect 3155 -2035 3205 -2005
rect 3235 -2035 3285 -2005
rect 3315 -2035 3365 -2005
rect 3395 -2035 3445 -2005
rect 3475 -2035 3525 -2005
rect 3555 -2035 3605 -2005
rect 3635 -2035 3685 -2005
rect 3715 -2035 3765 -2005
rect 3795 -2035 3845 -2005
rect 3875 -2035 3925 -2005
rect 3955 -2035 4005 -2005
rect 4035 -2035 4085 -2005
rect 4115 -2035 4165 -2005
rect 4195 -2035 4245 -2005
rect 4275 -2035 4325 -2005
rect 4355 -2035 4405 -2005
rect 4435 -2035 4485 -2005
rect 4515 -2035 4565 -2005
rect 4595 -2035 4645 -2005
rect 4675 -2035 4725 -2005
rect 4755 -2035 4805 -2005
rect 4835 -2035 4885 -2005
rect 4915 -2035 4965 -2005
rect 4995 -2035 5045 -2005
rect 5075 -2035 5125 -2005
rect 5155 -2035 5205 -2005
rect 5235 -2035 5285 -2005
rect 5315 -2035 5365 -2005
rect 5395 -2035 5445 -2005
rect 5475 -2035 5525 -2005
rect 5555 -2035 5605 -2005
rect 5635 -2035 5685 -2005
rect 5715 -2035 5765 -2005
rect 5795 -2035 5845 -2005
rect 5875 -2035 5925 -2005
rect 5955 -2035 6005 -2005
rect 6035 -2035 6085 -2005
rect 6115 -2035 6165 -2005
rect 6195 -2035 6245 -2005
rect 6275 -2035 6325 -2005
rect 6355 -2035 6405 -2005
rect 6435 -2035 6485 -2005
rect 6515 -2035 6565 -2005
rect 6595 -2035 6645 -2005
rect 6675 -2035 6725 -2005
rect 6755 -2035 6805 -2005
rect 6835 -2035 6885 -2005
rect 6915 -2035 6965 -2005
rect 6995 -2035 7045 -2005
rect 7075 -2035 7125 -2005
rect 7155 -2035 7205 -2005
rect 7235 -2035 7285 -2005
rect 7315 -2035 7365 -2005
rect 7395 -2035 7445 -2005
rect 7475 -2035 7525 -2005
rect 7555 -2035 7605 -2005
rect 7635 -2035 7685 -2005
rect 7715 -2035 7765 -2005
rect 7795 -2035 7845 -2005
rect 7875 -2035 7925 -2005
rect 7955 -2035 8005 -2005
rect 8035 -2035 8085 -2005
rect 8115 -2035 8165 -2005
rect 8195 -2035 8245 -2005
rect 8275 -2035 8325 -2005
rect 8355 -2035 8405 -2005
rect 8435 -2035 8485 -2005
rect 8515 -2035 8565 -2005
rect 8595 -2035 8645 -2005
rect 8675 -2035 8725 -2005
rect 8755 -2035 8805 -2005
rect 8835 -2035 8885 -2005
rect 8915 -2035 8965 -2005
rect 8995 -2035 9045 -2005
rect 9075 -2035 9125 -2005
rect 9155 -2035 9205 -2005
rect 9235 -2035 9285 -2005
rect 9315 -2035 9365 -2005
rect 9395 -2035 9445 -2005
rect 9475 -2035 9525 -2005
rect 9555 -2035 9605 -2005
rect 9635 -2035 9685 -2005
rect 9715 -2035 9765 -2005
rect 9795 -2035 9845 -2005
rect 9875 -2035 9925 -2005
rect 9955 -2035 10005 -2005
rect 10035 -2035 10085 -2005
rect 10115 -2035 10165 -2005
rect 10195 -2035 10245 -2005
rect 10275 -2035 10325 -2005
rect 10355 -2035 10405 -2005
rect 10435 -2035 10485 -2005
rect 10515 -2035 10565 -2005
rect 10595 -2035 10645 -2005
rect 10675 -2035 10805 -2005
rect 10835 -2035 10965 -2005
rect 10995 -2035 11000 -2005
rect -720 -2040 11000 -2035
rect -720 -2085 -360 -2080
rect -720 -2115 -715 -2085
rect -685 -2115 -555 -2085
rect -525 -2115 -395 -2085
rect -365 -2115 -360 -2085
rect -720 -2120 -360 -2115
rect -320 -2085 10920 -2080
rect -320 -2115 85 -2085
rect 115 -2115 245 -2085
rect 275 -2115 405 -2085
rect 435 -2115 725 -2085
rect 755 -2115 885 -2085
rect 915 -2115 1045 -2085
rect 1075 -2115 1205 -2085
rect 1235 -2115 1365 -2085
rect 1395 -2115 1525 -2085
rect 1555 -2115 1685 -2085
rect 1715 -2115 2005 -2085
rect 2035 -2115 2165 -2085
rect 2195 -2115 2325 -2085
rect 2355 -2115 2645 -2085
rect 2675 -2115 2805 -2085
rect 2835 -2115 2965 -2085
rect 2995 -2115 3285 -2085
rect 3315 -2115 3445 -2085
rect 3475 -2115 3605 -2085
rect 3635 -2115 3765 -2085
rect 3795 -2115 3925 -2085
rect 3955 -2115 4085 -2085
rect 4115 -2115 4245 -2085
rect 4275 -2115 4565 -2085
rect 4595 -2115 4725 -2085
rect 4755 -2115 4885 -2085
rect 4915 -2115 10885 -2085
rect 10915 -2115 10920 -2085
rect -320 -2120 10920 -2115
rect 10960 -2120 11000 -2080
rect -720 -2165 11000 -2160
rect -720 -2195 -715 -2165
rect -685 -2195 -555 -2165
rect -525 -2195 -395 -2165
rect -365 -2195 -235 -2165
rect -205 -2195 -155 -2165
rect -125 -2195 -75 -2165
rect -45 -2195 5 -2165
rect 35 -2195 85 -2165
rect 115 -2195 165 -2165
rect 195 -2195 245 -2165
rect 275 -2195 325 -2165
rect 355 -2195 405 -2165
rect 435 -2195 485 -2165
rect 515 -2195 565 -2165
rect 595 -2195 645 -2165
rect 675 -2195 725 -2165
rect 755 -2195 805 -2165
rect 835 -2195 885 -2165
rect 915 -2195 965 -2165
rect 995 -2195 1045 -2165
rect 1075 -2195 1125 -2165
rect 1155 -2195 1205 -2165
rect 1235 -2195 1285 -2165
rect 1315 -2195 1365 -2165
rect 1395 -2195 1445 -2165
rect 1475 -2195 1525 -2165
rect 1555 -2195 1605 -2165
rect 1635 -2195 1685 -2165
rect 1715 -2195 1765 -2165
rect 1795 -2195 1845 -2165
rect 1875 -2195 1925 -2165
rect 1955 -2195 2005 -2165
rect 2035 -2195 2085 -2165
rect 2115 -2195 2165 -2165
rect 2195 -2195 2245 -2165
rect 2275 -2195 2325 -2165
rect 2355 -2195 2405 -2165
rect 2435 -2195 2485 -2165
rect 2515 -2195 2565 -2165
rect 2595 -2195 2645 -2165
rect 2675 -2195 2725 -2165
rect 2755 -2195 2805 -2165
rect 2835 -2195 2885 -2165
rect 2915 -2195 2965 -2165
rect 2995 -2195 3045 -2165
rect 3075 -2195 3125 -2165
rect 3155 -2195 3205 -2165
rect 3235 -2195 3285 -2165
rect 3315 -2195 3365 -2165
rect 3395 -2195 3445 -2165
rect 3475 -2195 3525 -2165
rect 3555 -2195 3605 -2165
rect 3635 -2195 3685 -2165
rect 3715 -2195 3765 -2165
rect 3795 -2195 3845 -2165
rect 3875 -2195 3925 -2165
rect 3955 -2195 4005 -2165
rect 4035 -2195 4085 -2165
rect 4115 -2195 4165 -2165
rect 4195 -2195 4245 -2165
rect 4275 -2195 4325 -2165
rect 4355 -2195 4405 -2165
rect 4435 -2195 4485 -2165
rect 4515 -2195 4565 -2165
rect 4595 -2195 4645 -2165
rect 4675 -2195 4725 -2165
rect 4755 -2195 4805 -2165
rect 4835 -2195 4885 -2165
rect 4915 -2195 4965 -2165
rect 4995 -2195 5045 -2165
rect 5075 -2195 5125 -2165
rect 5155 -2195 5205 -2165
rect 5235 -2195 5285 -2165
rect 5315 -2195 5365 -2165
rect 5395 -2195 5445 -2165
rect 5475 -2195 5525 -2165
rect 5555 -2195 5605 -2165
rect 5635 -2195 5685 -2165
rect 5715 -2195 5765 -2165
rect 5795 -2195 5845 -2165
rect 5875 -2195 5925 -2165
rect 5955 -2195 6005 -2165
rect 6035 -2195 6085 -2165
rect 6115 -2195 6165 -2165
rect 6195 -2195 6245 -2165
rect 6275 -2195 6325 -2165
rect 6355 -2195 6405 -2165
rect 6435 -2195 6485 -2165
rect 6515 -2195 6565 -2165
rect 6595 -2195 6645 -2165
rect 6675 -2195 6725 -2165
rect 6755 -2195 6805 -2165
rect 6835 -2195 6885 -2165
rect 6915 -2195 6965 -2165
rect 6995 -2195 7045 -2165
rect 7075 -2195 7125 -2165
rect 7155 -2195 7205 -2165
rect 7235 -2195 7285 -2165
rect 7315 -2195 7365 -2165
rect 7395 -2195 7445 -2165
rect 7475 -2195 7525 -2165
rect 7555 -2195 7605 -2165
rect 7635 -2195 7685 -2165
rect 7715 -2195 7765 -2165
rect 7795 -2195 7845 -2165
rect 7875 -2195 7925 -2165
rect 7955 -2195 8005 -2165
rect 8035 -2195 8085 -2165
rect 8115 -2195 8165 -2165
rect 8195 -2195 8245 -2165
rect 8275 -2195 8325 -2165
rect 8355 -2195 8405 -2165
rect 8435 -2195 8485 -2165
rect 8515 -2195 8565 -2165
rect 8595 -2195 8645 -2165
rect 8675 -2195 8725 -2165
rect 8755 -2195 8805 -2165
rect 8835 -2195 8885 -2165
rect 8915 -2195 8965 -2165
rect 8995 -2195 9045 -2165
rect 9075 -2195 9125 -2165
rect 9155 -2195 9205 -2165
rect 9235 -2195 9285 -2165
rect 9315 -2195 9365 -2165
rect 9395 -2195 9445 -2165
rect 9475 -2195 9525 -2165
rect 9555 -2195 9605 -2165
rect 9635 -2195 9685 -2165
rect 9715 -2195 9765 -2165
rect 9795 -2195 9845 -2165
rect 9875 -2195 9925 -2165
rect 9955 -2195 10005 -2165
rect 10035 -2195 10085 -2165
rect 10115 -2195 10165 -2165
rect 10195 -2195 10245 -2165
rect 10275 -2195 10325 -2165
rect 10355 -2195 10405 -2165
rect 10435 -2195 10485 -2165
rect 10515 -2195 10565 -2165
rect 10595 -2195 10645 -2165
rect 10675 -2195 10805 -2165
rect 10835 -2195 10965 -2165
rect 10995 -2195 11000 -2165
rect -720 -2200 11000 -2195
rect -720 -2245 -360 -2240
rect -720 -2275 -715 -2245
rect -685 -2275 -555 -2245
rect -525 -2275 -395 -2245
rect -365 -2275 -360 -2245
rect -720 -2280 -360 -2275
rect -320 -2245 10760 -2240
rect -320 -2275 10 -2245
rect 190 -2275 330 -2245
rect 510 -2275 650 -2245
rect 830 -2275 970 -2245
rect 1150 -2275 1290 -2245
rect 1470 -2275 1610 -2245
rect 1790 -2275 1930 -2245
rect 2110 -2275 2250 -2245
rect 2430 -2275 2570 -2245
rect 2750 -2275 2890 -2245
rect 3070 -2275 3210 -2245
rect 3390 -2275 3530 -2245
rect 3710 -2275 3850 -2245
rect 4030 -2275 4170 -2245
rect 4350 -2275 4490 -2245
rect 4670 -2275 4810 -2245
rect 4990 -2275 5205 -2245
rect 5235 -2275 5290 -2245
rect 5470 -2275 5610 -2245
rect 5790 -2275 5930 -2245
rect 6110 -2275 6250 -2245
rect 6430 -2275 6485 -2245
rect 6515 -2275 6570 -2245
rect 6750 -2275 6890 -2245
rect 7070 -2275 7210 -2245
rect 7390 -2275 7530 -2245
rect 7710 -2275 7850 -2245
rect 8030 -2275 8170 -2245
rect 8350 -2275 8490 -2245
rect 8670 -2275 8810 -2245
rect 8990 -2275 9045 -2245
rect 9075 -2275 9130 -2245
rect 9310 -2275 9450 -2245
rect 9630 -2275 9770 -2245
rect 9950 -2275 10090 -2245
rect 10270 -2275 10725 -2245
rect 10755 -2275 10760 -2245
rect -320 -2280 10760 -2275
rect 10800 -2245 11000 -2240
rect 10800 -2275 10805 -2245
rect 10835 -2275 10965 -2245
rect 10995 -2275 11000 -2245
rect 10800 -2280 11000 -2275
rect -720 -2325 11000 -2320
rect -720 -2355 -715 -2325
rect -685 -2355 -555 -2325
rect -525 -2355 -395 -2325
rect -365 -2355 -235 -2325
rect -205 -2355 -155 -2325
rect -125 -2355 -75 -2325
rect -45 -2355 5 -2325
rect 35 -2355 85 -2325
rect 115 -2355 165 -2325
rect 195 -2355 245 -2325
rect 275 -2355 325 -2325
rect 355 -2355 405 -2325
rect 435 -2355 485 -2325
rect 515 -2355 565 -2325
rect 595 -2355 645 -2325
rect 675 -2355 725 -2325
rect 755 -2355 805 -2325
rect 835 -2355 885 -2325
rect 915 -2355 965 -2325
rect 995 -2355 1045 -2325
rect 1075 -2355 1125 -2325
rect 1155 -2355 1205 -2325
rect 1235 -2355 1285 -2325
rect 1315 -2355 1365 -2325
rect 1395 -2355 1445 -2325
rect 1475 -2355 1525 -2325
rect 1555 -2355 1605 -2325
rect 1635 -2355 1685 -2325
rect 1715 -2355 1765 -2325
rect 1795 -2355 1845 -2325
rect 1875 -2355 1925 -2325
rect 1955 -2355 2005 -2325
rect 2035 -2355 2085 -2325
rect 2115 -2355 2165 -2325
rect 2195 -2355 2245 -2325
rect 2275 -2355 2325 -2325
rect 2355 -2355 2405 -2325
rect 2435 -2355 2485 -2325
rect 2515 -2355 2565 -2325
rect 2595 -2355 2645 -2325
rect 2675 -2355 2725 -2325
rect 2755 -2355 2805 -2325
rect 2835 -2355 2885 -2325
rect 2915 -2355 2965 -2325
rect 2995 -2355 3045 -2325
rect 3075 -2355 3125 -2325
rect 3155 -2355 3205 -2325
rect 3235 -2355 3285 -2325
rect 3315 -2355 3365 -2325
rect 3395 -2355 3445 -2325
rect 3475 -2355 3525 -2325
rect 3555 -2355 3605 -2325
rect 3635 -2355 3685 -2325
rect 3715 -2355 3765 -2325
rect 3795 -2355 3845 -2325
rect 3875 -2355 3925 -2325
rect 3955 -2355 4005 -2325
rect 4035 -2355 4085 -2325
rect 4115 -2355 4165 -2325
rect 4195 -2355 4245 -2325
rect 4275 -2355 4325 -2325
rect 4355 -2355 4405 -2325
rect 4435 -2355 4485 -2325
rect 4515 -2355 4565 -2325
rect 4595 -2355 4645 -2325
rect 4675 -2355 4725 -2325
rect 4755 -2355 4805 -2325
rect 4835 -2355 4885 -2325
rect 4915 -2355 4965 -2325
rect 4995 -2355 5045 -2325
rect 5075 -2355 5125 -2325
rect 5155 -2355 5205 -2325
rect 5235 -2355 5285 -2325
rect 5315 -2355 5365 -2325
rect 5395 -2355 5445 -2325
rect 5475 -2355 5525 -2325
rect 5555 -2355 5605 -2325
rect 5635 -2355 5685 -2325
rect 5715 -2355 5765 -2325
rect 5795 -2355 5845 -2325
rect 5875 -2355 5925 -2325
rect 5955 -2355 6005 -2325
rect 6035 -2355 6085 -2325
rect 6115 -2355 6165 -2325
rect 6195 -2355 6245 -2325
rect 6275 -2355 6325 -2325
rect 6355 -2355 6405 -2325
rect 6435 -2355 6485 -2325
rect 6515 -2355 6565 -2325
rect 6595 -2355 6645 -2325
rect 6675 -2355 6725 -2325
rect 6755 -2355 6805 -2325
rect 6835 -2355 6885 -2325
rect 6915 -2355 6965 -2325
rect 6995 -2355 7045 -2325
rect 7075 -2355 7125 -2325
rect 7155 -2355 7205 -2325
rect 7235 -2355 7285 -2325
rect 7315 -2355 7365 -2325
rect 7395 -2355 7445 -2325
rect 7475 -2355 7525 -2325
rect 7555 -2355 7605 -2325
rect 7635 -2355 7685 -2325
rect 7715 -2355 7765 -2325
rect 7795 -2355 7845 -2325
rect 7875 -2355 7925 -2325
rect 7955 -2355 8005 -2325
rect 8035 -2355 8085 -2325
rect 8115 -2355 8165 -2325
rect 8195 -2355 8245 -2325
rect 8275 -2355 8325 -2325
rect 8355 -2355 8405 -2325
rect 8435 -2355 8485 -2325
rect 8515 -2355 8565 -2325
rect 8595 -2355 8645 -2325
rect 8675 -2355 8725 -2325
rect 8755 -2355 8805 -2325
rect 8835 -2355 8885 -2325
rect 8915 -2355 8965 -2325
rect 8995 -2355 9045 -2325
rect 9075 -2355 9125 -2325
rect 9155 -2355 9205 -2325
rect 9235 -2355 9285 -2325
rect 9315 -2355 9365 -2325
rect 9395 -2355 9445 -2325
rect 9475 -2355 9525 -2325
rect 9555 -2355 9605 -2325
rect 9635 -2355 9685 -2325
rect 9715 -2355 9765 -2325
rect 9795 -2355 9845 -2325
rect 9875 -2355 9925 -2325
rect 9955 -2355 10005 -2325
rect 10035 -2355 10085 -2325
rect 10115 -2355 10165 -2325
rect 10195 -2355 10245 -2325
rect 10275 -2355 10325 -2325
rect 10355 -2355 10405 -2325
rect 10435 -2355 10485 -2325
rect 10515 -2355 10565 -2325
rect 10595 -2355 10645 -2325
rect 10675 -2355 10805 -2325
rect 10835 -2355 10965 -2325
rect 10995 -2355 11000 -2325
rect -720 -2360 11000 -2355
rect -720 -2405 11000 -2400
rect -720 -2435 -715 -2405
rect -685 -2435 -555 -2405
rect -525 -2435 -395 -2405
rect -365 -2435 -235 -2405
rect -205 -2435 -155 -2405
rect -125 -2435 -75 -2405
rect -45 -2435 5 -2405
rect 35 -2435 85 -2405
rect 115 -2435 165 -2405
rect 195 -2435 245 -2405
rect 275 -2435 325 -2405
rect 355 -2435 405 -2405
rect 435 -2435 485 -2405
rect 515 -2435 565 -2405
rect 595 -2435 645 -2405
rect 675 -2435 725 -2405
rect 755 -2435 805 -2405
rect 835 -2435 885 -2405
rect 915 -2435 965 -2405
rect 995 -2435 1045 -2405
rect 1075 -2435 1125 -2405
rect 1155 -2435 1205 -2405
rect 1235 -2435 1285 -2405
rect 1315 -2435 1365 -2405
rect 1395 -2435 1445 -2405
rect 1475 -2435 1525 -2405
rect 1555 -2435 1605 -2405
rect 1635 -2435 1685 -2405
rect 1715 -2435 1765 -2405
rect 1795 -2435 1845 -2405
rect 1875 -2435 1925 -2405
rect 1955 -2435 2005 -2405
rect 2035 -2435 2085 -2405
rect 2115 -2435 2165 -2405
rect 2195 -2435 2245 -2405
rect 2275 -2435 2325 -2405
rect 2355 -2435 2405 -2405
rect 2435 -2435 2485 -2405
rect 2515 -2435 2565 -2405
rect 2595 -2435 2645 -2405
rect 2675 -2435 2725 -2405
rect 2755 -2435 2805 -2405
rect 2835 -2435 2885 -2405
rect 2915 -2435 2965 -2405
rect 2995 -2435 3045 -2405
rect 3075 -2435 3125 -2405
rect 3155 -2435 3205 -2405
rect 3235 -2435 3285 -2405
rect 3315 -2435 3365 -2405
rect 3395 -2435 3445 -2405
rect 3475 -2435 3525 -2405
rect 3555 -2435 3605 -2405
rect 3635 -2435 3685 -2405
rect 3715 -2435 3765 -2405
rect 3795 -2435 3845 -2405
rect 3875 -2435 3925 -2405
rect 3955 -2435 4005 -2405
rect 4035 -2435 4085 -2405
rect 4115 -2435 4165 -2405
rect 4195 -2435 4245 -2405
rect 4275 -2435 4325 -2405
rect 4355 -2435 4405 -2405
rect 4435 -2435 4485 -2405
rect 4515 -2435 4565 -2405
rect 4595 -2435 4645 -2405
rect 4675 -2435 4725 -2405
rect 4755 -2435 4805 -2405
rect 4835 -2435 4885 -2405
rect 4915 -2435 4965 -2405
rect 4995 -2435 5045 -2405
rect 5075 -2435 5125 -2405
rect 5155 -2435 5205 -2405
rect 5235 -2435 5285 -2405
rect 5315 -2435 5365 -2405
rect 5395 -2435 5445 -2405
rect 5475 -2435 5525 -2405
rect 5555 -2435 5605 -2405
rect 5635 -2435 5685 -2405
rect 5715 -2435 5765 -2405
rect 5795 -2435 5845 -2405
rect 5875 -2435 5925 -2405
rect 5955 -2435 6005 -2405
rect 6035 -2435 6085 -2405
rect 6115 -2435 6165 -2405
rect 6195 -2435 6245 -2405
rect 6275 -2435 6325 -2405
rect 6355 -2435 6405 -2405
rect 6435 -2435 6485 -2405
rect 6515 -2435 6565 -2405
rect 6595 -2435 6645 -2405
rect 6675 -2435 6725 -2405
rect 6755 -2435 6805 -2405
rect 6835 -2435 6885 -2405
rect 6915 -2435 6965 -2405
rect 6995 -2435 7045 -2405
rect 7075 -2435 7125 -2405
rect 7155 -2435 7205 -2405
rect 7235 -2435 7285 -2405
rect 7315 -2435 7365 -2405
rect 7395 -2435 7445 -2405
rect 7475 -2435 7525 -2405
rect 7555 -2435 7605 -2405
rect 7635 -2435 7685 -2405
rect 7715 -2435 7765 -2405
rect 7795 -2435 7845 -2405
rect 7875 -2435 7925 -2405
rect 7955 -2435 8005 -2405
rect 8035 -2435 8085 -2405
rect 8115 -2435 8165 -2405
rect 8195 -2435 8245 -2405
rect 8275 -2435 8325 -2405
rect 8355 -2435 8405 -2405
rect 8435 -2435 8485 -2405
rect 8515 -2435 8565 -2405
rect 8595 -2435 8645 -2405
rect 8675 -2435 8725 -2405
rect 8755 -2435 8805 -2405
rect 8835 -2435 8885 -2405
rect 8915 -2435 8965 -2405
rect 8995 -2435 9045 -2405
rect 9075 -2435 9125 -2405
rect 9155 -2435 9205 -2405
rect 9235 -2435 9285 -2405
rect 9315 -2435 9365 -2405
rect 9395 -2435 9445 -2405
rect 9475 -2435 9525 -2405
rect 9555 -2435 9605 -2405
rect 9635 -2435 9685 -2405
rect 9715 -2435 9765 -2405
rect 9795 -2435 9845 -2405
rect 9875 -2435 9925 -2405
rect 9955 -2435 10005 -2405
rect 10035 -2435 10085 -2405
rect 10115 -2435 10165 -2405
rect 10195 -2435 10245 -2405
rect 10275 -2435 10325 -2405
rect 10355 -2435 10405 -2405
rect 10435 -2435 10485 -2405
rect 10515 -2435 10565 -2405
rect 10595 -2435 10645 -2405
rect 10675 -2435 10805 -2405
rect 10835 -2435 10965 -2405
rect 10995 -2435 11000 -2405
rect -720 -2440 11000 -2435
rect -720 -2485 11000 -2480
rect -720 -2515 -715 -2485
rect -685 -2515 -555 -2485
rect -525 -2515 -395 -2485
rect -365 -2515 -235 -2485
rect -205 -2515 -155 -2485
rect -125 -2515 -75 -2485
rect -45 -2515 5 -2485
rect 35 -2515 85 -2485
rect 115 -2515 165 -2485
rect 195 -2515 245 -2485
rect 275 -2515 325 -2485
rect 355 -2515 405 -2485
rect 435 -2515 485 -2485
rect 515 -2515 565 -2485
rect 595 -2515 645 -2485
rect 675 -2515 725 -2485
rect 755 -2515 805 -2485
rect 835 -2515 885 -2485
rect 915 -2515 965 -2485
rect 995 -2515 1045 -2485
rect 1075 -2515 1125 -2485
rect 1155 -2515 1205 -2485
rect 1235 -2515 1285 -2485
rect 1315 -2515 1365 -2485
rect 1395 -2515 1445 -2485
rect 1475 -2515 1525 -2485
rect 1555 -2515 1605 -2485
rect 1635 -2515 1685 -2485
rect 1715 -2515 1765 -2485
rect 1795 -2515 1845 -2485
rect 1875 -2515 1925 -2485
rect 1955 -2515 2005 -2485
rect 2035 -2515 2085 -2485
rect 2115 -2515 2165 -2485
rect 2195 -2515 2245 -2485
rect 2275 -2515 2325 -2485
rect 2355 -2515 2405 -2485
rect 2435 -2515 2485 -2485
rect 2515 -2515 2565 -2485
rect 2595 -2515 2645 -2485
rect 2675 -2515 2725 -2485
rect 2755 -2515 2805 -2485
rect 2835 -2515 2885 -2485
rect 2915 -2515 2965 -2485
rect 2995 -2515 3045 -2485
rect 3075 -2515 3125 -2485
rect 3155 -2515 3205 -2485
rect 3235 -2515 3285 -2485
rect 3315 -2515 3365 -2485
rect 3395 -2515 3445 -2485
rect 3475 -2515 3525 -2485
rect 3555 -2515 3605 -2485
rect 3635 -2515 3685 -2485
rect 3715 -2515 3765 -2485
rect 3795 -2515 3845 -2485
rect 3875 -2515 3925 -2485
rect 3955 -2515 4005 -2485
rect 4035 -2515 4085 -2485
rect 4115 -2515 4165 -2485
rect 4195 -2515 4245 -2485
rect 4275 -2515 4325 -2485
rect 4355 -2515 4405 -2485
rect 4435 -2515 4485 -2485
rect 4515 -2515 4565 -2485
rect 4595 -2515 4645 -2485
rect 4675 -2515 4725 -2485
rect 4755 -2515 4805 -2485
rect 4835 -2515 4885 -2485
rect 4915 -2515 4965 -2485
rect 4995 -2515 5045 -2485
rect 5075 -2515 5125 -2485
rect 5155 -2515 5205 -2485
rect 5235 -2515 5285 -2485
rect 5315 -2515 5365 -2485
rect 5395 -2515 5445 -2485
rect 5475 -2515 5525 -2485
rect 5555 -2515 5605 -2485
rect 5635 -2515 5685 -2485
rect 5715 -2515 5765 -2485
rect 5795 -2515 5845 -2485
rect 5875 -2515 5925 -2485
rect 5955 -2515 6005 -2485
rect 6035 -2515 6085 -2485
rect 6115 -2515 6165 -2485
rect 6195 -2515 6245 -2485
rect 6275 -2515 6325 -2485
rect 6355 -2515 6405 -2485
rect 6435 -2515 6485 -2485
rect 6515 -2515 6565 -2485
rect 6595 -2515 6645 -2485
rect 6675 -2515 6725 -2485
rect 6755 -2515 6805 -2485
rect 6835 -2515 6885 -2485
rect 6915 -2515 6965 -2485
rect 6995 -2515 7045 -2485
rect 7075 -2515 7125 -2485
rect 7155 -2515 7205 -2485
rect 7235 -2515 7285 -2485
rect 7315 -2515 7365 -2485
rect 7395 -2515 7445 -2485
rect 7475 -2515 7525 -2485
rect 7555 -2515 7605 -2485
rect 7635 -2515 7685 -2485
rect 7715 -2515 7765 -2485
rect 7795 -2515 7845 -2485
rect 7875 -2515 7925 -2485
rect 7955 -2515 8005 -2485
rect 8035 -2515 8085 -2485
rect 8115 -2515 8165 -2485
rect 8195 -2515 8245 -2485
rect 8275 -2515 8325 -2485
rect 8355 -2515 8405 -2485
rect 8435 -2515 8485 -2485
rect 8515 -2515 8565 -2485
rect 8595 -2515 8645 -2485
rect 8675 -2515 8725 -2485
rect 8755 -2515 8805 -2485
rect 8835 -2515 8885 -2485
rect 8915 -2515 8965 -2485
rect 8995 -2515 9045 -2485
rect 9075 -2515 9125 -2485
rect 9155 -2515 9205 -2485
rect 9235 -2515 9285 -2485
rect 9315 -2515 9365 -2485
rect 9395 -2515 9445 -2485
rect 9475 -2515 9525 -2485
rect 9555 -2515 9605 -2485
rect 9635 -2515 9685 -2485
rect 9715 -2515 9765 -2485
rect 9795 -2515 9845 -2485
rect 9875 -2515 9925 -2485
rect 9955 -2515 10005 -2485
rect 10035 -2515 10085 -2485
rect 10115 -2515 10165 -2485
rect 10195 -2515 10245 -2485
rect 10275 -2515 10325 -2485
rect 10355 -2515 10405 -2485
rect 10435 -2515 10485 -2485
rect 10515 -2515 10565 -2485
rect 10595 -2515 10645 -2485
rect 10675 -2515 10805 -2485
rect 10835 -2515 10965 -2485
rect 10995 -2515 11000 -2485
rect -720 -2520 11000 -2515
rect -720 -2565 11000 -2560
rect -720 -2595 -715 -2565
rect -685 -2595 -555 -2565
rect -525 -2595 -395 -2565
rect -365 -2595 -315 -2565
rect -285 -2595 -235 -2565
rect -205 -2595 -155 -2565
rect -125 -2595 -75 -2565
rect -45 -2595 5 -2565
rect 35 -2595 85 -2565
rect 115 -2595 165 -2565
rect 195 -2595 245 -2565
rect 275 -2595 325 -2565
rect 355 -2595 405 -2565
rect 435 -2595 485 -2565
rect 515 -2595 565 -2565
rect 595 -2595 645 -2565
rect 675 -2595 725 -2565
rect 755 -2595 805 -2565
rect 835 -2595 885 -2565
rect 915 -2595 965 -2565
rect 995 -2595 1045 -2565
rect 1075 -2595 1125 -2565
rect 1155 -2595 1205 -2565
rect 1235 -2595 1285 -2565
rect 1315 -2595 1365 -2565
rect 1395 -2595 1445 -2565
rect 1475 -2595 1525 -2565
rect 1555 -2595 1605 -2565
rect 1635 -2595 1685 -2565
rect 1715 -2595 1765 -2565
rect 1795 -2595 1845 -2565
rect 1875 -2595 1925 -2565
rect 1955 -2595 2005 -2565
rect 2035 -2595 2085 -2565
rect 2115 -2595 2165 -2565
rect 2195 -2595 2245 -2565
rect 2275 -2595 2325 -2565
rect 2355 -2595 2405 -2565
rect 2435 -2595 2485 -2565
rect 2515 -2595 2565 -2565
rect 2595 -2595 2645 -2565
rect 2675 -2595 2725 -2565
rect 2755 -2595 2805 -2565
rect 2835 -2595 2885 -2565
rect 2915 -2595 2965 -2565
rect 2995 -2595 3045 -2565
rect 3075 -2595 3125 -2565
rect 3155 -2595 3205 -2565
rect 3235 -2595 3285 -2565
rect 3315 -2595 3365 -2565
rect 3395 -2595 3445 -2565
rect 3475 -2595 3525 -2565
rect 3555 -2595 3605 -2565
rect 3635 -2595 3685 -2565
rect 3715 -2595 3765 -2565
rect 3795 -2595 3845 -2565
rect 3875 -2595 3925 -2565
rect 3955 -2595 4005 -2565
rect 4035 -2595 4085 -2565
rect 4115 -2595 4165 -2565
rect 4195 -2595 4245 -2565
rect 4275 -2595 4325 -2565
rect 4355 -2595 4405 -2565
rect 4435 -2595 4485 -2565
rect 4515 -2595 4565 -2565
rect 4595 -2595 4645 -2565
rect 4675 -2595 4725 -2565
rect 4755 -2595 4805 -2565
rect 4835 -2595 4885 -2565
rect 4915 -2595 4965 -2565
rect 4995 -2595 5045 -2565
rect 5075 -2595 5125 -2565
rect 5155 -2595 5205 -2565
rect 5235 -2595 5285 -2565
rect 5315 -2595 5365 -2565
rect 5395 -2595 5445 -2565
rect 5475 -2595 5525 -2565
rect 5555 -2595 5605 -2565
rect 5635 -2595 5685 -2565
rect 5715 -2595 5765 -2565
rect 5795 -2595 5845 -2565
rect 5875 -2595 5925 -2565
rect 5955 -2595 6005 -2565
rect 6035 -2595 6085 -2565
rect 6115 -2595 6165 -2565
rect 6195 -2595 6245 -2565
rect 6275 -2595 6325 -2565
rect 6355 -2595 6405 -2565
rect 6435 -2595 6485 -2565
rect 6515 -2595 6565 -2565
rect 6595 -2595 6645 -2565
rect 6675 -2595 6725 -2565
rect 6755 -2595 6805 -2565
rect 6835 -2595 6885 -2565
rect 6915 -2595 6965 -2565
rect 6995 -2595 7045 -2565
rect 7075 -2595 7125 -2565
rect 7155 -2595 7205 -2565
rect 7235 -2595 7285 -2565
rect 7315 -2595 7365 -2565
rect 7395 -2595 7445 -2565
rect 7475 -2595 7525 -2565
rect 7555 -2595 7605 -2565
rect 7635 -2595 7685 -2565
rect 7715 -2595 7765 -2565
rect 7795 -2595 7845 -2565
rect 7875 -2595 7925 -2565
rect 7955 -2595 8005 -2565
rect 8035 -2595 8085 -2565
rect 8115 -2595 8165 -2565
rect 8195 -2595 8245 -2565
rect 8275 -2595 8325 -2565
rect 8355 -2595 8405 -2565
rect 8435 -2595 8485 -2565
rect 8515 -2595 8565 -2565
rect 8595 -2595 8645 -2565
rect 8675 -2595 8725 -2565
rect 8755 -2595 8805 -2565
rect 8835 -2595 8885 -2565
rect 8915 -2595 8965 -2565
rect 8995 -2595 9045 -2565
rect 9075 -2595 9125 -2565
rect 9155 -2595 9205 -2565
rect 9235 -2595 9285 -2565
rect 9315 -2595 9365 -2565
rect 9395 -2595 9445 -2565
rect 9475 -2595 9525 -2565
rect 9555 -2595 9605 -2565
rect 9635 -2595 9685 -2565
rect 9715 -2595 9765 -2565
rect 9795 -2595 9845 -2565
rect 9875 -2595 9925 -2565
rect 9955 -2595 10005 -2565
rect 10035 -2595 10085 -2565
rect 10115 -2595 10165 -2565
rect 10195 -2595 10245 -2565
rect 10275 -2595 10325 -2565
rect 10355 -2595 10405 -2565
rect 10435 -2595 10485 -2565
rect 10515 -2595 10645 -2565
rect 10675 -2595 10805 -2565
rect 10835 -2595 10965 -2565
rect 10995 -2595 11000 -2565
rect -720 -2600 11000 -2595
rect -720 -2645 11000 -2640
rect -720 -2675 -715 -2645
rect -685 -2675 -555 -2645
rect -525 -2675 -395 -2645
rect -365 -2675 -315 -2645
rect -285 -2675 -235 -2645
rect -205 -2675 -155 -2645
rect -125 -2675 -75 -2645
rect -45 -2675 5 -2645
rect 35 -2675 85 -2645
rect 115 -2675 165 -2645
rect 195 -2675 245 -2645
rect 275 -2675 325 -2645
rect 355 -2675 405 -2645
rect 435 -2675 485 -2645
rect 515 -2675 565 -2645
rect 595 -2675 645 -2645
rect 675 -2675 725 -2645
rect 755 -2675 805 -2645
rect 835 -2675 885 -2645
rect 915 -2675 965 -2645
rect 995 -2675 1045 -2645
rect 1075 -2675 1125 -2645
rect 1155 -2675 1205 -2645
rect 1235 -2675 1285 -2645
rect 1315 -2675 1365 -2645
rect 1395 -2675 1445 -2645
rect 1475 -2675 1525 -2645
rect 1555 -2675 1605 -2645
rect 1635 -2675 1685 -2645
rect 1715 -2675 1765 -2645
rect 1795 -2675 1845 -2645
rect 1875 -2675 1925 -2645
rect 1955 -2675 2005 -2645
rect 2035 -2675 2085 -2645
rect 2115 -2675 2165 -2645
rect 2195 -2675 2245 -2645
rect 2275 -2675 2325 -2645
rect 2355 -2675 2405 -2645
rect 2435 -2675 2485 -2645
rect 2515 -2675 2565 -2645
rect 2595 -2675 2645 -2645
rect 2675 -2675 2725 -2645
rect 2755 -2675 2805 -2645
rect 2835 -2675 2885 -2645
rect 2915 -2675 2965 -2645
rect 2995 -2675 3045 -2645
rect 3075 -2675 3125 -2645
rect 3155 -2675 3205 -2645
rect 3235 -2675 3285 -2645
rect 3315 -2675 3365 -2645
rect 3395 -2675 3445 -2645
rect 3475 -2675 3525 -2645
rect 3555 -2675 3605 -2645
rect 3635 -2675 3685 -2645
rect 3715 -2675 3765 -2645
rect 3795 -2675 3845 -2645
rect 3875 -2675 3925 -2645
rect 3955 -2675 4005 -2645
rect 4035 -2675 4085 -2645
rect 4115 -2675 4165 -2645
rect 4195 -2675 4245 -2645
rect 4275 -2675 4325 -2645
rect 4355 -2675 4405 -2645
rect 4435 -2675 4485 -2645
rect 4515 -2675 4565 -2645
rect 4595 -2675 4645 -2645
rect 4675 -2675 4725 -2645
rect 4755 -2675 4805 -2645
rect 4835 -2675 4885 -2645
rect 4915 -2675 4965 -2645
rect 4995 -2675 5045 -2645
rect 5075 -2675 5125 -2645
rect 5155 -2675 5205 -2645
rect 5235 -2675 5285 -2645
rect 5315 -2675 5365 -2645
rect 5395 -2675 5445 -2645
rect 5475 -2675 5525 -2645
rect 5555 -2675 5605 -2645
rect 5635 -2675 5685 -2645
rect 5715 -2675 5765 -2645
rect 5795 -2675 5845 -2645
rect 5875 -2675 5925 -2645
rect 5955 -2675 6005 -2645
rect 6035 -2675 6085 -2645
rect 6115 -2675 6165 -2645
rect 6195 -2675 6245 -2645
rect 6275 -2675 6325 -2645
rect 6355 -2675 6405 -2645
rect 6435 -2675 6485 -2645
rect 6515 -2675 6565 -2645
rect 6595 -2675 6645 -2645
rect 6675 -2675 6725 -2645
rect 6755 -2675 6805 -2645
rect 6835 -2675 6885 -2645
rect 6915 -2675 6965 -2645
rect 6995 -2675 7045 -2645
rect 7075 -2675 7125 -2645
rect 7155 -2675 7205 -2645
rect 7235 -2675 7285 -2645
rect 7315 -2675 7365 -2645
rect 7395 -2675 7445 -2645
rect 7475 -2675 7525 -2645
rect 7555 -2675 7605 -2645
rect 7635 -2675 7685 -2645
rect 7715 -2675 7765 -2645
rect 7795 -2675 7845 -2645
rect 7875 -2675 7925 -2645
rect 7955 -2675 8005 -2645
rect 8035 -2675 8085 -2645
rect 8115 -2675 8165 -2645
rect 8195 -2675 8245 -2645
rect 8275 -2675 8325 -2645
rect 8355 -2675 8405 -2645
rect 8435 -2675 8485 -2645
rect 8515 -2675 8565 -2645
rect 8595 -2675 8645 -2645
rect 8675 -2675 8725 -2645
rect 8755 -2675 8805 -2645
rect 8835 -2675 8885 -2645
rect 8915 -2675 8965 -2645
rect 8995 -2675 9045 -2645
rect 9075 -2675 9125 -2645
rect 9155 -2675 9205 -2645
rect 9235 -2675 9285 -2645
rect 9315 -2675 9365 -2645
rect 9395 -2675 9445 -2645
rect 9475 -2675 9525 -2645
rect 9555 -2675 9605 -2645
rect 9635 -2675 9685 -2645
rect 9715 -2675 9765 -2645
rect 9795 -2675 9845 -2645
rect 9875 -2675 9925 -2645
rect 9955 -2675 10005 -2645
rect 10035 -2675 10085 -2645
rect 10115 -2675 10165 -2645
rect 10195 -2675 10245 -2645
rect 10275 -2675 10325 -2645
rect 10355 -2675 10405 -2645
rect 10435 -2675 10485 -2645
rect 10515 -2675 10645 -2645
rect 10675 -2675 10805 -2645
rect 10835 -2675 10965 -2645
rect 10995 -2675 11000 -2645
rect -720 -2680 11000 -2675
rect -720 -2725 11000 -2720
rect -720 -2755 -715 -2725
rect -685 -2755 -555 -2725
rect -525 -2755 -395 -2725
rect -365 -2755 -315 -2725
rect -285 -2755 -235 -2725
rect -205 -2755 -155 -2725
rect -125 -2755 -75 -2725
rect -45 -2755 5 -2725
rect 35 -2755 85 -2725
rect 115 -2755 165 -2725
rect 195 -2755 245 -2725
rect 275 -2755 325 -2725
rect 355 -2755 405 -2725
rect 435 -2755 485 -2725
rect 515 -2755 565 -2725
rect 595 -2755 645 -2725
rect 675 -2755 725 -2725
rect 755 -2755 805 -2725
rect 835 -2755 885 -2725
rect 915 -2755 965 -2725
rect 995 -2755 1045 -2725
rect 1075 -2755 1125 -2725
rect 1155 -2755 1205 -2725
rect 1235 -2755 1285 -2725
rect 1315 -2755 1365 -2725
rect 1395 -2755 1445 -2725
rect 1475 -2755 1525 -2725
rect 1555 -2755 1605 -2725
rect 1635 -2755 1685 -2725
rect 1715 -2755 1765 -2725
rect 1795 -2755 1845 -2725
rect 1875 -2755 1925 -2725
rect 1955 -2755 2005 -2725
rect 2035 -2755 2085 -2725
rect 2115 -2755 2165 -2725
rect 2195 -2755 2245 -2725
rect 2275 -2755 2325 -2725
rect 2355 -2755 2405 -2725
rect 2435 -2755 2485 -2725
rect 2515 -2755 2565 -2725
rect 2595 -2755 2645 -2725
rect 2675 -2755 2725 -2725
rect 2755 -2755 2805 -2725
rect 2835 -2755 2885 -2725
rect 2915 -2755 2965 -2725
rect 2995 -2755 3045 -2725
rect 3075 -2755 3125 -2725
rect 3155 -2755 3205 -2725
rect 3235 -2755 3285 -2725
rect 3315 -2755 3365 -2725
rect 3395 -2755 3445 -2725
rect 3475 -2755 3525 -2725
rect 3555 -2755 3605 -2725
rect 3635 -2755 3685 -2725
rect 3715 -2755 3765 -2725
rect 3795 -2755 3845 -2725
rect 3875 -2755 3925 -2725
rect 3955 -2755 4005 -2725
rect 4035 -2755 4085 -2725
rect 4115 -2755 4165 -2725
rect 4195 -2755 4245 -2725
rect 4275 -2755 4325 -2725
rect 4355 -2755 4405 -2725
rect 4435 -2755 4485 -2725
rect 4515 -2755 4565 -2725
rect 4595 -2755 4645 -2725
rect 4675 -2755 4725 -2725
rect 4755 -2755 4805 -2725
rect 4835 -2755 4885 -2725
rect 4915 -2755 4965 -2725
rect 4995 -2755 5045 -2725
rect 5075 -2755 5125 -2725
rect 5155 -2755 5205 -2725
rect 5235 -2755 5285 -2725
rect 5315 -2755 5365 -2725
rect 5395 -2755 5445 -2725
rect 5475 -2755 5525 -2725
rect 5555 -2755 5605 -2725
rect 5635 -2755 5685 -2725
rect 5715 -2755 5765 -2725
rect 5795 -2755 5845 -2725
rect 5875 -2755 5925 -2725
rect 5955 -2755 6005 -2725
rect 6035 -2755 6085 -2725
rect 6115 -2755 6165 -2725
rect 6195 -2755 6245 -2725
rect 6275 -2755 6325 -2725
rect 6355 -2755 6405 -2725
rect 6435 -2755 6485 -2725
rect 6515 -2755 6565 -2725
rect 6595 -2755 6645 -2725
rect 6675 -2755 6725 -2725
rect 6755 -2755 6805 -2725
rect 6835 -2755 6885 -2725
rect 6915 -2755 6965 -2725
rect 6995 -2755 7045 -2725
rect 7075 -2755 7125 -2725
rect 7155 -2755 7205 -2725
rect 7235 -2755 7285 -2725
rect 7315 -2755 7365 -2725
rect 7395 -2755 7445 -2725
rect 7475 -2755 7525 -2725
rect 7555 -2755 7605 -2725
rect 7635 -2755 7685 -2725
rect 7715 -2755 7765 -2725
rect 7795 -2755 7845 -2725
rect 7875 -2755 7925 -2725
rect 7955 -2755 8005 -2725
rect 8035 -2755 8085 -2725
rect 8115 -2755 8165 -2725
rect 8195 -2755 8245 -2725
rect 8275 -2755 8325 -2725
rect 8355 -2755 8405 -2725
rect 8435 -2755 8485 -2725
rect 8515 -2755 8565 -2725
rect 8595 -2755 8645 -2725
rect 8675 -2755 8725 -2725
rect 8755 -2755 8805 -2725
rect 8835 -2755 8885 -2725
rect 8915 -2755 8965 -2725
rect 8995 -2755 9045 -2725
rect 9075 -2755 9125 -2725
rect 9155 -2755 9205 -2725
rect 9235 -2755 9285 -2725
rect 9315 -2755 9365 -2725
rect 9395 -2755 9445 -2725
rect 9475 -2755 9525 -2725
rect 9555 -2755 9605 -2725
rect 9635 -2755 9685 -2725
rect 9715 -2755 9765 -2725
rect 9795 -2755 9845 -2725
rect 9875 -2755 9925 -2725
rect 9955 -2755 10005 -2725
rect 10035 -2755 10085 -2725
rect 10115 -2755 10165 -2725
rect 10195 -2755 10245 -2725
rect 10275 -2755 10325 -2725
rect 10355 -2755 10405 -2725
rect 10435 -2755 10485 -2725
rect 10515 -2755 10645 -2725
rect 10675 -2755 10805 -2725
rect 10835 -2755 10965 -2725
rect 10995 -2755 11000 -2725
rect -720 -2760 11000 -2755
rect -720 -2805 -360 -2800
rect -720 -2835 -715 -2805
rect -685 -2835 -555 -2805
rect -525 -2835 -395 -2805
rect -365 -2835 -360 -2805
rect -720 -2840 -360 -2835
rect -320 -2805 10760 -2800
rect -320 -2835 10 -2805
rect 190 -2835 330 -2805
rect 510 -2835 650 -2805
rect 830 -2835 970 -2805
rect 1150 -2835 1205 -2805
rect 1235 -2835 1290 -2805
rect 1470 -2835 1610 -2805
rect 1790 -2835 1930 -2805
rect 2110 -2835 2250 -2805
rect 2430 -2835 2570 -2805
rect 2750 -2835 2890 -2805
rect 3070 -2835 3210 -2805
rect 3390 -2835 3530 -2805
rect 3710 -2835 3765 -2805
rect 3795 -2835 3850 -2805
rect 4030 -2835 4170 -2805
rect 4350 -2835 4490 -2805
rect 4670 -2835 4810 -2805
rect 4990 -2835 5045 -2805
rect 5075 -2835 5290 -2805
rect 5470 -2835 5610 -2805
rect 5790 -2835 5930 -2805
rect 6110 -2835 6250 -2805
rect 6430 -2835 6570 -2805
rect 6750 -2835 6890 -2805
rect 7070 -2835 7210 -2805
rect 7390 -2835 7530 -2805
rect 7710 -2835 7850 -2805
rect 8030 -2835 8170 -2805
rect 8350 -2835 8490 -2805
rect 8670 -2835 8810 -2805
rect 8990 -2835 9130 -2805
rect 9310 -2835 9450 -2805
rect 9630 -2835 9770 -2805
rect 9950 -2835 10090 -2805
rect 10270 -2835 10725 -2805
rect 10755 -2835 10760 -2805
rect -320 -2840 10760 -2835
rect 10800 -2805 11000 -2800
rect 10800 -2835 10805 -2805
rect 10835 -2835 10965 -2805
rect 10995 -2835 11000 -2805
rect 10800 -2840 11000 -2835
rect -720 -2885 11000 -2880
rect -720 -2915 -715 -2885
rect -685 -2915 -555 -2885
rect -525 -2915 -395 -2885
rect -365 -2915 -315 -2885
rect -285 -2915 -235 -2885
rect -205 -2915 -155 -2885
rect -125 -2915 -75 -2885
rect -45 -2915 5 -2885
rect 35 -2915 85 -2885
rect 115 -2915 165 -2885
rect 195 -2915 245 -2885
rect 275 -2915 325 -2885
rect 355 -2915 405 -2885
rect 435 -2915 485 -2885
rect 515 -2915 565 -2885
rect 595 -2915 645 -2885
rect 675 -2915 725 -2885
rect 755 -2915 805 -2885
rect 835 -2915 885 -2885
rect 915 -2915 965 -2885
rect 995 -2915 1045 -2885
rect 1075 -2915 1125 -2885
rect 1155 -2915 1205 -2885
rect 1235 -2915 1285 -2885
rect 1315 -2915 1365 -2885
rect 1395 -2915 1445 -2885
rect 1475 -2915 1525 -2885
rect 1555 -2915 1605 -2885
rect 1635 -2915 1685 -2885
rect 1715 -2915 1765 -2885
rect 1795 -2915 1845 -2885
rect 1875 -2915 1925 -2885
rect 1955 -2915 2005 -2885
rect 2035 -2915 2085 -2885
rect 2115 -2915 2165 -2885
rect 2195 -2915 2245 -2885
rect 2275 -2915 2325 -2885
rect 2355 -2915 2405 -2885
rect 2435 -2915 2485 -2885
rect 2515 -2915 2565 -2885
rect 2595 -2915 2645 -2885
rect 2675 -2915 2725 -2885
rect 2755 -2915 2805 -2885
rect 2835 -2915 2885 -2885
rect 2915 -2915 2965 -2885
rect 2995 -2915 3045 -2885
rect 3075 -2915 3125 -2885
rect 3155 -2915 3205 -2885
rect 3235 -2915 3285 -2885
rect 3315 -2915 3365 -2885
rect 3395 -2915 3445 -2885
rect 3475 -2915 3525 -2885
rect 3555 -2915 3605 -2885
rect 3635 -2915 3685 -2885
rect 3715 -2915 3765 -2885
rect 3795 -2915 3845 -2885
rect 3875 -2915 3925 -2885
rect 3955 -2915 4005 -2885
rect 4035 -2915 4085 -2885
rect 4115 -2915 4165 -2885
rect 4195 -2915 4245 -2885
rect 4275 -2915 4325 -2885
rect 4355 -2915 4405 -2885
rect 4435 -2915 4485 -2885
rect 4515 -2915 4565 -2885
rect 4595 -2915 4645 -2885
rect 4675 -2915 4725 -2885
rect 4755 -2915 4805 -2885
rect 4835 -2915 4885 -2885
rect 4915 -2915 4965 -2885
rect 4995 -2915 5045 -2885
rect 5075 -2915 5125 -2885
rect 5155 -2915 5205 -2885
rect 5235 -2915 5285 -2885
rect 5315 -2915 5365 -2885
rect 5395 -2915 5445 -2885
rect 5475 -2915 5525 -2885
rect 5555 -2915 5605 -2885
rect 5635 -2915 5685 -2885
rect 5715 -2915 5765 -2885
rect 5795 -2915 5845 -2885
rect 5875 -2915 5925 -2885
rect 5955 -2915 6005 -2885
rect 6035 -2915 6085 -2885
rect 6115 -2915 6165 -2885
rect 6195 -2915 6245 -2885
rect 6275 -2915 6325 -2885
rect 6355 -2915 6405 -2885
rect 6435 -2915 6485 -2885
rect 6515 -2915 6565 -2885
rect 6595 -2915 6645 -2885
rect 6675 -2915 6725 -2885
rect 6755 -2915 6805 -2885
rect 6835 -2915 6885 -2885
rect 6915 -2915 6965 -2885
rect 6995 -2915 7045 -2885
rect 7075 -2915 7125 -2885
rect 7155 -2915 7205 -2885
rect 7235 -2915 7285 -2885
rect 7315 -2915 7365 -2885
rect 7395 -2915 7445 -2885
rect 7475 -2915 7525 -2885
rect 7555 -2915 7605 -2885
rect 7635 -2915 7685 -2885
rect 7715 -2915 7765 -2885
rect 7795 -2915 7845 -2885
rect 7875 -2915 7925 -2885
rect 7955 -2915 8005 -2885
rect 8035 -2915 8085 -2885
rect 8115 -2915 8165 -2885
rect 8195 -2915 8245 -2885
rect 8275 -2915 8325 -2885
rect 8355 -2915 8405 -2885
rect 8435 -2915 8485 -2885
rect 8515 -2915 8565 -2885
rect 8595 -2915 8645 -2885
rect 8675 -2915 8725 -2885
rect 8755 -2915 8805 -2885
rect 8835 -2915 8885 -2885
rect 8915 -2915 8965 -2885
rect 8995 -2915 9045 -2885
rect 9075 -2915 9125 -2885
rect 9155 -2915 9205 -2885
rect 9235 -2915 9285 -2885
rect 9315 -2915 9365 -2885
rect 9395 -2915 9445 -2885
rect 9475 -2915 9525 -2885
rect 9555 -2915 9605 -2885
rect 9635 -2915 9685 -2885
rect 9715 -2915 9765 -2885
rect 9795 -2915 9845 -2885
rect 9875 -2915 9925 -2885
rect 9955 -2915 10005 -2885
rect 10035 -2915 10085 -2885
rect 10115 -2915 10165 -2885
rect 10195 -2915 10245 -2885
rect 10275 -2915 10325 -2885
rect 10355 -2915 10405 -2885
rect 10435 -2915 10485 -2885
rect 10515 -2915 10645 -2885
rect 10675 -2915 10805 -2885
rect 10835 -2915 10965 -2885
rect 10995 -2915 11000 -2885
rect -720 -2920 11000 -2915
rect -720 -2965 -360 -2960
rect -720 -2995 -715 -2965
rect -685 -2995 -555 -2965
rect -525 -2995 -395 -2965
rect -365 -2995 -360 -2965
rect -720 -3000 -360 -2995
rect -320 -2965 10920 -2960
rect -320 -2995 5365 -2965
rect 5395 -2995 5525 -2965
rect 5555 -2995 5685 -2965
rect 5715 -2995 6005 -2965
rect 6035 -2995 6165 -2965
rect 6195 -2995 6325 -2965
rect 6355 -2995 6485 -2965
rect 6515 -2995 6645 -2965
rect 6675 -2995 6805 -2965
rect 6835 -2995 6965 -2965
rect 6995 -2995 7285 -2965
rect 7315 -2995 7445 -2965
rect 7475 -2995 7605 -2965
rect 7635 -2995 7925 -2965
rect 7955 -2995 8085 -2965
rect 8115 -2995 8245 -2965
rect 8275 -2995 8565 -2965
rect 8595 -2995 8725 -2965
rect 8755 -2995 8885 -2965
rect 8915 -2995 9045 -2965
rect 9075 -2995 9205 -2965
rect 9235 -2995 9365 -2965
rect 9395 -2995 9525 -2965
rect 9555 -2995 9845 -2965
rect 9875 -2995 10005 -2965
rect 10035 -2995 10165 -2965
rect 10195 -2995 10885 -2965
rect 10915 -2995 10920 -2965
rect -320 -3000 10920 -2995
rect 10960 -3000 11000 -2960
rect -720 -3045 11000 -3040
rect -720 -3075 -715 -3045
rect -685 -3075 -555 -3045
rect -525 -3075 -395 -3045
rect -365 -3075 -315 -3045
rect -285 -3075 -235 -3045
rect -205 -3075 -155 -3045
rect -125 -3075 -75 -3045
rect -45 -3075 5 -3045
rect 35 -3075 85 -3045
rect 115 -3075 165 -3045
rect 195 -3075 245 -3045
rect 275 -3075 325 -3045
rect 355 -3075 405 -3045
rect 435 -3075 485 -3045
rect 515 -3075 565 -3045
rect 595 -3075 645 -3045
rect 675 -3075 725 -3045
rect 755 -3075 805 -3045
rect 835 -3075 885 -3045
rect 915 -3075 965 -3045
rect 995 -3075 1045 -3045
rect 1075 -3075 1125 -3045
rect 1155 -3075 1205 -3045
rect 1235 -3075 1285 -3045
rect 1315 -3075 1365 -3045
rect 1395 -3075 1445 -3045
rect 1475 -3075 1525 -3045
rect 1555 -3075 1605 -3045
rect 1635 -3075 1685 -3045
rect 1715 -3075 1765 -3045
rect 1795 -3075 1845 -3045
rect 1875 -3075 1925 -3045
rect 1955 -3075 2005 -3045
rect 2035 -3075 2085 -3045
rect 2115 -3075 2165 -3045
rect 2195 -3075 2245 -3045
rect 2275 -3075 2325 -3045
rect 2355 -3075 2405 -3045
rect 2435 -3075 2485 -3045
rect 2515 -3075 2565 -3045
rect 2595 -3075 2645 -3045
rect 2675 -3075 2725 -3045
rect 2755 -3075 2805 -3045
rect 2835 -3075 2885 -3045
rect 2915 -3075 2965 -3045
rect 2995 -3075 3045 -3045
rect 3075 -3075 3125 -3045
rect 3155 -3075 3205 -3045
rect 3235 -3075 3285 -3045
rect 3315 -3075 3365 -3045
rect 3395 -3075 3445 -3045
rect 3475 -3075 3525 -3045
rect 3555 -3075 3605 -3045
rect 3635 -3075 3685 -3045
rect 3715 -3075 3765 -3045
rect 3795 -3075 3845 -3045
rect 3875 -3075 3925 -3045
rect 3955 -3075 4005 -3045
rect 4035 -3075 4085 -3045
rect 4115 -3075 4165 -3045
rect 4195 -3075 4245 -3045
rect 4275 -3075 4325 -3045
rect 4355 -3075 4405 -3045
rect 4435 -3075 4485 -3045
rect 4515 -3075 4565 -3045
rect 4595 -3075 4645 -3045
rect 4675 -3075 4725 -3045
rect 4755 -3075 4805 -3045
rect 4835 -3075 4885 -3045
rect 4915 -3075 4965 -3045
rect 4995 -3075 5045 -3045
rect 5075 -3075 5125 -3045
rect 5155 -3075 5205 -3045
rect 5235 -3075 5285 -3045
rect 5315 -3075 5365 -3045
rect 5395 -3075 5445 -3045
rect 5475 -3075 5525 -3045
rect 5555 -3075 5605 -3045
rect 5635 -3075 5685 -3045
rect 5715 -3075 5765 -3045
rect 5795 -3075 5845 -3045
rect 5875 -3075 5925 -3045
rect 5955 -3075 6005 -3045
rect 6035 -3075 6085 -3045
rect 6115 -3075 6165 -3045
rect 6195 -3075 6245 -3045
rect 6275 -3075 6325 -3045
rect 6355 -3075 6405 -3045
rect 6435 -3075 6485 -3045
rect 6515 -3075 6565 -3045
rect 6595 -3075 6645 -3045
rect 6675 -3075 6725 -3045
rect 6755 -3075 6805 -3045
rect 6835 -3075 6885 -3045
rect 6915 -3075 6965 -3045
rect 6995 -3075 7045 -3045
rect 7075 -3075 7125 -3045
rect 7155 -3075 7205 -3045
rect 7235 -3075 7285 -3045
rect 7315 -3075 7365 -3045
rect 7395 -3075 7445 -3045
rect 7475 -3075 7525 -3045
rect 7555 -3075 7605 -3045
rect 7635 -3075 7685 -3045
rect 7715 -3075 7765 -3045
rect 7795 -3075 7845 -3045
rect 7875 -3075 7925 -3045
rect 7955 -3075 8005 -3045
rect 8035 -3075 8085 -3045
rect 8115 -3075 8165 -3045
rect 8195 -3075 8245 -3045
rect 8275 -3075 8325 -3045
rect 8355 -3075 8405 -3045
rect 8435 -3075 8485 -3045
rect 8515 -3075 8565 -3045
rect 8595 -3075 8645 -3045
rect 8675 -3075 8725 -3045
rect 8755 -3075 8805 -3045
rect 8835 -3075 8885 -3045
rect 8915 -3075 8965 -3045
rect 8995 -3075 9045 -3045
rect 9075 -3075 9125 -3045
rect 9155 -3075 9205 -3045
rect 9235 -3075 9285 -3045
rect 9315 -3075 9365 -3045
rect 9395 -3075 9445 -3045
rect 9475 -3075 9525 -3045
rect 9555 -3075 9605 -3045
rect 9635 -3075 9685 -3045
rect 9715 -3075 9765 -3045
rect 9795 -3075 9845 -3045
rect 9875 -3075 9925 -3045
rect 9955 -3075 10005 -3045
rect 10035 -3075 10085 -3045
rect 10115 -3075 10165 -3045
rect 10195 -3075 10245 -3045
rect 10275 -3075 10325 -3045
rect 10355 -3075 10405 -3045
rect 10435 -3075 10485 -3045
rect 10515 -3075 10645 -3045
rect 10675 -3075 10805 -3045
rect 10835 -3075 10965 -3045
rect 10995 -3075 11000 -3045
rect -720 -3080 11000 -3075
rect -720 -3125 -520 -3120
rect -720 -3155 -715 -3125
rect -685 -3155 -555 -3125
rect -525 -3155 -520 -3125
rect -720 -3160 -520 -3155
rect -480 -3125 10600 -3120
rect -480 -3155 -475 -3125
rect -445 -3155 85 -3125
rect 115 -3155 405 -3125
rect 435 -3155 725 -3125
rect 755 -3155 1045 -3125
rect 1075 -3155 1365 -3125
rect 1395 -3155 1685 -3125
rect 1715 -3155 2005 -3125
rect 2035 -3155 2325 -3125
rect 2355 -3155 2645 -3125
rect 2675 -3155 2965 -3125
rect 2995 -3155 3285 -3125
rect 3315 -3155 3605 -3125
rect 3635 -3155 3925 -3125
rect 3955 -3155 4245 -3125
rect 4275 -3155 4565 -3125
rect 4595 -3155 4885 -3125
rect 4915 -3155 10600 -3125
rect -480 -3160 10600 -3155
rect 10640 -3125 11000 -3120
rect 10640 -3155 10645 -3125
rect 10675 -3155 10805 -3125
rect 10835 -3155 10965 -3125
rect 10995 -3155 11000 -3125
rect 10640 -3160 11000 -3155
rect -720 -3205 11000 -3200
rect -720 -3235 -715 -3205
rect -685 -3235 -555 -3205
rect -525 -3235 -395 -3205
rect -365 -3235 -315 -3205
rect -285 -3235 -235 -3205
rect -205 -3235 -155 -3205
rect -125 -3235 -75 -3205
rect -45 -3235 5 -3205
rect 35 -3235 85 -3205
rect 115 -3235 165 -3205
rect 195 -3235 245 -3205
rect 275 -3235 325 -3205
rect 355 -3235 405 -3205
rect 435 -3235 485 -3205
rect 515 -3235 565 -3205
rect 595 -3235 645 -3205
rect 675 -3235 725 -3205
rect 755 -3235 805 -3205
rect 835 -3235 885 -3205
rect 915 -3235 965 -3205
rect 995 -3235 1045 -3205
rect 1075 -3235 1125 -3205
rect 1155 -3235 1205 -3205
rect 1235 -3235 1285 -3205
rect 1315 -3235 1365 -3205
rect 1395 -3235 1445 -3205
rect 1475 -3235 1525 -3205
rect 1555 -3235 1605 -3205
rect 1635 -3235 1685 -3205
rect 1715 -3235 1765 -3205
rect 1795 -3235 1845 -3205
rect 1875 -3235 1925 -3205
rect 1955 -3235 2005 -3205
rect 2035 -3235 2085 -3205
rect 2115 -3235 2165 -3205
rect 2195 -3235 2245 -3205
rect 2275 -3235 2325 -3205
rect 2355 -3235 2405 -3205
rect 2435 -3235 2485 -3205
rect 2515 -3235 2565 -3205
rect 2595 -3235 2645 -3205
rect 2675 -3235 2725 -3205
rect 2755 -3235 2805 -3205
rect 2835 -3235 2885 -3205
rect 2915 -3235 2965 -3205
rect 2995 -3235 3045 -3205
rect 3075 -3235 3125 -3205
rect 3155 -3235 3205 -3205
rect 3235 -3235 3285 -3205
rect 3315 -3235 3365 -3205
rect 3395 -3235 3445 -3205
rect 3475 -3235 3525 -3205
rect 3555 -3235 3605 -3205
rect 3635 -3235 3685 -3205
rect 3715 -3235 3765 -3205
rect 3795 -3235 3845 -3205
rect 3875 -3235 3925 -3205
rect 3955 -3235 4005 -3205
rect 4035 -3235 4085 -3205
rect 4115 -3235 4165 -3205
rect 4195 -3235 4245 -3205
rect 4275 -3235 4325 -3205
rect 4355 -3235 4405 -3205
rect 4435 -3235 4485 -3205
rect 4515 -3235 4565 -3205
rect 4595 -3235 4645 -3205
rect 4675 -3235 4725 -3205
rect 4755 -3235 4805 -3205
rect 4835 -3235 4885 -3205
rect 4915 -3235 4965 -3205
rect 4995 -3235 5045 -3205
rect 5075 -3235 5125 -3205
rect 5155 -3235 5205 -3205
rect 5235 -3235 5285 -3205
rect 5315 -3235 5365 -3205
rect 5395 -3235 5445 -3205
rect 5475 -3235 5525 -3205
rect 5555 -3235 5605 -3205
rect 5635 -3235 5685 -3205
rect 5715 -3235 5765 -3205
rect 5795 -3235 5845 -3205
rect 5875 -3235 5925 -3205
rect 5955 -3235 6005 -3205
rect 6035 -3235 6085 -3205
rect 6115 -3235 6165 -3205
rect 6195 -3235 6245 -3205
rect 6275 -3235 6325 -3205
rect 6355 -3235 6405 -3205
rect 6435 -3235 6485 -3205
rect 6515 -3235 6565 -3205
rect 6595 -3235 6645 -3205
rect 6675 -3235 6725 -3205
rect 6755 -3235 6805 -3205
rect 6835 -3235 6885 -3205
rect 6915 -3235 6965 -3205
rect 6995 -3235 7045 -3205
rect 7075 -3235 7125 -3205
rect 7155 -3235 7205 -3205
rect 7235 -3235 7285 -3205
rect 7315 -3235 7365 -3205
rect 7395 -3235 7445 -3205
rect 7475 -3235 7525 -3205
rect 7555 -3235 7605 -3205
rect 7635 -3235 7685 -3205
rect 7715 -3235 7765 -3205
rect 7795 -3235 7845 -3205
rect 7875 -3235 7925 -3205
rect 7955 -3235 8005 -3205
rect 8035 -3235 8085 -3205
rect 8115 -3235 8165 -3205
rect 8195 -3235 8245 -3205
rect 8275 -3235 8325 -3205
rect 8355 -3235 8405 -3205
rect 8435 -3235 8485 -3205
rect 8515 -3235 8565 -3205
rect 8595 -3235 8645 -3205
rect 8675 -3235 8725 -3205
rect 8755 -3235 8805 -3205
rect 8835 -3235 8885 -3205
rect 8915 -3235 8965 -3205
rect 8995 -3235 9045 -3205
rect 9075 -3235 9125 -3205
rect 9155 -3235 9205 -3205
rect 9235 -3235 9285 -3205
rect 9315 -3235 9365 -3205
rect 9395 -3235 9445 -3205
rect 9475 -3235 9525 -3205
rect 9555 -3235 9605 -3205
rect 9635 -3235 9685 -3205
rect 9715 -3235 9765 -3205
rect 9795 -3235 9845 -3205
rect 9875 -3235 9925 -3205
rect 9955 -3235 10005 -3205
rect 10035 -3235 10085 -3205
rect 10115 -3235 10165 -3205
rect 10195 -3235 10245 -3205
rect 10275 -3235 10325 -3205
rect 10355 -3235 10405 -3205
rect 10435 -3235 10485 -3205
rect 10515 -3235 10645 -3205
rect 10675 -3235 10805 -3205
rect 10835 -3235 10965 -3205
rect 10995 -3235 11000 -3205
rect -720 -3240 11000 -3235
rect -720 -3285 11000 -3280
rect -720 -3315 -715 -3285
rect -685 -3315 -555 -3285
rect -525 -3315 -395 -3285
rect -365 -3315 -315 -3285
rect -285 -3315 -235 -3285
rect -205 -3315 -155 -3285
rect -125 -3315 -75 -3285
rect -45 -3315 5 -3285
rect 35 -3315 85 -3285
rect 115 -3315 165 -3285
rect 195 -3315 245 -3285
rect 275 -3315 325 -3285
rect 355 -3315 405 -3285
rect 435 -3315 485 -3285
rect 515 -3315 565 -3285
rect 595 -3315 645 -3285
rect 675 -3315 725 -3285
rect 755 -3315 805 -3285
rect 835 -3315 885 -3285
rect 915 -3315 965 -3285
rect 995 -3315 1045 -3285
rect 1075 -3315 1125 -3285
rect 1155 -3315 1205 -3285
rect 1235 -3315 1285 -3285
rect 1315 -3315 1365 -3285
rect 1395 -3315 1445 -3285
rect 1475 -3315 1525 -3285
rect 1555 -3315 1605 -3285
rect 1635 -3315 1685 -3285
rect 1715 -3315 1765 -3285
rect 1795 -3315 1845 -3285
rect 1875 -3315 1925 -3285
rect 1955 -3315 2005 -3285
rect 2035 -3315 2085 -3285
rect 2115 -3315 2165 -3285
rect 2195 -3315 2245 -3285
rect 2275 -3315 2325 -3285
rect 2355 -3315 2405 -3285
rect 2435 -3315 2485 -3285
rect 2515 -3315 2565 -3285
rect 2595 -3315 2645 -3285
rect 2675 -3315 2725 -3285
rect 2755 -3315 2805 -3285
rect 2835 -3315 2885 -3285
rect 2915 -3315 2965 -3285
rect 2995 -3315 3045 -3285
rect 3075 -3315 3125 -3285
rect 3155 -3315 3205 -3285
rect 3235 -3315 3285 -3285
rect 3315 -3315 3365 -3285
rect 3395 -3315 3445 -3285
rect 3475 -3315 3525 -3285
rect 3555 -3315 3605 -3285
rect 3635 -3315 3685 -3285
rect 3715 -3315 3765 -3285
rect 3795 -3315 3845 -3285
rect 3875 -3315 3925 -3285
rect 3955 -3315 4005 -3285
rect 4035 -3315 4085 -3285
rect 4115 -3315 4165 -3285
rect 4195 -3315 4245 -3285
rect 4275 -3315 4325 -3285
rect 4355 -3315 4405 -3285
rect 4435 -3315 4485 -3285
rect 4515 -3315 4565 -3285
rect 4595 -3315 4645 -3285
rect 4675 -3315 4725 -3285
rect 4755 -3315 4805 -3285
rect 4835 -3315 4885 -3285
rect 4915 -3315 4965 -3285
rect 4995 -3315 5045 -3285
rect 5075 -3315 5125 -3285
rect 5155 -3315 5205 -3285
rect 5235 -3315 5285 -3285
rect 5315 -3315 5365 -3285
rect 5395 -3315 5445 -3285
rect 5475 -3315 5525 -3285
rect 5555 -3315 5605 -3285
rect 5635 -3315 5685 -3285
rect 5715 -3315 5765 -3285
rect 5795 -3315 5845 -3285
rect 5875 -3315 5925 -3285
rect 5955 -3315 6005 -3285
rect 6035 -3315 6085 -3285
rect 6115 -3315 6165 -3285
rect 6195 -3315 6245 -3285
rect 6275 -3315 6325 -3285
rect 6355 -3315 6405 -3285
rect 6435 -3315 6485 -3285
rect 6515 -3315 6565 -3285
rect 6595 -3315 6645 -3285
rect 6675 -3315 6725 -3285
rect 6755 -3315 6805 -3285
rect 6835 -3315 6885 -3285
rect 6915 -3315 6965 -3285
rect 6995 -3315 7045 -3285
rect 7075 -3315 7125 -3285
rect 7155 -3315 7205 -3285
rect 7235 -3315 7285 -3285
rect 7315 -3315 7365 -3285
rect 7395 -3315 7445 -3285
rect 7475 -3315 7525 -3285
rect 7555 -3315 7605 -3285
rect 7635 -3315 7685 -3285
rect 7715 -3315 7765 -3285
rect 7795 -3315 7845 -3285
rect 7875 -3315 7925 -3285
rect 7955 -3315 8005 -3285
rect 8035 -3315 8085 -3285
rect 8115 -3315 8165 -3285
rect 8195 -3315 8245 -3285
rect 8275 -3315 8325 -3285
rect 8355 -3315 8405 -3285
rect 8435 -3315 8485 -3285
rect 8515 -3315 8565 -3285
rect 8595 -3315 8645 -3285
rect 8675 -3315 8725 -3285
rect 8755 -3315 8805 -3285
rect 8835 -3315 8885 -3285
rect 8915 -3315 8965 -3285
rect 8995 -3315 9045 -3285
rect 9075 -3315 9125 -3285
rect 9155 -3315 9205 -3285
rect 9235 -3315 9285 -3285
rect 9315 -3315 9365 -3285
rect 9395 -3315 9445 -3285
rect 9475 -3315 9525 -3285
rect 9555 -3315 9605 -3285
rect 9635 -3315 9685 -3285
rect 9715 -3315 9765 -3285
rect 9795 -3315 9845 -3285
rect 9875 -3315 9925 -3285
rect 9955 -3315 10005 -3285
rect 10035 -3315 10085 -3285
rect 10115 -3315 10165 -3285
rect 10195 -3315 10245 -3285
rect 10275 -3315 10325 -3285
rect 10355 -3315 10405 -3285
rect 10435 -3315 10485 -3285
rect 10515 -3315 10645 -3285
rect 10675 -3315 10805 -3285
rect 10835 -3315 10965 -3285
rect 10995 -3315 11000 -3285
rect -720 -3320 11000 -3315
rect -640 -3365 10600 -3360
rect -640 -3395 -635 -3365
rect -605 -3395 -75 -3365
rect -45 -3395 5205 -3365
rect 5235 -3395 5845 -3365
rect 5875 -3395 6485 -3365
rect 6515 -3395 7125 -3365
rect 7155 -3395 7765 -3365
rect 7795 -3395 8405 -3365
rect 8435 -3395 9045 -3365
rect 9075 -3395 9685 -3365
rect 9715 -3395 10325 -3365
rect 10355 -3395 10600 -3365
rect -640 -3400 10600 -3395
rect 10640 -3365 11000 -3360
rect 10640 -3395 10645 -3365
rect 10675 -3395 10805 -3365
rect 10835 -3395 10965 -3365
rect 10995 -3395 11000 -3365
rect 10640 -3400 11000 -3395
rect -640 -3445 10600 -3440
rect -640 -3475 -635 -3445
rect -605 -3475 -75 -3445
rect -45 -3475 5205 -3445
rect 5235 -3475 5845 -3445
rect 5875 -3475 6485 -3445
rect 6515 -3475 7125 -3445
rect 7155 -3475 7765 -3445
rect 7795 -3475 8405 -3445
rect 8435 -3475 9045 -3445
rect 9075 -3475 9685 -3445
rect 9715 -3475 10325 -3445
rect 10355 -3475 10600 -3445
rect -640 -3480 10600 -3475
rect 10640 -3445 11000 -3440
rect 10640 -3475 10645 -3445
rect 10675 -3475 10805 -3445
rect 10835 -3475 10965 -3445
rect 10995 -3475 11000 -3445
rect 10640 -3480 11000 -3475
rect -720 -3525 11000 -3520
rect -720 -3555 -715 -3525
rect -685 -3555 -555 -3525
rect -525 -3555 -395 -3525
rect -365 -3555 -315 -3525
rect -285 -3555 -235 -3525
rect -205 -3555 -155 -3525
rect -125 -3555 -75 -3525
rect -45 -3555 5 -3525
rect 35 -3555 85 -3525
rect 115 -3555 165 -3525
rect 195 -3555 245 -3525
rect 275 -3555 325 -3525
rect 355 -3555 405 -3525
rect 435 -3555 485 -3525
rect 515 -3555 565 -3525
rect 595 -3555 645 -3525
rect 675 -3555 725 -3525
rect 755 -3555 805 -3525
rect 835 -3555 885 -3525
rect 915 -3555 965 -3525
rect 995 -3555 1045 -3525
rect 1075 -3555 1125 -3525
rect 1155 -3555 1205 -3525
rect 1235 -3555 1285 -3525
rect 1315 -3555 1365 -3525
rect 1395 -3555 1445 -3525
rect 1475 -3555 1525 -3525
rect 1555 -3555 1605 -3525
rect 1635 -3555 1685 -3525
rect 1715 -3555 1765 -3525
rect 1795 -3555 1845 -3525
rect 1875 -3555 1925 -3525
rect 1955 -3555 2005 -3525
rect 2035 -3555 2085 -3525
rect 2115 -3555 2165 -3525
rect 2195 -3555 2245 -3525
rect 2275 -3555 2325 -3525
rect 2355 -3555 2405 -3525
rect 2435 -3555 2485 -3525
rect 2515 -3555 2565 -3525
rect 2595 -3555 2645 -3525
rect 2675 -3555 2725 -3525
rect 2755 -3555 2805 -3525
rect 2835 -3555 2885 -3525
rect 2915 -3555 2965 -3525
rect 2995 -3555 3045 -3525
rect 3075 -3555 3125 -3525
rect 3155 -3555 3205 -3525
rect 3235 -3555 3285 -3525
rect 3315 -3555 3365 -3525
rect 3395 -3555 3445 -3525
rect 3475 -3555 3525 -3525
rect 3555 -3555 3605 -3525
rect 3635 -3555 3685 -3525
rect 3715 -3555 3765 -3525
rect 3795 -3555 3845 -3525
rect 3875 -3555 3925 -3525
rect 3955 -3555 4005 -3525
rect 4035 -3555 4085 -3525
rect 4115 -3555 4165 -3525
rect 4195 -3555 4245 -3525
rect 4275 -3555 4325 -3525
rect 4355 -3555 4405 -3525
rect 4435 -3555 4485 -3525
rect 4515 -3555 4565 -3525
rect 4595 -3555 4645 -3525
rect 4675 -3555 4725 -3525
rect 4755 -3555 4805 -3525
rect 4835 -3555 4885 -3525
rect 4915 -3555 4965 -3525
rect 4995 -3555 5045 -3525
rect 5075 -3555 5125 -3525
rect 5155 -3555 5205 -3525
rect 5235 -3555 5285 -3525
rect 5315 -3555 5365 -3525
rect 5395 -3555 5445 -3525
rect 5475 -3555 5525 -3525
rect 5555 -3555 5605 -3525
rect 5635 -3555 5685 -3525
rect 5715 -3555 5765 -3525
rect 5795 -3555 5845 -3525
rect 5875 -3555 5925 -3525
rect 5955 -3555 6005 -3525
rect 6035 -3555 6085 -3525
rect 6115 -3555 6165 -3525
rect 6195 -3555 6245 -3525
rect 6275 -3555 6325 -3525
rect 6355 -3555 6405 -3525
rect 6435 -3555 6485 -3525
rect 6515 -3555 6565 -3525
rect 6595 -3555 6645 -3525
rect 6675 -3555 6725 -3525
rect 6755 -3555 6805 -3525
rect 6835 -3555 6885 -3525
rect 6915 -3555 6965 -3525
rect 6995 -3555 7045 -3525
rect 7075 -3555 7125 -3525
rect 7155 -3555 7205 -3525
rect 7235 -3555 7285 -3525
rect 7315 -3555 7365 -3525
rect 7395 -3555 7445 -3525
rect 7475 -3555 7525 -3525
rect 7555 -3555 7605 -3525
rect 7635 -3555 7685 -3525
rect 7715 -3555 7765 -3525
rect 7795 -3555 7845 -3525
rect 7875 -3555 7925 -3525
rect 7955 -3555 8005 -3525
rect 8035 -3555 8085 -3525
rect 8115 -3555 8165 -3525
rect 8195 -3555 8245 -3525
rect 8275 -3555 8325 -3525
rect 8355 -3555 8405 -3525
rect 8435 -3555 8485 -3525
rect 8515 -3555 8565 -3525
rect 8595 -3555 8645 -3525
rect 8675 -3555 8725 -3525
rect 8755 -3555 8805 -3525
rect 8835 -3555 8885 -3525
rect 8915 -3555 8965 -3525
rect 8995 -3555 9045 -3525
rect 9075 -3555 9125 -3525
rect 9155 -3555 9205 -3525
rect 9235 -3555 9285 -3525
rect 9315 -3555 9365 -3525
rect 9395 -3555 9445 -3525
rect 9475 -3555 9525 -3525
rect 9555 -3555 9605 -3525
rect 9635 -3555 9685 -3525
rect 9715 -3555 9765 -3525
rect 9795 -3555 9845 -3525
rect 9875 -3555 9925 -3525
rect 9955 -3555 10005 -3525
rect 10035 -3555 10085 -3525
rect 10115 -3555 10165 -3525
rect 10195 -3555 10245 -3525
rect 10275 -3555 10325 -3525
rect 10355 -3555 10405 -3525
rect 10435 -3555 10485 -3525
rect 10515 -3555 10645 -3525
rect 10675 -3555 10805 -3525
rect 10835 -3555 10965 -3525
rect 10995 -3555 11000 -3525
rect -720 -3560 11000 -3555
rect -720 -3605 11000 -3600
rect -720 -3635 -715 -3605
rect -685 -3635 -555 -3605
rect -525 -3635 -395 -3605
rect -365 -3635 -315 -3605
rect -285 -3635 -235 -3605
rect -205 -3635 -155 -3605
rect -125 -3635 -75 -3605
rect -45 -3635 5 -3605
rect 35 -3635 85 -3605
rect 115 -3635 165 -3605
rect 195 -3635 245 -3605
rect 275 -3635 325 -3605
rect 355 -3635 405 -3605
rect 435 -3635 485 -3605
rect 515 -3635 565 -3605
rect 595 -3635 645 -3605
rect 675 -3635 725 -3605
rect 755 -3635 805 -3605
rect 835 -3635 885 -3605
rect 915 -3635 965 -3605
rect 995 -3635 1045 -3605
rect 1075 -3635 1125 -3605
rect 1155 -3635 1205 -3605
rect 1235 -3635 1285 -3605
rect 1315 -3635 1365 -3605
rect 1395 -3635 1445 -3605
rect 1475 -3635 1525 -3605
rect 1555 -3635 1605 -3605
rect 1635 -3635 1685 -3605
rect 1715 -3635 1765 -3605
rect 1795 -3635 1845 -3605
rect 1875 -3635 1925 -3605
rect 1955 -3635 2005 -3605
rect 2035 -3635 2085 -3605
rect 2115 -3635 2165 -3605
rect 2195 -3635 2245 -3605
rect 2275 -3635 2325 -3605
rect 2355 -3635 2405 -3605
rect 2435 -3635 2485 -3605
rect 2515 -3635 2565 -3605
rect 2595 -3635 2645 -3605
rect 2675 -3635 2725 -3605
rect 2755 -3635 2805 -3605
rect 2835 -3635 2885 -3605
rect 2915 -3635 2965 -3605
rect 2995 -3635 3045 -3605
rect 3075 -3635 3125 -3605
rect 3155 -3635 3205 -3605
rect 3235 -3635 3285 -3605
rect 3315 -3635 3365 -3605
rect 3395 -3635 3445 -3605
rect 3475 -3635 3525 -3605
rect 3555 -3635 3605 -3605
rect 3635 -3635 3685 -3605
rect 3715 -3635 3765 -3605
rect 3795 -3635 3845 -3605
rect 3875 -3635 3925 -3605
rect 3955 -3635 4005 -3605
rect 4035 -3635 4085 -3605
rect 4115 -3635 4165 -3605
rect 4195 -3635 4245 -3605
rect 4275 -3635 4325 -3605
rect 4355 -3635 4405 -3605
rect 4435 -3635 4485 -3605
rect 4515 -3635 4565 -3605
rect 4595 -3635 4645 -3605
rect 4675 -3635 4725 -3605
rect 4755 -3635 4805 -3605
rect 4835 -3635 4885 -3605
rect 4915 -3635 4965 -3605
rect 4995 -3635 5045 -3605
rect 5075 -3635 5125 -3605
rect 5155 -3635 5205 -3605
rect 5235 -3635 5285 -3605
rect 5315 -3635 5365 -3605
rect 5395 -3635 5445 -3605
rect 5475 -3635 5525 -3605
rect 5555 -3635 5605 -3605
rect 5635 -3635 5685 -3605
rect 5715 -3635 5765 -3605
rect 5795 -3635 5845 -3605
rect 5875 -3635 5925 -3605
rect 5955 -3635 6005 -3605
rect 6035 -3635 6085 -3605
rect 6115 -3635 6165 -3605
rect 6195 -3635 6245 -3605
rect 6275 -3635 6325 -3605
rect 6355 -3635 6405 -3605
rect 6435 -3635 6485 -3605
rect 6515 -3635 6565 -3605
rect 6595 -3635 6645 -3605
rect 6675 -3635 6725 -3605
rect 6755 -3635 6805 -3605
rect 6835 -3635 6885 -3605
rect 6915 -3635 6965 -3605
rect 6995 -3635 7045 -3605
rect 7075 -3635 7125 -3605
rect 7155 -3635 7205 -3605
rect 7235 -3635 7285 -3605
rect 7315 -3635 7365 -3605
rect 7395 -3635 7445 -3605
rect 7475 -3635 7525 -3605
rect 7555 -3635 7605 -3605
rect 7635 -3635 7685 -3605
rect 7715 -3635 7765 -3605
rect 7795 -3635 7845 -3605
rect 7875 -3635 7925 -3605
rect 7955 -3635 8005 -3605
rect 8035 -3635 8085 -3605
rect 8115 -3635 8165 -3605
rect 8195 -3635 8245 -3605
rect 8275 -3635 8325 -3605
rect 8355 -3635 8405 -3605
rect 8435 -3635 8485 -3605
rect 8515 -3635 8565 -3605
rect 8595 -3635 8645 -3605
rect 8675 -3635 8725 -3605
rect 8755 -3635 8805 -3605
rect 8835 -3635 8885 -3605
rect 8915 -3635 8965 -3605
rect 8995 -3635 9045 -3605
rect 9075 -3635 9125 -3605
rect 9155 -3635 9205 -3605
rect 9235 -3635 9285 -3605
rect 9315 -3635 9365 -3605
rect 9395 -3635 9445 -3605
rect 9475 -3635 9525 -3605
rect 9555 -3635 9605 -3605
rect 9635 -3635 9685 -3605
rect 9715 -3635 9765 -3605
rect 9795 -3635 9845 -3605
rect 9875 -3635 9925 -3605
rect 9955 -3635 10005 -3605
rect 10035 -3635 10085 -3605
rect 10115 -3635 10165 -3605
rect 10195 -3635 10245 -3605
rect 10275 -3635 10325 -3605
rect 10355 -3635 10405 -3605
rect 10435 -3635 10485 -3605
rect 10515 -3635 10645 -3605
rect 10675 -3635 10805 -3605
rect 10835 -3635 10965 -3605
rect 10995 -3635 11000 -3605
rect -720 -3640 11000 -3635
rect -720 -3685 11000 -3680
rect -720 -3715 -715 -3685
rect -685 -3715 -555 -3685
rect -525 -3715 -395 -3685
rect -365 -3715 -315 -3685
rect -285 -3715 -235 -3685
rect -205 -3715 -155 -3685
rect -125 -3715 -75 -3685
rect -45 -3715 5 -3685
rect 35 -3715 85 -3685
rect 115 -3715 165 -3685
rect 195 -3715 245 -3685
rect 275 -3715 325 -3685
rect 355 -3715 405 -3685
rect 435 -3715 485 -3685
rect 515 -3715 565 -3685
rect 595 -3715 645 -3685
rect 675 -3715 725 -3685
rect 755 -3715 805 -3685
rect 835 -3715 885 -3685
rect 915 -3715 965 -3685
rect 995 -3715 1045 -3685
rect 1075 -3715 1125 -3685
rect 1155 -3715 1205 -3685
rect 1235 -3715 1285 -3685
rect 1315 -3715 1365 -3685
rect 1395 -3715 1445 -3685
rect 1475 -3715 1525 -3685
rect 1555 -3715 1605 -3685
rect 1635 -3715 1685 -3685
rect 1715 -3715 1765 -3685
rect 1795 -3715 1845 -3685
rect 1875 -3715 1925 -3685
rect 1955 -3715 2005 -3685
rect 2035 -3715 2085 -3685
rect 2115 -3715 2165 -3685
rect 2195 -3715 2245 -3685
rect 2275 -3715 2325 -3685
rect 2355 -3715 2405 -3685
rect 2435 -3715 2485 -3685
rect 2515 -3715 2565 -3685
rect 2595 -3715 2645 -3685
rect 2675 -3715 2725 -3685
rect 2755 -3715 2805 -3685
rect 2835 -3715 2885 -3685
rect 2915 -3715 2965 -3685
rect 2995 -3715 3045 -3685
rect 3075 -3715 3125 -3685
rect 3155 -3715 3205 -3685
rect 3235 -3715 3285 -3685
rect 3315 -3715 3365 -3685
rect 3395 -3715 3445 -3685
rect 3475 -3715 3525 -3685
rect 3555 -3715 3605 -3685
rect 3635 -3715 3685 -3685
rect 3715 -3715 3765 -3685
rect 3795 -3715 3845 -3685
rect 3875 -3715 3925 -3685
rect 3955 -3715 4005 -3685
rect 4035 -3715 4085 -3685
rect 4115 -3715 4165 -3685
rect 4195 -3715 4245 -3685
rect 4275 -3715 4325 -3685
rect 4355 -3715 4405 -3685
rect 4435 -3715 4485 -3685
rect 4515 -3715 4565 -3685
rect 4595 -3715 4645 -3685
rect 4675 -3715 4725 -3685
rect 4755 -3715 4805 -3685
rect 4835 -3715 4885 -3685
rect 4915 -3715 4965 -3685
rect 4995 -3715 5045 -3685
rect 5075 -3715 5125 -3685
rect 5155 -3715 5205 -3685
rect 5235 -3715 5285 -3685
rect 5315 -3715 5365 -3685
rect 5395 -3715 5445 -3685
rect 5475 -3715 5525 -3685
rect 5555 -3715 5605 -3685
rect 5635 -3715 5685 -3685
rect 5715 -3715 5765 -3685
rect 5795 -3715 5845 -3685
rect 5875 -3715 5925 -3685
rect 5955 -3715 6005 -3685
rect 6035 -3715 6085 -3685
rect 6115 -3715 6165 -3685
rect 6195 -3715 6245 -3685
rect 6275 -3715 6325 -3685
rect 6355 -3715 6405 -3685
rect 6435 -3715 6485 -3685
rect 6515 -3715 6565 -3685
rect 6595 -3715 6645 -3685
rect 6675 -3715 6725 -3685
rect 6755 -3715 6805 -3685
rect 6835 -3715 6885 -3685
rect 6915 -3715 6965 -3685
rect 6995 -3715 7045 -3685
rect 7075 -3715 7125 -3685
rect 7155 -3715 7205 -3685
rect 7235 -3715 7285 -3685
rect 7315 -3715 7365 -3685
rect 7395 -3715 7445 -3685
rect 7475 -3715 7525 -3685
rect 7555 -3715 7605 -3685
rect 7635 -3715 7685 -3685
rect 7715 -3715 7765 -3685
rect 7795 -3715 7845 -3685
rect 7875 -3715 7925 -3685
rect 7955 -3715 8005 -3685
rect 8035 -3715 8085 -3685
rect 8115 -3715 8165 -3685
rect 8195 -3715 8245 -3685
rect 8275 -3715 8325 -3685
rect 8355 -3715 8405 -3685
rect 8435 -3715 8485 -3685
rect 8515 -3715 8565 -3685
rect 8595 -3715 8645 -3685
rect 8675 -3715 8725 -3685
rect 8755 -3715 8805 -3685
rect 8835 -3715 8885 -3685
rect 8915 -3715 8965 -3685
rect 8995 -3715 9045 -3685
rect 9075 -3715 9125 -3685
rect 9155 -3715 9205 -3685
rect 9235 -3715 9285 -3685
rect 9315 -3715 9365 -3685
rect 9395 -3715 9445 -3685
rect 9475 -3715 9525 -3685
rect 9555 -3715 9605 -3685
rect 9635 -3715 9685 -3685
rect 9715 -3715 9765 -3685
rect 9795 -3715 9845 -3685
rect 9875 -3715 9925 -3685
rect 9955 -3715 10005 -3685
rect 10035 -3715 10085 -3685
rect 10115 -3715 10165 -3685
rect 10195 -3715 10245 -3685
rect 10275 -3715 10325 -3685
rect 10355 -3715 10405 -3685
rect 10435 -3715 10485 -3685
rect 10515 -3715 10645 -3685
rect 10675 -3715 10805 -3685
rect 10835 -3715 10965 -3685
rect 10995 -3715 11000 -3685
rect -720 -3720 11000 -3715
<< via2 >>
rect -715 1005 -685 1035
rect -555 1005 -525 1035
rect -395 1005 -365 1035
rect -315 1005 -285 1035
rect -235 1005 -205 1035
rect -155 1005 -125 1035
rect -75 1005 -45 1035
rect 5 1005 35 1035
rect 85 1005 115 1035
rect 165 1005 195 1035
rect 245 1005 275 1035
rect 325 1005 355 1035
rect 405 1005 435 1035
rect 485 1005 515 1035
rect 565 1005 595 1035
rect 645 1005 675 1035
rect 725 1005 755 1035
rect 805 1005 835 1035
rect 885 1005 915 1035
rect 965 1005 995 1035
rect 1045 1005 1075 1035
rect 1125 1005 1155 1035
rect 1205 1005 1235 1035
rect 1285 1005 1315 1035
rect 1365 1005 1395 1035
rect 1445 1005 1475 1035
rect 1525 1005 1555 1035
rect 1605 1005 1635 1035
rect 1685 1005 1715 1035
rect 1765 1005 1795 1035
rect 1845 1005 1875 1035
rect 1925 1005 1955 1035
rect 2005 1005 2035 1035
rect 2085 1005 2115 1035
rect 2165 1005 2195 1035
rect 2245 1005 2275 1035
rect 2325 1005 2355 1035
rect 2405 1005 2435 1035
rect 2485 1005 2515 1035
rect 2565 1005 2595 1035
rect 2645 1005 2675 1035
rect 2725 1005 2755 1035
rect 2805 1005 2835 1035
rect 2885 1005 2915 1035
rect 2965 1005 2995 1035
rect 3045 1005 3075 1035
rect 3125 1005 3155 1035
rect 3205 1005 3235 1035
rect 3285 1005 3315 1035
rect 3365 1005 3395 1035
rect 3445 1005 3475 1035
rect 3525 1005 3555 1035
rect 3605 1005 3635 1035
rect 3685 1005 3715 1035
rect 3765 1005 3795 1035
rect 3845 1005 3875 1035
rect 3925 1005 3955 1035
rect 4005 1005 4035 1035
rect 4085 1005 4115 1035
rect 4165 1005 4195 1035
rect 4245 1005 4275 1035
rect 4325 1005 4355 1035
rect 4405 1005 4435 1035
rect 4485 1005 4515 1035
rect 4565 1005 4595 1035
rect 4645 1005 4675 1035
rect 4725 1005 4755 1035
rect 4805 1005 4835 1035
rect 4885 1005 4915 1035
rect 4965 1005 4995 1035
rect 5045 1005 5075 1035
rect 5125 1005 5155 1035
rect 5205 1005 5235 1035
rect 5285 1005 5315 1035
rect 5365 1005 5395 1035
rect 5445 1005 5475 1035
rect 5525 1005 5555 1035
rect 5605 1005 5635 1035
rect 5685 1005 5715 1035
rect 5765 1005 5795 1035
rect 5845 1005 5875 1035
rect 5925 1005 5955 1035
rect 6005 1005 6035 1035
rect 6085 1005 6115 1035
rect 6165 1005 6195 1035
rect 6245 1005 6275 1035
rect 6325 1005 6355 1035
rect 6405 1005 6435 1035
rect 6485 1005 6515 1035
rect 6565 1005 6595 1035
rect 6645 1005 6675 1035
rect 6725 1005 6755 1035
rect 6805 1005 6835 1035
rect 6885 1005 6915 1035
rect 6965 1005 6995 1035
rect 7045 1005 7075 1035
rect 7125 1005 7155 1035
rect 7205 1005 7235 1035
rect 7285 1005 7315 1035
rect 7365 1005 7395 1035
rect 7445 1005 7475 1035
rect 7525 1005 7555 1035
rect 7605 1005 7635 1035
rect 7685 1005 7715 1035
rect 7765 1005 7795 1035
rect 7845 1005 7875 1035
rect 7925 1005 7955 1035
rect 8005 1005 8035 1035
rect 8085 1005 8115 1035
rect 8165 1005 8195 1035
rect 8245 1005 8275 1035
rect 8325 1005 8355 1035
rect 8405 1005 8435 1035
rect 8485 1005 8515 1035
rect 8565 1005 8595 1035
rect 8645 1005 8675 1035
rect 8725 1005 8755 1035
rect 8805 1005 8835 1035
rect 8885 1005 8915 1035
rect 8965 1005 8995 1035
rect 9045 1005 9075 1035
rect 9125 1005 9155 1035
rect 9205 1005 9235 1035
rect 9285 1005 9315 1035
rect 9365 1005 9395 1035
rect 9445 1005 9475 1035
rect 9525 1005 9555 1035
rect 9605 1005 9635 1035
rect 9685 1005 9715 1035
rect 9765 1005 9795 1035
rect 9845 1005 9875 1035
rect 9925 1005 9955 1035
rect 10005 1005 10035 1035
rect 10085 1005 10115 1035
rect 10165 1005 10195 1035
rect 10245 1005 10275 1035
rect 10325 1005 10355 1035
rect 10405 1005 10435 1035
rect 10485 1005 10515 1035
rect 10645 1005 10675 1035
rect 10805 1005 10835 1035
rect 10965 1005 10995 1035
rect -715 925 -685 955
rect -555 925 -525 955
rect -395 925 -365 955
rect -315 925 -285 955
rect -235 925 -205 955
rect -155 925 -125 955
rect -75 925 -45 955
rect 5 925 35 955
rect 85 925 115 955
rect 165 925 195 955
rect 245 925 275 955
rect 325 925 355 955
rect 405 925 435 955
rect 485 925 515 955
rect 565 925 595 955
rect 645 925 675 955
rect 725 925 755 955
rect 805 925 835 955
rect 885 925 915 955
rect 965 925 995 955
rect 1045 925 1075 955
rect 1125 925 1155 955
rect 1205 925 1235 955
rect 1285 925 1315 955
rect 1365 925 1395 955
rect 1445 925 1475 955
rect 1525 925 1555 955
rect 1605 925 1635 955
rect 1685 925 1715 955
rect 1765 925 1795 955
rect 1845 925 1875 955
rect 1925 925 1955 955
rect 2005 925 2035 955
rect 2085 925 2115 955
rect 2165 925 2195 955
rect 2245 925 2275 955
rect 2325 925 2355 955
rect 2405 925 2435 955
rect 2485 925 2515 955
rect 2565 925 2595 955
rect 2645 925 2675 955
rect 2725 925 2755 955
rect 2805 925 2835 955
rect 2885 925 2915 955
rect 2965 925 2995 955
rect 3045 925 3075 955
rect 3125 925 3155 955
rect 3205 925 3235 955
rect 3285 925 3315 955
rect 3365 925 3395 955
rect 3445 925 3475 955
rect 3525 925 3555 955
rect 3605 925 3635 955
rect 3685 925 3715 955
rect 3765 925 3795 955
rect 3845 925 3875 955
rect 3925 925 3955 955
rect 4005 925 4035 955
rect 4085 925 4115 955
rect 4165 925 4195 955
rect 4245 925 4275 955
rect 4325 925 4355 955
rect 4405 925 4435 955
rect 4485 925 4515 955
rect 4565 925 4595 955
rect 4645 925 4675 955
rect 4725 925 4755 955
rect 4805 925 4835 955
rect 4885 925 4915 955
rect 4965 925 4995 955
rect 5045 925 5075 955
rect 5125 925 5155 955
rect 5205 925 5235 955
rect 5285 925 5315 955
rect 5365 925 5395 955
rect 5445 925 5475 955
rect 5525 925 5555 955
rect 5605 925 5635 955
rect 5685 925 5715 955
rect 5765 925 5795 955
rect 5845 925 5875 955
rect 5925 925 5955 955
rect 6005 925 6035 955
rect 6085 925 6115 955
rect 6165 925 6195 955
rect 6245 925 6275 955
rect 6325 925 6355 955
rect 6405 925 6435 955
rect 6485 925 6515 955
rect 6565 925 6595 955
rect 6645 925 6675 955
rect 6725 925 6755 955
rect 6805 925 6835 955
rect 6885 925 6915 955
rect 6965 925 6995 955
rect 7045 925 7075 955
rect 7125 925 7155 955
rect 7205 925 7235 955
rect 7285 925 7315 955
rect 7365 925 7395 955
rect 7445 925 7475 955
rect 7525 925 7555 955
rect 7605 925 7635 955
rect 7685 925 7715 955
rect 7765 925 7795 955
rect 7845 925 7875 955
rect 7925 925 7955 955
rect 8005 925 8035 955
rect 8085 925 8115 955
rect 8165 925 8195 955
rect 8245 925 8275 955
rect 8325 925 8355 955
rect 8405 925 8435 955
rect 8485 925 8515 955
rect 8565 925 8595 955
rect 8645 925 8675 955
rect 8725 925 8755 955
rect 8805 925 8835 955
rect 8885 925 8915 955
rect 8965 925 8995 955
rect 9045 925 9075 955
rect 9125 925 9155 955
rect 9205 925 9235 955
rect 9285 925 9315 955
rect 9365 925 9395 955
rect 9445 925 9475 955
rect 9525 925 9555 955
rect 9605 925 9635 955
rect 9685 925 9715 955
rect 9765 925 9795 955
rect 9845 925 9875 955
rect 9925 925 9955 955
rect 10005 925 10035 955
rect 10085 925 10115 955
rect 10165 925 10195 955
rect 10245 925 10275 955
rect 10325 925 10355 955
rect 10405 925 10435 955
rect 10485 925 10515 955
rect 10645 925 10675 955
rect 10805 925 10835 955
rect 10965 925 10995 955
rect -715 845 -685 875
rect -555 845 -525 875
rect -395 845 -365 875
rect -315 845 -285 875
rect -235 845 -205 875
rect -155 845 -125 875
rect -75 845 -45 875
rect 5 845 35 875
rect 85 845 115 875
rect 165 845 195 875
rect 245 845 275 875
rect 325 845 355 875
rect 405 845 435 875
rect 485 845 515 875
rect 565 845 595 875
rect 645 845 675 875
rect 725 845 755 875
rect 805 845 835 875
rect 885 845 915 875
rect 965 845 995 875
rect 1045 845 1075 875
rect 1125 845 1155 875
rect 1205 845 1235 875
rect 1285 845 1315 875
rect 1365 845 1395 875
rect 1445 845 1475 875
rect 1525 845 1555 875
rect 1605 845 1635 875
rect 1685 845 1715 875
rect 1765 845 1795 875
rect 1845 845 1875 875
rect 1925 845 1955 875
rect 2005 845 2035 875
rect 2085 845 2115 875
rect 2165 845 2195 875
rect 2245 845 2275 875
rect 2325 845 2355 875
rect 2405 845 2435 875
rect 2485 845 2515 875
rect 2565 845 2595 875
rect 2645 845 2675 875
rect 2725 845 2755 875
rect 2805 845 2835 875
rect 2885 845 2915 875
rect 2965 845 2995 875
rect 3045 845 3075 875
rect 3125 845 3155 875
rect 3205 845 3235 875
rect 3285 845 3315 875
rect 3365 845 3395 875
rect 3445 845 3475 875
rect 3525 845 3555 875
rect 3605 845 3635 875
rect 3685 845 3715 875
rect 3765 845 3795 875
rect 3845 845 3875 875
rect 3925 845 3955 875
rect 4005 845 4035 875
rect 4085 845 4115 875
rect 4165 845 4195 875
rect 4245 845 4275 875
rect 4325 845 4355 875
rect 4405 845 4435 875
rect 4485 845 4515 875
rect 4565 845 4595 875
rect 4645 845 4675 875
rect 4725 845 4755 875
rect 4805 845 4835 875
rect 4885 845 4915 875
rect 4965 845 4995 875
rect 5045 845 5075 875
rect 5125 845 5155 875
rect 5205 845 5235 875
rect 5285 845 5315 875
rect 5365 845 5395 875
rect 5445 845 5475 875
rect 5525 845 5555 875
rect 5605 845 5635 875
rect 5685 845 5715 875
rect 5765 845 5795 875
rect 5845 845 5875 875
rect 5925 845 5955 875
rect 6005 845 6035 875
rect 6085 845 6115 875
rect 6165 845 6195 875
rect 6245 845 6275 875
rect 6325 845 6355 875
rect 6405 845 6435 875
rect 6485 845 6515 875
rect 6565 845 6595 875
rect 6645 845 6675 875
rect 6725 845 6755 875
rect 6805 845 6835 875
rect 6885 845 6915 875
rect 6965 845 6995 875
rect 7045 845 7075 875
rect 7125 845 7155 875
rect 7205 845 7235 875
rect 7285 845 7315 875
rect 7365 845 7395 875
rect 7445 845 7475 875
rect 7525 845 7555 875
rect 7605 845 7635 875
rect 7685 845 7715 875
rect 7765 845 7795 875
rect 7845 845 7875 875
rect 7925 845 7955 875
rect 8005 845 8035 875
rect 8085 845 8115 875
rect 8165 845 8195 875
rect 8245 845 8275 875
rect 8325 845 8355 875
rect 8405 845 8435 875
rect 8485 845 8515 875
rect 8565 845 8595 875
rect 8645 845 8675 875
rect 8725 845 8755 875
rect 8805 845 8835 875
rect 8885 845 8915 875
rect 8965 845 8995 875
rect 9045 845 9075 875
rect 9125 845 9155 875
rect 9205 845 9235 875
rect 9285 845 9315 875
rect 9365 845 9395 875
rect 9445 845 9475 875
rect 9525 845 9555 875
rect 9605 845 9635 875
rect 9685 845 9715 875
rect 9765 845 9795 875
rect 9845 845 9875 875
rect 9925 845 9955 875
rect 10005 845 10035 875
rect 10085 845 10115 875
rect 10165 845 10195 875
rect 10245 845 10275 875
rect 10325 845 10355 875
rect 10405 845 10435 875
rect 10485 845 10515 875
rect 10645 845 10675 875
rect 10805 845 10835 875
rect 10965 845 10995 875
rect -635 765 -605 795
rect 10645 765 10675 795
rect 10805 765 10835 795
rect 10965 765 10995 795
rect -635 685 -605 715
rect 10645 685 10675 715
rect 10805 685 10835 715
rect 10965 685 10995 715
rect -715 605 -685 635
rect -555 605 -525 635
rect -395 605 -365 635
rect -315 605 -285 635
rect -235 605 -205 635
rect -155 605 -125 635
rect -75 605 -45 635
rect 5 605 35 635
rect 85 605 115 635
rect 165 605 195 635
rect 245 605 275 635
rect 325 605 355 635
rect 405 605 435 635
rect 485 605 515 635
rect 565 605 595 635
rect 645 605 675 635
rect 725 605 755 635
rect 805 605 835 635
rect 885 605 915 635
rect 965 605 995 635
rect 1045 605 1075 635
rect 1125 605 1155 635
rect 1205 605 1235 635
rect 1285 605 1315 635
rect 1365 605 1395 635
rect 1445 605 1475 635
rect 1525 605 1555 635
rect 1605 605 1635 635
rect 1685 605 1715 635
rect 1765 605 1795 635
rect 1845 605 1875 635
rect 1925 605 1955 635
rect 2005 605 2035 635
rect 2085 605 2115 635
rect 2165 605 2195 635
rect 2245 605 2275 635
rect 2325 605 2355 635
rect 2405 605 2435 635
rect 2485 605 2515 635
rect 2565 605 2595 635
rect 2645 605 2675 635
rect 2725 605 2755 635
rect 2805 605 2835 635
rect 2885 605 2915 635
rect 2965 605 2995 635
rect 3045 605 3075 635
rect 3125 605 3155 635
rect 3205 605 3235 635
rect 3285 605 3315 635
rect 3365 605 3395 635
rect 3445 605 3475 635
rect 3525 605 3555 635
rect 3605 605 3635 635
rect 3685 605 3715 635
rect 3765 605 3795 635
rect 3845 605 3875 635
rect 3925 605 3955 635
rect 4005 605 4035 635
rect 4085 605 4115 635
rect 4165 605 4195 635
rect 4245 605 4275 635
rect 4325 605 4355 635
rect 4405 605 4435 635
rect 4485 605 4515 635
rect 4565 605 4595 635
rect 4645 605 4675 635
rect 4725 605 4755 635
rect 4805 605 4835 635
rect 4885 605 4915 635
rect 4965 605 4995 635
rect 5045 605 5075 635
rect 5125 605 5155 635
rect 5205 605 5235 635
rect 5285 605 5315 635
rect 5365 605 5395 635
rect 5445 605 5475 635
rect 5525 605 5555 635
rect 5605 605 5635 635
rect 5685 605 5715 635
rect 5765 605 5795 635
rect 5845 605 5875 635
rect 5925 605 5955 635
rect 6005 605 6035 635
rect 6085 605 6115 635
rect 6165 605 6195 635
rect 6245 605 6275 635
rect 6325 605 6355 635
rect 6405 605 6435 635
rect 6485 605 6515 635
rect 6565 605 6595 635
rect 6645 605 6675 635
rect 6725 605 6755 635
rect 6805 605 6835 635
rect 6885 605 6915 635
rect 6965 605 6995 635
rect 7045 605 7075 635
rect 7125 605 7155 635
rect 7205 605 7235 635
rect 7285 605 7315 635
rect 7365 605 7395 635
rect 7445 605 7475 635
rect 7525 605 7555 635
rect 7605 605 7635 635
rect 7685 605 7715 635
rect 7765 605 7795 635
rect 7845 605 7875 635
rect 7925 605 7955 635
rect 8005 605 8035 635
rect 8085 605 8115 635
rect 8165 605 8195 635
rect 8245 605 8275 635
rect 8325 605 8355 635
rect 8405 605 8435 635
rect 8485 605 8515 635
rect 8565 605 8595 635
rect 8645 605 8675 635
rect 8725 605 8755 635
rect 8805 605 8835 635
rect 8885 605 8915 635
rect 8965 605 8995 635
rect 9045 605 9075 635
rect 9125 605 9155 635
rect 9205 605 9235 635
rect 9285 605 9315 635
rect 9365 605 9395 635
rect 9445 605 9475 635
rect 9525 605 9555 635
rect 9605 605 9635 635
rect 9685 605 9715 635
rect 9765 605 9795 635
rect 9845 605 9875 635
rect 9925 605 9955 635
rect 10005 605 10035 635
rect 10085 605 10115 635
rect 10165 605 10195 635
rect 10245 605 10275 635
rect 10325 605 10355 635
rect 10405 605 10435 635
rect 10485 605 10515 635
rect 10645 605 10675 635
rect 10805 605 10835 635
rect 10965 605 10995 635
rect -715 525 -685 555
rect -555 525 -525 555
rect -395 525 -365 555
rect -315 525 -285 555
rect -235 525 -205 555
rect -155 525 -125 555
rect -75 525 -45 555
rect 5 525 35 555
rect 85 525 115 555
rect 165 525 195 555
rect 245 525 275 555
rect 325 525 355 555
rect 405 525 435 555
rect 485 525 515 555
rect 565 525 595 555
rect 645 525 675 555
rect 725 525 755 555
rect 805 525 835 555
rect 885 525 915 555
rect 965 525 995 555
rect 1045 525 1075 555
rect 1125 525 1155 555
rect 1205 525 1235 555
rect 1285 525 1315 555
rect 1365 525 1395 555
rect 1445 525 1475 555
rect 1525 525 1555 555
rect 1605 525 1635 555
rect 1685 525 1715 555
rect 1765 525 1795 555
rect 1845 525 1875 555
rect 1925 525 1955 555
rect 2005 525 2035 555
rect 2085 525 2115 555
rect 2165 525 2195 555
rect 2245 525 2275 555
rect 2325 525 2355 555
rect 2405 525 2435 555
rect 2485 525 2515 555
rect 2565 525 2595 555
rect 2645 525 2675 555
rect 2725 525 2755 555
rect 2805 525 2835 555
rect 2885 525 2915 555
rect 2965 525 2995 555
rect 3045 525 3075 555
rect 3125 525 3155 555
rect 3205 525 3235 555
rect 3285 525 3315 555
rect 3365 525 3395 555
rect 3445 525 3475 555
rect 3525 525 3555 555
rect 3605 525 3635 555
rect 3685 525 3715 555
rect 3765 525 3795 555
rect 3845 525 3875 555
rect 3925 525 3955 555
rect 4005 525 4035 555
rect 4085 525 4115 555
rect 4165 525 4195 555
rect 4245 525 4275 555
rect 4325 525 4355 555
rect 4405 525 4435 555
rect 4485 525 4515 555
rect 4565 525 4595 555
rect 4645 525 4675 555
rect 4725 525 4755 555
rect 4805 525 4835 555
rect 4885 525 4915 555
rect 4965 525 4995 555
rect 5045 525 5075 555
rect 5125 525 5155 555
rect 5205 525 5235 555
rect 5285 525 5315 555
rect 5365 525 5395 555
rect 5445 525 5475 555
rect 5525 525 5555 555
rect 5605 525 5635 555
rect 5685 525 5715 555
rect 5765 525 5795 555
rect 5845 525 5875 555
rect 5925 525 5955 555
rect 6005 525 6035 555
rect 6085 525 6115 555
rect 6165 525 6195 555
rect 6245 525 6275 555
rect 6325 525 6355 555
rect 6405 525 6435 555
rect 6485 525 6515 555
rect 6565 525 6595 555
rect 6645 525 6675 555
rect 6725 525 6755 555
rect 6805 525 6835 555
rect 6885 525 6915 555
rect 6965 525 6995 555
rect 7045 525 7075 555
rect 7125 525 7155 555
rect 7205 525 7235 555
rect 7285 525 7315 555
rect 7365 525 7395 555
rect 7445 525 7475 555
rect 7525 525 7555 555
rect 7605 525 7635 555
rect 7685 525 7715 555
rect 7765 525 7795 555
rect 7845 525 7875 555
rect 7925 525 7955 555
rect 8005 525 8035 555
rect 8085 525 8115 555
rect 8165 525 8195 555
rect 8245 525 8275 555
rect 8325 525 8355 555
rect 8405 525 8435 555
rect 8485 525 8515 555
rect 8565 525 8595 555
rect 8645 525 8675 555
rect 8725 525 8755 555
rect 8805 525 8835 555
rect 8885 525 8915 555
rect 8965 525 8995 555
rect 9045 525 9075 555
rect 9125 525 9155 555
rect 9205 525 9235 555
rect 9285 525 9315 555
rect 9365 525 9395 555
rect 9445 525 9475 555
rect 9525 525 9555 555
rect 9605 525 9635 555
rect 9685 525 9715 555
rect 9765 525 9795 555
rect 9845 525 9875 555
rect 9925 525 9955 555
rect 10005 525 10035 555
rect 10085 525 10115 555
rect 10165 525 10195 555
rect 10245 525 10275 555
rect 10325 525 10355 555
rect 10405 525 10435 555
rect 10485 525 10515 555
rect 10645 525 10675 555
rect 10805 525 10835 555
rect 10965 525 10995 555
rect -715 445 -685 475
rect -555 445 -525 475
rect -475 445 -445 475
rect 10645 445 10675 475
rect 10805 445 10835 475
rect 10965 445 10995 475
rect -715 365 -685 395
rect -555 365 -525 395
rect -395 365 -365 395
rect -315 365 -285 395
rect -235 365 -205 395
rect -155 365 -125 395
rect -75 365 -45 395
rect 5 365 35 395
rect 85 365 115 395
rect 165 365 195 395
rect 245 365 275 395
rect 325 365 355 395
rect 405 365 435 395
rect 485 365 515 395
rect 565 365 595 395
rect 645 365 675 395
rect 725 365 755 395
rect 805 365 835 395
rect 885 365 915 395
rect 965 365 995 395
rect 1045 365 1075 395
rect 1125 365 1155 395
rect 1205 365 1235 395
rect 1285 365 1315 395
rect 1365 365 1395 395
rect 1445 365 1475 395
rect 1525 365 1555 395
rect 1605 365 1635 395
rect 1685 365 1715 395
rect 1765 365 1795 395
rect 1845 365 1875 395
rect 1925 365 1955 395
rect 2005 365 2035 395
rect 2085 365 2115 395
rect 2165 365 2195 395
rect 2245 365 2275 395
rect 2325 365 2355 395
rect 2405 365 2435 395
rect 2485 365 2515 395
rect 2565 365 2595 395
rect 2645 365 2675 395
rect 2725 365 2755 395
rect 2805 365 2835 395
rect 2885 365 2915 395
rect 2965 365 2995 395
rect 3045 365 3075 395
rect 3125 365 3155 395
rect 3205 365 3235 395
rect 3285 365 3315 395
rect 3365 365 3395 395
rect 3445 365 3475 395
rect 3525 365 3555 395
rect 3605 365 3635 395
rect 3685 365 3715 395
rect 3765 365 3795 395
rect 3845 365 3875 395
rect 3925 365 3955 395
rect 4005 365 4035 395
rect 4085 365 4115 395
rect 4165 365 4195 395
rect 4245 365 4275 395
rect 4325 365 4355 395
rect 4405 365 4435 395
rect 4485 365 4515 395
rect 4565 365 4595 395
rect 4645 365 4675 395
rect 4725 365 4755 395
rect 4805 365 4835 395
rect 4885 365 4915 395
rect 4965 365 4995 395
rect 5045 365 5075 395
rect 5125 365 5155 395
rect 5205 365 5235 395
rect 5285 365 5315 395
rect 5365 365 5395 395
rect 5445 365 5475 395
rect 5525 365 5555 395
rect 5605 365 5635 395
rect 5685 365 5715 395
rect 5765 365 5795 395
rect 5845 365 5875 395
rect 5925 365 5955 395
rect 6005 365 6035 395
rect 6085 365 6115 395
rect 6165 365 6195 395
rect 6245 365 6275 395
rect 6325 365 6355 395
rect 6405 365 6435 395
rect 6485 365 6515 395
rect 6565 365 6595 395
rect 6645 365 6675 395
rect 6725 365 6755 395
rect 6805 365 6835 395
rect 6885 365 6915 395
rect 6965 365 6995 395
rect 7045 365 7075 395
rect 7125 365 7155 395
rect 7205 365 7235 395
rect 7285 365 7315 395
rect 7365 365 7395 395
rect 7445 365 7475 395
rect 7525 365 7555 395
rect 7605 365 7635 395
rect 7685 365 7715 395
rect 7765 365 7795 395
rect 7845 365 7875 395
rect 7925 365 7955 395
rect 8005 365 8035 395
rect 8085 365 8115 395
rect 8165 365 8195 395
rect 8245 365 8275 395
rect 8325 365 8355 395
rect 8405 365 8435 395
rect 8485 365 8515 395
rect 8565 365 8595 395
rect 8645 365 8675 395
rect 8725 365 8755 395
rect 8805 365 8835 395
rect 8885 365 8915 395
rect 8965 365 8995 395
rect 9045 365 9075 395
rect 9125 365 9155 395
rect 9205 365 9235 395
rect 9285 365 9315 395
rect 9365 365 9395 395
rect 9445 365 9475 395
rect 9525 365 9555 395
rect 9605 365 9635 395
rect 9685 365 9715 395
rect 9765 365 9795 395
rect 9845 365 9875 395
rect 9925 365 9955 395
rect 10005 365 10035 395
rect 10085 365 10115 395
rect 10165 365 10195 395
rect 10245 365 10275 395
rect 10325 365 10355 395
rect 10405 365 10435 395
rect 10485 365 10515 395
rect 10645 365 10675 395
rect 10805 365 10835 395
rect 10965 365 10995 395
rect -715 285 -685 315
rect -555 285 -525 315
rect -395 285 -365 315
rect 10885 285 10915 315
rect -715 205 -685 235
rect -555 205 -525 235
rect -395 205 -365 235
rect -315 205 -285 235
rect -235 205 -205 235
rect -155 205 -125 235
rect -75 205 -45 235
rect 5 205 35 235
rect 85 205 115 235
rect 165 205 195 235
rect 245 205 275 235
rect 325 205 355 235
rect 405 205 435 235
rect 485 205 515 235
rect 565 205 595 235
rect 645 205 675 235
rect 725 205 755 235
rect 805 205 835 235
rect 885 205 915 235
rect 965 205 995 235
rect 1045 205 1075 235
rect 1125 205 1155 235
rect 1205 205 1235 235
rect 1285 205 1315 235
rect 1365 205 1395 235
rect 1445 205 1475 235
rect 1525 205 1555 235
rect 1605 205 1635 235
rect 1685 205 1715 235
rect 1765 205 1795 235
rect 1845 205 1875 235
rect 1925 205 1955 235
rect 2005 205 2035 235
rect 2085 205 2115 235
rect 2165 205 2195 235
rect 2245 205 2275 235
rect 2325 205 2355 235
rect 2405 205 2435 235
rect 2485 205 2515 235
rect 2565 205 2595 235
rect 2645 205 2675 235
rect 2725 205 2755 235
rect 2805 205 2835 235
rect 2885 205 2915 235
rect 2965 205 2995 235
rect 3045 205 3075 235
rect 3125 205 3155 235
rect 3205 205 3235 235
rect 3285 205 3315 235
rect 3365 205 3395 235
rect 3445 205 3475 235
rect 3525 205 3555 235
rect 3605 205 3635 235
rect 3685 205 3715 235
rect 3765 205 3795 235
rect 3845 205 3875 235
rect 3925 205 3955 235
rect 4005 205 4035 235
rect 4085 205 4115 235
rect 4165 205 4195 235
rect 4245 205 4275 235
rect 4325 205 4355 235
rect 4405 205 4435 235
rect 4485 205 4515 235
rect 4565 205 4595 235
rect 4645 205 4675 235
rect 4725 205 4755 235
rect 4805 205 4835 235
rect 4885 205 4915 235
rect 4965 205 4995 235
rect 5045 205 5075 235
rect 5125 205 5155 235
rect 5205 205 5235 235
rect 5285 205 5315 235
rect 5365 205 5395 235
rect 5445 205 5475 235
rect 5525 205 5555 235
rect 5605 205 5635 235
rect 5685 205 5715 235
rect 5765 205 5795 235
rect 5845 205 5875 235
rect 5925 205 5955 235
rect 6005 205 6035 235
rect 6085 205 6115 235
rect 6165 205 6195 235
rect 6245 205 6275 235
rect 6325 205 6355 235
rect 6405 205 6435 235
rect 6485 205 6515 235
rect 6565 205 6595 235
rect 6645 205 6675 235
rect 6725 205 6755 235
rect 6805 205 6835 235
rect 6885 205 6915 235
rect 6965 205 6995 235
rect 7045 205 7075 235
rect 7125 205 7155 235
rect 7205 205 7235 235
rect 7285 205 7315 235
rect 7365 205 7395 235
rect 7445 205 7475 235
rect 7525 205 7555 235
rect 7605 205 7635 235
rect 7685 205 7715 235
rect 7765 205 7795 235
rect 7845 205 7875 235
rect 7925 205 7955 235
rect 8005 205 8035 235
rect 8085 205 8115 235
rect 8165 205 8195 235
rect 8245 205 8275 235
rect 8325 205 8355 235
rect 8405 205 8435 235
rect 8485 205 8515 235
rect 8565 205 8595 235
rect 8645 205 8675 235
rect 8725 205 8755 235
rect 8805 205 8835 235
rect 8885 205 8915 235
rect 8965 205 8995 235
rect 9045 205 9075 235
rect 9125 205 9155 235
rect 9205 205 9235 235
rect 9285 205 9315 235
rect 9365 205 9395 235
rect 9445 205 9475 235
rect 9525 205 9555 235
rect 9605 205 9635 235
rect 9685 205 9715 235
rect 9765 205 9795 235
rect 9845 205 9875 235
rect 9925 205 9955 235
rect 10005 205 10035 235
rect 10085 205 10115 235
rect 10165 205 10195 235
rect 10245 205 10275 235
rect 10325 205 10355 235
rect 10405 205 10435 235
rect 10485 205 10515 235
rect 10645 205 10675 235
rect 10805 205 10835 235
rect 10965 205 10995 235
rect -715 125 -685 155
rect -555 125 -525 155
rect -395 125 -365 155
rect 10725 125 10755 155
rect 10805 125 10835 155
rect 10965 125 10995 155
rect -715 45 -685 75
rect -555 45 -525 75
rect -395 45 -365 75
rect -315 45 -285 75
rect -235 45 -205 75
rect -155 45 -125 75
rect -75 45 -45 75
rect 5 45 35 75
rect 85 45 115 75
rect 165 45 195 75
rect 245 45 275 75
rect 325 45 355 75
rect 405 45 435 75
rect 485 45 515 75
rect 565 45 595 75
rect 645 45 675 75
rect 725 45 755 75
rect 805 45 835 75
rect 885 45 915 75
rect 965 45 995 75
rect 1045 45 1075 75
rect 1125 45 1155 75
rect 1205 45 1235 75
rect 1285 45 1315 75
rect 1365 45 1395 75
rect 1445 45 1475 75
rect 1525 45 1555 75
rect 1605 45 1635 75
rect 1685 45 1715 75
rect 1765 45 1795 75
rect 1845 45 1875 75
rect 1925 45 1955 75
rect 2005 45 2035 75
rect 2085 45 2115 75
rect 2165 45 2195 75
rect 2245 45 2275 75
rect 2325 45 2355 75
rect 2405 45 2435 75
rect 2485 45 2515 75
rect 2565 45 2595 75
rect 2645 45 2675 75
rect 2725 45 2755 75
rect 2805 45 2835 75
rect 2885 45 2915 75
rect 2965 45 2995 75
rect 3045 45 3075 75
rect 3125 45 3155 75
rect 3205 45 3235 75
rect 3285 45 3315 75
rect 3365 45 3395 75
rect 3445 45 3475 75
rect 3525 45 3555 75
rect 3605 45 3635 75
rect 3685 45 3715 75
rect 3765 45 3795 75
rect 3845 45 3875 75
rect 3925 45 3955 75
rect 4005 45 4035 75
rect 4085 45 4115 75
rect 4165 45 4195 75
rect 4245 45 4275 75
rect 4325 45 4355 75
rect 4405 45 4435 75
rect 4485 45 4515 75
rect 4565 45 4595 75
rect 4645 45 4675 75
rect 4725 45 4755 75
rect 4805 45 4835 75
rect 4885 45 4915 75
rect 4965 45 4995 75
rect 5045 45 5075 75
rect 5125 45 5155 75
rect 5205 45 5235 75
rect 5285 45 5315 75
rect 5365 45 5395 75
rect 5445 45 5475 75
rect 5525 45 5555 75
rect 5605 45 5635 75
rect 5685 45 5715 75
rect 5765 45 5795 75
rect 5845 45 5875 75
rect 5925 45 5955 75
rect 6005 45 6035 75
rect 6085 45 6115 75
rect 6165 45 6195 75
rect 6245 45 6275 75
rect 6325 45 6355 75
rect 6405 45 6435 75
rect 6485 45 6515 75
rect 6565 45 6595 75
rect 6645 45 6675 75
rect 6725 45 6755 75
rect 6805 45 6835 75
rect 6885 45 6915 75
rect 6965 45 6995 75
rect 7045 45 7075 75
rect 7125 45 7155 75
rect 7205 45 7235 75
rect 7285 45 7315 75
rect 7365 45 7395 75
rect 7445 45 7475 75
rect 7525 45 7555 75
rect 7605 45 7635 75
rect 7685 45 7715 75
rect 7765 45 7795 75
rect 7845 45 7875 75
rect 7925 45 7955 75
rect 8005 45 8035 75
rect 8085 45 8115 75
rect 8165 45 8195 75
rect 8245 45 8275 75
rect 8325 45 8355 75
rect 8405 45 8435 75
rect 8485 45 8515 75
rect 8565 45 8595 75
rect 8645 45 8675 75
rect 8725 45 8755 75
rect 8805 45 8835 75
rect 8885 45 8915 75
rect 8965 45 8995 75
rect 9045 45 9075 75
rect 9125 45 9155 75
rect 9205 45 9235 75
rect 9285 45 9315 75
rect 9365 45 9395 75
rect 9445 45 9475 75
rect 9525 45 9555 75
rect 9605 45 9635 75
rect 9685 45 9715 75
rect 9765 45 9795 75
rect 9845 45 9875 75
rect 9925 45 9955 75
rect 10005 45 10035 75
rect 10085 45 10115 75
rect 10165 45 10195 75
rect 10245 45 10275 75
rect 10325 45 10355 75
rect 10405 45 10435 75
rect 10485 45 10515 75
rect 10645 45 10675 75
rect 10805 45 10835 75
rect 10965 45 10995 75
rect -715 -35 -685 -5
rect -555 -35 -525 -5
rect -395 -35 -365 -5
rect -315 -35 -285 -5
rect -235 -35 -205 -5
rect -155 -35 -125 -5
rect -75 -35 -45 -5
rect 5 -35 35 -5
rect 85 -35 115 -5
rect 165 -35 195 -5
rect 245 -35 275 -5
rect 325 -35 355 -5
rect 405 -35 435 -5
rect 485 -35 515 -5
rect 565 -35 595 -5
rect 645 -35 675 -5
rect 725 -35 755 -5
rect 805 -35 835 -5
rect 885 -35 915 -5
rect 965 -35 995 -5
rect 1045 -35 1075 -5
rect 1125 -35 1155 -5
rect 1205 -35 1235 -5
rect 1285 -35 1315 -5
rect 1365 -35 1395 -5
rect 1445 -35 1475 -5
rect 1525 -35 1555 -5
rect 1605 -35 1635 -5
rect 1685 -35 1715 -5
rect 1765 -35 1795 -5
rect 1845 -35 1875 -5
rect 1925 -35 1955 -5
rect 2005 -35 2035 -5
rect 2085 -35 2115 -5
rect 2165 -35 2195 -5
rect 2245 -35 2275 -5
rect 2325 -35 2355 -5
rect 2405 -35 2435 -5
rect 2485 -35 2515 -5
rect 2565 -35 2595 -5
rect 2645 -35 2675 -5
rect 2725 -35 2755 -5
rect 2805 -35 2835 -5
rect 2885 -35 2915 -5
rect 2965 -35 2995 -5
rect 3045 -35 3075 -5
rect 3125 -35 3155 -5
rect 3205 -35 3235 -5
rect 3285 -35 3315 -5
rect 3365 -35 3395 -5
rect 3445 -35 3475 -5
rect 3525 -35 3555 -5
rect 3605 -35 3635 -5
rect 3685 -35 3715 -5
rect 3765 -35 3795 -5
rect 3845 -35 3875 -5
rect 3925 -35 3955 -5
rect 4005 -35 4035 -5
rect 4085 -35 4115 -5
rect 4165 -35 4195 -5
rect 4245 -35 4275 -5
rect 4325 -35 4355 -5
rect 4405 -35 4435 -5
rect 4485 -35 4515 -5
rect 4565 -35 4595 -5
rect 4645 -35 4675 -5
rect 4725 -35 4755 -5
rect 4805 -35 4835 -5
rect 4885 -35 4915 -5
rect 4965 -35 4995 -5
rect 5045 -35 5075 -5
rect 5125 -35 5155 -5
rect 5205 -35 5235 -5
rect 5285 -35 5315 -5
rect 5365 -35 5395 -5
rect 5445 -35 5475 -5
rect 5525 -35 5555 -5
rect 5605 -35 5635 -5
rect 5685 -35 5715 -5
rect 5765 -35 5795 -5
rect 5845 -35 5875 -5
rect 5925 -35 5955 -5
rect 6005 -35 6035 -5
rect 6085 -35 6115 -5
rect 6165 -35 6195 -5
rect 6245 -35 6275 -5
rect 6325 -35 6355 -5
rect 6405 -35 6435 -5
rect 6485 -35 6515 -5
rect 6565 -35 6595 -5
rect 6645 -35 6675 -5
rect 6725 -35 6755 -5
rect 6805 -35 6835 -5
rect 6885 -35 6915 -5
rect 6965 -35 6995 -5
rect 7045 -35 7075 -5
rect 7125 -35 7155 -5
rect 7205 -35 7235 -5
rect 7285 -35 7315 -5
rect 7365 -35 7395 -5
rect 7445 -35 7475 -5
rect 7525 -35 7555 -5
rect 7605 -35 7635 -5
rect 7685 -35 7715 -5
rect 7765 -35 7795 -5
rect 7845 -35 7875 -5
rect 7925 -35 7955 -5
rect 8005 -35 8035 -5
rect 8085 -35 8115 -5
rect 8165 -35 8195 -5
rect 8245 -35 8275 -5
rect 8325 -35 8355 -5
rect 8405 -35 8435 -5
rect 8485 -35 8515 -5
rect 8565 -35 8595 -5
rect 8645 -35 8675 -5
rect 8725 -35 8755 -5
rect 8805 -35 8835 -5
rect 8885 -35 8915 -5
rect 8965 -35 8995 -5
rect 9045 -35 9075 -5
rect 9125 -35 9155 -5
rect 9205 -35 9235 -5
rect 9285 -35 9315 -5
rect 9365 -35 9395 -5
rect 9445 -35 9475 -5
rect 9525 -35 9555 -5
rect 9605 -35 9635 -5
rect 9685 -35 9715 -5
rect 9765 -35 9795 -5
rect 9845 -35 9875 -5
rect 9925 -35 9955 -5
rect 10005 -35 10035 -5
rect 10085 -35 10115 -5
rect 10165 -35 10195 -5
rect 10245 -35 10275 -5
rect 10325 -35 10355 -5
rect 10405 -35 10435 -5
rect 10485 -35 10515 -5
rect 10645 -35 10675 -5
rect 10805 -35 10835 -5
rect 10965 -35 10995 -5
rect -715 -115 -685 -85
rect -555 -115 -525 -85
rect -395 -115 -365 -85
rect -315 -115 -285 -85
rect -235 -115 -205 -85
rect -155 -115 -125 -85
rect -75 -115 -45 -85
rect 5 -115 35 -85
rect 85 -115 115 -85
rect 165 -115 195 -85
rect 245 -115 275 -85
rect 325 -115 355 -85
rect 405 -115 435 -85
rect 485 -115 515 -85
rect 565 -115 595 -85
rect 645 -115 675 -85
rect 725 -115 755 -85
rect 805 -115 835 -85
rect 885 -115 915 -85
rect 965 -115 995 -85
rect 1045 -115 1075 -85
rect 1125 -115 1155 -85
rect 1205 -115 1235 -85
rect 1285 -115 1315 -85
rect 1365 -115 1395 -85
rect 1445 -115 1475 -85
rect 1525 -115 1555 -85
rect 1605 -115 1635 -85
rect 1685 -115 1715 -85
rect 1765 -115 1795 -85
rect 1845 -115 1875 -85
rect 1925 -115 1955 -85
rect 2005 -115 2035 -85
rect 2085 -115 2115 -85
rect 2165 -115 2195 -85
rect 2245 -115 2275 -85
rect 2325 -115 2355 -85
rect 2405 -115 2435 -85
rect 2485 -115 2515 -85
rect 2565 -115 2595 -85
rect 2645 -115 2675 -85
rect 2725 -115 2755 -85
rect 2805 -115 2835 -85
rect 2885 -115 2915 -85
rect 2965 -115 2995 -85
rect 3045 -115 3075 -85
rect 3125 -115 3155 -85
rect 3205 -115 3235 -85
rect 3285 -115 3315 -85
rect 3365 -115 3395 -85
rect 3445 -115 3475 -85
rect 3525 -115 3555 -85
rect 3605 -115 3635 -85
rect 3685 -115 3715 -85
rect 3765 -115 3795 -85
rect 3845 -115 3875 -85
rect 3925 -115 3955 -85
rect 4005 -115 4035 -85
rect 4085 -115 4115 -85
rect 4165 -115 4195 -85
rect 4245 -115 4275 -85
rect 4325 -115 4355 -85
rect 4405 -115 4435 -85
rect 4485 -115 4515 -85
rect 4565 -115 4595 -85
rect 4645 -115 4675 -85
rect 4725 -115 4755 -85
rect 4805 -115 4835 -85
rect 4885 -115 4915 -85
rect 4965 -115 4995 -85
rect 5045 -115 5075 -85
rect 5125 -115 5155 -85
rect 5205 -115 5235 -85
rect 5285 -115 5315 -85
rect 5365 -115 5395 -85
rect 5445 -115 5475 -85
rect 5525 -115 5555 -85
rect 5605 -115 5635 -85
rect 5685 -115 5715 -85
rect 5765 -115 5795 -85
rect 5845 -115 5875 -85
rect 5925 -115 5955 -85
rect 6005 -115 6035 -85
rect 6085 -115 6115 -85
rect 6165 -115 6195 -85
rect 6245 -115 6275 -85
rect 6325 -115 6355 -85
rect 6405 -115 6435 -85
rect 6485 -115 6515 -85
rect 6565 -115 6595 -85
rect 6645 -115 6675 -85
rect 6725 -115 6755 -85
rect 6805 -115 6835 -85
rect 6885 -115 6915 -85
rect 6965 -115 6995 -85
rect 7045 -115 7075 -85
rect 7125 -115 7155 -85
rect 7205 -115 7235 -85
rect 7285 -115 7315 -85
rect 7365 -115 7395 -85
rect 7445 -115 7475 -85
rect 7525 -115 7555 -85
rect 7605 -115 7635 -85
rect 7685 -115 7715 -85
rect 7765 -115 7795 -85
rect 7845 -115 7875 -85
rect 7925 -115 7955 -85
rect 8005 -115 8035 -85
rect 8085 -115 8115 -85
rect 8165 -115 8195 -85
rect 8245 -115 8275 -85
rect 8325 -115 8355 -85
rect 8405 -115 8435 -85
rect 8485 -115 8515 -85
rect 8565 -115 8595 -85
rect 8645 -115 8675 -85
rect 8725 -115 8755 -85
rect 8805 -115 8835 -85
rect 8885 -115 8915 -85
rect 8965 -115 8995 -85
rect 9045 -115 9075 -85
rect 9125 -115 9155 -85
rect 9205 -115 9235 -85
rect 9285 -115 9315 -85
rect 9365 -115 9395 -85
rect 9445 -115 9475 -85
rect 9525 -115 9555 -85
rect 9605 -115 9635 -85
rect 9685 -115 9715 -85
rect 9765 -115 9795 -85
rect 9845 -115 9875 -85
rect 9925 -115 9955 -85
rect 10005 -115 10035 -85
rect 10085 -115 10115 -85
rect 10165 -115 10195 -85
rect 10245 -115 10275 -85
rect 10325 -115 10355 -85
rect 10405 -115 10435 -85
rect 10485 -115 10515 -85
rect 10645 -115 10675 -85
rect 10805 -115 10835 -85
rect 10965 -115 10995 -85
rect -715 -195 -685 -165
rect -555 -195 -525 -165
rect -395 -195 -365 -165
rect -235 -195 -205 -165
rect -155 -195 -125 -165
rect -75 -195 -45 -165
rect 5 -195 35 -165
rect 85 -195 115 -165
rect 165 -195 195 -165
rect 245 -195 275 -165
rect 325 -195 355 -165
rect 405 -195 435 -165
rect 485 -195 515 -165
rect 565 -195 595 -165
rect 645 -195 675 -165
rect 725 -195 755 -165
rect 805 -195 835 -165
rect 885 -195 915 -165
rect 965 -195 995 -165
rect 1045 -195 1075 -165
rect 1125 -195 1155 -165
rect 1205 -195 1235 -165
rect 1285 -195 1315 -165
rect 1365 -195 1395 -165
rect 1445 -195 1475 -165
rect 1525 -195 1555 -165
rect 1605 -195 1635 -165
rect 1685 -195 1715 -165
rect 1765 -195 1795 -165
rect 1845 -195 1875 -165
rect 1925 -195 1955 -165
rect 2005 -195 2035 -165
rect 2085 -195 2115 -165
rect 2165 -195 2195 -165
rect 2245 -195 2275 -165
rect 2325 -195 2355 -165
rect 2405 -195 2435 -165
rect 2485 -195 2515 -165
rect 2565 -195 2595 -165
rect 2645 -195 2675 -165
rect 2725 -195 2755 -165
rect 2805 -195 2835 -165
rect 2885 -195 2915 -165
rect 2965 -195 2995 -165
rect 3045 -195 3075 -165
rect 3125 -195 3155 -165
rect 3205 -195 3235 -165
rect 3285 -195 3315 -165
rect 3365 -195 3395 -165
rect 3445 -195 3475 -165
rect 3525 -195 3555 -165
rect 3605 -195 3635 -165
rect 3685 -195 3715 -165
rect 3765 -195 3795 -165
rect 3845 -195 3875 -165
rect 3925 -195 3955 -165
rect 4005 -195 4035 -165
rect 4085 -195 4115 -165
rect 4165 -195 4195 -165
rect 4245 -195 4275 -165
rect 4325 -195 4355 -165
rect 4405 -195 4435 -165
rect 4485 -195 4515 -165
rect 4565 -195 4595 -165
rect 4645 -195 4675 -165
rect 4725 -195 4755 -165
rect 4805 -195 4835 -165
rect 4885 -195 4915 -165
rect 4965 -195 4995 -165
rect 5045 -195 5075 -165
rect 5125 -195 5155 -165
rect 5205 -195 5235 -165
rect 5285 -195 5315 -165
rect 5365 -195 5395 -165
rect 5445 -195 5475 -165
rect 5525 -195 5555 -165
rect 5605 -195 5635 -165
rect 5685 -195 5715 -165
rect 5765 -195 5795 -165
rect 5845 -195 5875 -165
rect 5925 -195 5955 -165
rect 6005 -195 6035 -165
rect 6085 -195 6115 -165
rect 6165 -195 6195 -165
rect 6245 -195 6275 -165
rect 6325 -195 6355 -165
rect 6405 -195 6435 -165
rect 6485 -195 6515 -165
rect 6565 -195 6595 -165
rect 6645 -195 6675 -165
rect 6725 -195 6755 -165
rect 6805 -195 6835 -165
rect 6885 -195 6915 -165
rect 6965 -195 6995 -165
rect 7045 -195 7075 -165
rect 7125 -195 7155 -165
rect 7205 -195 7235 -165
rect 7285 -195 7315 -165
rect 7365 -195 7395 -165
rect 7445 -195 7475 -165
rect 7525 -195 7555 -165
rect 7605 -195 7635 -165
rect 7685 -195 7715 -165
rect 7765 -195 7795 -165
rect 7845 -195 7875 -165
rect 7925 -195 7955 -165
rect 8005 -195 8035 -165
rect 8085 -195 8115 -165
rect 8165 -195 8195 -165
rect 8245 -195 8275 -165
rect 8325 -195 8355 -165
rect 8405 -195 8435 -165
rect 8485 -195 8515 -165
rect 8565 -195 8595 -165
rect 8645 -195 8675 -165
rect 8725 -195 8755 -165
rect 8805 -195 8835 -165
rect 8885 -195 8915 -165
rect 8965 -195 8995 -165
rect 9045 -195 9075 -165
rect 9125 -195 9155 -165
rect 9205 -195 9235 -165
rect 9285 -195 9315 -165
rect 9365 -195 9395 -165
rect 9445 -195 9475 -165
rect 9525 -195 9555 -165
rect 9605 -195 9635 -165
rect 9685 -195 9715 -165
rect 9765 -195 9795 -165
rect 9845 -195 9875 -165
rect 9925 -195 9955 -165
rect 10005 -195 10035 -165
rect 10085 -195 10115 -165
rect 10165 -195 10195 -165
rect 10245 -195 10275 -165
rect 10325 -195 10355 -165
rect 10405 -195 10435 -165
rect 10485 -195 10515 -165
rect 10565 -195 10595 -165
rect 10645 -195 10675 -165
rect 10805 -195 10835 -165
rect 10965 -195 10995 -165
rect -715 -275 -685 -245
rect -555 -275 -525 -245
rect -395 -275 -365 -245
rect -235 -275 -205 -245
rect -155 -275 -125 -245
rect -75 -275 -45 -245
rect 5 -275 35 -245
rect 85 -275 115 -245
rect 165 -275 195 -245
rect 245 -275 275 -245
rect 325 -275 355 -245
rect 405 -275 435 -245
rect 485 -275 515 -245
rect 565 -275 595 -245
rect 645 -275 675 -245
rect 725 -275 755 -245
rect 805 -275 835 -245
rect 885 -275 915 -245
rect 965 -275 995 -245
rect 1045 -275 1075 -245
rect 1125 -275 1155 -245
rect 1205 -275 1235 -245
rect 1285 -275 1315 -245
rect 1365 -275 1395 -245
rect 1445 -275 1475 -245
rect 1525 -275 1555 -245
rect 1605 -275 1635 -245
rect 1685 -275 1715 -245
rect 1765 -275 1795 -245
rect 1845 -275 1875 -245
rect 1925 -275 1955 -245
rect 2005 -275 2035 -245
rect 2085 -275 2115 -245
rect 2165 -275 2195 -245
rect 2245 -275 2275 -245
rect 2325 -275 2355 -245
rect 2405 -275 2435 -245
rect 2485 -275 2515 -245
rect 2565 -275 2595 -245
rect 2645 -275 2675 -245
rect 2725 -275 2755 -245
rect 2805 -275 2835 -245
rect 2885 -275 2915 -245
rect 2965 -275 2995 -245
rect 3045 -275 3075 -245
rect 3125 -275 3155 -245
rect 3205 -275 3235 -245
rect 3285 -275 3315 -245
rect 3365 -275 3395 -245
rect 3445 -275 3475 -245
rect 3525 -275 3555 -245
rect 3605 -275 3635 -245
rect 3685 -275 3715 -245
rect 3765 -275 3795 -245
rect 3845 -275 3875 -245
rect 3925 -275 3955 -245
rect 4005 -275 4035 -245
rect 4085 -275 4115 -245
rect 4165 -275 4195 -245
rect 4245 -275 4275 -245
rect 4325 -275 4355 -245
rect 4405 -275 4435 -245
rect 4485 -275 4515 -245
rect 4565 -275 4595 -245
rect 4645 -275 4675 -245
rect 4725 -275 4755 -245
rect 4805 -275 4835 -245
rect 4885 -275 4915 -245
rect 4965 -275 4995 -245
rect 5045 -275 5075 -245
rect 5125 -275 5155 -245
rect 5205 -275 5235 -245
rect 5285 -275 5315 -245
rect 5365 -275 5395 -245
rect 5445 -275 5475 -245
rect 5525 -275 5555 -245
rect 5605 -275 5635 -245
rect 5685 -275 5715 -245
rect 5765 -275 5795 -245
rect 5845 -275 5875 -245
rect 5925 -275 5955 -245
rect 6005 -275 6035 -245
rect 6085 -275 6115 -245
rect 6165 -275 6195 -245
rect 6245 -275 6275 -245
rect 6325 -275 6355 -245
rect 6405 -275 6435 -245
rect 6485 -275 6515 -245
rect 6565 -275 6595 -245
rect 6645 -275 6675 -245
rect 6725 -275 6755 -245
rect 6805 -275 6835 -245
rect 6885 -275 6915 -245
rect 6965 -275 6995 -245
rect 7045 -275 7075 -245
rect 7125 -275 7155 -245
rect 7205 -275 7235 -245
rect 7285 -275 7315 -245
rect 7365 -275 7395 -245
rect 7445 -275 7475 -245
rect 7525 -275 7555 -245
rect 7605 -275 7635 -245
rect 7685 -275 7715 -245
rect 7765 -275 7795 -245
rect 7845 -275 7875 -245
rect 7925 -275 7955 -245
rect 8005 -275 8035 -245
rect 8085 -275 8115 -245
rect 8165 -275 8195 -245
rect 8245 -275 8275 -245
rect 8325 -275 8355 -245
rect 8405 -275 8435 -245
rect 8485 -275 8515 -245
rect 8565 -275 8595 -245
rect 8645 -275 8675 -245
rect 8725 -275 8755 -245
rect 8805 -275 8835 -245
rect 8885 -275 8915 -245
rect 8965 -275 8995 -245
rect 9045 -275 9075 -245
rect 9125 -275 9155 -245
rect 9205 -275 9235 -245
rect 9285 -275 9315 -245
rect 9365 -275 9395 -245
rect 9445 -275 9475 -245
rect 9525 -275 9555 -245
rect 9605 -275 9635 -245
rect 9685 -275 9715 -245
rect 9765 -275 9795 -245
rect 9845 -275 9875 -245
rect 9925 -275 9955 -245
rect 10005 -275 10035 -245
rect 10085 -275 10115 -245
rect 10165 -275 10195 -245
rect 10245 -275 10275 -245
rect 10325 -275 10355 -245
rect 10405 -275 10435 -245
rect 10485 -275 10515 -245
rect 10565 -275 10595 -245
rect 10645 -275 10675 -245
rect 10805 -275 10835 -245
rect 10965 -275 10995 -245
rect -715 -355 -685 -325
rect -555 -355 -525 -325
rect -395 -355 -365 -325
rect -235 -355 -205 -325
rect -155 -355 -125 -325
rect -75 -355 -45 -325
rect 5 -355 35 -325
rect 85 -355 115 -325
rect 165 -355 195 -325
rect 245 -355 275 -325
rect 325 -355 355 -325
rect 405 -355 435 -325
rect 485 -355 515 -325
rect 565 -355 595 -325
rect 645 -355 675 -325
rect 725 -355 755 -325
rect 805 -355 835 -325
rect 885 -355 915 -325
rect 965 -355 995 -325
rect 1045 -355 1075 -325
rect 1125 -355 1155 -325
rect 1205 -355 1235 -325
rect 1285 -355 1315 -325
rect 1365 -355 1395 -325
rect 1445 -355 1475 -325
rect 1525 -355 1555 -325
rect 1605 -355 1635 -325
rect 1685 -355 1715 -325
rect 1765 -355 1795 -325
rect 1845 -355 1875 -325
rect 1925 -355 1955 -325
rect 2005 -355 2035 -325
rect 2085 -355 2115 -325
rect 2165 -355 2195 -325
rect 2245 -355 2275 -325
rect 2325 -355 2355 -325
rect 2405 -355 2435 -325
rect 2485 -355 2515 -325
rect 2565 -355 2595 -325
rect 2645 -355 2675 -325
rect 2725 -355 2755 -325
rect 2805 -355 2835 -325
rect 2885 -355 2915 -325
rect 2965 -355 2995 -325
rect 3045 -355 3075 -325
rect 3125 -355 3155 -325
rect 3205 -355 3235 -325
rect 3285 -355 3315 -325
rect 3365 -355 3395 -325
rect 3445 -355 3475 -325
rect 3525 -355 3555 -325
rect 3605 -355 3635 -325
rect 3685 -355 3715 -325
rect 3765 -355 3795 -325
rect 3845 -355 3875 -325
rect 3925 -355 3955 -325
rect 4005 -355 4035 -325
rect 4085 -355 4115 -325
rect 4165 -355 4195 -325
rect 4245 -355 4275 -325
rect 4325 -355 4355 -325
rect 4405 -355 4435 -325
rect 4485 -355 4515 -325
rect 4565 -355 4595 -325
rect 4645 -355 4675 -325
rect 4725 -355 4755 -325
rect 4805 -355 4835 -325
rect 4885 -355 4915 -325
rect 4965 -355 4995 -325
rect 5045 -355 5075 -325
rect 5125 -355 5155 -325
rect 5205 -355 5235 -325
rect 5285 -355 5315 -325
rect 5365 -355 5395 -325
rect 5445 -355 5475 -325
rect 5525 -355 5555 -325
rect 5605 -355 5635 -325
rect 5685 -355 5715 -325
rect 5765 -355 5795 -325
rect 5845 -355 5875 -325
rect 5925 -355 5955 -325
rect 6005 -355 6035 -325
rect 6085 -355 6115 -325
rect 6165 -355 6195 -325
rect 6245 -355 6275 -325
rect 6325 -355 6355 -325
rect 6405 -355 6435 -325
rect 6485 -355 6515 -325
rect 6565 -355 6595 -325
rect 6645 -355 6675 -325
rect 6725 -355 6755 -325
rect 6805 -355 6835 -325
rect 6885 -355 6915 -325
rect 6965 -355 6995 -325
rect 7045 -355 7075 -325
rect 7125 -355 7155 -325
rect 7205 -355 7235 -325
rect 7285 -355 7315 -325
rect 7365 -355 7395 -325
rect 7445 -355 7475 -325
rect 7525 -355 7555 -325
rect 7605 -355 7635 -325
rect 7685 -355 7715 -325
rect 7765 -355 7795 -325
rect 7845 -355 7875 -325
rect 7925 -355 7955 -325
rect 8005 -355 8035 -325
rect 8085 -355 8115 -325
rect 8165 -355 8195 -325
rect 8245 -355 8275 -325
rect 8325 -355 8355 -325
rect 8405 -355 8435 -325
rect 8485 -355 8515 -325
rect 8565 -355 8595 -325
rect 8645 -355 8675 -325
rect 8725 -355 8755 -325
rect 8805 -355 8835 -325
rect 8885 -355 8915 -325
rect 8965 -355 8995 -325
rect 9045 -355 9075 -325
rect 9125 -355 9155 -325
rect 9205 -355 9235 -325
rect 9285 -355 9315 -325
rect 9365 -355 9395 -325
rect 9445 -355 9475 -325
rect 9525 -355 9555 -325
rect 9605 -355 9635 -325
rect 9685 -355 9715 -325
rect 9765 -355 9795 -325
rect 9845 -355 9875 -325
rect 9925 -355 9955 -325
rect 10005 -355 10035 -325
rect 10085 -355 10115 -325
rect 10165 -355 10195 -325
rect 10245 -355 10275 -325
rect 10325 -355 10355 -325
rect 10405 -355 10435 -325
rect 10485 -355 10515 -325
rect 10565 -355 10595 -325
rect 10645 -355 10675 -325
rect 10805 -355 10835 -325
rect 10965 -355 10995 -325
rect -715 -435 -685 -405
rect -555 -435 -525 -405
rect -395 -435 -365 -405
rect 10725 -435 10755 -405
rect 10805 -435 10835 -405
rect 10965 -435 10995 -405
rect -715 -515 -685 -485
rect -555 -515 -525 -485
rect -395 -515 -365 -485
rect -235 -515 -205 -485
rect -155 -515 -125 -485
rect -75 -515 -45 -485
rect 5 -515 35 -485
rect 85 -515 115 -485
rect 165 -515 195 -485
rect 245 -515 275 -485
rect 325 -515 355 -485
rect 405 -515 435 -485
rect 485 -515 515 -485
rect 565 -515 595 -485
rect 645 -515 675 -485
rect 725 -515 755 -485
rect 805 -515 835 -485
rect 885 -515 915 -485
rect 965 -515 995 -485
rect 1045 -515 1075 -485
rect 1125 -515 1155 -485
rect 1205 -515 1235 -485
rect 1285 -515 1315 -485
rect 1365 -515 1395 -485
rect 1445 -515 1475 -485
rect 1525 -515 1555 -485
rect 1605 -515 1635 -485
rect 1685 -515 1715 -485
rect 1765 -515 1795 -485
rect 1845 -515 1875 -485
rect 1925 -515 1955 -485
rect 2005 -515 2035 -485
rect 2085 -515 2115 -485
rect 2165 -515 2195 -485
rect 2245 -515 2275 -485
rect 2325 -515 2355 -485
rect 2405 -515 2435 -485
rect 2485 -515 2515 -485
rect 2565 -515 2595 -485
rect 2645 -515 2675 -485
rect 2725 -515 2755 -485
rect 2805 -515 2835 -485
rect 2885 -515 2915 -485
rect 2965 -515 2995 -485
rect 3045 -515 3075 -485
rect 3125 -515 3155 -485
rect 3205 -515 3235 -485
rect 3285 -515 3315 -485
rect 3365 -515 3395 -485
rect 3445 -515 3475 -485
rect 3525 -515 3555 -485
rect 3605 -515 3635 -485
rect 3685 -515 3715 -485
rect 3765 -515 3795 -485
rect 3845 -515 3875 -485
rect 3925 -515 3955 -485
rect 4005 -515 4035 -485
rect 4085 -515 4115 -485
rect 4165 -515 4195 -485
rect 4245 -515 4275 -485
rect 4325 -515 4355 -485
rect 4405 -515 4435 -485
rect 4485 -515 4515 -485
rect 4565 -515 4595 -485
rect 4645 -515 4675 -485
rect 4725 -515 4755 -485
rect 4805 -515 4835 -485
rect 4885 -515 4915 -485
rect 4965 -515 4995 -485
rect 5045 -515 5075 -485
rect 5125 -515 5155 -485
rect 5205 -515 5235 -485
rect 5285 -515 5315 -485
rect 5365 -515 5395 -485
rect 5445 -515 5475 -485
rect 5525 -515 5555 -485
rect 5605 -515 5635 -485
rect 5685 -515 5715 -485
rect 5765 -515 5795 -485
rect 5845 -515 5875 -485
rect 5925 -515 5955 -485
rect 6005 -515 6035 -485
rect 6085 -515 6115 -485
rect 6165 -515 6195 -485
rect 6245 -515 6275 -485
rect 6325 -515 6355 -485
rect 6405 -515 6435 -485
rect 6485 -515 6515 -485
rect 6565 -515 6595 -485
rect 6645 -515 6675 -485
rect 6725 -515 6755 -485
rect 6805 -515 6835 -485
rect 6885 -515 6915 -485
rect 6965 -515 6995 -485
rect 7045 -515 7075 -485
rect 7125 -515 7155 -485
rect 7205 -515 7235 -485
rect 7285 -515 7315 -485
rect 7365 -515 7395 -485
rect 7445 -515 7475 -485
rect 7525 -515 7555 -485
rect 7605 -515 7635 -485
rect 7685 -515 7715 -485
rect 7765 -515 7795 -485
rect 7845 -515 7875 -485
rect 7925 -515 7955 -485
rect 8005 -515 8035 -485
rect 8085 -515 8115 -485
rect 8165 -515 8195 -485
rect 8245 -515 8275 -485
rect 8325 -515 8355 -485
rect 8405 -515 8435 -485
rect 8485 -515 8515 -485
rect 8565 -515 8595 -485
rect 8645 -515 8675 -485
rect 8725 -515 8755 -485
rect 8805 -515 8835 -485
rect 8885 -515 8915 -485
rect 8965 -515 8995 -485
rect 9045 -515 9075 -485
rect 9125 -515 9155 -485
rect 9205 -515 9235 -485
rect 9285 -515 9315 -485
rect 9365 -515 9395 -485
rect 9445 -515 9475 -485
rect 9525 -515 9555 -485
rect 9605 -515 9635 -485
rect 9685 -515 9715 -485
rect 9765 -515 9795 -485
rect 9845 -515 9875 -485
rect 9925 -515 9955 -485
rect 10005 -515 10035 -485
rect 10085 -515 10115 -485
rect 10165 -515 10195 -485
rect 10245 -515 10275 -485
rect 10325 -515 10355 -485
rect 10405 -515 10435 -485
rect 10485 -515 10515 -485
rect 10565 -515 10595 -485
rect 10645 -515 10675 -485
rect 10805 -515 10835 -485
rect 10965 -515 10995 -485
rect -715 -595 -685 -565
rect -555 -595 -525 -565
rect -395 -595 -365 -565
rect 10885 -595 10915 -565
rect -715 -675 -685 -645
rect -555 -675 -525 -645
rect -395 -675 -365 -645
rect -235 -675 -205 -645
rect -155 -675 -125 -645
rect -75 -675 -45 -645
rect 5 -675 35 -645
rect 85 -675 115 -645
rect 165 -675 195 -645
rect 245 -675 275 -645
rect 325 -675 355 -645
rect 405 -675 435 -645
rect 485 -675 515 -645
rect 565 -675 595 -645
rect 645 -675 675 -645
rect 725 -675 755 -645
rect 805 -675 835 -645
rect 885 -675 915 -645
rect 965 -675 995 -645
rect 1045 -675 1075 -645
rect 1125 -675 1155 -645
rect 1205 -675 1235 -645
rect 1285 -675 1315 -645
rect 1365 -675 1395 -645
rect 1445 -675 1475 -645
rect 1525 -675 1555 -645
rect 1605 -675 1635 -645
rect 1685 -675 1715 -645
rect 1765 -675 1795 -645
rect 1845 -675 1875 -645
rect 1925 -675 1955 -645
rect 2005 -675 2035 -645
rect 2085 -675 2115 -645
rect 2165 -675 2195 -645
rect 2245 -675 2275 -645
rect 2325 -675 2355 -645
rect 2405 -675 2435 -645
rect 2485 -675 2515 -645
rect 2565 -675 2595 -645
rect 2645 -675 2675 -645
rect 2725 -675 2755 -645
rect 2805 -675 2835 -645
rect 2885 -675 2915 -645
rect 2965 -675 2995 -645
rect 3045 -675 3075 -645
rect 3125 -675 3155 -645
rect 3205 -675 3235 -645
rect 3285 -675 3315 -645
rect 3365 -675 3395 -645
rect 3445 -675 3475 -645
rect 3525 -675 3555 -645
rect 3605 -675 3635 -645
rect 3685 -675 3715 -645
rect 3765 -675 3795 -645
rect 3845 -675 3875 -645
rect 3925 -675 3955 -645
rect 4005 -675 4035 -645
rect 4085 -675 4115 -645
rect 4165 -675 4195 -645
rect 4245 -675 4275 -645
rect 4325 -675 4355 -645
rect 4405 -675 4435 -645
rect 4485 -675 4515 -645
rect 4565 -675 4595 -645
rect 4645 -675 4675 -645
rect 4725 -675 4755 -645
rect 4805 -675 4835 -645
rect 4885 -675 4915 -645
rect 4965 -675 4995 -645
rect 5045 -675 5075 -645
rect 5125 -675 5155 -645
rect 5205 -675 5235 -645
rect 5285 -675 5315 -645
rect 5365 -675 5395 -645
rect 5445 -675 5475 -645
rect 5525 -675 5555 -645
rect 5605 -675 5635 -645
rect 5685 -675 5715 -645
rect 5765 -675 5795 -645
rect 5845 -675 5875 -645
rect 5925 -675 5955 -645
rect 6005 -675 6035 -645
rect 6085 -675 6115 -645
rect 6165 -675 6195 -645
rect 6245 -675 6275 -645
rect 6325 -675 6355 -645
rect 6405 -675 6435 -645
rect 6485 -675 6515 -645
rect 6565 -675 6595 -645
rect 6645 -675 6675 -645
rect 6725 -675 6755 -645
rect 6805 -675 6835 -645
rect 6885 -675 6915 -645
rect 6965 -675 6995 -645
rect 7045 -675 7075 -645
rect 7125 -675 7155 -645
rect 7205 -675 7235 -645
rect 7285 -675 7315 -645
rect 7365 -675 7395 -645
rect 7445 -675 7475 -645
rect 7525 -675 7555 -645
rect 7605 -675 7635 -645
rect 7685 -675 7715 -645
rect 7765 -675 7795 -645
rect 7845 -675 7875 -645
rect 7925 -675 7955 -645
rect 8005 -675 8035 -645
rect 8085 -675 8115 -645
rect 8165 -675 8195 -645
rect 8245 -675 8275 -645
rect 8325 -675 8355 -645
rect 8405 -675 8435 -645
rect 8485 -675 8515 -645
rect 8565 -675 8595 -645
rect 8645 -675 8675 -645
rect 8725 -675 8755 -645
rect 8805 -675 8835 -645
rect 8885 -675 8915 -645
rect 8965 -675 8995 -645
rect 9045 -675 9075 -645
rect 9125 -675 9155 -645
rect 9205 -675 9235 -645
rect 9285 -675 9315 -645
rect 9365 -675 9395 -645
rect 9445 -675 9475 -645
rect 9525 -675 9555 -645
rect 9605 -675 9635 -645
rect 9685 -675 9715 -645
rect 9765 -675 9795 -645
rect 9845 -675 9875 -645
rect 9925 -675 9955 -645
rect 10005 -675 10035 -645
rect 10085 -675 10115 -645
rect 10165 -675 10195 -645
rect 10245 -675 10275 -645
rect 10325 -675 10355 -645
rect 10405 -675 10435 -645
rect 10485 -675 10515 -645
rect 10565 -675 10595 -645
rect 10645 -675 10675 -645
rect 10805 -675 10835 -645
rect 10965 -675 10995 -645
rect -715 -755 -685 -725
rect -555 -755 -525 -725
rect -475 -755 -445 -725
rect 10645 -755 10675 -725
rect 10805 -755 10835 -725
rect 10965 -755 10995 -725
rect -715 -835 -685 -805
rect -555 -835 -525 -805
rect -395 -835 -365 -805
rect -235 -835 -205 -805
rect -155 -835 -125 -805
rect -75 -835 -45 -805
rect 5 -835 35 -805
rect 85 -835 115 -805
rect 165 -835 195 -805
rect 245 -835 275 -805
rect 325 -835 355 -805
rect 405 -835 435 -805
rect 485 -835 515 -805
rect 565 -835 595 -805
rect 645 -835 675 -805
rect 725 -835 755 -805
rect 805 -835 835 -805
rect 885 -835 915 -805
rect 965 -835 995 -805
rect 1045 -835 1075 -805
rect 1125 -835 1155 -805
rect 1205 -835 1235 -805
rect 1285 -835 1315 -805
rect 1365 -835 1395 -805
rect 1445 -835 1475 -805
rect 1525 -835 1555 -805
rect 1605 -835 1635 -805
rect 1685 -835 1715 -805
rect 1765 -835 1795 -805
rect 1845 -835 1875 -805
rect 1925 -835 1955 -805
rect 2005 -835 2035 -805
rect 2085 -835 2115 -805
rect 2165 -835 2195 -805
rect 2245 -835 2275 -805
rect 2325 -835 2355 -805
rect 2405 -835 2435 -805
rect 2485 -835 2515 -805
rect 2565 -835 2595 -805
rect 2645 -835 2675 -805
rect 2725 -835 2755 -805
rect 2805 -835 2835 -805
rect 2885 -835 2915 -805
rect 2965 -835 2995 -805
rect 3045 -835 3075 -805
rect 3125 -835 3155 -805
rect 3205 -835 3235 -805
rect 3285 -835 3315 -805
rect 3365 -835 3395 -805
rect 3445 -835 3475 -805
rect 3525 -835 3555 -805
rect 3605 -835 3635 -805
rect 3685 -835 3715 -805
rect 3765 -835 3795 -805
rect 3845 -835 3875 -805
rect 3925 -835 3955 -805
rect 4005 -835 4035 -805
rect 4085 -835 4115 -805
rect 4165 -835 4195 -805
rect 4245 -835 4275 -805
rect 4325 -835 4355 -805
rect 4405 -835 4435 -805
rect 4485 -835 4515 -805
rect 4565 -835 4595 -805
rect 4645 -835 4675 -805
rect 4725 -835 4755 -805
rect 4805 -835 4835 -805
rect 4885 -835 4915 -805
rect 4965 -835 4995 -805
rect 5045 -835 5075 -805
rect 5125 -835 5155 -805
rect 5205 -835 5235 -805
rect 5285 -835 5315 -805
rect 5365 -835 5395 -805
rect 5445 -835 5475 -805
rect 5525 -835 5555 -805
rect 5605 -835 5635 -805
rect 5685 -835 5715 -805
rect 5765 -835 5795 -805
rect 5845 -835 5875 -805
rect 5925 -835 5955 -805
rect 6005 -835 6035 -805
rect 6085 -835 6115 -805
rect 6165 -835 6195 -805
rect 6245 -835 6275 -805
rect 6325 -835 6355 -805
rect 6405 -835 6435 -805
rect 6485 -835 6515 -805
rect 6565 -835 6595 -805
rect 6645 -835 6675 -805
rect 6725 -835 6755 -805
rect 6805 -835 6835 -805
rect 6885 -835 6915 -805
rect 6965 -835 6995 -805
rect 7045 -835 7075 -805
rect 7125 -835 7155 -805
rect 7205 -835 7235 -805
rect 7285 -835 7315 -805
rect 7365 -835 7395 -805
rect 7445 -835 7475 -805
rect 7525 -835 7555 -805
rect 7605 -835 7635 -805
rect 7685 -835 7715 -805
rect 7765 -835 7795 -805
rect 7845 -835 7875 -805
rect 7925 -835 7955 -805
rect 8005 -835 8035 -805
rect 8085 -835 8115 -805
rect 8165 -835 8195 -805
rect 8245 -835 8275 -805
rect 8325 -835 8355 -805
rect 8405 -835 8435 -805
rect 8485 -835 8515 -805
rect 8565 -835 8595 -805
rect 8645 -835 8675 -805
rect 8725 -835 8755 -805
rect 8805 -835 8835 -805
rect 8885 -835 8915 -805
rect 8965 -835 8995 -805
rect 9045 -835 9075 -805
rect 9125 -835 9155 -805
rect 9205 -835 9235 -805
rect 9285 -835 9315 -805
rect 9365 -835 9395 -805
rect 9445 -835 9475 -805
rect 9525 -835 9555 -805
rect 9605 -835 9635 -805
rect 9685 -835 9715 -805
rect 9765 -835 9795 -805
rect 9845 -835 9875 -805
rect 9925 -835 9955 -805
rect 10005 -835 10035 -805
rect 10085 -835 10115 -805
rect 10165 -835 10195 -805
rect 10245 -835 10275 -805
rect 10325 -835 10355 -805
rect 10405 -835 10435 -805
rect 10485 -835 10515 -805
rect 10565 -835 10595 -805
rect 10645 -835 10675 -805
rect 10805 -835 10835 -805
rect 10965 -835 10995 -805
rect -715 -915 -685 -885
rect -555 -915 -525 -885
rect -395 -915 -365 -885
rect -235 -915 -205 -885
rect -155 -915 -125 -885
rect -75 -915 -45 -885
rect 5 -915 35 -885
rect 85 -915 115 -885
rect 165 -915 195 -885
rect 245 -915 275 -885
rect 325 -915 355 -885
rect 405 -915 435 -885
rect 485 -915 515 -885
rect 565 -915 595 -885
rect 645 -915 675 -885
rect 725 -915 755 -885
rect 805 -915 835 -885
rect 885 -915 915 -885
rect 965 -915 995 -885
rect 1045 -915 1075 -885
rect 1125 -915 1155 -885
rect 1205 -915 1235 -885
rect 1285 -915 1315 -885
rect 1365 -915 1395 -885
rect 1445 -915 1475 -885
rect 1525 -915 1555 -885
rect 1605 -915 1635 -885
rect 1685 -915 1715 -885
rect 1765 -915 1795 -885
rect 1845 -915 1875 -885
rect 1925 -915 1955 -885
rect 2005 -915 2035 -885
rect 2085 -915 2115 -885
rect 2165 -915 2195 -885
rect 2245 -915 2275 -885
rect 2325 -915 2355 -885
rect 2405 -915 2435 -885
rect 2485 -915 2515 -885
rect 2565 -915 2595 -885
rect 2645 -915 2675 -885
rect 2725 -915 2755 -885
rect 2805 -915 2835 -885
rect 2885 -915 2915 -885
rect 2965 -915 2995 -885
rect 3045 -915 3075 -885
rect 3125 -915 3155 -885
rect 3205 -915 3235 -885
rect 3285 -915 3315 -885
rect 3365 -915 3395 -885
rect 3445 -915 3475 -885
rect 3525 -915 3555 -885
rect 3605 -915 3635 -885
rect 3685 -915 3715 -885
rect 3765 -915 3795 -885
rect 3845 -915 3875 -885
rect 3925 -915 3955 -885
rect 4005 -915 4035 -885
rect 4085 -915 4115 -885
rect 4165 -915 4195 -885
rect 4245 -915 4275 -885
rect 4325 -915 4355 -885
rect 4405 -915 4435 -885
rect 4485 -915 4515 -885
rect 4565 -915 4595 -885
rect 4645 -915 4675 -885
rect 4725 -915 4755 -885
rect 4805 -915 4835 -885
rect 4885 -915 4915 -885
rect 4965 -915 4995 -885
rect 5045 -915 5075 -885
rect 5125 -915 5155 -885
rect 5205 -915 5235 -885
rect 5285 -915 5315 -885
rect 5365 -915 5395 -885
rect 5445 -915 5475 -885
rect 5525 -915 5555 -885
rect 5605 -915 5635 -885
rect 5685 -915 5715 -885
rect 5765 -915 5795 -885
rect 5845 -915 5875 -885
rect 5925 -915 5955 -885
rect 6005 -915 6035 -885
rect 6085 -915 6115 -885
rect 6165 -915 6195 -885
rect 6245 -915 6275 -885
rect 6325 -915 6355 -885
rect 6405 -915 6435 -885
rect 6485 -915 6515 -885
rect 6565 -915 6595 -885
rect 6645 -915 6675 -885
rect 6725 -915 6755 -885
rect 6805 -915 6835 -885
rect 6885 -915 6915 -885
rect 6965 -915 6995 -885
rect 7045 -915 7075 -885
rect 7125 -915 7155 -885
rect 7205 -915 7235 -885
rect 7285 -915 7315 -885
rect 7365 -915 7395 -885
rect 7445 -915 7475 -885
rect 7525 -915 7555 -885
rect 7605 -915 7635 -885
rect 7685 -915 7715 -885
rect 7765 -915 7795 -885
rect 7845 -915 7875 -885
rect 7925 -915 7955 -885
rect 8005 -915 8035 -885
rect 8085 -915 8115 -885
rect 8165 -915 8195 -885
rect 8245 -915 8275 -885
rect 8325 -915 8355 -885
rect 8405 -915 8435 -885
rect 8485 -915 8515 -885
rect 8565 -915 8595 -885
rect 8645 -915 8675 -885
rect 8725 -915 8755 -885
rect 8805 -915 8835 -885
rect 8885 -915 8915 -885
rect 8965 -915 8995 -885
rect 9045 -915 9075 -885
rect 9125 -915 9155 -885
rect 9205 -915 9235 -885
rect 9285 -915 9315 -885
rect 9365 -915 9395 -885
rect 9445 -915 9475 -885
rect 9525 -915 9555 -885
rect 9605 -915 9635 -885
rect 9685 -915 9715 -885
rect 9765 -915 9795 -885
rect 9845 -915 9875 -885
rect 9925 -915 9955 -885
rect 10005 -915 10035 -885
rect 10085 -915 10115 -885
rect 10165 -915 10195 -885
rect 10245 -915 10275 -885
rect 10325 -915 10355 -885
rect 10405 -915 10435 -885
rect 10485 -915 10515 -885
rect 10565 -915 10595 -885
rect 10645 -915 10675 -885
rect 10805 -915 10835 -885
rect 10965 -915 10995 -885
rect -635 -995 -605 -965
rect 10645 -995 10675 -965
rect 10805 -995 10835 -965
rect 10965 -995 10995 -965
rect -635 -1075 -605 -1045
rect 10645 -1075 10675 -1045
rect 10805 -1075 10835 -1045
rect 10965 -1075 10995 -1045
rect -715 -1155 -685 -1125
rect -555 -1155 -525 -1125
rect -395 -1155 -365 -1125
rect -235 -1155 -205 -1125
rect -155 -1155 -125 -1125
rect -75 -1155 -45 -1125
rect 5 -1155 35 -1125
rect 85 -1155 115 -1125
rect 165 -1155 195 -1125
rect 245 -1155 275 -1125
rect 325 -1155 355 -1125
rect 405 -1155 435 -1125
rect 485 -1155 515 -1125
rect 565 -1155 595 -1125
rect 645 -1155 675 -1125
rect 725 -1155 755 -1125
rect 805 -1155 835 -1125
rect 885 -1155 915 -1125
rect 965 -1155 995 -1125
rect 1045 -1155 1075 -1125
rect 1125 -1155 1155 -1125
rect 1205 -1155 1235 -1125
rect 1285 -1155 1315 -1125
rect 1365 -1155 1395 -1125
rect 1445 -1155 1475 -1125
rect 1525 -1155 1555 -1125
rect 1605 -1155 1635 -1125
rect 1685 -1155 1715 -1125
rect 1765 -1155 1795 -1125
rect 1845 -1155 1875 -1125
rect 1925 -1155 1955 -1125
rect 2005 -1155 2035 -1125
rect 2085 -1155 2115 -1125
rect 2165 -1155 2195 -1125
rect 2245 -1155 2275 -1125
rect 2325 -1155 2355 -1125
rect 2405 -1155 2435 -1125
rect 2485 -1155 2515 -1125
rect 2565 -1155 2595 -1125
rect 2645 -1155 2675 -1125
rect 2725 -1155 2755 -1125
rect 2805 -1155 2835 -1125
rect 2885 -1155 2915 -1125
rect 2965 -1155 2995 -1125
rect 3045 -1155 3075 -1125
rect 3125 -1155 3155 -1125
rect 3205 -1155 3235 -1125
rect 3285 -1155 3315 -1125
rect 3365 -1155 3395 -1125
rect 3445 -1155 3475 -1125
rect 3525 -1155 3555 -1125
rect 3605 -1155 3635 -1125
rect 3685 -1155 3715 -1125
rect 3765 -1155 3795 -1125
rect 3845 -1155 3875 -1125
rect 3925 -1155 3955 -1125
rect 4005 -1155 4035 -1125
rect 4085 -1155 4115 -1125
rect 4165 -1155 4195 -1125
rect 4245 -1155 4275 -1125
rect 4325 -1155 4355 -1125
rect 4405 -1155 4435 -1125
rect 4485 -1155 4515 -1125
rect 4565 -1155 4595 -1125
rect 4645 -1155 4675 -1125
rect 4725 -1155 4755 -1125
rect 4805 -1155 4835 -1125
rect 4885 -1155 4915 -1125
rect 4965 -1155 4995 -1125
rect 5045 -1155 5075 -1125
rect 5125 -1155 5155 -1125
rect 5205 -1155 5235 -1125
rect 5285 -1155 5315 -1125
rect 5365 -1155 5395 -1125
rect 5445 -1155 5475 -1125
rect 5525 -1155 5555 -1125
rect 5605 -1155 5635 -1125
rect 5685 -1155 5715 -1125
rect 5765 -1155 5795 -1125
rect 5845 -1155 5875 -1125
rect 5925 -1155 5955 -1125
rect 6005 -1155 6035 -1125
rect 6085 -1155 6115 -1125
rect 6165 -1155 6195 -1125
rect 6245 -1155 6275 -1125
rect 6325 -1155 6355 -1125
rect 6405 -1155 6435 -1125
rect 6485 -1155 6515 -1125
rect 6565 -1155 6595 -1125
rect 6645 -1155 6675 -1125
rect 6725 -1155 6755 -1125
rect 6805 -1155 6835 -1125
rect 6885 -1155 6915 -1125
rect 6965 -1155 6995 -1125
rect 7045 -1155 7075 -1125
rect 7125 -1155 7155 -1125
rect 7205 -1155 7235 -1125
rect 7285 -1155 7315 -1125
rect 7365 -1155 7395 -1125
rect 7445 -1155 7475 -1125
rect 7525 -1155 7555 -1125
rect 7605 -1155 7635 -1125
rect 7685 -1155 7715 -1125
rect 7765 -1155 7795 -1125
rect 7845 -1155 7875 -1125
rect 7925 -1155 7955 -1125
rect 8005 -1155 8035 -1125
rect 8085 -1155 8115 -1125
rect 8165 -1155 8195 -1125
rect 8245 -1155 8275 -1125
rect 8325 -1155 8355 -1125
rect 8405 -1155 8435 -1125
rect 8485 -1155 8515 -1125
rect 8565 -1155 8595 -1125
rect 8645 -1155 8675 -1125
rect 8725 -1155 8755 -1125
rect 8805 -1155 8835 -1125
rect 8885 -1155 8915 -1125
rect 8965 -1155 8995 -1125
rect 9045 -1155 9075 -1125
rect 9125 -1155 9155 -1125
rect 9205 -1155 9235 -1125
rect 9285 -1155 9315 -1125
rect 9365 -1155 9395 -1125
rect 9445 -1155 9475 -1125
rect 9525 -1155 9555 -1125
rect 9605 -1155 9635 -1125
rect 9685 -1155 9715 -1125
rect 9765 -1155 9795 -1125
rect 9845 -1155 9875 -1125
rect 9925 -1155 9955 -1125
rect 10005 -1155 10035 -1125
rect 10085 -1155 10115 -1125
rect 10165 -1155 10195 -1125
rect 10245 -1155 10275 -1125
rect 10325 -1155 10355 -1125
rect 10405 -1155 10435 -1125
rect 10485 -1155 10515 -1125
rect 10565 -1155 10595 -1125
rect 10645 -1155 10675 -1125
rect 10805 -1155 10835 -1125
rect 10965 -1155 10995 -1125
rect -715 -1235 -685 -1205
rect -555 -1235 -525 -1205
rect -395 -1235 -365 -1205
rect -235 -1235 -205 -1205
rect -155 -1235 -125 -1205
rect -75 -1235 -45 -1205
rect 5 -1235 35 -1205
rect 85 -1235 115 -1205
rect 165 -1235 195 -1205
rect 245 -1235 275 -1205
rect 325 -1235 355 -1205
rect 405 -1235 435 -1205
rect 485 -1235 515 -1205
rect 565 -1235 595 -1205
rect 645 -1235 675 -1205
rect 725 -1235 755 -1205
rect 805 -1235 835 -1205
rect 885 -1235 915 -1205
rect 965 -1235 995 -1205
rect 1045 -1235 1075 -1205
rect 1125 -1235 1155 -1205
rect 1205 -1235 1235 -1205
rect 1285 -1235 1315 -1205
rect 1365 -1235 1395 -1205
rect 1445 -1235 1475 -1205
rect 1525 -1235 1555 -1205
rect 1605 -1235 1635 -1205
rect 1685 -1235 1715 -1205
rect 1765 -1235 1795 -1205
rect 1845 -1235 1875 -1205
rect 1925 -1235 1955 -1205
rect 2005 -1235 2035 -1205
rect 2085 -1235 2115 -1205
rect 2165 -1235 2195 -1205
rect 2245 -1235 2275 -1205
rect 2325 -1235 2355 -1205
rect 2405 -1235 2435 -1205
rect 2485 -1235 2515 -1205
rect 2565 -1235 2595 -1205
rect 2645 -1235 2675 -1205
rect 2725 -1235 2755 -1205
rect 2805 -1235 2835 -1205
rect 2885 -1235 2915 -1205
rect 2965 -1235 2995 -1205
rect 3045 -1235 3075 -1205
rect 3125 -1235 3155 -1205
rect 3205 -1235 3235 -1205
rect 3285 -1235 3315 -1205
rect 3365 -1235 3395 -1205
rect 3445 -1235 3475 -1205
rect 3525 -1235 3555 -1205
rect 3605 -1235 3635 -1205
rect 3685 -1235 3715 -1205
rect 3765 -1235 3795 -1205
rect 3845 -1235 3875 -1205
rect 3925 -1235 3955 -1205
rect 4005 -1235 4035 -1205
rect 4085 -1235 4115 -1205
rect 4165 -1235 4195 -1205
rect 4245 -1235 4275 -1205
rect 4325 -1235 4355 -1205
rect 4405 -1235 4435 -1205
rect 4485 -1235 4515 -1205
rect 4565 -1235 4595 -1205
rect 4645 -1235 4675 -1205
rect 4725 -1235 4755 -1205
rect 4805 -1235 4835 -1205
rect 4885 -1235 4915 -1205
rect 4965 -1235 4995 -1205
rect 5045 -1235 5075 -1205
rect 5125 -1235 5155 -1205
rect 5205 -1235 5235 -1205
rect 5285 -1235 5315 -1205
rect 5365 -1235 5395 -1205
rect 5445 -1235 5475 -1205
rect 5525 -1235 5555 -1205
rect 5605 -1235 5635 -1205
rect 5685 -1235 5715 -1205
rect 5765 -1235 5795 -1205
rect 5845 -1235 5875 -1205
rect 5925 -1235 5955 -1205
rect 6005 -1235 6035 -1205
rect 6085 -1235 6115 -1205
rect 6165 -1235 6195 -1205
rect 6245 -1235 6275 -1205
rect 6325 -1235 6355 -1205
rect 6405 -1235 6435 -1205
rect 6485 -1235 6515 -1205
rect 6565 -1235 6595 -1205
rect 6645 -1235 6675 -1205
rect 6725 -1235 6755 -1205
rect 6805 -1235 6835 -1205
rect 6885 -1235 6915 -1205
rect 6965 -1235 6995 -1205
rect 7045 -1235 7075 -1205
rect 7125 -1235 7155 -1205
rect 7205 -1235 7235 -1205
rect 7285 -1235 7315 -1205
rect 7365 -1235 7395 -1205
rect 7445 -1235 7475 -1205
rect 7525 -1235 7555 -1205
rect 7605 -1235 7635 -1205
rect 7685 -1235 7715 -1205
rect 7765 -1235 7795 -1205
rect 7845 -1235 7875 -1205
rect 7925 -1235 7955 -1205
rect 8005 -1235 8035 -1205
rect 8085 -1235 8115 -1205
rect 8165 -1235 8195 -1205
rect 8245 -1235 8275 -1205
rect 8325 -1235 8355 -1205
rect 8405 -1235 8435 -1205
rect 8485 -1235 8515 -1205
rect 8565 -1235 8595 -1205
rect 8645 -1235 8675 -1205
rect 8725 -1235 8755 -1205
rect 8805 -1235 8835 -1205
rect 8885 -1235 8915 -1205
rect 8965 -1235 8995 -1205
rect 9045 -1235 9075 -1205
rect 9125 -1235 9155 -1205
rect 9205 -1235 9235 -1205
rect 9285 -1235 9315 -1205
rect 9365 -1235 9395 -1205
rect 9445 -1235 9475 -1205
rect 9525 -1235 9555 -1205
rect 9605 -1235 9635 -1205
rect 9685 -1235 9715 -1205
rect 9765 -1235 9795 -1205
rect 9845 -1235 9875 -1205
rect 9925 -1235 9955 -1205
rect 10005 -1235 10035 -1205
rect 10085 -1235 10115 -1205
rect 10165 -1235 10195 -1205
rect 10245 -1235 10275 -1205
rect 10325 -1235 10355 -1205
rect 10405 -1235 10435 -1205
rect 10485 -1235 10515 -1205
rect 10565 -1235 10595 -1205
rect 10645 -1235 10675 -1205
rect 10805 -1235 10835 -1205
rect 10965 -1235 10995 -1205
rect -715 -1315 -685 -1285
rect -555 -1315 -525 -1285
rect -395 -1315 -365 -1285
rect -235 -1315 -205 -1285
rect -155 -1315 -125 -1285
rect -75 -1315 -45 -1285
rect 5 -1315 35 -1285
rect 85 -1315 115 -1285
rect 165 -1315 195 -1285
rect 245 -1315 275 -1285
rect 325 -1315 355 -1285
rect 405 -1315 435 -1285
rect 485 -1315 515 -1285
rect 565 -1315 595 -1285
rect 645 -1315 675 -1285
rect 725 -1315 755 -1285
rect 805 -1315 835 -1285
rect 885 -1315 915 -1285
rect 965 -1315 995 -1285
rect 1045 -1315 1075 -1285
rect 1125 -1315 1155 -1285
rect 1205 -1315 1235 -1285
rect 1285 -1315 1315 -1285
rect 1365 -1315 1395 -1285
rect 1445 -1315 1475 -1285
rect 1525 -1315 1555 -1285
rect 1605 -1315 1635 -1285
rect 1685 -1315 1715 -1285
rect 1765 -1315 1795 -1285
rect 1845 -1315 1875 -1285
rect 1925 -1315 1955 -1285
rect 2005 -1315 2035 -1285
rect 2085 -1315 2115 -1285
rect 2165 -1315 2195 -1285
rect 2245 -1315 2275 -1285
rect 2325 -1315 2355 -1285
rect 2405 -1315 2435 -1285
rect 2485 -1315 2515 -1285
rect 2565 -1315 2595 -1285
rect 2645 -1315 2675 -1285
rect 2725 -1315 2755 -1285
rect 2805 -1315 2835 -1285
rect 2885 -1315 2915 -1285
rect 2965 -1315 2995 -1285
rect 3045 -1315 3075 -1285
rect 3125 -1315 3155 -1285
rect 3205 -1315 3235 -1285
rect 3285 -1315 3315 -1285
rect 3365 -1315 3395 -1285
rect 3445 -1315 3475 -1285
rect 3525 -1315 3555 -1285
rect 3605 -1315 3635 -1285
rect 3685 -1315 3715 -1285
rect 3765 -1315 3795 -1285
rect 3845 -1315 3875 -1285
rect 3925 -1315 3955 -1285
rect 4005 -1315 4035 -1285
rect 4085 -1315 4115 -1285
rect 4165 -1315 4195 -1285
rect 4245 -1315 4275 -1285
rect 4325 -1315 4355 -1285
rect 4405 -1315 4435 -1285
rect 4485 -1315 4515 -1285
rect 4565 -1315 4595 -1285
rect 4645 -1315 4675 -1285
rect 4725 -1315 4755 -1285
rect 4805 -1315 4835 -1285
rect 4885 -1315 4915 -1285
rect 4965 -1315 4995 -1285
rect 5045 -1315 5075 -1285
rect 5125 -1315 5155 -1285
rect 5205 -1315 5235 -1285
rect 5285 -1315 5315 -1285
rect 5365 -1315 5395 -1285
rect 5445 -1315 5475 -1285
rect 5525 -1315 5555 -1285
rect 5605 -1315 5635 -1285
rect 5685 -1315 5715 -1285
rect 5765 -1315 5795 -1285
rect 5845 -1315 5875 -1285
rect 5925 -1315 5955 -1285
rect 6005 -1315 6035 -1285
rect 6085 -1315 6115 -1285
rect 6165 -1315 6195 -1285
rect 6245 -1315 6275 -1285
rect 6325 -1315 6355 -1285
rect 6405 -1315 6435 -1285
rect 6485 -1315 6515 -1285
rect 6565 -1315 6595 -1285
rect 6645 -1315 6675 -1285
rect 6725 -1315 6755 -1285
rect 6805 -1315 6835 -1285
rect 6885 -1315 6915 -1285
rect 6965 -1315 6995 -1285
rect 7045 -1315 7075 -1285
rect 7125 -1315 7155 -1285
rect 7205 -1315 7235 -1285
rect 7285 -1315 7315 -1285
rect 7365 -1315 7395 -1285
rect 7445 -1315 7475 -1285
rect 7525 -1315 7555 -1285
rect 7605 -1315 7635 -1285
rect 7685 -1315 7715 -1285
rect 7765 -1315 7795 -1285
rect 7845 -1315 7875 -1285
rect 7925 -1315 7955 -1285
rect 8005 -1315 8035 -1285
rect 8085 -1315 8115 -1285
rect 8165 -1315 8195 -1285
rect 8245 -1315 8275 -1285
rect 8325 -1315 8355 -1285
rect 8405 -1315 8435 -1285
rect 8485 -1315 8515 -1285
rect 8565 -1315 8595 -1285
rect 8645 -1315 8675 -1285
rect 8725 -1315 8755 -1285
rect 8805 -1315 8835 -1285
rect 8885 -1315 8915 -1285
rect 8965 -1315 8995 -1285
rect 9045 -1315 9075 -1285
rect 9125 -1315 9155 -1285
rect 9205 -1315 9235 -1285
rect 9285 -1315 9315 -1285
rect 9365 -1315 9395 -1285
rect 9445 -1315 9475 -1285
rect 9525 -1315 9555 -1285
rect 9605 -1315 9635 -1285
rect 9685 -1315 9715 -1285
rect 9765 -1315 9795 -1285
rect 9845 -1315 9875 -1285
rect 9925 -1315 9955 -1285
rect 10005 -1315 10035 -1285
rect 10085 -1315 10115 -1285
rect 10165 -1315 10195 -1285
rect 10245 -1315 10275 -1285
rect 10325 -1315 10355 -1285
rect 10405 -1315 10435 -1285
rect 10485 -1315 10515 -1285
rect 10565 -1315 10595 -1285
rect 10645 -1315 10675 -1285
rect 10805 -1315 10835 -1285
rect 10965 -1315 10995 -1285
rect -715 -1395 -685 -1365
rect -555 -1395 -525 -1365
rect -395 -1395 -365 -1365
rect -235 -1395 -205 -1365
rect -155 -1395 -125 -1365
rect -75 -1395 -45 -1365
rect 5 -1395 35 -1365
rect 85 -1395 115 -1365
rect 165 -1395 195 -1365
rect 245 -1395 275 -1365
rect 325 -1395 355 -1365
rect 405 -1395 435 -1365
rect 485 -1395 515 -1365
rect 565 -1395 595 -1365
rect 645 -1395 675 -1365
rect 725 -1395 755 -1365
rect 805 -1395 835 -1365
rect 885 -1395 915 -1365
rect 965 -1395 995 -1365
rect 1045 -1395 1075 -1365
rect 1125 -1395 1155 -1365
rect 1205 -1395 1235 -1365
rect 1285 -1395 1315 -1365
rect 1365 -1395 1395 -1365
rect 1445 -1395 1475 -1365
rect 1525 -1395 1555 -1365
rect 1605 -1395 1635 -1365
rect 1685 -1395 1715 -1365
rect 1765 -1395 1795 -1365
rect 1845 -1395 1875 -1365
rect 1925 -1395 1955 -1365
rect 2005 -1395 2035 -1365
rect 2085 -1395 2115 -1365
rect 2165 -1395 2195 -1365
rect 2245 -1395 2275 -1365
rect 2325 -1395 2355 -1365
rect 2405 -1395 2435 -1365
rect 2485 -1395 2515 -1365
rect 2565 -1395 2595 -1365
rect 2645 -1395 2675 -1365
rect 2725 -1395 2755 -1365
rect 2805 -1395 2835 -1365
rect 2885 -1395 2915 -1365
rect 2965 -1395 2995 -1365
rect 3045 -1395 3075 -1365
rect 3125 -1395 3155 -1365
rect 3205 -1395 3235 -1365
rect 3285 -1395 3315 -1365
rect 3365 -1395 3395 -1365
rect 3445 -1395 3475 -1365
rect 3525 -1395 3555 -1365
rect 3605 -1395 3635 -1365
rect 3685 -1395 3715 -1365
rect 3765 -1395 3795 -1365
rect 3845 -1395 3875 -1365
rect 3925 -1395 3955 -1365
rect 4005 -1395 4035 -1365
rect 4085 -1395 4115 -1365
rect 4165 -1395 4195 -1365
rect 4245 -1395 4275 -1365
rect 4325 -1395 4355 -1365
rect 4405 -1395 4435 -1365
rect 4485 -1395 4515 -1365
rect 4565 -1395 4595 -1365
rect 4645 -1395 4675 -1365
rect 4725 -1395 4755 -1365
rect 4805 -1395 4835 -1365
rect 4885 -1395 4915 -1365
rect 4965 -1395 4995 -1365
rect 5045 -1395 5075 -1365
rect 5125 -1395 5155 -1365
rect 5205 -1395 5235 -1365
rect 5285 -1395 5315 -1365
rect 5365 -1395 5395 -1365
rect 5445 -1395 5475 -1365
rect 5525 -1395 5555 -1365
rect 5605 -1395 5635 -1365
rect 5685 -1395 5715 -1365
rect 5765 -1395 5795 -1365
rect 5845 -1395 5875 -1365
rect 5925 -1395 5955 -1365
rect 6005 -1395 6035 -1365
rect 6085 -1395 6115 -1365
rect 6165 -1395 6195 -1365
rect 6245 -1395 6275 -1365
rect 6325 -1395 6355 -1365
rect 6405 -1395 6435 -1365
rect 6485 -1395 6515 -1365
rect 6565 -1395 6595 -1365
rect 6645 -1395 6675 -1365
rect 6725 -1395 6755 -1365
rect 6805 -1395 6835 -1365
rect 6885 -1395 6915 -1365
rect 6965 -1395 6995 -1365
rect 7045 -1395 7075 -1365
rect 7125 -1395 7155 -1365
rect 7205 -1395 7235 -1365
rect 7285 -1395 7315 -1365
rect 7365 -1395 7395 -1365
rect 7445 -1395 7475 -1365
rect 7525 -1395 7555 -1365
rect 7605 -1395 7635 -1365
rect 7685 -1395 7715 -1365
rect 7765 -1395 7795 -1365
rect 7845 -1395 7875 -1365
rect 7925 -1395 7955 -1365
rect 8005 -1395 8035 -1365
rect 8085 -1395 8115 -1365
rect 8165 -1395 8195 -1365
rect 8245 -1395 8275 -1365
rect 8325 -1395 8355 -1365
rect 8405 -1395 8435 -1365
rect 8485 -1395 8515 -1365
rect 8565 -1395 8595 -1365
rect 8645 -1395 8675 -1365
rect 8725 -1395 8755 -1365
rect 8805 -1395 8835 -1365
rect 8885 -1395 8915 -1365
rect 8965 -1395 8995 -1365
rect 9045 -1395 9075 -1365
rect 9125 -1395 9155 -1365
rect 9205 -1395 9235 -1365
rect 9285 -1395 9315 -1365
rect 9365 -1395 9395 -1365
rect 9445 -1395 9475 -1365
rect 9525 -1395 9555 -1365
rect 9605 -1395 9635 -1365
rect 9685 -1395 9715 -1365
rect 9765 -1395 9795 -1365
rect 9845 -1395 9875 -1365
rect 9925 -1395 9955 -1365
rect 10005 -1395 10035 -1365
rect 10085 -1395 10115 -1365
rect 10165 -1395 10195 -1365
rect 10245 -1395 10275 -1365
rect 10325 -1395 10355 -1365
rect 10405 -1395 10435 -1365
rect 10485 -1395 10515 -1365
rect 10565 -1395 10595 -1365
rect 10645 -1395 10675 -1365
rect 10805 -1395 10835 -1365
rect 10965 -1395 10995 -1365
rect -715 -1475 -685 -1445
rect -555 -1475 -525 -1445
rect -395 -1475 -365 -1445
rect -235 -1475 -205 -1445
rect -155 -1475 -125 -1445
rect -75 -1475 -45 -1445
rect 5 -1475 35 -1445
rect 85 -1475 115 -1445
rect 165 -1475 195 -1445
rect 245 -1475 275 -1445
rect 325 -1475 355 -1445
rect 405 -1475 435 -1445
rect 485 -1475 515 -1445
rect 565 -1475 595 -1445
rect 645 -1475 675 -1445
rect 725 -1475 755 -1445
rect 805 -1475 835 -1445
rect 885 -1475 915 -1445
rect 965 -1475 995 -1445
rect 1045 -1475 1075 -1445
rect 1125 -1475 1155 -1445
rect 1205 -1475 1235 -1445
rect 1285 -1475 1315 -1445
rect 1365 -1475 1395 -1445
rect 1445 -1475 1475 -1445
rect 1525 -1475 1555 -1445
rect 1605 -1475 1635 -1445
rect 1685 -1475 1715 -1445
rect 1765 -1475 1795 -1445
rect 1845 -1475 1875 -1445
rect 1925 -1475 1955 -1445
rect 2005 -1475 2035 -1445
rect 2085 -1475 2115 -1445
rect 2165 -1475 2195 -1445
rect 2245 -1475 2275 -1445
rect 2325 -1475 2355 -1445
rect 2405 -1475 2435 -1445
rect 2485 -1475 2515 -1445
rect 2565 -1475 2595 -1445
rect 2645 -1475 2675 -1445
rect 2725 -1475 2755 -1445
rect 2805 -1475 2835 -1445
rect 2885 -1475 2915 -1445
rect 2965 -1475 2995 -1445
rect 3045 -1475 3075 -1445
rect 3125 -1475 3155 -1445
rect 3205 -1475 3235 -1445
rect 3285 -1475 3315 -1445
rect 3365 -1475 3395 -1445
rect 3445 -1475 3475 -1445
rect 3525 -1475 3555 -1445
rect 3605 -1475 3635 -1445
rect 3685 -1475 3715 -1445
rect 3765 -1475 3795 -1445
rect 3845 -1475 3875 -1445
rect 3925 -1475 3955 -1445
rect 4005 -1475 4035 -1445
rect 4085 -1475 4115 -1445
rect 4165 -1475 4195 -1445
rect 4245 -1475 4275 -1445
rect 4325 -1475 4355 -1445
rect 4405 -1475 4435 -1445
rect 4485 -1475 4515 -1445
rect 4565 -1475 4595 -1445
rect 4645 -1475 4675 -1445
rect 4725 -1475 4755 -1445
rect 4805 -1475 4835 -1445
rect 4885 -1475 4915 -1445
rect 4965 -1475 4995 -1445
rect 5045 -1475 5075 -1445
rect 5125 -1475 5155 -1445
rect 5205 -1475 5235 -1445
rect 5285 -1475 5315 -1445
rect 5365 -1475 5395 -1445
rect 5445 -1475 5475 -1445
rect 5525 -1475 5555 -1445
rect 5605 -1475 5635 -1445
rect 5685 -1475 5715 -1445
rect 5765 -1475 5795 -1445
rect 5845 -1475 5875 -1445
rect 5925 -1475 5955 -1445
rect 6005 -1475 6035 -1445
rect 6085 -1475 6115 -1445
rect 6165 -1475 6195 -1445
rect 6245 -1475 6275 -1445
rect 6325 -1475 6355 -1445
rect 6405 -1475 6435 -1445
rect 6485 -1475 6515 -1445
rect 6565 -1475 6595 -1445
rect 6645 -1475 6675 -1445
rect 6725 -1475 6755 -1445
rect 6805 -1475 6835 -1445
rect 6885 -1475 6915 -1445
rect 6965 -1475 6995 -1445
rect 7045 -1475 7075 -1445
rect 7125 -1475 7155 -1445
rect 7205 -1475 7235 -1445
rect 7285 -1475 7315 -1445
rect 7365 -1475 7395 -1445
rect 7445 -1475 7475 -1445
rect 7525 -1475 7555 -1445
rect 7605 -1475 7635 -1445
rect 7685 -1475 7715 -1445
rect 7765 -1475 7795 -1445
rect 7845 -1475 7875 -1445
rect 7925 -1475 7955 -1445
rect 8005 -1475 8035 -1445
rect 8085 -1475 8115 -1445
rect 8165 -1475 8195 -1445
rect 8245 -1475 8275 -1445
rect 8325 -1475 8355 -1445
rect 8405 -1475 8435 -1445
rect 8485 -1475 8515 -1445
rect 8565 -1475 8595 -1445
rect 8645 -1475 8675 -1445
rect 8725 -1475 8755 -1445
rect 8805 -1475 8835 -1445
rect 8885 -1475 8915 -1445
rect 8965 -1475 8995 -1445
rect 9045 -1475 9075 -1445
rect 9125 -1475 9155 -1445
rect 9205 -1475 9235 -1445
rect 9285 -1475 9315 -1445
rect 9365 -1475 9395 -1445
rect 9445 -1475 9475 -1445
rect 9525 -1475 9555 -1445
rect 9605 -1475 9635 -1445
rect 9685 -1475 9715 -1445
rect 9765 -1475 9795 -1445
rect 9845 -1475 9875 -1445
rect 9925 -1475 9955 -1445
rect 10005 -1475 10035 -1445
rect 10085 -1475 10115 -1445
rect 10165 -1475 10195 -1445
rect 10245 -1475 10275 -1445
rect 10325 -1475 10355 -1445
rect 10405 -1475 10435 -1445
rect 10485 -1475 10515 -1445
rect 10565 -1475 10595 -1445
rect 10645 -1475 10675 -1445
rect 10805 -1475 10835 -1445
rect 10965 -1475 10995 -1445
rect -715 -1555 -685 -1525
rect -555 -1555 -525 -1525
rect -395 -1555 -365 -1525
rect -235 -1555 -205 -1525
rect -155 -1555 -125 -1525
rect -75 -1555 -45 -1525
rect 5 -1555 35 -1525
rect 85 -1555 115 -1525
rect 165 -1555 195 -1525
rect 245 -1555 275 -1525
rect 325 -1555 355 -1525
rect 405 -1555 435 -1525
rect 485 -1555 515 -1525
rect 565 -1555 595 -1525
rect 645 -1555 675 -1525
rect 725 -1555 755 -1525
rect 805 -1555 835 -1525
rect 885 -1555 915 -1525
rect 965 -1555 995 -1525
rect 1045 -1555 1075 -1525
rect 1125 -1555 1155 -1525
rect 1205 -1555 1235 -1525
rect 1285 -1555 1315 -1525
rect 1365 -1555 1395 -1525
rect 1445 -1555 1475 -1525
rect 1525 -1555 1555 -1525
rect 1605 -1555 1635 -1525
rect 1685 -1555 1715 -1525
rect 1765 -1555 1795 -1525
rect 1845 -1555 1875 -1525
rect 1925 -1555 1955 -1525
rect 2005 -1555 2035 -1525
rect 2085 -1555 2115 -1525
rect 2165 -1555 2195 -1525
rect 2245 -1555 2275 -1525
rect 2325 -1555 2355 -1525
rect 2405 -1555 2435 -1525
rect 2485 -1555 2515 -1525
rect 2565 -1555 2595 -1525
rect 2645 -1555 2675 -1525
rect 2725 -1555 2755 -1525
rect 2805 -1555 2835 -1525
rect 2885 -1555 2915 -1525
rect 2965 -1555 2995 -1525
rect 3045 -1555 3075 -1525
rect 3125 -1555 3155 -1525
rect 3205 -1555 3235 -1525
rect 3285 -1555 3315 -1525
rect 3365 -1555 3395 -1525
rect 3445 -1555 3475 -1525
rect 3525 -1555 3555 -1525
rect 3605 -1555 3635 -1525
rect 3685 -1555 3715 -1525
rect 3765 -1555 3795 -1525
rect 3845 -1555 3875 -1525
rect 3925 -1555 3955 -1525
rect 4005 -1555 4035 -1525
rect 4085 -1555 4115 -1525
rect 4165 -1555 4195 -1525
rect 4245 -1555 4275 -1525
rect 4325 -1555 4355 -1525
rect 4405 -1555 4435 -1525
rect 4485 -1555 4515 -1525
rect 4565 -1555 4595 -1525
rect 4645 -1555 4675 -1525
rect 4725 -1555 4755 -1525
rect 4805 -1555 4835 -1525
rect 4885 -1555 4915 -1525
rect 4965 -1555 4995 -1525
rect 5045 -1555 5075 -1525
rect 5125 -1555 5155 -1525
rect 5205 -1555 5235 -1525
rect 5285 -1555 5315 -1525
rect 5365 -1555 5395 -1525
rect 5445 -1555 5475 -1525
rect 5525 -1555 5555 -1525
rect 5605 -1555 5635 -1525
rect 5685 -1555 5715 -1525
rect 5765 -1555 5795 -1525
rect 5845 -1555 5875 -1525
rect 5925 -1555 5955 -1525
rect 6005 -1555 6035 -1525
rect 6085 -1555 6115 -1525
rect 6165 -1555 6195 -1525
rect 6245 -1555 6275 -1525
rect 6325 -1555 6355 -1525
rect 6405 -1555 6435 -1525
rect 6485 -1555 6515 -1525
rect 6565 -1555 6595 -1525
rect 6645 -1555 6675 -1525
rect 6725 -1555 6755 -1525
rect 6805 -1555 6835 -1525
rect 6885 -1555 6915 -1525
rect 6965 -1555 6995 -1525
rect 7045 -1555 7075 -1525
rect 7125 -1555 7155 -1525
rect 7205 -1555 7235 -1525
rect 7285 -1555 7315 -1525
rect 7365 -1555 7395 -1525
rect 7445 -1555 7475 -1525
rect 7525 -1555 7555 -1525
rect 7605 -1555 7635 -1525
rect 7685 -1555 7715 -1525
rect 7765 -1555 7795 -1525
rect 7845 -1555 7875 -1525
rect 7925 -1555 7955 -1525
rect 8005 -1555 8035 -1525
rect 8085 -1555 8115 -1525
rect 8165 -1555 8195 -1525
rect 8245 -1555 8275 -1525
rect 8325 -1555 8355 -1525
rect 8405 -1555 8435 -1525
rect 8485 -1555 8515 -1525
rect 8565 -1555 8595 -1525
rect 8645 -1555 8675 -1525
rect 8725 -1555 8755 -1525
rect 8805 -1555 8835 -1525
rect 8885 -1555 8915 -1525
rect 8965 -1555 8995 -1525
rect 9045 -1555 9075 -1525
rect 9125 -1555 9155 -1525
rect 9205 -1555 9235 -1525
rect 9285 -1555 9315 -1525
rect 9365 -1555 9395 -1525
rect 9445 -1555 9475 -1525
rect 9525 -1555 9555 -1525
rect 9605 -1555 9635 -1525
rect 9685 -1555 9715 -1525
rect 9765 -1555 9795 -1525
rect 9845 -1555 9875 -1525
rect 9925 -1555 9955 -1525
rect 10005 -1555 10035 -1525
rect 10085 -1555 10115 -1525
rect 10165 -1555 10195 -1525
rect 10245 -1555 10275 -1525
rect 10325 -1555 10355 -1525
rect 10405 -1555 10435 -1525
rect 10485 -1555 10515 -1525
rect 10565 -1555 10595 -1525
rect 10645 -1555 10675 -1525
rect 10805 -1555 10835 -1525
rect 10965 -1555 10995 -1525
rect -635 -1635 -605 -1605
rect 10645 -1635 10675 -1605
rect 10805 -1635 10835 -1605
rect 10965 -1635 10995 -1605
rect -635 -1715 -605 -1685
rect 10645 -1715 10675 -1685
rect 10805 -1715 10835 -1685
rect 10965 -1715 10995 -1685
rect -715 -1795 -685 -1765
rect -555 -1795 -525 -1765
rect -395 -1795 -365 -1765
rect -235 -1795 -205 -1765
rect -155 -1795 -125 -1765
rect -75 -1795 -45 -1765
rect 5 -1795 35 -1765
rect 85 -1795 115 -1765
rect 165 -1795 195 -1765
rect 245 -1795 275 -1765
rect 325 -1795 355 -1765
rect 405 -1795 435 -1765
rect 485 -1795 515 -1765
rect 565 -1795 595 -1765
rect 645 -1795 675 -1765
rect 725 -1795 755 -1765
rect 805 -1795 835 -1765
rect 885 -1795 915 -1765
rect 965 -1795 995 -1765
rect 1045 -1795 1075 -1765
rect 1125 -1795 1155 -1765
rect 1205 -1795 1235 -1765
rect 1285 -1795 1315 -1765
rect 1365 -1795 1395 -1765
rect 1445 -1795 1475 -1765
rect 1525 -1795 1555 -1765
rect 1605 -1795 1635 -1765
rect 1685 -1795 1715 -1765
rect 1765 -1795 1795 -1765
rect 1845 -1795 1875 -1765
rect 1925 -1795 1955 -1765
rect 2005 -1795 2035 -1765
rect 2085 -1795 2115 -1765
rect 2165 -1795 2195 -1765
rect 2245 -1795 2275 -1765
rect 2325 -1795 2355 -1765
rect 2405 -1795 2435 -1765
rect 2485 -1795 2515 -1765
rect 2565 -1795 2595 -1765
rect 2645 -1795 2675 -1765
rect 2725 -1795 2755 -1765
rect 2805 -1795 2835 -1765
rect 2885 -1795 2915 -1765
rect 2965 -1795 2995 -1765
rect 3045 -1795 3075 -1765
rect 3125 -1795 3155 -1765
rect 3205 -1795 3235 -1765
rect 3285 -1795 3315 -1765
rect 3365 -1795 3395 -1765
rect 3445 -1795 3475 -1765
rect 3525 -1795 3555 -1765
rect 3605 -1795 3635 -1765
rect 3685 -1795 3715 -1765
rect 3765 -1795 3795 -1765
rect 3845 -1795 3875 -1765
rect 3925 -1795 3955 -1765
rect 4005 -1795 4035 -1765
rect 4085 -1795 4115 -1765
rect 4165 -1795 4195 -1765
rect 4245 -1795 4275 -1765
rect 4325 -1795 4355 -1765
rect 4405 -1795 4435 -1765
rect 4485 -1795 4515 -1765
rect 4565 -1795 4595 -1765
rect 4645 -1795 4675 -1765
rect 4725 -1795 4755 -1765
rect 4805 -1795 4835 -1765
rect 4885 -1795 4915 -1765
rect 4965 -1795 4995 -1765
rect 5045 -1795 5075 -1765
rect 5125 -1795 5155 -1765
rect 5205 -1795 5235 -1765
rect 5285 -1795 5315 -1765
rect 5365 -1795 5395 -1765
rect 5445 -1795 5475 -1765
rect 5525 -1795 5555 -1765
rect 5605 -1795 5635 -1765
rect 5685 -1795 5715 -1765
rect 5765 -1795 5795 -1765
rect 5845 -1795 5875 -1765
rect 5925 -1795 5955 -1765
rect 6005 -1795 6035 -1765
rect 6085 -1795 6115 -1765
rect 6165 -1795 6195 -1765
rect 6245 -1795 6275 -1765
rect 6325 -1795 6355 -1765
rect 6405 -1795 6435 -1765
rect 6485 -1795 6515 -1765
rect 6565 -1795 6595 -1765
rect 6645 -1795 6675 -1765
rect 6725 -1795 6755 -1765
rect 6805 -1795 6835 -1765
rect 6885 -1795 6915 -1765
rect 6965 -1795 6995 -1765
rect 7045 -1795 7075 -1765
rect 7125 -1795 7155 -1765
rect 7205 -1795 7235 -1765
rect 7285 -1795 7315 -1765
rect 7365 -1795 7395 -1765
rect 7445 -1795 7475 -1765
rect 7525 -1795 7555 -1765
rect 7605 -1795 7635 -1765
rect 7685 -1795 7715 -1765
rect 7765 -1795 7795 -1765
rect 7845 -1795 7875 -1765
rect 7925 -1795 7955 -1765
rect 8005 -1795 8035 -1765
rect 8085 -1795 8115 -1765
rect 8165 -1795 8195 -1765
rect 8245 -1795 8275 -1765
rect 8325 -1795 8355 -1765
rect 8405 -1795 8435 -1765
rect 8485 -1795 8515 -1765
rect 8565 -1795 8595 -1765
rect 8645 -1795 8675 -1765
rect 8725 -1795 8755 -1765
rect 8805 -1795 8835 -1765
rect 8885 -1795 8915 -1765
rect 8965 -1795 8995 -1765
rect 9045 -1795 9075 -1765
rect 9125 -1795 9155 -1765
rect 9205 -1795 9235 -1765
rect 9285 -1795 9315 -1765
rect 9365 -1795 9395 -1765
rect 9445 -1795 9475 -1765
rect 9525 -1795 9555 -1765
rect 9605 -1795 9635 -1765
rect 9685 -1795 9715 -1765
rect 9765 -1795 9795 -1765
rect 9845 -1795 9875 -1765
rect 9925 -1795 9955 -1765
rect 10005 -1795 10035 -1765
rect 10085 -1795 10115 -1765
rect 10165 -1795 10195 -1765
rect 10245 -1795 10275 -1765
rect 10325 -1795 10355 -1765
rect 10405 -1795 10435 -1765
rect 10485 -1795 10515 -1765
rect 10565 -1795 10595 -1765
rect 10645 -1795 10675 -1765
rect 10805 -1795 10835 -1765
rect 10965 -1795 10995 -1765
rect -715 -1875 -685 -1845
rect -555 -1875 -525 -1845
rect -395 -1875 -365 -1845
rect -235 -1875 -205 -1845
rect -155 -1875 -125 -1845
rect -75 -1875 -45 -1845
rect 5 -1875 35 -1845
rect 85 -1875 115 -1845
rect 165 -1875 195 -1845
rect 245 -1875 275 -1845
rect 325 -1875 355 -1845
rect 405 -1875 435 -1845
rect 485 -1875 515 -1845
rect 565 -1875 595 -1845
rect 645 -1875 675 -1845
rect 725 -1875 755 -1845
rect 805 -1875 835 -1845
rect 885 -1875 915 -1845
rect 965 -1875 995 -1845
rect 1045 -1875 1075 -1845
rect 1125 -1875 1155 -1845
rect 1205 -1875 1235 -1845
rect 1285 -1875 1315 -1845
rect 1365 -1875 1395 -1845
rect 1445 -1875 1475 -1845
rect 1525 -1875 1555 -1845
rect 1605 -1875 1635 -1845
rect 1685 -1875 1715 -1845
rect 1765 -1875 1795 -1845
rect 1845 -1875 1875 -1845
rect 1925 -1875 1955 -1845
rect 2005 -1875 2035 -1845
rect 2085 -1875 2115 -1845
rect 2165 -1875 2195 -1845
rect 2245 -1875 2275 -1845
rect 2325 -1875 2355 -1845
rect 2405 -1875 2435 -1845
rect 2485 -1875 2515 -1845
rect 2565 -1875 2595 -1845
rect 2645 -1875 2675 -1845
rect 2725 -1875 2755 -1845
rect 2805 -1875 2835 -1845
rect 2885 -1875 2915 -1845
rect 2965 -1875 2995 -1845
rect 3045 -1875 3075 -1845
rect 3125 -1875 3155 -1845
rect 3205 -1875 3235 -1845
rect 3285 -1875 3315 -1845
rect 3365 -1875 3395 -1845
rect 3445 -1875 3475 -1845
rect 3525 -1875 3555 -1845
rect 3605 -1875 3635 -1845
rect 3685 -1875 3715 -1845
rect 3765 -1875 3795 -1845
rect 3845 -1875 3875 -1845
rect 3925 -1875 3955 -1845
rect 4005 -1875 4035 -1845
rect 4085 -1875 4115 -1845
rect 4165 -1875 4195 -1845
rect 4245 -1875 4275 -1845
rect 4325 -1875 4355 -1845
rect 4405 -1875 4435 -1845
rect 4485 -1875 4515 -1845
rect 4565 -1875 4595 -1845
rect 4645 -1875 4675 -1845
rect 4725 -1875 4755 -1845
rect 4805 -1875 4835 -1845
rect 4885 -1875 4915 -1845
rect 4965 -1875 4995 -1845
rect 5045 -1875 5075 -1845
rect 5125 -1875 5155 -1845
rect 5205 -1875 5235 -1845
rect 5285 -1875 5315 -1845
rect 5365 -1875 5395 -1845
rect 5445 -1875 5475 -1845
rect 5525 -1875 5555 -1845
rect 5605 -1875 5635 -1845
rect 5685 -1875 5715 -1845
rect 5765 -1875 5795 -1845
rect 5845 -1875 5875 -1845
rect 5925 -1875 5955 -1845
rect 6005 -1875 6035 -1845
rect 6085 -1875 6115 -1845
rect 6165 -1875 6195 -1845
rect 6245 -1875 6275 -1845
rect 6325 -1875 6355 -1845
rect 6405 -1875 6435 -1845
rect 6485 -1875 6515 -1845
rect 6565 -1875 6595 -1845
rect 6645 -1875 6675 -1845
rect 6725 -1875 6755 -1845
rect 6805 -1875 6835 -1845
rect 6885 -1875 6915 -1845
rect 6965 -1875 6995 -1845
rect 7045 -1875 7075 -1845
rect 7125 -1875 7155 -1845
rect 7205 -1875 7235 -1845
rect 7285 -1875 7315 -1845
rect 7365 -1875 7395 -1845
rect 7445 -1875 7475 -1845
rect 7525 -1875 7555 -1845
rect 7605 -1875 7635 -1845
rect 7685 -1875 7715 -1845
rect 7765 -1875 7795 -1845
rect 7845 -1875 7875 -1845
rect 7925 -1875 7955 -1845
rect 8005 -1875 8035 -1845
rect 8085 -1875 8115 -1845
rect 8165 -1875 8195 -1845
rect 8245 -1875 8275 -1845
rect 8325 -1875 8355 -1845
rect 8405 -1875 8435 -1845
rect 8485 -1875 8515 -1845
rect 8565 -1875 8595 -1845
rect 8645 -1875 8675 -1845
rect 8725 -1875 8755 -1845
rect 8805 -1875 8835 -1845
rect 8885 -1875 8915 -1845
rect 8965 -1875 8995 -1845
rect 9045 -1875 9075 -1845
rect 9125 -1875 9155 -1845
rect 9205 -1875 9235 -1845
rect 9285 -1875 9315 -1845
rect 9365 -1875 9395 -1845
rect 9445 -1875 9475 -1845
rect 9525 -1875 9555 -1845
rect 9605 -1875 9635 -1845
rect 9685 -1875 9715 -1845
rect 9765 -1875 9795 -1845
rect 9845 -1875 9875 -1845
rect 9925 -1875 9955 -1845
rect 10005 -1875 10035 -1845
rect 10085 -1875 10115 -1845
rect 10165 -1875 10195 -1845
rect 10245 -1875 10275 -1845
rect 10325 -1875 10355 -1845
rect 10405 -1875 10435 -1845
rect 10485 -1875 10515 -1845
rect 10565 -1875 10595 -1845
rect 10645 -1875 10675 -1845
rect 10805 -1875 10835 -1845
rect 10965 -1875 10995 -1845
rect -715 -1955 -685 -1925
rect -555 -1955 -525 -1925
rect -475 -1955 -445 -1925
rect 10645 -1955 10675 -1925
rect 10805 -1955 10835 -1925
rect 10965 -1955 10995 -1925
rect -715 -2035 -685 -2005
rect -555 -2035 -525 -2005
rect -395 -2035 -365 -2005
rect -235 -2035 -205 -2005
rect -155 -2035 -125 -2005
rect -75 -2035 -45 -2005
rect 5 -2035 35 -2005
rect 85 -2035 115 -2005
rect 165 -2035 195 -2005
rect 245 -2035 275 -2005
rect 325 -2035 355 -2005
rect 405 -2035 435 -2005
rect 485 -2035 515 -2005
rect 565 -2035 595 -2005
rect 645 -2035 675 -2005
rect 725 -2035 755 -2005
rect 805 -2035 835 -2005
rect 885 -2035 915 -2005
rect 965 -2035 995 -2005
rect 1045 -2035 1075 -2005
rect 1125 -2035 1155 -2005
rect 1205 -2035 1235 -2005
rect 1285 -2035 1315 -2005
rect 1365 -2035 1395 -2005
rect 1445 -2035 1475 -2005
rect 1525 -2035 1555 -2005
rect 1605 -2035 1635 -2005
rect 1685 -2035 1715 -2005
rect 1765 -2035 1795 -2005
rect 1845 -2035 1875 -2005
rect 1925 -2035 1955 -2005
rect 2005 -2035 2035 -2005
rect 2085 -2035 2115 -2005
rect 2165 -2035 2195 -2005
rect 2245 -2035 2275 -2005
rect 2325 -2035 2355 -2005
rect 2405 -2035 2435 -2005
rect 2485 -2035 2515 -2005
rect 2565 -2035 2595 -2005
rect 2645 -2035 2675 -2005
rect 2725 -2035 2755 -2005
rect 2805 -2035 2835 -2005
rect 2885 -2035 2915 -2005
rect 2965 -2035 2995 -2005
rect 3045 -2035 3075 -2005
rect 3125 -2035 3155 -2005
rect 3205 -2035 3235 -2005
rect 3285 -2035 3315 -2005
rect 3365 -2035 3395 -2005
rect 3445 -2035 3475 -2005
rect 3525 -2035 3555 -2005
rect 3605 -2035 3635 -2005
rect 3685 -2035 3715 -2005
rect 3765 -2035 3795 -2005
rect 3845 -2035 3875 -2005
rect 3925 -2035 3955 -2005
rect 4005 -2035 4035 -2005
rect 4085 -2035 4115 -2005
rect 4165 -2035 4195 -2005
rect 4245 -2035 4275 -2005
rect 4325 -2035 4355 -2005
rect 4405 -2035 4435 -2005
rect 4485 -2035 4515 -2005
rect 4565 -2035 4595 -2005
rect 4645 -2035 4675 -2005
rect 4725 -2035 4755 -2005
rect 4805 -2035 4835 -2005
rect 4885 -2035 4915 -2005
rect 4965 -2035 4995 -2005
rect 5045 -2035 5075 -2005
rect 5125 -2035 5155 -2005
rect 5205 -2035 5235 -2005
rect 5285 -2035 5315 -2005
rect 5365 -2035 5395 -2005
rect 5445 -2035 5475 -2005
rect 5525 -2035 5555 -2005
rect 5605 -2035 5635 -2005
rect 5685 -2035 5715 -2005
rect 5765 -2035 5795 -2005
rect 5845 -2035 5875 -2005
rect 5925 -2035 5955 -2005
rect 6005 -2035 6035 -2005
rect 6085 -2035 6115 -2005
rect 6165 -2035 6195 -2005
rect 6245 -2035 6275 -2005
rect 6325 -2035 6355 -2005
rect 6405 -2035 6435 -2005
rect 6485 -2035 6515 -2005
rect 6565 -2035 6595 -2005
rect 6645 -2035 6675 -2005
rect 6725 -2035 6755 -2005
rect 6805 -2035 6835 -2005
rect 6885 -2035 6915 -2005
rect 6965 -2035 6995 -2005
rect 7045 -2035 7075 -2005
rect 7125 -2035 7155 -2005
rect 7205 -2035 7235 -2005
rect 7285 -2035 7315 -2005
rect 7365 -2035 7395 -2005
rect 7445 -2035 7475 -2005
rect 7525 -2035 7555 -2005
rect 7605 -2035 7635 -2005
rect 7685 -2035 7715 -2005
rect 7765 -2035 7795 -2005
rect 7845 -2035 7875 -2005
rect 7925 -2035 7955 -2005
rect 8005 -2035 8035 -2005
rect 8085 -2035 8115 -2005
rect 8165 -2035 8195 -2005
rect 8245 -2035 8275 -2005
rect 8325 -2035 8355 -2005
rect 8405 -2035 8435 -2005
rect 8485 -2035 8515 -2005
rect 8565 -2035 8595 -2005
rect 8645 -2035 8675 -2005
rect 8725 -2035 8755 -2005
rect 8805 -2035 8835 -2005
rect 8885 -2035 8915 -2005
rect 8965 -2035 8995 -2005
rect 9045 -2035 9075 -2005
rect 9125 -2035 9155 -2005
rect 9205 -2035 9235 -2005
rect 9285 -2035 9315 -2005
rect 9365 -2035 9395 -2005
rect 9445 -2035 9475 -2005
rect 9525 -2035 9555 -2005
rect 9605 -2035 9635 -2005
rect 9685 -2035 9715 -2005
rect 9765 -2035 9795 -2005
rect 9845 -2035 9875 -2005
rect 9925 -2035 9955 -2005
rect 10005 -2035 10035 -2005
rect 10085 -2035 10115 -2005
rect 10165 -2035 10195 -2005
rect 10245 -2035 10275 -2005
rect 10325 -2035 10355 -2005
rect 10405 -2035 10435 -2005
rect 10485 -2035 10515 -2005
rect 10565 -2035 10595 -2005
rect 10645 -2035 10675 -2005
rect 10805 -2035 10835 -2005
rect 10965 -2035 10995 -2005
rect -715 -2115 -685 -2085
rect -555 -2115 -525 -2085
rect -395 -2115 -365 -2085
rect 10885 -2115 10915 -2085
rect -715 -2195 -685 -2165
rect -555 -2195 -525 -2165
rect -395 -2195 -365 -2165
rect -235 -2195 -205 -2165
rect -155 -2195 -125 -2165
rect -75 -2195 -45 -2165
rect 5 -2195 35 -2165
rect 85 -2195 115 -2165
rect 165 -2195 195 -2165
rect 245 -2195 275 -2165
rect 325 -2195 355 -2165
rect 405 -2195 435 -2165
rect 485 -2195 515 -2165
rect 565 -2195 595 -2165
rect 645 -2195 675 -2165
rect 725 -2195 755 -2165
rect 805 -2195 835 -2165
rect 885 -2195 915 -2165
rect 965 -2195 995 -2165
rect 1045 -2195 1075 -2165
rect 1125 -2195 1155 -2165
rect 1205 -2195 1235 -2165
rect 1285 -2195 1315 -2165
rect 1365 -2195 1395 -2165
rect 1445 -2195 1475 -2165
rect 1525 -2195 1555 -2165
rect 1605 -2195 1635 -2165
rect 1685 -2195 1715 -2165
rect 1765 -2195 1795 -2165
rect 1845 -2195 1875 -2165
rect 1925 -2195 1955 -2165
rect 2005 -2195 2035 -2165
rect 2085 -2195 2115 -2165
rect 2165 -2195 2195 -2165
rect 2245 -2195 2275 -2165
rect 2325 -2195 2355 -2165
rect 2405 -2195 2435 -2165
rect 2485 -2195 2515 -2165
rect 2565 -2195 2595 -2165
rect 2645 -2195 2675 -2165
rect 2725 -2195 2755 -2165
rect 2805 -2195 2835 -2165
rect 2885 -2195 2915 -2165
rect 2965 -2195 2995 -2165
rect 3045 -2195 3075 -2165
rect 3125 -2195 3155 -2165
rect 3205 -2195 3235 -2165
rect 3285 -2195 3315 -2165
rect 3365 -2195 3395 -2165
rect 3445 -2195 3475 -2165
rect 3525 -2195 3555 -2165
rect 3605 -2195 3635 -2165
rect 3685 -2195 3715 -2165
rect 3765 -2195 3795 -2165
rect 3845 -2195 3875 -2165
rect 3925 -2195 3955 -2165
rect 4005 -2195 4035 -2165
rect 4085 -2195 4115 -2165
rect 4165 -2195 4195 -2165
rect 4245 -2195 4275 -2165
rect 4325 -2195 4355 -2165
rect 4405 -2195 4435 -2165
rect 4485 -2195 4515 -2165
rect 4565 -2195 4595 -2165
rect 4645 -2195 4675 -2165
rect 4725 -2195 4755 -2165
rect 4805 -2195 4835 -2165
rect 4885 -2195 4915 -2165
rect 4965 -2195 4995 -2165
rect 5045 -2195 5075 -2165
rect 5125 -2195 5155 -2165
rect 5205 -2195 5235 -2165
rect 5285 -2195 5315 -2165
rect 5365 -2195 5395 -2165
rect 5445 -2195 5475 -2165
rect 5525 -2195 5555 -2165
rect 5605 -2195 5635 -2165
rect 5685 -2195 5715 -2165
rect 5765 -2195 5795 -2165
rect 5845 -2195 5875 -2165
rect 5925 -2195 5955 -2165
rect 6005 -2195 6035 -2165
rect 6085 -2195 6115 -2165
rect 6165 -2195 6195 -2165
rect 6245 -2195 6275 -2165
rect 6325 -2195 6355 -2165
rect 6405 -2195 6435 -2165
rect 6485 -2195 6515 -2165
rect 6565 -2195 6595 -2165
rect 6645 -2195 6675 -2165
rect 6725 -2195 6755 -2165
rect 6805 -2195 6835 -2165
rect 6885 -2195 6915 -2165
rect 6965 -2195 6995 -2165
rect 7045 -2195 7075 -2165
rect 7125 -2195 7155 -2165
rect 7205 -2195 7235 -2165
rect 7285 -2195 7315 -2165
rect 7365 -2195 7395 -2165
rect 7445 -2195 7475 -2165
rect 7525 -2195 7555 -2165
rect 7605 -2195 7635 -2165
rect 7685 -2195 7715 -2165
rect 7765 -2195 7795 -2165
rect 7845 -2195 7875 -2165
rect 7925 -2195 7955 -2165
rect 8005 -2195 8035 -2165
rect 8085 -2195 8115 -2165
rect 8165 -2195 8195 -2165
rect 8245 -2195 8275 -2165
rect 8325 -2195 8355 -2165
rect 8405 -2195 8435 -2165
rect 8485 -2195 8515 -2165
rect 8565 -2195 8595 -2165
rect 8645 -2195 8675 -2165
rect 8725 -2195 8755 -2165
rect 8805 -2195 8835 -2165
rect 8885 -2195 8915 -2165
rect 8965 -2195 8995 -2165
rect 9045 -2195 9075 -2165
rect 9125 -2195 9155 -2165
rect 9205 -2195 9235 -2165
rect 9285 -2195 9315 -2165
rect 9365 -2195 9395 -2165
rect 9445 -2195 9475 -2165
rect 9525 -2195 9555 -2165
rect 9605 -2195 9635 -2165
rect 9685 -2195 9715 -2165
rect 9765 -2195 9795 -2165
rect 9845 -2195 9875 -2165
rect 9925 -2195 9955 -2165
rect 10005 -2195 10035 -2165
rect 10085 -2195 10115 -2165
rect 10165 -2195 10195 -2165
rect 10245 -2195 10275 -2165
rect 10325 -2195 10355 -2165
rect 10405 -2195 10435 -2165
rect 10485 -2195 10515 -2165
rect 10565 -2195 10595 -2165
rect 10645 -2195 10675 -2165
rect 10805 -2195 10835 -2165
rect 10965 -2195 10995 -2165
rect -715 -2275 -685 -2245
rect -555 -2275 -525 -2245
rect -395 -2275 -365 -2245
rect 10725 -2275 10755 -2245
rect 10805 -2275 10835 -2245
rect 10965 -2275 10995 -2245
rect -715 -2355 -685 -2325
rect -555 -2355 -525 -2325
rect -395 -2355 -365 -2325
rect -235 -2355 -205 -2325
rect -155 -2355 -125 -2325
rect -75 -2355 -45 -2325
rect 5 -2355 35 -2325
rect 85 -2355 115 -2325
rect 165 -2355 195 -2325
rect 245 -2355 275 -2325
rect 325 -2355 355 -2325
rect 405 -2355 435 -2325
rect 485 -2355 515 -2325
rect 565 -2355 595 -2325
rect 645 -2355 675 -2325
rect 725 -2355 755 -2325
rect 805 -2355 835 -2325
rect 885 -2355 915 -2325
rect 965 -2355 995 -2325
rect 1045 -2355 1075 -2325
rect 1125 -2355 1155 -2325
rect 1205 -2355 1235 -2325
rect 1285 -2355 1315 -2325
rect 1365 -2355 1395 -2325
rect 1445 -2355 1475 -2325
rect 1525 -2355 1555 -2325
rect 1605 -2355 1635 -2325
rect 1685 -2355 1715 -2325
rect 1765 -2355 1795 -2325
rect 1845 -2355 1875 -2325
rect 1925 -2355 1955 -2325
rect 2005 -2355 2035 -2325
rect 2085 -2355 2115 -2325
rect 2165 -2355 2195 -2325
rect 2245 -2355 2275 -2325
rect 2325 -2355 2355 -2325
rect 2405 -2355 2435 -2325
rect 2485 -2355 2515 -2325
rect 2565 -2355 2595 -2325
rect 2645 -2355 2675 -2325
rect 2725 -2355 2755 -2325
rect 2805 -2355 2835 -2325
rect 2885 -2355 2915 -2325
rect 2965 -2355 2995 -2325
rect 3045 -2355 3075 -2325
rect 3125 -2355 3155 -2325
rect 3205 -2355 3235 -2325
rect 3285 -2355 3315 -2325
rect 3365 -2355 3395 -2325
rect 3445 -2355 3475 -2325
rect 3525 -2355 3555 -2325
rect 3605 -2355 3635 -2325
rect 3685 -2355 3715 -2325
rect 3765 -2355 3795 -2325
rect 3845 -2355 3875 -2325
rect 3925 -2355 3955 -2325
rect 4005 -2355 4035 -2325
rect 4085 -2355 4115 -2325
rect 4165 -2355 4195 -2325
rect 4245 -2355 4275 -2325
rect 4325 -2355 4355 -2325
rect 4405 -2355 4435 -2325
rect 4485 -2355 4515 -2325
rect 4565 -2355 4595 -2325
rect 4645 -2355 4675 -2325
rect 4725 -2355 4755 -2325
rect 4805 -2355 4835 -2325
rect 4885 -2355 4915 -2325
rect 4965 -2355 4995 -2325
rect 5045 -2355 5075 -2325
rect 5125 -2355 5155 -2325
rect 5205 -2355 5235 -2325
rect 5285 -2355 5315 -2325
rect 5365 -2355 5395 -2325
rect 5445 -2355 5475 -2325
rect 5525 -2355 5555 -2325
rect 5605 -2355 5635 -2325
rect 5685 -2355 5715 -2325
rect 5765 -2355 5795 -2325
rect 5845 -2355 5875 -2325
rect 5925 -2355 5955 -2325
rect 6005 -2355 6035 -2325
rect 6085 -2355 6115 -2325
rect 6165 -2355 6195 -2325
rect 6245 -2355 6275 -2325
rect 6325 -2355 6355 -2325
rect 6405 -2355 6435 -2325
rect 6485 -2355 6515 -2325
rect 6565 -2355 6595 -2325
rect 6645 -2355 6675 -2325
rect 6725 -2355 6755 -2325
rect 6805 -2355 6835 -2325
rect 6885 -2355 6915 -2325
rect 6965 -2355 6995 -2325
rect 7045 -2355 7075 -2325
rect 7125 -2355 7155 -2325
rect 7205 -2355 7235 -2325
rect 7285 -2355 7315 -2325
rect 7365 -2355 7395 -2325
rect 7445 -2355 7475 -2325
rect 7525 -2355 7555 -2325
rect 7605 -2355 7635 -2325
rect 7685 -2355 7715 -2325
rect 7765 -2355 7795 -2325
rect 7845 -2355 7875 -2325
rect 7925 -2355 7955 -2325
rect 8005 -2355 8035 -2325
rect 8085 -2355 8115 -2325
rect 8165 -2355 8195 -2325
rect 8245 -2355 8275 -2325
rect 8325 -2355 8355 -2325
rect 8405 -2355 8435 -2325
rect 8485 -2355 8515 -2325
rect 8565 -2355 8595 -2325
rect 8645 -2355 8675 -2325
rect 8725 -2355 8755 -2325
rect 8805 -2355 8835 -2325
rect 8885 -2355 8915 -2325
rect 8965 -2355 8995 -2325
rect 9045 -2355 9075 -2325
rect 9125 -2355 9155 -2325
rect 9205 -2355 9235 -2325
rect 9285 -2355 9315 -2325
rect 9365 -2355 9395 -2325
rect 9445 -2355 9475 -2325
rect 9525 -2355 9555 -2325
rect 9605 -2355 9635 -2325
rect 9685 -2355 9715 -2325
rect 9765 -2355 9795 -2325
rect 9845 -2355 9875 -2325
rect 9925 -2355 9955 -2325
rect 10005 -2355 10035 -2325
rect 10085 -2355 10115 -2325
rect 10165 -2355 10195 -2325
rect 10245 -2355 10275 -2325
rect 10325 -2355 10355 -2325
rect 10405 -2355 10435 -2325
rect 10485 -2355 10515 -2325
rect 10565 -2355 10595 -2325
rect 10645 -2355 10675 -2325
rect 10805 -2355 10835 -2325
rect 10965 -2355 10995 -2325
rect -715 -2435 -685 -2405
rect -555 -2435 -525 -2405
rect -395 -2435 -365 -2405
rect -235 -2435 -205 -2405
rect -155 -2435 -125 -2405
rect -75 -2435 -45 -2405
rect 5 -2435 35 -2405
rect 85 -2435 115 -2405
rect 165 -2435 195 -2405
rect 245 -2435 275 -2405
rect 325 -2435 355 -2405
rect 405 -2435 435 -2405
rect 485 -2435 515 -2405
rect 565 -2435 595 -2405
rect 645 -2435 675 -2405
rect 725 -2435 755 -2405
rect 805 -2435 835 -2405
rect 885 -2435 915 -2405
rect 965 -2435 995 -2405
rect 1045 -2435 1075 -2405
rect 1125 -2435 1155 -2405
rect 1205 -2435 1235 -2405
rect 1285 -2435 1315 -2405
rect 1365 -2435 1395 -2405
rect 1445 -2435 1475 -2405
rect 1525 -2435 1555 -2405
rect 1605 -2435 1635 -2405
rect 1685 -2435 1715 -2405
rect 1765 -2435 1795 -2405
rect 1845 -2435 1875 -2405
rect 1925 -2435 1955 -2405
rect 2005 -2435 2035 -2405
rect 2085 -2435 2115 -2405
rect 2165 -2435 2195 -2405
rect 2245 -2435 2275 -2405
rect 2325 -2435 2355 -2405
rect 2405 -2435 2435 -2405
rect 2485 -2435 2515 -2405
rect 2565 -2435 2595 -2405
rect 2645 -2435 2675 -2405
rect 2725 -2435 2755 -2405
rect 2805 -2435 2835 -2405
rect 2885 -2435 2915 -2405
rect 2965 -2435 2995 -2405
rect 3045 -2435 3075 -2405
rect 3125 -2435 3155 -2405
rect 3205 -2435 3235 -2405
rect 3285 -2435 3315 -2405
rect 3365 -2435 3395 -2405
rect 3445 -2435 3475 -2405
rect 3525 -2435 3555 -2405
rect 3605 -2435 3635 -2405
rect 3685 -2435 3715 -2405
rect 3765 -2435 3795 -2405
rect 3845 -2435 3875 -2405
rect 3925 -2435 3955 -2405
rect 4005 -2435 4035 -2405
rect 4085 -2435 4115 -2405
rect 4165 -2435 4195 -2405
rect 4245 -2435 4275 -2405
rect 4325 -2435 4355 -2405
rect 4405 -2435 4435 -2405
rect 4485 -2435 4515 -2405
rect 4565 -2435 4595 -2405
rect 4645 -2435 4675 -2405
rect 4725 -2435 4755 -2405
rect 4805 -2435 4835 -2405
rect 4885 -2435 4915 -2405
rect 4965 -2435 4995 -2405
rect 5045 -2435 5075 -2405
rect 5125 -2435 5155 -2405
rect 5205 -2435 5235 -2405
rect 5285 -2435 5315 -2405
rect 5365 -2435 5395 -2405
rect 5445 -2435 5475 -2405
rect 5525 -2435 5555 -2405
rect 5605 -2435 5635 -2405
rect 5685 -2435 5715 -2405
rect 5765 -2435 5795 -2405
rect 5845 -2435 5875 -2405
rect 5925 -2435 5955 -2405
rect 6005 -2435 6035 -2405
rect 6085 -2435 6115 -2405
rect 6165 -2435 6195 -2405
rect 6245 -2435 6275 -2405
rect 6325 -2435 6355 -2405
rect 6405 -2435 6435 -2405
rect 6485 -2435 6515 -2405
rect 6565 -2435 6595 -2405
rect 6645 -2435 6675 -2405
rect 6725 -2435 6755 -2405
rect 6805 -2435 6835 -2405
rect 6885 -2435 6915 -2405
rect 6965 -2435 6995 -2405
rect 7045 -2435 7075 -2405
rect 7125 -2435 7155 -2405
rect 7205 -2435 7235 -2405
rect 7285 -2435 7315 -2405
rect 7365 -2435 7395 -2405
rect 7445 -2435 7475 -2405
rect 7525 -2435 7555 -2405
rect 7605 -2435 7635 -2405
rect 7685 -2435 7715 -2405
rect 7765 -2435 7795 -2405
rect 7845 -2435 7875 -2405
rect 7925 -2435 7955 -2405
rect 8005 -2435 8035 -2405
rect 8085 -2435 8115 -2405
rect 8165 -2435 8195 -2405
rect 8245 -2435 8275 -2405
rect 8325 -2435 8355 -2405
rect 8405 -2435 8435 -2405
rect 8485 -2435 8515 -2405
rect 8565 -2435 8595 -2405
rect 8645 -2435 8675 -2405
rect 8725 -2435 8755 -2405
rect 8805 -2435 8835 -2405
rect 8885 -2435 8915 -2405
rect 8965 -2435 8995 -2405
rect 9045 -2435 9075 -2405
rect 9125 -2435 9155 -2405
rect 9205 -2435 9235 -2405
rect 9285 -2435 9315 -2405
rect 9365 -2435 9395 -2405
rect 9445 -2435 9475 -2405
rect 9525 -2435 9555 -2405
rect 9605 -2435 9635 -2405
rect 9685 -2435 9715 -2405
rect 9765 -2435 9795 -2405
rect 9845 -2435 9875 -2405
rect 9925 -2435 9955 -2405
rect 10005 -2435 10035 -2405
rect 10085 -2435 10115 -2405
rect 10165 -2435 10195 -2405
rect 10245 -2435 10275 -2405
rect 10325 -2435 10355 -2405
rect 10405 -2435 10435 -2405
rect 10485 -2435 10515 -2405
rect 10565 -2435 10595 -2405
rect 10645 -2435 10675 -2405
rect 10805 -2435 10835 -2405
rect 10965 -2435 10995 -2405
rect -715 -2515 -685 -2485
rect -555 -2515 -525 -2485
rect -395 -2515 -365 -2485
rect -235 -2515 -205 -2485
rect -155 -2515 -125 -2485
rect -75 -2515 -45 -2485
rect 5 -2515 35 -2485
rect 85 -2515 115 -2485
rect 165 -2515 195 -2485
rect 245 -2515 275 -2485
rect 325 -2515 355 -2485
rect 405 -2515 435 -2485
rect 485 -2515 515 -2485
rect 565 -2515 595 -2485
rect 645 -2515 675 -2485
rect 725 -2515 755 -2485
rect 805 -2515 835 -2485
rect 885 -2515 915 -2485
rect 965 -2515 995 -2485
rect 1045 -2515 1075 -2485
rect 1125 -2515 1155 -2485
rect 1205 -2515 1235 -2485
rect 1285 -2515 1315 -2485
rect 1365 -2515 1395 -2485
rect 1445 -2515 1475 -2485
rect 1525 -2515 1555 -2485
rect 1605 -2515 1635 -2485
rect 1685 -2515 1715 -2485
rect 1765 -2515 1795 -2485
rect 1845 -2515 1875 -2485
rect 1925 -2515 1955 -2485
rect 2005 -2515 2035 -2485
rect 2085 -2515 2115 -2485
rect 2165 -2515 2195 -2485
rect 2245 -2515 2275 -2485
rect 2325 -2515 2355 -2485
rect 2405 -2515 2435 -2485
rect 2485 -2515 2515 -2485
rect 2565 -2515 2595 -2485
rect 2645 -2515 2675 -2485
rect 2725 -2515 2755 -2485
rect 2805 -2515 2835 -2485
rect 2885 -2515 2915 -2485
rect 2965 -2515 2995 -2485
rect 3045 -2515 3075 -2485
rect 3125 -2515 3155 -2485
rect 3205 -2515 3235 -2485
rect 3285 -2515 3315 -2485
rect 3365 -2515 3395 -2485
rect 3445 -2515 3475 -2485
rect 3525 -2515 3555 -2485
rect 3605 -2515 3635 -2485
rect 3685 -2515 3715 -2485
rect 3765 -2515 3795 -2485
rect 3845 -2515 3875 -2485
rect 3925 -2515 3955 -2485
rect 4005 -2515 4035 -2485
rect 4085 -2515 4115 -2485
rect 4165 -2515 4195 -2485
rect 4245 -2515 4275 -2485
rect 4325 -2515 4355 -2485
rect 4405 -2515 4435 -2485
rect 4485 -2515 4515 -2485
rect 4565 -2515 4595 -2485
rect 4645 -2515 4675 -2485
rect 4725 -2515 4755 -2485
rect 4805 -2515 4835 -2485
rect 4885 -2515 4915 -2485
rect 4965 -2515 4995 -2485
rect 5045 -2515 5075 -2485
rect 5125 -2515 5155 -2485
rect 5205 -2515 5235 -2485
rect 5285 -2515 5315 -2485
rect 5365 -2515 5395 -2485
rect 5445 -2515 5475 -2485
rect 5525 -2515 5555 -2485
rect 5605 -2515 5635 -2485
rect 5685 -2515 5715 -2485
rect 5765 -2515 5795 -2485
rect 5845 -2515 5875 -2485
rect 5925 -2515 5955 -2485
rect 6005 -2515 6035 -2485
rect 6085 -2515 6115 -2485
rect 6165 -2515 6195 -2485
rect 6245 -2515 6275 -2485
rect 6325 -2515 6355 -2485
rect 6405 -2515 6435 -2485
rect 6485 -2515 6515 -2485
rect 6565 -2515 6595 -2485
rect 6645 -2515 6675 -2485
rect 6725 -2515 6755 -2485
rect 6805 -2515 6835 -2485
rect 6885 -2515 6915 -2485
rect 6965 -2515 6995 -2485
rect 7045 -2515 7075 -2485
rect 7125 -2515 7155 -2485
rect 7205 -2515 7235 -2485
rect 7285 -2515 7315 -2485
rect 7365 -2515 7395 -2485
rect 7445 -2515 7475 -2485
rect 7525 -2515 7555 -2485
rect 7605 -2515 7635 -2485
rect 7685 -2515 7715 -2485
rect 7765 -2515 7795 -2485
rect 7845 -2515 7875 -2485
rect 7925 -2515 7955 -2485
rect 8005 -2515 8035 -2485
rect 8085 -2515 8115 -2485
rect 8165 -2515 8195 -2485
rect 8245 -2515 8275 -2485
rect 8325 -2515 8355 -2485
rect 8405 -2515 8435 -2485
rect 8485 -2515 8515 -2485
rect 8565 -2515 8595 -2485
rect 8645 -2515 8675 -2485
rect 8725 -2515 8755 -2485
rect 8805 -2515 8835 -2485
rect 8885 -2515 8915 -2485
rect 8965 -2515 8995 -2485
rect 9045 -2515 9075 -2485
rect 9125 -2515 9155 -2485
rect 9205 -2515 9235 -2485
rect 9285 -2515 9315 -2485
rect 9365 -2515 9395 -2485
rect 9445 -2515 9475 -2485
rect 9525 -2515 9555 -2485
rect 9605 -2515 9635 -2485
rect 9685 -2515 9715 -2485
rect 9765 -2515 9795 -2485
rect 9845 -2515 9875 -2485
rect 9925 -2515 9955 -2485
rect 10005 -2515 10035 -2485
rect 10085 -2515 10115 -2485
rect 10165 -2515 10195 -2485
rect 10245 -2515 10275 -2485
rect 10325 -2515 10355 -2485
rect 10405 -2515 10435 -2485
rect 10485 -2515 10515 -2485
rect 10565 -2515 10595 -2485
rect 10645 -2515 10675 -2485
rect 10805 -2515 10835 -2485
rect 10965 -2515 10995 -2485
rect -715 -2595 -685 -2565
rect -555 -2595 -525 -2565
rect -395 -2595 -365 -2565
rect -315 -2595 -285 -2565
rect -235 -2595 -205 -2565
rect -155 -2595 -125 -2565
rect -75 -2595 -45 -2565
rect 5 -2595 35 -2565
rect 85 -2595 115 -2565
rect 165 -2595 195 -2565
rect 245 -2595 275 -2565
rect 325 -2595 355 -2565
rect 405 -2595 435 -2565
rect 485 -2595 515 -2565
rect 565 -2595 595 -2565
rect 645 -2595 675 -2565
rect 725 -2595 755 -2565
rect 805 -2595 835 -2565
rect 885 -2595 915 -2565
rect 965 -2595 995 -2565
rect 1045 -2595 1075 -2565
rect 1125 -2595 1155 -2565
rect 1205 -2595 1235 -2565
rect 1285 -2595 1315 -2565
rect 1365 -2595 1395 -2565
rect 1445 -2595 1475 -2565
rect 1525 -2595 1555 -2565
rect 1605 -2595 1635 -2565
rect 1685 -2595 1715 -2565
rect 1765 -2595 1795 -2565
rect 1845 -2595 1875 -2565
rect 1925 -2595 1955 -2565
rect 2005 -2595 2035 -2565
rect 2085 -2595 2115 -2565
rect 2165 -2595 2195 -2565
rect 2245 -2595 2275 -2565
rect 2325 -2595 2355 -2565
rect 2405 -2595 2435 -2565
rect 2485 -2595 2515 -2565
rect 2565 -2595 2595 -2565
rect 2645 -2595 2675 -2565
rect 2725 -2595 2755 -2565
rect 2805 -2595 2835 -2565
rect 2885 -2595 2915 -2565
rect 2965 -2595 2995 -2565
rect 3045 -2595 3075 -2565
rect 3125 -2595 3155 -2565
rect 3205 -2595 3235 -2565
rect 3285 -2595 3315 -2565
rect 3365 -2595 3395 -2565
rect 3445 -2595 3475 -2565
rect 3525 -2595 3555 -2565
rect 3605 -2595 3635 -2565
rect 3685 -2595 3715 -2565
rect 3765 -2595 3795 -2565
rect 3845 -2595 3875 -2565
rect 3925 -2595 3955 -2565
rect 4005 -2595 4035 -2565
rect 4085 -2595 4115 -2565
rect 4165 -2595 4195 -2565
rect 4245 -2595 4275 -2565
rect 4325 -2595 4355 -2565
rect 4405 -2595 4435 -2565
rect 4485 -2595 4515 -2565
rect 4565 -2595 4595 -2565
rect 4645 -2595 4675 -2565
rect 4725 -2595 4755 -2565
rect 4805 -2595 4835 -2565
rect 4885 -2595 4915 -2565
rect 4965 -2595 4995 -2565
rect 5045 -2595 5075 -2565
rect 5125 -2595 5155 -2565
rect 5205 -2595 5235 -2565
rect 5285 -2595 5315 -2565
rect 5365 -2595 5395 -2565
rect 5445 -2595 5475 -2565
rect 5525 -2595 5555 -2565
rect 5605 -2595 5635 -2565
rect 5685 -2595 5715 -2565
rect 5765 -2595 5795 -2565
rect 5845 -2595 5875 -2565
rect 5925 -2595 5955 -2565
rect 6005 -2595 6035 -2565
rect 6085 -2595 6115 -2565
rect 6165 -2595 6195 -2565
rect 6245 -2595 6275 -2565
rect 6325 -2595 6355 -2565
rect 6405 -2595 6435 -2565
rect 6485 -2595 6515 -2565
rect 6565 -2595 6595 -2565
rect 6645 -2595 6675 -2565
rect 6725 -2595 6755 -2565
rect 6805 -2595 6835 -2565
rect 6885 -2595 6915 -2565
rect 6965 -2595 6995 -2565
rect 7045 -2595 7075 -2565
rect 7125 -2595 7155 -2565
rect 7205 -2595 7235 -2565
rect 7285 -2595 7315 -2565
rect 7365 -2595 7395 -2565
rect 7445 -2595 7475 -2565
rect 7525 -2595 7555 -2565
rect 7605 -2595 7635 -2565
rect 7685 -2595 7715 -2565
rect 7765 -2595 7795 -2565
rect 7845 -2595 7875 -2565
rect 7925 -2595 7955 -2565
rect 8005 -2595 8035 -2565
rect 8085 -2595 8115 -2565
rect 8165 -2595 8195 -2565
rect 8245 -2595 8275 -2565
rect 8325 -2595 8355 -2565
rect 8405 -2595 8435 -2565
rect 8485 -2595 8515 -2565
rect 8565 -2595 8595 -2565
rect 8645 -2595 8675 -2565
rect 8725 -2595 8755 -2565
rect 8805 -2595 8835 -2565
rect 8885 -2595 8915 -2565
rect 8965 -2595 8995 -2565
rect 9045 -2595 9075 -2565
rect 9125 -2595 9155 -2565
rect 9205 -2595 9235 -2565
rect 9285 -2595 9315 -2565
rect 9365 -2595 9395 -2565
rect 9445 -2595 9475 -2565
rect 9525 -2595 9555 -2565
rect 9605 -2595 9635 -2565
rect 9685 -2595 9715 -2565
rect 9765 -2595 9795 -2565
rect 9845 -2595 9875 -2565
rect 9925 -2595 9955 -2565
rect 10005 -2595 10035 -2565
rect 10085 -2595 10115 -2565
rect 10165 -2595 10195 -2565
rect 10245 -2595 10275 -2565
rect 10325 -2595 10355 -2565
rect 10405 -2595 10435 -2565
rect 10485 -2595 10515 -2565
rect 10645 -2595 10675 -2565
rect 10805 -2595 10835 -2565
rect 10965 -2595 10995 -2565
rect -715 -2675 -685 -2645
rect -555 -2675 -525 -2645
rect -395 -2675 -365 -2645
rect -315 -2675 -285 -2645
rect -235 -2675 -205 -2645
rect -155 -2675 -125 -2645
rect -75 -2675 -45 -2645
rect 5 -2675 35 -2645
rect 85 -2675 115 -2645
rect 165 -2675 195 -2645
rect 245 -2675 275 -2645
rect 325 -2675 355 -2645
rect 405 -2675 435 -2645
rect 485 -2675 515 -2645
rect 565 -2675 595 -2645
rect 645 -2675 675 -2645
rect 725 -2675 755 -2645
rect 805 -2675 835 -2645
rect 885 -2675 915 -2645
rect 965 -2675 995 -2645
rect 1045 -2675 1075 -2645
rect 1125 -2675 1155 -2645
rect 1205 -2675 1235 -2645
rect 1285 -2675 1315 -2645
rect 1365 -2675 1395 -2645
rect 1445 -2675 1475 -2645
rect 1525 -2675 1555 -2645
rect 1605 -2675 1635 -2645
rect 1685 -2675 1715 -2645
rect 1765 -2675 1795 -2645
rect 1845 -2675 1875 -2645
rect 1925 -2675 1955 -2645
rect 2005 -2675 2035 -2645
rect 2085 -2675 2115 -2645
rect 2165 -2675 2195 -2645
rect 2245 -2675 2275 -2645
rect 2325 -2675 2355 -2645
rect 2405 -2675 2435 -2645
rect 2485 -2675 2515 -2645
rect 2565 -2675 2595 -2645
rect 2645 -2675 2675 -2645
rect 2725 -2675 2755 -2645
rect 2805 -2675 2835 -2645
rect 2885 -2675 2915 -2645
rect 2965 -2675 2995 -2645
rect 3045 -2675 3075 -2645
rect 3125 -2675 3155 -2645
rect 3205 -2675 3235 -2645
rect 3285 -2675 3315 -2645
rect 3365 -2675 3395 -2645
rect 3445 -2675 3475 -2645
rect 3525 -2675 3555 -2645
rect 3605 -2675 3635 -2645
rect 3685 -2675 3715 -2645
rect 3765 -2675 3795 -2645
rect 3845 -2675 3875 -2645
rect 3925 -2675 3955 -2645
rect 4005 -2675 4035 -2645
rect 4085 -2675 4115 -2645
rect 4165 -2675 4195 -2645
rect 4245 -2675 4275 -2645
rect 4325 -2675 4355 -2645
rect 4405 -2675 4435 -2645
rect 4485 -2675 4515 -2645
rect 4565 -2675 4595 -2645
rect 4645 -2675 4675 -2645
rect 4725 -2675 4755 -2645
rect 4805 -2675 4835 -2645
rect 4885 -2675 4915 -2645
rect 4965 -2675 4995 -2645
rect 5045 -2675 5075 -2645
rect 5125 -2675 5155 -2645
rect 5205 -2675 5235 -2645
rect 5285 -2675 5315 -2645
rect 5365 -2675 5395 -2645
rect 5445 -2675 5475 -2645
rect 5525 -2675 5555 -2645
rect 5605 -2675 5635 -2645
rect 5685 -2675 5715 -2645
rect 5765 -2675 5795 -2645
rect 5845 -2675 5875 -2645
rect 5925 -2675 5955 -2645
rect 6005 -2675 6035 -2645
rect 6085 -2675 6115 -2645
rect 6165 -2675 6195 -2645
rect 6245 -2675 6275 -2645
rect 6325 -2675 6355 -2645
rect 6405 -2675 6435 -2645
rect 6485 -2675 6515 -2645
rect 6565 -2675 6595 -2645
rect 6645 -2675 6675 -2645
rect 6725 -2675 6755 -2645
rect 6805 -2675 6835 -2645
rect 6885 -2675 6915 -2645
rect 6965 -2675 6995 -2645
rect 7045 -2675 7075 -2645
rect 7125 -2675 7155 -2645
rect 7205 -2675 7235 -2645
rect 7285 -2675 7315 -2645
rect 7365 -2675 7395 -2645
rect 7445 -2675 7475 -2645
rect 7525 -2675 7555 -2645
rect 7605 -2675 7635 -2645
rect 7685 -2675 7715 -2645
rect 7765 -2675 7795 -2645
rect 7845 -2675 7875 -2645
rect 7925 -2675 7955 -2645
rect 8005 -2675 8035 -2645
rect 8085 -2675 8115 -2645
rect 8165 -2675 8195 -2645
rect 8245 -2675 8275 -2645
rect 8325 -2675 8355 -2645
rect 8405 -2675 8435 -2645
rect 8485 -2675 8515 -2645
rect 8565 -2675 8595 -2645
rect 8645 -2675 8675 -2645
rect 8725 -2675 8755 -2645
rect 8805 -2675 8835 -2645
rect 8885 -2675 8915 -2645
rect 8965 -2675 8995 -2645
rect 9045 -2675 9075 -2645
rect 9125 -2675 9155 -2645
rect 9205 -2675 9235 -2645
rect 9285 -2675 9315 -2645
rect 9365 -2675 9395 -2645
rect 9445 -2675 9475 -2645
rect 9525 -2675 9555 -2645
rect 9605 -2675 9635 -2645
rect 9685 -2675 9715 -2645
rect 9765 -2675 9795 -2645
rect 9845 -2675 9875 -2645
rect 9925 -2675 9955 -2645
rect 10005 -2675 10035 -2645
rect 10085 -2675 10115 -2645
rect 10165 -2675 10195 -2645
rect 10245 -2675 10275 -2645
rect 10325 -2675 10355 -2645
rect 10405 -2675 10435 -2645
rect 10485 -2675 10515 -2645
rect 10645 -2675 10675 -2645
rect 10805 -2675 10835 -2645
rect 10965 -2675 10995 -2645
rect -715 -2755 -685 -2725
rect -555 -2755 -525 -2725
rect -395 -2755 -365 -2725
rect -315 -2755 -285 -2725
rect -235 -2755 -205 -2725
rect -155 -2755 -125 -2725
rect -75 -2755 -45 -2725
rect 5 -2755 35 -2725
rect 85 -2755 115 -2725
rect 165 -2755 195 -2725
rect 245 -2755 275 -2725
rect 325 -2755 355 -2725
rect 405 -2755 435 -2725
rect 485 -2755 515 -2725
rect 565 -2755 595 -2725
rect 645 -2755 675 -2725
rect 725 -2755 755 -2725
rect 805 -2755 835 -2725
rect 885 -2755 915 -2725
rect 965 -2755 995 -2725
rect 1045 -2755 1075 -2725
rect 1125 -2755 1155 -2725
rect 1205 -2755 1235 -2725
rect 1285 -2755 1315 -2725
rect 1365 -2755 1395 -2725
rect 1445 -2755 1475 -2725
rect 1525 -2755 1555 -2725
rect 1605 -2755 1635 -2725
rect 1685 -2755 1715 -2725
rect 1765 -2755 1795 -2725
rect 1845 -2755 1875 -2725
rect 1925 -2755 1955 -2725
rect 2005 -2755 2035 -2725
rect 2085 -2755 2115 -2725
rect 2165 -2755 2195 -2725
rect 2245 -2755 2275 -2725
rect 2325 -2755 2355 -2725
rect 2405 -2755 2435 -2725
rect 2485 -2755 2515 -2725
rect 2565 -2755 2595 -2725
rect 2645 -2755 2675 -2725
rect 2725 -2755 2755 -2725
rect 2805 -2755 2835 -2725
rect 2885 -2755 2915 -2725
rect 2965 -2755 2995 -2725
rect 3045 -2755 3075 -2725
rect 3125 -2755 3155 -2725
rect 3205 -2755 3235 -2725
rect 3285 -2755 3315 -2725
rect 3365 -2755 3395 -2725
rect 3445 -2755 3475 -2725
rect 3525 -2755 3555 -2725
rect 3605 -2755 3635 -2725
rect 3685 -2755 3715 -2725
rect 3765 -2755 3795 -2725
rect 3845 -2755 3875 -2725
rect 3925 -2755 3955 -2725
rect 4005 -2755 4035 -2725
rect 4085 -2755 4115 -2725
rect 4165 -2755 4195 -2725
rect 4245 -2755 4275 -2725
rect 4325 -2755 4355 -2725
rect 4405 -2755 4435 -2725
rect 4485 -2755 4515 -2725
rect 4565 -2755 4595 -2725
rect 4645 -2755 4675 -2725
rect 4725 -2755 4755 -2725
rect 4805 -2755 4835 -2725
rect 4885 -2755 4915 -2725
rect 4965 -2755 4995 -2725
rect 5045 -2755 5075 -2725
rect 5125 -2755 5155 -2725
rect 5205 -2755 5235 -2725
rect 5285 -2755 5315 -2725
rect 5365 -2755 5395 -2725
rect 5445 -2755 5475 -2725
rect 5525 -2755 5555 -2725
rect 5605 -2755 5635 -2725
rect 5685 -2755 5715 -2725
rect 5765 -2755 5795 -2725
rect 5845 -2755 5875 -2725
rect 5925 -2755 5955 -2725
rect 6005 -2755 6035 -2725
rect 6085 -2755 6115 -2725
rect 6165 -2755 6195 -2725
rect 6245 -2755 6275 -2725
rect 6325 -2755 6355 -2725
rect 6405 -2755 6435 -2725
rect 6485 -2755 6515 -2725
rect 6565 -2755 6595 -2725
rect 6645 -2755 6675 -2725
rect 6725 -2755 6755 -2725
rect 6805 -2755 6835 -2725
rect 6885 -2755 6915 -2725
rect 6965 -2755 6995 -2725
rect 7045 -2755 7075 -2725
rect 7125 -2755 7155 -2725
rect 7205 -2755 7235 -2725
rect 7285 -2755 7315 -2725
rect 7365 -2755 7395 -2725
rect 7445 -2755 7475 -2725
rect 7525 -2755 7555 -2725
rect 7605 -2755 7635 -2725
rect 7685 -2755 7715 -2725
rect 7765 -2755 7795 -2725
rect 7845 -2755 7875 -2725
rect 7925 -2755 7955 -2725
rect 8005 -2755 8035 -2725
rect 8085 -2755 8115 -2725
rect 8165 -2755 8195 -2725
rect 8245 -2755 8275 -2725
rect 8325 -2755 8355 -2725
rect 8405 -2755 8435 -2725
rect 8485 -2755 8515 -2725
rect 8565 -2755 8595 -2725
rect 8645 -2755 8675 -2725
rect 8725 -2755 8755 -2725
rect 8805 -2755 8835 -2725
rect 8885 -2755 8915 -2725
rect 8965 -2755 8995 -2725
rect 9045 -2755 9075 -2725
rect 9125 -2755 9155 -2725
rect 9205 -2755 9235 -2725
rect 9285 -2755 9315 -2725
rect 9365 -2755 9395 -2725
rect 9445 -2755 9475 -2725
rect 9525 -2755 9555 -2725
rect 9605 -2755 9635 -2725
rect 9685 -2755 9715 -2725
rect 9765 -2755 9795 -2725
rect 9845 -2755 9875 -2725
rect 9925 -2755 9955 -2725
rect 10005 -2755 10035 -2725
rect 10085 -2755 10115 -2725
rect 10165 -2755 10195 -2725
rect 10245 -2755 10275 -2725
rect 10325 -2755 10355 -2725
rect 10405 -2755 10435 -2725
rect 10485 -2755 10515 -2725
rect 10645 -2755 10675 -2725
rect 10805 -2755 10835 -2725
rect 10965 -2755 10995 -2725
rect -715 -2835 -685 -2805
rect -555 -2835 -525 -2805
rect -395 -2835 -365 -2805
rect 10725 -2835 10755 -2805
rect 10805 -2835 10835 -2805
rect 10965 -2835 10995 -2805
rect -715 -2915 -685 -2885
rect -555 -2915 -525 -2885
rect -395 -2915 -365 -2885
rect -315 -2915 -285 -2885
rect -235 -2915 -205 -2885
rect -155 -2915 -125 -2885
rect -75 -2915 -45 -2885
rect 5 -2915 35 -2885
rect 85 -2915 115 -2885
rect 165 -2915 195 -2885
rect 245 -2915 275 -2885
rect 325 -2915 355 -2885
rect 405 -2915 435 -2885
rect 485 -2915 515 -2885
rect 565 -2915 595 -2885
rect 645 -2915 675 -2885
rect 725 -2915 755 -2885
rect 805 -2915 835 -2885
rect 885 -2915 915 -2885
rect 965 -2915 995 -2885
rect 1045 -2915 1075 -2885
rect 1125 -2915 1155 -2885
rect 1205 -2915 1235 -2885
rect 1285 -2915 1315 -2885
rect 1365 -2915 1395 -2885
rect 1445 -2915 1475 -2885
rect 1525 -2915 1555 -2885
rect 1605 -2915 1635 -2885
rect 1685 -2915 1715 -2885
rect 1765 -2915 1795 -2885
rect 1845 -2915 1875 -2885
rect 1925 -2915 1955 -2885
rect 2005 -2915 2035 -2885
rect 2085 -2915 2115 -2885
rect 2165 -2915 2195 -2885
rect 2245 -2915 2275 -2885
rect 2325 -2915 2355 -2885
rect 2405 -2915 2435 -2885
rect 2485 -2915 2515 -2885
rect 2565 -2915 2595 -2885
rect 2645 -2915 2675 -2885
rect 2725 -2915 2755 -2885
rect 2805 -2915 2835 -2885
rect 2885 -2915 2915 -2885
rect 2965 -2915 2995 -2885
rect 3045 -2915 3075 -2885
rect 3125 -2915 3155 -2885
rect 3205 -2915 3235 -2885
rect 3285 -2915 3315 -2885
rect 3365 -2915 3395 -2885
rect 3445 -2915 3475 -2885
rect 3525 -2915 3555 -2885
rect 3605 -2915 3635 -2885
rect 3685 -2915 3715 -2885
rect 3765 -2915 3795 -2885
rect 3845 -2915 3875 -2885
rect 3925 -2915 3955 -2885
rect 4005 -2915 4035 -2885
rect 4085 -2915 4115 -2885
rect 4165 -2915 4195 -2885
rect 4245 -2915 4275 -2885
rect 4325 -2915 4355 -2885
rect 4405 -2915 4435 -2885
rect 4485 -2915 4515 -2885
rect 4565 -2915 4595 -2885
rect 4645 -2915 4675 -2885
rect 4725 -2915 4755 -2885
rect 4805 -2915 4835 -2885
rect 4885 -2915 4915 -2885
rect 4965 -2915 4995 -2885
rect 5045 -2915 5075 -2885
rect 5125 -2915 5155 -2885
rect 5205 -2915 5235 -2885
rect 5285 -2915 5315 -2885
rect 5365 -2915 5395 -2885
rect 5445 -2915 5475 -2885
rect 5525 -2915 5555 -2885
rect 5605 -2915 5635 -2885
rect 5685 -2915 5715 -2885
rect 5765 -2915 5795 -2885
rect 5845 -2915 5875 -2885
rect 5925 -2915 5955 -2885
rect 6005 -2915 6035 -2885
rect 6085 -2915 6115 -2885
rect 6165 -2915 6195 -2885
rect 6245 -2915 6275 -2885
rect 6325 -2915 6355 -2885
rect 6405 -2915 6435 -2885
rect 6485 -2915 6515 -2885
rect 6565 -2915 6595 -2885
rect 6645 -2915 6675 -2885
rect 6725 -2915 6755 -2885
rect 6805 -2915 6835 -2885
rect 6885 -2915 6915 -2885
rect 6965 -2915 6995 -2885
rect 7045 -2915 7075 -2885
rect 7125 -2915 7155 -2885
rect 7205 -2915 7235 -2885
rect 7285 -2915 7315 -2885
rect 7365 -2915 7395 -2885
rect 7445 -2915 7475 -2885
rect 7525 -2915 7555 -2885
rect 7605 -2915 7635 -2885
rect 7685 -2915 7715 -2885
rect 7765 -2915 7795 -2885
rect 7845 -2915 7875 -2885
rect 7925 -2915 7955 -2885
rect 8005 -2915 8035 -2885
rect 8085 -2915 8115 -2885
rect 8165 -2915 8195 -2885
rect 8245 -2915 8275 -2885
rect 8325 -2915 8355 -2885
rect 8405 -2915 8435 -2885
rect 8485 -2915 8515 -2885
rect 8565 -2915 8595 -2885
rect 8645 -2915 8675 -2885
rect 8725 -2915 8755 -2885
rect 8805 -2915 8835 -2885
rect 8885 -2915 8915 -2885
rect 8965 -2915 8995 -2885
rect 9045 -2915 9075 -2885
rect 9125 -2915 9155 -2885
rect 9205 -2915 9235 -2885
rect 9285 -2915 9315 -2885
rect 9365 -2915 9395 -2885
rect 9445 -2915 9475 -2885
rect 9525 -2915 9555 -2885
rect 9605 -2915 9635 -2885
rect 9685 -2915 9715 -2885
rect 9765 -2915 9795 -2885
rect 9845 -2915 9875 -2885
rect 9925 -2915 9955 -2885
rect 10005 -2915 10035 -2885
rect 10085 -2915 10115 -2885
rect 10165 -2915 10195 -2885
rect 10245 -2915 10275 -2885
rect 10325 -2915 10355 -2885
rect 10405 -2915 10435 -2885
rect 10485 -2915 10515 -2885
rect 10645 -2915 10675 -2885
rect 10805 -2915 10835 -2885
rect 10965 -2915 10995 -2885
rect -715 -2995 -685 -2965
rect -555 -2995 -525 -2965
rect -395 -2995 -365 -2965
rect 10885 -2995 10915 -2965
rect -715 -3075 -685 -3045
rect -555 -3075 -525 -3045
rect -395 -3075 -365 -3045
rect -315 -3075 -285 -3045
rect -235 -3075 -205 -3045
rect -155 -3075 -125 -3045
rect -75 -3075 -45 -3045
rect 5 -3075 35 -3045
rect 85 -3075 115 -3045
rect 165 -3075 195 -3045
rect 245 -3075 275 -3045
rect 325 -3075 355 -3045
rect 405 -3075 435 -3045
rect 485 -3075 515 -3045
rect 565 -3075 595 -3045
rect 645 -3075 675 -3045
rect 725 -3075 755 -3045
rect 805 -3075 835 -3045
rect 885 -3075 915 -3045
rect 965 -3075 995 -3045
rect 1045 -3075 1075 -3045
rect 1125 -3075 1155 -3045
rect 1205 -3075 1235 -3045
rect 1285 -3075 1315 -3045
rect 1365 -3075 1395 -3045
rect 1445 -3075 1475 -3045
rect 1525 -3075 1555 -3045
rect 1605 -3075 1635 -3045
rect 1685 -3075 1715 -3045
rect 1765 -3075 1795 -3045
rect 1845 -3075 1875 -3045
rect 1925 -3075 1955 -3045
rect 2005 -3075 2035 -3045
rect 2085 -3075 2115 -3045
rect 2165 -3075 2195 -3045
rect 2245 -3075 2275 -3045
rect 2325 -3075 2355 -3045
rect 2405 -3075 2435 -3045
rect 2485 -3075 2515 -3045
rect 2565 -3075 2595 -3045
rect 2645 -3075 2675 -3045
rect 2725 -3075 2755 -3045
rect 2805 -3075 2835 -3045
rect 2885 -3075 2915 -3045
rect 2965 -3075 2995 -3045
rect 3045 -3075 3075 -3045
rect 3125 -3075 3155 -3045
rect 3205 -3075 3235 -3045
rect 3285 -3075 3315 -3045
rect 3365 -3075 3395 -3045
rect 3445 -3075 3475 -3045
rect 3525 -3075 3555 -3045
rect 3605 -3075 3635 -3045
rect 3685 -3075 3715 -3045
rect 3765 -3075 3795 -3045
rect 3845 -3075 3875 -3045
rect 3925 -3075 3955 -3045
rect 4005 -3075 4035 -3045
rect 4085 -3075 4115 -3045
rect 4165 -3075 4195 -3045
rect 4245 -3075 4275 -3045
rect 4325 -3075 4355 -3045
rect 4405 -3075 4435 -3045
rect 4485 -3075 4515 -3045
rect 4565 -3075 4595 -3045
rect 4645 -3075 4675 -3045
rect 4725 -3075 4755 -3045
rect 4805 -3075 4835 -3045
rect 4885 -3075 4915 -3045
rect 4965 -3075 4995 -3045
rect 5045 -3075 5075 -3045
rect 5125 -3075 5155 -3045
rect 5205 -3075 5235 -3045
rect 5285 -3075 5315 -3045
rect 5365 -3075 5395 -3045
rect 5445 -3075 5475 -3045
rect 5525 -3075 5555 -3045
rect 5605 -3075 5635 -3045
rect 5685 -3075 5715 -3045
rect 5765 -3075 5795 -3045
rect 5845 -3075 5875 -3045
rect 5925 -3075 5955 -3045
rect 6005 -3075 6035 -3045
rect 6085 -3075 6115 -3045
rect 6165 -3075 6195 -3045
rect 6245 -3075 6275 -3045
rect 6325 -3075 6355 -3045
rect 6405 -3075 6435 -3045
rect 6485 -3075 6515 -3045
rect 6565 -3075 6595 -3045
rect 6645 -3075 6675 -3045
rect 6725 -3075 6755 -3045
rect 6805 -3075 6835 -3045
rect 6885 -3075 6915 -3045
rect 6965 -3075 6995 -3045
rect 7045 -3075 7075 -3045
rect 7125 -3075 7155 -3045
rect 7205 -3075 7235 -3045
rect 7285 -3075 7315 -3045
rect 7365 -3075 7395 -3045
rect 7445 -3075 7475 -3045
rect 7525 -3075 7555 -3045
rect 7605 -3075 7635 -3045
rect 7685 -3075 7715 -3045
rect 7765 -3075 7795 -3045
rect 7845 -3075 7875 -3045
rect 7925 -3075 7955 -3045
rect 8005 -3075 8035 -3045
rect 8085 -3075 8115 -3045
rect 8165 -3075 8195 -3045
rect 8245 -3075 8275 -3045
rect 8325 -3075 8355 -3045
rect 8405 -3075 8435 -3045
rect 8485 -3075 8515 -3045
rect 8565 -3075 8595 -3045
rect 8645 -3075 8675 -3045
rect 8725 -3075 8755 -3045
rect 8805 -3075 8835 -3045
rect 8885 -3075 8915 -3045
rect 8965 -3075 8995 -3045
rect 9045 -3075 9075 -3045
rect 9125 -3075 9155 -3045
rect 9205 -3075 9235 -3045
rect 9285 -3075 9315 -3045
rect 9365 -3075 9395 -3045
rect 9445 -3075 9475 -3045
rect 9525 -3075 9555 -3045
rect 9605 -3075 9635 -3045
rect 9685 -3075 9715 -3045
rect 9765 -3075 9795 -3045
rect 9845 -3075 9875 -3045
rect 9925 -3075 9955 -3045
rect 10005 -3075 10035 -3045
rect 10085 -3075 10115 -3045
rect 10165 -3075 10195 -3045
rect 10245 -3075 10275 -3045
rect 10325 -3075 10355 -3045
rect 10405 -3075 10435 -3045
rect 10485 -3075 10515 -3045
rect 10645 -3075 10675 -3045
rect 10805 -3075 10835 -3045
rect 10965 -3075 10995 -3045
rect -715 -3155 -685 -3125
rect -555 -3155 -525 -3125
rect -475 -3155 -445 -3125
rect 10645 -3155 10675 -3125
rect 10805 -3155 10835 -3125
rect 10965 -3155 10995 -3125
rect -715 -3235 -685 -3205
rect -555 -3235 -525 -3205
rect -395 -3235 -365 -3205
rect -315 -3235 -285 -3205
rect -235 -3235 -205 -3205
rect -155 -3235 -125 -3205
rect -75 -3235 -45 -3205
rect 5 -3235 35 -3205
rect 85 -3235 115 -3205
rect 165 -3235 195 -3205
rect 245 -3235 275 -3205
rect 325 -3235 355 -3205
rect 405 -3235 435 -3205
rect 485 -3235 515 -3205
rect 565 -3235 595 -3205
rect 645 -3235 675 -3205
rect 725 -3235 755 -3205
rect 805 -3235 835 -3205
rect 885 -3235 915 -3205
rect 965 -3235 995 -3205
rect 1045 -3235 1075 -3205
rect 1125 -3235 1155 -3205
rect 1205 -3235 1235 -3205
rect 1285 -3235 1315 -3205
rect 1365 -3235 1395 -3205
rect 1445 -3235 1475 -3205
rect 1525 -3235 1555 -3205
rect 1605 -3235 1635 -3205
rect 1685 -3235 1715 -3205
rect 1765 -3235 1795 -3205
rect 1845 -3235 1875 -3205
rect 1925 -3235 1955 -3205
rect 2005 -3235 2035 -3205
rect 2085 -3235 2115 -3205
rect 2165 -3235 2195 -3205
rect 2245 -3235 2275 -3205
rect 2325 -3235 2355 -3205
rect 2405 -3235 2435 -3205
rect 2485 -3235 2515 -3205
rect 2565 -3235 2595 -3205
rect 2645 -3235 2675 -3205
rect 2725 -3235 2755 -3205
rect 2805 -3235 2835 -3205
rect 2885 -3235 2915 -3205
rect 2965 -3235 2995 -3205
rect 3045 -3235 3075 -3205
rect 3125 -3235 3155 -3205
rect 3205 -3235 3235 -3205
rect 3285 -3235 3315 -3205
rect 3365 -3235 3395 -3205
rect 3445 -3235 3475 -3205
rect 3525 -3235 3555 -3205
rect 3605 -3235 3635 -3205
rect 3685 -3235 3715 -3205
rect 3765 -3235 3795 -3205
rect 3845 -3235 3875 -3205
rect 3925 -3235 3955 -3205
rect 4005 -3235 4035 -3205
rect 4085 -3235 4115 -3205
rect 4165 -3235 4195 -3205
rect 4245 -3235 4275 -3205
rect 4325 -3235 4355 -3205
rect 4405 -3235 4435 -3205
rect 4485 -3235 4515 -3205
rect 4565 -3235 4595 -3205
rect 4645 -3235 4675 -3205
rect 4725 -3235 4755 -3205
rect 4805 -3235 4835 -3205
rect 4885 -3235 4915 -3205
rect 4965 -3235 4995 -3205
rect 5045 -3235 5075 -3205
rect 5125 -3235 5155 -3205
rect 5205 -3235 5235 -3205
rect 5285 -3235 5315 -3205
rect 5365 -3235 5395 -3205
rect 5445 -3235 5475 -3205
rect 5525 -3235 5555 -3205
rect 5605 -3235 5635 -3205
rect 5685 -3235 5715 -3205
rect 5765 -3235 5795 -3205
rect 5845 -3235 5875 -3205
rect 5925 -3235 5955 -3205
rect 6005 -3235 6035 -3205
rect 6085 -3235 6115 -3205
rect 6165 -3235 6195 -3205
rect 6245 -3235 6275 -3205
rect 6325 -3235 6355 -3205
rect 6405 -3235 6435 -3205
rect 6485 -3235 6515 -3205
rect 6565 -3235 6595 -3205
rect 6645 -3235 6675 -3205
rect 6725 -3235 6755 -3205
rect 6805 -3235 6835 -3205
rect 6885 -3235 6915 -3205
rect 6965 -3235 6995 -3205
rect 7045 -3235 7075 -3205
rect 7125 -3235 7155 -3205
rect 7205 -3235 7235 -3205
rect 7285 -3235 7315 -3205
rect 7365 -3235 7395 -3205
rect 7445 -3235 7475 -3205
rect 7525 -3235 7555 -3205
rect 7605 -3235 7635 -3205
rect 7685 -3235 7715 -3205
rect 7765 -3235 7795 -3205
rect 7845 -3235 7875 -3205
rect 7925 -3235 7955 -3205
rect 8005 -3235 8035 -3205
rect 8085 -3235 8115 -3205
rect 8165 -3235 8195 -3205
rect 8245 -3235 8275 -3205
rect 8325 -3235 8355 -3205
rect 8405 -3235 8435 -3205
rect 8485 -3235 8515 -3205
rect 8565 -3235 8595 -3205
rect 8645 -3235 8675 -3205
rect 8725 -3235 8755 -3205
rect 8805 -3235 8835 -3205
rect 8885 -3235 8915 -3205
rect 8965 -3235 8995 -3205
rect 9045 -3235 9075 -3205
rect 9125 -3235 9155 -3205
rect 9205 -3235 9235 -3205
rect 9285 -3235 9315 -3205
rect 9365 -3235 9395 -3205
rect 9445 -3235 9475 -3205
rect 9525 -3235 9555 -3205
rect 9605 -3235 9635 -3205
rect 9685 -3235 9715 -3205
rect 9765 -3235 9795 -3205
rect 9845 -3235 9875 -3205
rect 9925 -3235 9955 -3205
rect 10005 -3235 10035 -3205
rect 10085 -3235 10115 -3205
rect 10165 -3235 10195 -3205
rect 10245 -3235 10275 -3205
rect 10325 -3235 10355 -3205
rect 10405 -3235 10435 -3205
rect 10485 -3235 10515 -3205
rect 10645 -3235 10675 -3205
rect 10805 -3235 10835 -3205
rect 10965 -3235 10995 -3205
rect -715 -3315 -685 -3285
rect -555 -3315 -525 -3285
rect -395 -3315 -365 -3285
rect -315 -3315 -285 -3285
rect -235 -3315 -205 -3285
rect -155 -3315 -125 -3285
rect -75 -3315 -45 -3285
rect 5 -3315 35 -3285
rect 85 -3315 115 -3285
rect 165 -3315 195 -3285
rect 245 -3315 275 -3285
rect 325 -3315 355 -3285
rect 405 -3315 435 -3285
rect 485 -3315 515 -3285
rect 565 -3315 595 -3285
rect 645 -3315 675 -3285
rect 725 -3315 755 -3285
rect 805 -3315 835 -3285
rect 885 -3315 915 -3285
rect 965 -3315 995 -3285
rect 1045 -3315 1075 -3285
rect 1125 -3315 1155 -3285
rect 1205 -3315 1235 -3285
rect 1285 -3315 1315 -3285
rect 1365 -3315 1395 -3285
rect 1445 -3315 1475 -3285
rect 1525 -3315 1555 -3285
rect 1605 -3315 1635 -3285
rect 1685 -3315 1715 -3285
rect 1765 -3315 1795 -3285
rect 1845 -3315 1875 -3285
rect 1925 -3315 1955 -3285
rect 2005 -3315 2035 -3285
rect 2085 -3315 2115 -3285
rect 2165 -3315 2195 -3285
rect 2245 -3315 2275 -3285
rect 2325 -3315 2355 -3285
rect 2405 -3315 2435 -3285
rect 2485 -3315 2515 -3285
rect 2565 -3315 2595 -3285
rect 2645 -3315 2675 -3285
rect 2725 -3315 2755 -3285
rect 2805 -3315 2835 -3285
rect 2885 -3315 2915 -3285
rect 2965 -3315 2995 -3285
rect 3045 -3315 3075 -3285
rect 3125 -3315 3155 -3285
rect 3205 -3315 3235 -3285
rect 3285 -3315 3315 -3285
rect 3365 -3315 3395 -3285
rect 3445 -3315 3475 -3285
rect 3525 -3315 3555 -3285
rect 3605 -3315 3635 -3285
rect 3685 -3315 3715 -3285
rect 3765 -3315 3795 -3285
rect 3845 -3315 3875 -3285
rect 3925 -3315 3955 -3285
rect 4005 -3315 4035 -3285
rect 4085 -3315 4115 -3285
rect 4165 -3315 4195 -3285
rect 4245 -3315 4275 -3285
rect 4325 -3315 4355 -3285
rect 4405 -3315 4435 -3285
rect 4485 -3315 4515 -3285
rect 4565 -3315 4595 -3285
rect 4645 -3315 4675 -3285
rect 4725 -3315 4755 -3285
rect 4805 -3315 4835 -3285
rect 4885 -3315 4915 -3285
rect 4965 -3315 4995 -3285
rect 5045 -3315 5075 -3285
rect 5125 -3315 5155 -3285
rect 5205 -3315 5235 -3285
rect 5285 -3315 5315 -3285
rect 5365 -3315 5395 -3285
rect 5445 -3315 5475 -3285
rect 5525 -3315 5555 -3285
rect 5605 -3315 5635 -3285
rect 5685 -3315 5715 -3285
rect 5765 -3315 5795 -3285
rect 5845 -3315 5875 -3285
rect 5925 -3315 5955 -3285
rect 6005 -3315 6035 -3285
rect 6085 -3315 6115 -3285
rect 6165 -3315 6195 -3285
rect 6245 -3315 6275 -3285
rect 6325 -3315 6355 -3285
rect 6405 -3315 6435 -3285
rect 6485 -3315 6515 -3285
rect 6565 -3315 6595 -3285
rect 6645 -3315 6675 -3285
rect 6725 -3315 6755 -3285
rect 6805 -3315 6835 -3285
rect 6885 -3315 6915 -3285
rect 6965 -3315 6995 -3285
rect 7045 -3315 7075 -3285
rect 7125 -3315 7155 -3285
rect 7205 -3315 7235 -3285
rect 7285 -3315 7315 -3285
rect 7365 -3315 7395 -3285
rect 7445 -3315 7475 -3285
rect 7525 -3315 7555 -3285
rect 7605 -3315 7635 -3285
rect 7685 -3315 7715 -3285
rect 7765 -3315 7795 -3285
rect 7845 -3315 7875 -3285
rect 7925 -3315 7955 -3285
rect 8005 -3315 8035 -3285
rect 8085 -3315 8115 -3285
rect 8165 -3315 8195 -3285
rect 8245 -3315 8275 -3285
rect 8325 -3315 8355 -3285
rect 8405 -3315 8435 -3285
rect 8485 -3315 8515 -3285
rect 8565 -3315 8595 -3285
rect 8645 -3315 8675 -3285
rect 8725 -3315 8755 -3285
rect 8805 -3315 8835 -3285
rect 8885 -3315 8915 -3285
rect 8965 -3315 8995 -3285
rect 9045 -3315 9075 -3285
rect 9125 -3315 9155 -3285
rect 9205 -3315 9235 -3285
rect 9285 -3315 9315 -3285
rect 9365 -3315 9395 -3285
rect 9445 -3315 9475 -3285
rect 9525 -3315 9555 -3285
rect 9605 -3315 9635 -3285
rect 9685 -3315 9715 -3285
rect 9765 -3315 9795 -3285
rect 9845 -3315 9875 -3285
rect 9925 -3315 9955 -3285
rect 10005 -3315 10035 -3285
rect 10085 -3315 10115 -3285
rect 10165 -3315 10195 -3285
rect 10245 -3315 10275 -3285
rect 10325 -3315 10355 -3285
rect 10405 -3315 10435 -3285
rect 10485 -3315 10515 -3285
rect 10645 -3315 10675 -3285
rect 10805 -3315 10835 -3285
rect 10965 -3315 10995 -3285
rect -635 -3395 -605 -3365
rect 10645 -3395 10675 -3365
rect 10805 -3395 10835 -3365
rect 10965 -3395 10995 -3365
rect -635 -3475 -605 -3445
rect 10645 -3475 10675 -3445
rect 10805 -3475 10835 -3445
rect 10965 -3475 10995 -3445
rect -715 -3555 -685 -3525
rect -555 -3555 -525 -3525
rect -395 -3555 -365 -3525
rect -315 -3555 -285 -3525
rect -235 -3555 -205 -3525
rect -155 -3555 -125 -3525
rect -75 -3555 -45 -3525
rect 5 -3555 35 -3525
rect 85 -3555 115 -3525
rect 165 -3555 195 -3525
rect 245 -3555 275 -3525
rect 325 -3555 355 -3525
rect 405 -3555 435 -3525
rect 485 -3555 515 -3525
rect 565 -3555 595 -3525
rect 645 -3555 675 -3525
rect 725 -3555 755 -3525
rect 805 -3555 835 -3525
rect 885 -3555 915 -3525
rect 965 -3555 995 -3525
rect 1045 -3555 1075 -3525
rect 1125 -3555 1155 -3525
rect 1205 -3555 1235 -3525
rect 1285 -3555 1315 -3525
rect 1365 -3555 1395 -3525
rect 1445 -3555 1475 -3525
rect 1525 -3555 1555 -3525
rect 1605 -3555 1635 -3525
rect 1685 -3555 1715 -3525
rect 1765 -3555 1795 -3525
rect 1845 -3555 1875 -3525
rect 1925 -3555 1955 -3525
rect 2005 -3555 2035 -3525
rect 2085 -3555 2115 -3525
rect 2165 -3555 2195 -3525
rect 2245 -3555 2275 -3525
rect 2325 -3555 2355 -3525
rect 2405 -3555 2435 -3525
rect 2485 -3555 2515 -3525
rect 2565 -3555 2595 -3525
rect 2645 -3555 2675 -3525
rect 2725 -3555 2755 -3525
rect 2805 -3555 2835 -3525
rect 2885 -3555 2915 -3525
rect 2965 -3555 2995 -3525
rect 3045 -3555 3075 -3525
rect 3125 -3555 3155 -3525
rect 3205 -3555 3235 -3525
rect 3285 -3555 3315 -3525
rect 3365 -3555 3395 -3525
rect 3445 -3555 3475 -3525
rect 3525 -3555 3555 -3525
rect 3605 -3555 3635 -3525
rect 3685 -3555 3715 -3525
rect 3765 -3555 3795 -3525
rect 3845 -3555 3875 -3525
rect 3925 -3555 3955 -3525
rect 4005 -3555 4035 -3525
rect 4085 -3555 4115 -3525
rect 4165 -3555 4195 -3525
rect 4245 -3555 4275 -3525
rect 4325 -3555 4355 -3525
rect 4405 -3555 4435 -3525
rect 4485 -3555 4515 -3525
rect 4565 -3555 4595 -3525
rect 4645 -3555 4675 -3525
rect 4725 -3555 4755 -3525
rect 4805 -3555 4835 -3525
rect 4885 -3555 4915 -3525
rect 4965 -3555 4995 -3525
rect 5045 -3555 5075 -3525
rect 5125 -3555 5155 -3525
rect 5205 -3555 5235 -3525
rect 5285 -3555 5315 -3525
rect 5365 -3555 5395 -3525
rect 5445 -3555 5475 -3525
rect 5525 -3555 5555 -3525
rect 5605 -3555 5635 -3525
rect 5685 -3555 5715 -3525
rect 5765 -3555 5795 -3525
rect 5845 -3555 5875 -3525
rect 5925 -3555 5955 -3525
rect 6005 -3555 6035 -3525
rect 6085 -3555 6115 -3525
rect 6165 -3555 6195 -3525
rect 6245 -3555 6275 -3525
rect 6325 -3555 6355 -3525
rect 6405 -3555 6435 -3525
rect 6485 -3555 6515 -3525
rect 6565 -3555 6595 -3525
rect 6645 -3555 6675 -3525
rect 6725 -3555 6755 -3525
rect 6805 -3555 6835 -3525
rect 6885 -3555 6915 -3525
rect 6965 -3555 6995 -3525
rect 7045 -3555 7075 -3525
rect 7125 -3555 7155 -3525
rect 7205 -3555 7235 -3525
rect 7285 -3555 7315 -3525
rect 7365 -3555 7395 -3525
rect 7445 -3555 7475 -3525
rect 7525 -3555 7555 -3525
rect 7605 -3555 7635 -3525
rect 7685 -3555 7715 -3525
rect 7765 -3555 7795 -3525
rect 7845 -3555 7875 -3525
rect 7925 -3555 7955 -3525
rect 8005 -3555 8035 -3525
rect 8085 -3555 8115 -3525
rect 8165 -3555 8195 -3525
rect 8245 -3555 8275 -3525
rect 8325 -3555 8355 -3525
rect 8405 -3555 8435 -3525
rect 8485 -3555 8515 -3525
rect 8565 -3555 8595 -3525
rect 8645 -3555 8675 -3525
rect 8725 -3555 8755 -3525
rect 8805 -3555 8835 -3525
rect 8885 -3555 8915 -3525
rect 8965 -3555 8995 -3525
rect 9045 -3555 9075 -3525
rect 9125 -3555 9155 -3525
rect 9205 -3555 9235 -3525
rect 9285 -3555 9315 -3525
rect 9365 -3555 9395 -3525
rect 9445 -3555 9475 -3525
rect 9525 -3555 9555 -3525
rect 9605 -3555 9635 -3525
rect 9685 -3555 9715 -3525
rect 9765 -3555 9795 -3525
rect 9845 -3555 9875 -3525
rect 9925 -3555 9955 -3525
rect 10005 -3555 10035 -3525
rect 10085 -3555 10115 -3525
rect 10165 -3555 10195 -3525
rect 10245 -3555 10275 -3525
rect 10325 -3555 10355 -3525
rect 10405 -3555 10435 -3525
rect 10485 -3555 10515 -3525
rect 10645 -3555 10675 -3525
rect 10805 -3555 10835 -3525
rect 10965 -3555 10995 -3525
rect -715 -3635 -685 -3605
rect -555 -3635 -525 -3605
rect -395 -3635 -365 -3605
rect -315 -3635 -285 -3605
rect -235 -3635 -205 -3605
rect -155 -3635 -125 -3605
rect -75 -3635 -45 -3605
rect 5 -3635 35 -3605
rect 85 -3635 115 -3605
rect 165 -3635 195 -3605
rect 245 -3635 275 -3605
rect 325 -3635 355 -3605
rect 405 -3635 435 -3605
rect 485 -3635 515 -3605
rect 565 -3635 595 -3605
rect 645 -3635 675 -3605
rect 725 -3635 755 -3605
rect 805 -3635 835 -3605
rect 885 -3635 915 -3605
rect 965 -3635 995 -3605
rect 1045 -3635 1075 -3605
rect 1125 -3635 1155 -3605
rect 1205 -3635 1235 -3605
rect 1285 -3635 1315 -3605
rect 1365 -3635 1395 -3605
rect 1445 -3635 1475 -3605
rect 1525 -3635 1555 -3605
rect 1605 -3635 1635 -3605
rect 1685 -3635 1715 -3605
rect 1765 -3635 1795 -3605
rect 1845 -3635 1875 -3605
rect 1925 -3635 1955 -3605
rect 2005 -3635 2035 -3605
rect 2085 -3635 2115 -3605
rect 2165 -3635 2195 -3605
rect 2245 -3635 2275 -3605
rect 2325 -3635 2355 -3605
rect 2405 -3635 2435 -3605
rect 2485 -3635 2515 -3605
rect 2565 -3635 2595 -3605
rect 2645 -3635 2675 -3605
rect 2725 -3635 2755 -3605
rect 2805 -3635 2835 -3605
rect 2885 -3635 2915 -3605
rect 2965 -3635 2995 -3605
rect 3045 -3635 3075 -3605
rect 3125 -3635 3155 -3605
rect 3205 -3635 3235 -3605
rect 3285 -3635 3315 -3605
rect 3365 -3635 3395 -3605
rect 3445 -3635 3475 -3605
rect 3525 -3635 3555 -3605
rect 3605 -3635 3635 -3605
rect 3685 -3635 3715 -3605
rect 3765 -3635 3795 -3605
rect 3845 -3635 3875 -3605
rect 3925 -3635 3955 -3605
rect 4005 -3635 4035 -3605
rect 4085 -3635 4115 -3605
rect 4165 -3635 4195 -3605
rect 4245 -3635 4275 -3605
rect 4325 -3635 4355 -3605
rect 4405 -3635 4435 -3605
rect 4485 -3635 4515 -3605
rect 4565 -3635 4595 -3605
rect 4645 -3635 4675 -3605
rect 4725 -3635 4755 -3605
rect 4805 -3635 4835 -3605
rect 4885 -3635 4915 -3605
rect 4965 -3635 4995 -3605
rect 5045 -3635 5075 -3605
rect 5125 -3635 5155 -3605
rect 5205 -3635 5235 -3605
rect 5285 -3635 5315 -3605
rect 5365 -3635 5395 -3605
rect 5445 -3635 5475 -3605
rect 5525 -3635 5555 -3605
rect 5605 -3635 5635 -3605
rect 5685 -3635 5715 -3605
rect 5765 -3635 5795 -3605
rect 5845 -3635 5875 -3605
rect 5925 -3635 5955 -3605
rect 6005 -3635 6035 -3605
rect 6085 -3635 6115 -3605
rect 6165 -3635 6195 -3605
rect 6245 -3635 6275 -3605
rect 6325 -3635 6355 -3605
rect 6405 -3635 6435 -3605
rect 6485 -3635 6515 -3605
rect 6565 -3635 6595 -3605
rect 6645 -3635 6675 -3605
rect 6725 -3635 6755 -3605
rect 6805 -3635 6835 -3605
rect 6885 -3635 6915 -3605
rect 6965 -3635 6995 -3605
rect 7045 -3635 7075 -3605
rect 7125 -3635 7155 -3605
rect 7205 -3635 7235 -3605
rect 7285 -3635 7315 -3605
rect 7365 -3635 7395 -3605
rect 7445 -3635 7475 -3605
rect 7525 -3635 7555 -3605
rect 7605 -3635 7635 -3605
rect 7685 -3635 7715 -3605
rect 7765 -3635 7795 -3605
rect 7845 -3635 7875 -3605
rect 7925 -3635 7955 -3605
rect 8005 -3635 8035 -3605
rect 8085 -3635 8115 -3605
rect 8165 -3635 8195 -3605
rect 8245 -3635 8275 -3605
rect 8325 -3635 8355 -3605
rect 8405 -3635 8435 -3605
rect 8485 -3635 8515 -3605
rect 8565 -3635 8595 -3605
rect 8645 -3635 8675 -3605
rect 8725 -3635 8755 -3605
rect 8805 -3635 8835 -3605
rect 8885 -3635 8915 -3605
rect 8965 -3635 8995 -3605
rect 9045 -3635 9075 -3605
rect 9125 -3635 9155 -3605
rect 9205 -3635 9235 -3605
rect 9285 -3635 9315 -3605
rect 9365 -3635 9395 -3605
rect 9445 -3635 9475 -3605
rect 9525 -3635 9555 -3605
rect 9605 -3635 9635 -3605
rect 9685 -3635 9715 -3605
rect 9765 -3635 9795 -3605
rect 9845 -3635 9875 -3605
rect 9925 -3635 9955 -3605
rect 10005 -3635 10035 -3605
rect 10085 -3635 10115 -3605
rect 10165 -3635 10195 -3605
rect 10245 -3635 10275 -3605
rect 10325 -3635 10355 -3605
rect 10405 -3635 10435 -3605
rect 10485 -3635 10515 -3605
rect 10645 -3635 10675 -3605
rect 10805 -3635 10835 -3605
rect 10965 -3635 10995 -3605
rect -715 -3715 -685 -3685
rect -555 -3715 -525 -3685
rect -395 -3715 -365 -3685
rect -315 -3715 -285 -3685
rect -235 -3715 -205 -3685
rect -155 -3715 -125 -3685
rect -75 -3715 -45 -3685
rect 5 -3715 35 -3685
rect 85 -3715 115 -3685
rect 165 -3715 195 -3685
rect 245 -3715 275 -3685
rect 325 -3715 355 -3685
rect 405 -3715 435 -3685
rect 485 -3715 515 -3685
rect 565 -3715 595 -3685
rect 645 -3715 675 -3685
rect 725 -3715 755 -3685
rect 805 -3715 835 -3685
rect 885 -3715 915 -3685
rect 965 -3715 995 -3685
rect 1045 -3715 1075 -3685
rect 1125 -3715 1155 -3685
rect 1205 -3715 1235 -3685
rect 1285 -3715 1315 -3685
rect 1365 -3715 1395 -3685
rect 1445 -3715 1475 -3685
rect 1525 -3715 1555 -3685
rect 1605 -3715 1635 -3685
rect 1685 -3715 1715 -3685
rect 1765 -3715 1795 -3685
rect 1845 -3715 1875 -3685
rect 1925 -3715 1955 -3685
rect 2005 -3715 2035 -3685
rect 2085 -3715 2115 -3685
rect 2165 -3715 2195 -3685
rect 2245 -3715 2275 -3685
rect 2325 -3715 2355 -3685
rect 2405 -3715 2435 -3685
rect 2485 -3715 2515 -3685
rect 2565 -3715 2595 -3685
rect 2645 -3715 2675 -3685
rect 2725 -3715 2755 -3685
rect 2805 -3715 2835 -3685
rect 2885 -3715 2915 -3685
rect 2965 -3715 2995 -3685
rect 3045 -3715 3075 -3685
rect 3125 -3715 3155 -3685
rect 3205 -3715 3235 -3685
rect 3285 -3715 3315 -3685
rect 3365 -3715 3395 -3685
rect 3445 -3715 3475 -3685
rect 3525 -3715 3555 -3685
rect 3605 -3715 3635 -3685
rect 3685 -3715 3715 -3685
rect 3765 -3715 3795 -3685
rect 3845 -3715 3875 -3685
rect 3925 -3715 3955 -3685
rect 4005 -3715 4035 -3685
rect 4085 -3715 4115 -3685
rect 4165 -3715 4195 -3685
rect 4245 -3715 4275 -3685
rect 4325 -3715 4355 -3685
rect 4405 -3715 4435 -3685
rect 4485 -3715 4515 -3685
rect 4565 -3715 4595 -3685
rect 4645 -3715 4675 -3685
rect 4725 -3715 4755 -3685
rect 4805 -3715 4835 -3685
rect 4885 -3715 4915 -3685
rect 4965 -3715 4995 -3685
rect 5045 -3715 5075 -3685
rect 5125 -3715 5155 -3685
rect 5205 -3715 5235 -3685
rect 5285 -3715 5315 -3685
rect 5365 -3715 5395 -3685
rect 5445 -3715 5475 -3685
rect 5525 -3715 5555 -3685
rect 5605 -3715 5635 -3685
rect 5685 -3715 5715 -3685
rect 5765 -3715 5795 -3685
rect 5845 -3715 5875 -3685
rect 5925 -3715 5955 -3685
rect 6005 -3715 6035 -3685
rect 6085 -3715 6115 -3685
rect 6165 -3715 6195 -3685
rect 6245 -3715 6275 -3685
rect 6325 -3715 6355 -3685
rect 6405 -3715 6435 -3685
rect 6485 -3715 6515 -3685
rect 6565 -3715 6595 -3685
rect 6645 -3715 6675 -3685
rect 6725 -3715 6755 -3685
rect 6805 -3715 6835 -3685
rect 6885 -3715 6915 -3685
rect 6965 -3715 6995 -3685
rect 7045 -3715 7075 -3685
rect 7125 -3715 7155 -3685
rect 7205 -3715 7235 -3685
rect 7285 -3715 7315 -3685
rect 7365 -3715 7395 -3685
rect 7445 -3715 7475 -3685
rect 7525 -3715 7555 -3685
rect 7605 -3715 7635 -3685
rect 7685 -3715 7715 -3685
rect 7765 -3715 7795 -3685
rect 7845 -3715 7875 -3685
rect 7925 -3715 7955 -3685
rect 8005 -3715 8035 -3685
rect 8085 -3715 8115 -3685
rect 8165 -3715 8195 -3685
rect 8245 -3715 8275 -3685
rect 8325 -3715 8355 -3685
rect 8405 -3715 8435 -3685
rect 8485 -3715 8515 -3685
rect 8565 -3715 8595 -3685
rect 8645 -3715 8675 -3685
rect 8725 -3715 8755 -3685
rect 8805 -3715 8835 -3685
rect 8885 -3715 8915 -3685
rect 8965 -3715 8995 -3685
rect 9045 -3715 9075 -3685
rect 9125 -3715 9155 -3685
rect 9205 -3715 9235 -3685
rect 9285 -3715 9315 -3685
rect 9365 -3715 9395 -3685
rect 9445 -3715 9475 -3685
rect 9525 -3715 9555 -3685
rect 9605 -3715 9635 -3685
rect 9685 -3715 9715 -3685
rect 9765 -3715 9795 -3685
rect 9845 -3715 9875 -3685
rect 9925 -3715 9955 -3685
rect 10005 -3715 10035 -3685
rect 10085 -3715 10115 -3685
rect 10165 -3715 10195 -3685
rect 10245 -3715 10275 -3685
rect 10325 -3715 10355 -3685
rect 10405 -3715 10435 -3685
rect 10485 -3715 10515 -3685
rect 10645 -3715 10675 -3685
rect 10805 -3715 10835 -3685
rect 10965 -3715 10995 -3685
<< metal3 >>
rect -720 1036 -680 1040
rect -720 1004 -716 1036
rect -684 1004 -680 1036
rect -720 956 -680 1004
rect -720 924 -716 956
rect -684 924 -680 956
rect -720 876 -680 924
rect -720 844 -716 876
rect -684 844 -680 876
rect -720 796 -680 844
rect -720 764 -716 796
rect -684 764 -680 796
rect -720 716 -680 764
rect -720 684 -716 716
rect -684 684 -680 716
rect -720 636 -680 684
rect -720 604 -716 636
rect -684 604 -680 636
rect -720 556 -680 604
rect -720 524 -716 556
rect -684 524 -680 556
rect -720 476 -680 524
rect -720 444 -716 476
rect -684 444 -680 476
rect -720 396 -680 444
rect -720 364 -716 396
rect -684 364 -680 396
rect -720 316 -680 364
rect -720 284 -716 316
rect -684 284 -680 316
rect -720 236 -680 284
rect -720 204 -716 236
rect -684 204 -680 236
rect -720 156 -680 204
rect -720 124 -716 156
rect -684 124 -680 156
rect -720 76 -680 124
rect -720 44 -716 76
rect -684 44 -680 76
rect -720 -4 -680 44
rect -720 -36 -716 -4
rect -684 -36 -680 -4
rect -720 -84 -680 -36
rect -720 -116 -716 -84
rect -684 -116 -680 -84
rect -720 -164 -680 -116
rect -720 -196 -716 -164
rect -684 -196 -680 -164
rect -720 -244 -680 -196
rect -720 -276 -716 -244
rect -684 -276 -680 -244
rect -720 -324 -680 -276
rect -720 -356 -716 -324
rect -684 -356 -680 -324
rect -720 -404 -680 -356
rect -720 -436 -716 -404
rect -684 -436 -680 -404
rect -720 -484 -680 -436
rect -720 -516 -716 -484
rect -684 -516 -680 -484
rect -720 -564 -680 -516
rect -720 -596 -716 -564
rect -684 -596 -680 -564
rect -720 -644 -680 -596
rect -720 -676 -716 -644
rect -684 -676 -680 -644
rect -720 -724 -680 -676
rect -720 -756 -716 -724
rect -684 -756 -680 -724
rect -720 -804 -680 -756
rect -720 -836 -716 -804
rect -684 -836 -680 -804
rect -720 -884 -680 -836
rect -720 -916 -716 -884
rect -684 -916 -680 -884
rect -720 -964 -680 -916
rect -720 -996 -716 -964
rect -684 -996 -680 -964
rect -720 -1044 -680 -996
rect -720 -1076 -716 -1044
rect -684 -1076 -680 -1044
rect -720 -1124 -680 -1076
rect -720 -1156 -716 -1124
rect -684 -1156 -680 -1124
rect -720 -1204 -680 -1156
rect -720 -1236 -716 -1204
rect -684 -1236 -680 -1204
rect -720 -1284 -680 -1236
rect -720 -1316 -716 -1284
rect -684 -1316 -680 -1284
rect -720 -1364 -680 -1316
rect -720 -1396 -716 -1364
rect -684 -1396 -680 -1364
rect -720 -1444 -680 -1396
rect -720 -1476 -716 -1444
rect -684 -1476 -680 -1444
rect -720 -1524 -680 -1476
rect -720 -1556 -716 -1524
rect -684 -1556 -680 -1524
rect -720 -1604 -680 -1556
rect -720 -1636 -716 -1604
rect -684 -1636 -680 -1604
rect -720 -1684 -680 -1636
rect -720 -1716 -716 -1684
rect -684 -1716 -680 -1684
rect -720 -1764 -680 -1716
rect -720 -1796 -716 -1764
rect -684 -1796 -680 -1764
rect -720 -1844 -680 -1796
rect -720 -1876 -716 -1844
rect -684 -1876 -680 -1844
rect -720 -1924 -680 -1876
rect -720 -1956 -716 -1924
rect -684 -1956 -680 -1924
rect -720 -2004 -680 -1956
rect -720 -2036 -716 -2004
rect -684 -2036 -680 -2004
rect -720 -2084 -680 -2036
rect -720 -2116 -716 -2084
rect -684 -2116 -680 -2084
rect -720 -2164 -680 -2116
rect -720 -2196 -716 -2164
rect -684 -2196 -680 -2164
rect -720 -2244 -680 -2196
rect -720 -2276 -716 -2244
rect -684 -2276 -680 -2244
rect -720 -2324 -680 -2276
rect -720 -2356 -716 -2324
rect -684 -2356 -680 -2324
rect -720 -2404 -680 -2356
rect -720 -2436 -716 -2404
rect -684 -2436 -680 -2404
rect -720 -2484 -680 -2436
rect -720 -2516 -716 -2484
rect -684 -2516 -680 -2484
rect -720 -2564 -680 -2516
rect -720 -2596 -716 -2564
rect -684 -2596 -680 -2564
rect -720 -2644 -680 -2596
rect -720 -2676 -716 -2644
rect -684 -2676 -680 -2644
rect -720 -2724 -680 -2676
rect -720 -2756 -716 -2724
rect -684 -2756 -680 -2724
rect -720 -2804 -680 -2756
rect -720 -2836 -716 -2804
rect -684 -2836 -680 -2804
rect -720 -2884 -680 -2836
rect -720 -2916 -716 -2884
rect -684 -2916 -680 -2884
rect -720 -2964 -680 -2916
rect -720 -2996 -716 -2964
rect -684 -2996 -680 -2964
rect -720 -3044 -680 -2996
rect -720 -3076 -716 -3044
rect -684 -3076 -680 -3044
rect -720 -3124 -680 -3076
rect -720 -3156 -716 -3124
rect -684 -3156 -680 -3124
rect -720 -3204 -680 -3156
rect -720 -3236 -716 -3204
rect -684 -3236 -680 -3204
rect -720 -3284 -680 -3236
rect -720 -3316 -716 -3284
rect -684 -3316 -680 -3284
rect -720 -3364 -680 -3316
rect -720 -3396 -716 -3364
rect -684 -3396 -680 -3364
rect -720 -3444 -680 -3396
rect -720 -3476 -716 -3444
rect -684 -3476 -680 -3444
rect -720 -3524 -680 -3476
rect -720 -3556 -716 -3524
rect -684 -3556 -680 -3524
rect -720 -3604 -680 -3556
rect -720 -3636 -716 -3604
rect -684 -3636 -680 -3604
rect -720 -3684 -680 -3636
rect -720 -3716 -716 -3684
rect -684 -3716 -680 -3684
rect -720 -3720 -680 -3716
rect -640 795 -600 1080
rect -640 765 -635 795
rect -605 765 -600 795
rect -640 715 -600 765
rect -640 685 -635 715
rect -605 685 -600 715
rect -640 -965 -600 685
rect -640 -995 -635 -965
rect -605 -995 -600 -965
rect -640 -1045 -600 -995
rect -640 -1075 -635 -1045
rect -605 -1075 -600 -1045
rect -640 -1605 -600 -1075
rect -640 -1635 -635 -1605
rect -605 -1635 -600 -1605
rect -640 -1685 -600 -1635
rect -640 -1715 -635 -1685
rect -605 -1715 -600 -1685
rect -640 -3365 -600 -1715
rect -640 -3395 -635 -3365
rect -605 -3395 -600 -3365
rect -640 -3445 -600 -3395
rect -640 -3475 -635 -3445
rect -605 -3475 -600 -3445
rect -640 -3720 -600 -3475
rect -560 1036 -520 1040
rect -560 1004 -556 1036
rect -524 1004 -520 1036
rect -560 956 -520 1004
rect -560 924 -556 956
rect -524 924 -520 956
rect -560 876 -520 924
rect -560 844 -556 876
rect -524 844 -520 876
rect -560 796 -520 844
rect -560 764 -556 796
rect -524 764 -520 796
rect -560 716 -520 764
rect -560 684 -556 716
rect -524 684 -520 716
rect -560 636 -520 684
rect -560 604 -556 636
rect -524 604 -520 636
rect -560 556 -520 604
rect -560 524 -556 556
rect -524 524 -520 556
rect -560 476 -520 524
rect -560 444 -556 476
rect -524 444 -520 476
rect -560 396 -520 444
rect -560 364 -556 396
rect -524 364 -520 396
rect -560 316 -520 364
rect -560 284 -556 316
rect -524 284 -520 316
rect -560 236 -520 284
rect -560 204 -556 236
rect -524 204 -520 236
rect -560 156 -520 204
rect -560 124 -556 156
rect -524 124 -520 156
rect -560 76 -520 124
rect -560 44 -556 76
rect -524 44 -520 76
rect -560 -4 -520 44
rect -560 -36 -556 -4
rect -524 -36 -520 -4
rect -560 -84 -520 -36
rect -560 -116 -556 -84
rect -524 -116 -520 -84
rect -560 -164 -520 -116
rect -560 -196 -556 -164
rect -524 -196 -520 -164
rect -560 -244 -520 -196
rect -560 -276 -556 -244
rect -524 -276 -520 -244
rect -560 -324 -520 -276
rect -560 -356 -556 -324
rect -524 -356 -520 -324
rect -560 -404 -520 -356
rect -560 -436 -556 -404
rect -524 -436 -520 -404
rect -560 -484 -520 -436
rect -560 -516 -556 -484
rect -524 -516 -520 -484
rect -560 -564 -520 -516
rect -560 -596 -556 -564
rect -524 -596 -520 -564
rect -560 -644 -520 -596
rect -560 -676 -556 -644
rect -524 -676 -520 -644
rect -560 -724 -520 -676
rect -560 -756 -556 -724
rect -524 -756 -520 -724
rect -560 -804 -520 -756
rect -560 -836 -556 -804
rect -524 -836 -520 -804
rect -560 -884 -520 -836
rect -560 -916 -556 -884
rect -524 -916 -520 -884
rect -560 -964 -520 -916
rect -560 -996 -556 -964
rect -524 -996 -520 -964
rect -560 -1044 -520 -996
rect -560 -1076 -556 -1044
rect -524 -1076 -520 -1044
rect -560 -1124 -520 -1076
rect -560 -1156 -556 -1124
rect -524 -1156 -520 -1124
rect -560 -1204 -520 -1156
rect -560 -1236 -556 -1204
rect -524 -1236 -520 -1204
rect -560 -1284 -520 -1236
rect -560 -1316 -556 -1284
rect -524 -1316 -520 -1284
rect -560 -1364 -520 -1316
rect -560 -1396 -556 -1364
rect -524 -1396 -520 -1364
rect -560 -1444 -520 -1396
rect -560 -1476 -556 -1444
rect -524 -1476 -520 -1444
rect -560 -1524 -520 -1476
rect -560 -1556 -556 -1524
rect -524 -1556 -520 -1524
rect -560 -1604 -520 -1556
rect -560 -1636 -556 -1604
rect -524 -1636 -520 -1604
rect -560 -1684 -520 -1636
rect -560 -1716 -556 -1684
rect -524 -1716 -520 -1684
rect -560 -1764 -520 -1716
rect -560 -1796 -556 -1764
rect -524 -1796 -520 -1764
rect -560 -1844 -520 -1796
rect -560 -1876 -556 -1844
rect -524 -1876 -520 -1844
rect -560 -1924 -520 -1876
rect -560 -1956 -556 -1924
rect -524 -1956 -520 -1924
rect -560 -2004 -520 -1956
rect -560 -2036 -556 -2004
rect -524 -2036 -520 -2004
rect -560 -2084 -520 -2036
rect -560 -2116 -556 -2084
rect -524 -2116 -520 -2084
rect -560 -2164 -520 -2116
rect -560 -2196 -556 -2164
rect -524 -2196 -520 -2164
rect -560 -2244 -520 -2196
rect -560 -2276 -556 -2244
rect -524 -2276 -520 -2244
rect -560 -2324 -520 -2276
rect -560 -2356 -556 -2324
rect -524 -2356 -520 -2324
rect -560 -2404 -520 -2356
rect -560 -2436 -556 -2404
rect -524 -2436 -520 -2404
rect -560 -2484 -520 -2436
rect -560 -2516 -556 -2484
rect -524 -2516 -520 -2484
rect -560 -2564 -520 -2516
rect -560 -2596 -556 -2564
rect -524 -2596 -520 -2564
rect -560 -2644 -520 -2596
rect -560 -2676 -556 -2644
rect -524 -2676 -520 -2644
rect -560 -2724 -520 -2676
rect -560 -2756 -556 -2724
rect -524 -2756 -520 -2724
rect -560 -2804 -520 -2756
rect -560 -2836 -556 -2804
rect -524 -2836 -520 -2804
rect -560 -2884 -520 -2836
rect -560 -2916 -556 -2884
rect -524 -2916 -520 -2884
rect -560 -2964 -520 -2916
rect -560 -2996 -556 -2964
rect -524 -2996 -520 -2964
rect -560 -3044 -520 -2996
rect -560 -3076 -556 -3044
rect -524 -3076 -520 -3044
rect -560 -3124 -520 -3076
rect -560 -3156 -556 -3124
rect -524 -3156 -520 -3124
rect -560 -3204 -520 -3156
rect -560 -3236 -556 -3204
rect -524 -3236 -520 -3204
rect -560 -3284 -520 -3236
rect -560 -3316 -556 -3284
rect -524 -3316 -520 -3284
rect -560 -3364 -520 -3316
rect -560 -3396 -556 -3364
rect -524 -3396 -520 -3364
rect -560 -3444 -520 -3396
rect -560 -3476 -556 -3444
rect -524 -3476 -520 -3444
rect -560 -3524 -520 -3476
rect -560 -3556 -556 -3524
rect -524 -3556 -520 -3524
rect -560 -3604 -520 -3556
rect -560 -3636 -556 -3604
rect -524 -3636 -520 -3604
rect -560 -3684 -520 -3636
rect -560 -3716 -556 -3684
rect -524 -3716 -520 -3684
rect -560 -3720 -520 -3716
rect -480 475 -440 1080
rect -480 445 -475 475
rect -445 445 -440 475
rect -480 -725 -440 445
rect -480 -755 -475 -725
rect -445 -755 -440 -725
rect -480 -1925 -440 -755
rect -480 -1955 -475 -1925
rect -445 -1955 -440 -1925
rect -480 -3125 -440 -1955
rect -480 -3155 -475 -3125
rect -445 -3155 -440 -3125
rect -480 -3720 -440 -3155
rect -400 1036 -360 1040
rect -400 1004 -396 1036
rect -364 1004 -360 1036
rect -400 956 -360 1004
rect -400 924 -396 956
rect -364 924 -360 956
rect -400 876 -360 924
rect -400 844 -396 876
rect -364 844 -360 876
rect -400 796 -360 844
rect -400 764 -396 796
rect -364 764 -360 796
rect -400 716 -360 764
rect -400 684 -396 716
rect -364 684 -360 716
rect -400 636 -360 684
rect -400 604 -396 636
rect -364 604 -360 636
rect -400 556 -360 604
rect -400 524 -396 556
rect -364 524 -360 556
rect -400 476 -360 524
rect -400 444 -396 476
rect -364 444 -360 476
rect -400 396 -360 444
rect -400 364 -396 396
rect -364 364 -360 396
rect -400 316 -360 364
rect -400 284 -396 316
rect -364 284 -360 316
rect -400 236 -360 284
rect -400 204 -396 236
rect -364 204 -360 236
rect -400 156 -360 204
rect -400 124 -396 156
rect -364 124 -360 156
rect -400 76 -360 124
rect -400 44 -396 76
rect -364 44 -360 76
rect -400 -4 -360 44
rect -400 -36 -396 -4
rect -364 -36 -360 -4
rect -400 -84 -360 -36
rect -400 -116 -396 -84
rect -364 -116 -360 -84
rect -400 -164 -360 -116
rect -400 -196 -396 -164
rect -364 -196 -360 -164
rect -400 -244 -360 -196
rect -400 -276 -396 -244
rect -364 -276 -360 -244
rect -400 -324 -360 -276
rect -400 -356 -396 -324
rect -364 -356 -360 -324
rect -400 -404 -360 -356
rect -400 -436 -396 -404
rect -364 -436 -360 -404
rect -400 -484 -360 -436
rect -400 -516 -396 -484
rect -364 -516 -360 -484
rect -400 -564 -360 -516
rect -400 -596 -396 -564
rect -364 -596 -360 -564
rect -400 -644 -360 -596
rect -400 -676 -396 -644
rect -364 -676 -360 -644
rect -400 -724 -360 -676
rect -400 -756 -396 -724
rect -364 -756 -360 -724
rect -400 -804 -360 -756
rect -400 -836 -396 -804
rect -364 -836 -360 -804
rect -400 -884 -360 -836
rect -400 -916 -396 -884
rect -364 -916 -360 -884
rect -400 -964 -360 -916
rect -400 -996 -396 -964
rect -364 -996 -360 -964
rect -400 -1044 -360 -996
rect -400 -1076 -396 -1044
rect -364 -1076 -360 -1044
rect -400 -1124 -360 -1076
rect -400 -1156 -396 -1124
rect -364 -1156 -360 -1124
rect -400 -1204 -360 -1156
rect -400 -1236 -396 -1204
rect -364 -1236 -360 -1204
rect -400 -1284 -360 -1236
rect -400 -1316 -396 -1284
rect -364 -1316 -360 -1284
rect -400 -1364 -360 -1316
rect -400 -1396 -396 -1364
rect -364 -1396 -360 -1364
rect -400 -1444 -360 -1396
rect -400 -1476 -396 -1444
rect -364 -1476 -360 -1444
rect -400 -1524 -360 -1476
rect -400 -1556 -396 -1524
rect -364 -1556 -360 -1524
rect -400 -1604 -360 -1556
rect -400 -1636 -396 -1604
rect -364 -1636 -360 -1604
rect -400 -1684 -360 -1636
rect -400 -1716 -396 -1684
rect -364 -1716 -360 -1684
rect -400 -1764 -360 -1716
rect -400 -1796 -396 -1764
rect -364 -1796 -360 -1764
rect -400 -1844 -360 -1796
rect -400 -1876 -396 -1844
rect -364 -1876 -360 -1844
rect -400 -1924 -360 -1876
rect -400 -1956 -396 -1924
rect -364 -1956 -360 -1924
rect -400 -2004 -360 -1956
rect -400 -2036 -396 -2004
rect -364 -2036 -360 -2004
rect -400 -2084 -360 -2036
rect -400 -2116 -396 -2084
rect -364 -2116 -360 -2084
rect -400 -2164 -360 -2116
rect -400 -2196 -396 -2164
rect -364 -2196 -360 -2164
rect -400 -2244 -360 -2196
rect -400 -2276 -396 -2244
rect -364 -2276 -360 -2244
rect -400 -2324 -360 -2276
rect -400 -2356 -396 -2324
rect -364 -2356 -360 -2324
rect -400 -2404 -360 -2356
rect -400 -2436 -396 -2404
rect -364 -2436 -360 -2404
rect -400 -2484 -360 -2436
rect -400 -2516 -396 -2484
rect -364 -2516 -360 -2484
rect -400 -2564 -360 -2516
rect -400 -2596 -396 -2564
rect -364 -2596 -360 -2564
rect -400 -2644 -360 -2596
rect -400 -2676 -396 -2644
rect -364 -2676 -360 -2644
rect -400 -2724 -360 -2676
rect -400 -2756 -396 -2724
rect -364 -2756 -360 -2724
rect -400 -2804 -360 -2756
rect -400 -2836 -396 -2804
rect -364 -2836 -360 -2804
rect -400 -2884 -360 -2836
rect -400 -2916 -396 -2884
rect -364 -2916 -360 -2884
rect -400 -2964 -360 -2916
rect -400 -2996 -396 -2964
rect -364 -2996 -360 -2964
rect -400 -3044 -360 -2996
rect -400 -3076 -396 -3044
rect -364 -3076 -360 -3044
rect -400 -3124 -360 -3076
rect -400 -3156 -396 -3124
rect -364 -3156 -360 -3124
rect -400 -3204 -360 -3156
rect -400 -3236 -396 -3204
rect -364 -3236 -360 -3204
rect -400 -3284 -360 -3236
rect -400 -3316 -396 -3284
rect -364 -3316 -360 -3284
rect -400 -3364 -360 -3316
rect -400 -3396 -396 -3364
rect -364 -3396 -360 -3364
rect -400 -3444 -360 -3396
rect -400 -3476 -396 -3444
rect -364 -3476 -360 -3444
rect -400 -3524 -360 -3476
rect -400 -3556 -396 -3524
rect -364 -3556 -360 -3524
rect -400 -3604 -360 -3556
rect -400 -3636 -396 -3604
rect -364 -3636 -360 -3604
rect -400 -3684 -360 -3636
rect -400 -3716 -396 -3684
rect -364 -3716 -360 -3684
rect -400 -3720 -360 -3716
rect -320 1036 -280 1040
rect -320 1004 -316 1036
rect -284 1004 -280 1036
rect -320 956 -280 1004
rect -320 924 -316 956
rect -284 924 -280 956
rect -320 876 -280 924
rect -320 844 -316 876
rect -284 844 -280 876
rect -320 796 -280 844
rect -320 764 -316 796
rect -284 764 -280 796
rect -320 716 -280 764
rect -320 684 -316 716
rect -284 684 -280 716
rect -320 636 -280 684
rect -320 604 -316 636
rect -284 604 -280 636
rect -320 556 -280 604
rect -320 524 -316 556
rect -284 524 -280 556
rect -320 476 -280 524
rect -320 444 -316 476
rect -284 444 -280 476
rect -320 396 -280 444
rect -320 364 -316 396
rect -284 364 -280 396
rect -320 316 -280 364
rect -320 284 -316 316
rect -284 284 -280 316
rect -320 236 -280 284
rect -320 204 -316 236
rect -284 204 -280 236
rect -320 156 -280 204
rect -320 124 -316 156
rect -284 124 -280 156
rect -320 76 -280 124
rect -320 44 -316 76
rect -284 44 -280 76
rect -320 -4 -280 44
rect -320 -36 -316 -4
rect -284 -36 -280 -4
rect -320 -84 -280 -36
rect -320 -116 -316 -84
rect -284 -116 -280 -84
rect -320 -2564 -280 -116
rect -320 -2596 -316 -2564
rect -284 -2596 -280 -2564
rect -320 -2644 -280 -2596
rect -320 -2676 -316 -2644
rect -284 -2676 -280 -2644
rect -320 -2724 -280 -2676
rect -320 -2756 -316 -2724
rect -284 -2756 -280 -2724
rect -320 -2804 -280 -2756
rect -320 -2836 -316 -2804
rect -284 -2836 -280 -2804
rect -320 -2884 -280 -2836
rect -320 -2916 -316 -2884
rect -284 -2916 -280 -2884
rect -320 -2964 -280 -2916
rect -320 -2996 -316 -2964
rect -284 -2996 -280 -2964
rect -320 -3044 -280 -2996
rect -320 -3076 -316 -3044
rect -284 -3076 -280 -3044
rect -320 -3124 -280 -3076
rect -320 -3156 -316 -3124
rect -284 -3156 -280 -3124
rect -320 -3204 -280 -3156
rect -320 -3236 -316 -3204
rect -284 -3236 -280 -3204
rect -320 -3284 -280 -3236
rect -320 -3316 -316 -3284
rect -284 -3316 -280 -3284
rect -320 -3364 -280 -3316
rect -320 -3396 -316 -3364
rect -284 -3396 -280 -3364
rect -320 -3444 -280 -3396
rect -320 -3476 -316 -3444
rect -284 -3476 -280 -3444
rect -320 -3524 -280 -3476
rect -320 -3556 -316 -3524
rect -284 -3556 -280 -3524
rect -320 -3604 -280 -3556
rect -320 -3636 -316 -3604
rect -284 -3636 -280 -3604
rect -320 -3684 -280 -3636
rect -320 -3716 -316 -3684
rect -284 -3716 -280 -3684
rect -320 -3720 -280 -3716
rect -240 1036 -200 1040
rect -240 1004 -236 1036
rect -204 1004 -200 1036
rect -240 956 -200 1004
rect -240 924 -236 956
rect -204 924 -200 956
rect -240 876 -200 924
rect -240 844 -236 876
rect -204 844 -200 876
rect -240 796 -200 844
rect -240 764 -236 796
rect -204 764 -200 796
rect -240 716 -200 764
rect -240 684 -236 716
rect -204 684 -200 716
rect -240 636 -200 684
rect -240 604 -236 636
rect -204 604 -200 636
rect -240 556 -200 604
rect -240 524 -236 556
rect -204 524 -200 556
rect -240 476 -200 524
rect -240 444 -236 476
rect -204 444 -200 476
rect -240 396 -200 444
rect -240 364 -236 396
rect -204 364 -200 396
rect -240 316 -200 364
rect -240 284 -236 316
rect -204 284 -200 316
rect -240 236 -200 284
rect -240 204 -236 236
rect -204 204 -200 236
rect -240 156 -200 204
rect -240 124 -236 156
rect -204 124 -200 156
rect -240 76 -200 124
rect -240 44 -236 76
rect -204 44 -200 76
rect -240 -4 -200 44
rect -240 -36 -236 -4
rect -204 -36 -200 -4
rect -240 -84 -200 -36
rect -240 -116 -236 -84
rect -204 -116 -200 -84
rect -240 -164 -200 -116
rect -240 -196 -236 -164
rect -204 -196 -200 -164
rect -240 -244 -200 -196
rect -240 -276 -236 -244
rect -204 -276 -200 -244
rect -240 -324 -200 -276
rect -240 -356 -236 -324
rect -204 -356 -200 -324
rect -240 -404 -200 -356
rect -240 -436 -236 -404
rect -204 -436 -200 -404
rect -240 -484 -200 -436
rect -240 -516 -236 -484
rect -204 -516 -200 -484
rect -240 -564 -200 -516
rect -240 -596 -236 -564
rect -204 -596 -200 -564
rect -240 -644 -200 -596
rect -240 -676 -236 -644
rect -204 -676 -200 -644
rect -240 -724 -200 -676
rect -240 -756 -236 -724
rect -204 -756 -200 -724
rect -240 -804 -200 -756
rect -240 -836 -236 -804
rect -204 -836 -200 -804
rect -240 -884 -200 -836
rect -240 -916 -236 -884
rect -204 -916 -200 -884
rect -240 -964 -200 -916
rect -240 -996 -236 -964
rect -204 -996 -200 -964
rect -240 -1044 -200 -996
rect -240 -1076 -236 -1044
rect -204 -1076 -200 -1044
rect -240 -1124 -200 -1076
rect -240 -1156 -236 -1124
rect -204 -1156 -200 -1124
rect -240 -1204 -200 -1156
rect -240 -1236 -236 -1204
rect -204 -1236 -200 -1204
rect -240 -1284 -200 -1236
rect -240 -1316 -236 -1284
rect -204 -1316 -200 -1284
rect -240 -1364 -200 -1316
rect -240 -1396 -236 -1364
rect -204 -1396 -200 -1364
rect -240 -1444 -200 -1396
rect -240 -1476 -236 -1444
rect -204 -1476 -200 -1444
rect -240 -1524 -200 -1476
rect -240 -1556 -236 -1524
rect -204 -1556 -200 -1524
rect -240 -1604 -200 -1556
rect -240 -1636 -236 -1604
rect -204 -1636 -200 -1604
rect -240 -1684 -200 -1636
rect -240 -1716 -236 -1684
rect -204 -1716 -200 -1684
rect -240 -1764 -200 -1716
rect -240 -1796 -236 -1764
rect -204 -1796 -200 -1764
rect -240 -1844 -200 -1796
rect -240 -1876 -236 -1844
rect -204 -1876 -200 -1844
rect -240 -1924 -200 -1876
rect -240 -1956 -236 -1924
rect -204 -1956 -200 -1924
rect -240 -2004 -200 -1956
rect -240 -2036 -236 -2004
rect -204 -2036 -200 -2004
rect -240 -2084 -200 -2036
rect -240 -2116 -236 -2084
rect -204 -2116 -200 -2084
rect -240 -2164 -200 -2116
rect -240 -2196 -236 -2164
rect -204 -2196 -200 -2164
rect -240 -2244 -200 -2196
rect -240 -2276 -236 -2244
rect -204 -2276 -200 -2244
rect -240 -2324 -200 -2276
rect -240 -2356 -236 -2324
rect -204 -2356 -200 -2324
rect -240 -2404 -200 -2356
rect -240 -2436 -236 -2404
rect -204 -2436 -200 -2404
rect -240 -2484 -200 -2436
rect -240 -2516 -236 -2484
rect -204 -2516 -200 -2484
rect -240 -2564 -200 -2516
rect -240 -2596 -236 -2564
rect -204 -2596 -200 -2564
rect -240 -2644 -200 -2596
rect -240 -2676 -236 -2644
rect -204 -2676 -200 -2644
rect -240 -2724 -200 -2676
rect -240 -2756 -236 -2724
rect -204 -2756 -200 -2724
rect -240 -2804 -200 -2756
rect -240 -2836 -236 -2804
rect -204 -2836 -200 -2804
rect -240 -2884 -200 -2836
rect -240 -2916 -236 -2884
rect -204 -2916 -200 -2884
rect -240 -2964 -200 -2916
rect -240 -2996 -236 -2964
rect -204 -2996 -200 -2964
rect -240 -3044 -200 -2996
rect -240 -3076 -236 -3044
rect -204 -3076 -200 -3044
rect -240 -3124 -200 -3076
rect -240 -3156 -236 -3124
rect -204 -3156 -200 -3124
rect -240 -3204 -200 -3156
rect -240 -3236 -236 -3204
rect -204 -3236 -200 -3204
rect -240 -3284 -200 -3236
rect -240 -3316 -236 -3284
rect -204 -3316 -200 -3284
rect -240 -3364 -200 -3316
rect -240 -3396 -236 -3364
rect -204 -3396 -200 -3364
rect -240 -3444 -200 -3396
rect -240 -3476 -236 -3444
rect -204 -3476 -200 -3444
rect -240 -3524 -200 -3476
rect -240 -3556 -236 -3524
rect -204 -3556 -200 -3524
rect -240 -3604 -200 -3556
rect -240 -3636 -236 -3604
rect -204 -3636 -200 -3604
rect -240 -3684 -200 -3636
rect -240 -3716 -236 -3684
rect -204 -3716 -200 -3684
rect -240 -3720 -200 -3716
rect -160 1036 -120 1040
rect -160 1004 -156 1036
rect -124 1004 -120 1036
rect -160 956 -120 1004
rect -160 924 -156 956
rect -124 924 -120 956
rect -160 876 -120 924
rect -160 844 -156 876
rect -124 844 -120 876
rect -160 796 -120 844
rect -160 764 -156 796
rect -124 764 -120 796
rect -160 716 -120 764
rect -160 684 -156 716
rect -124 684 -120 716
rect -160 636 -120 684
rect -160 604 -156 636
rect -124 604 -120 636
rect -160 556 -120 604
rect -160 524 -156 556
rect -124 524 -120 556
rect -160 476 -120 524
rect -160 444 -156 476
rect -124 444 -120 476
rect -160 396 -120 444
rect -160 364 -156 396
rect -124 364 -120 396
rect -160 316 -120 364
rect -160 284 -156 316
rect -124 284 -120 316
rect -160 236 -120 284
rect -160 204 -156 236
rect -124 204 -120 236
rect -160 156 -120 204
rect -160 124 -156 156
rect -124 124 -120 156
rect -160 76 -120 124
rect -160 44 -156 76
rect -124 44 -120 76
rect -160 -4 -120 44
rect -160 -36 -156 -4
rect -124 -36 -120 -4
rect -160 -84 -120 -36
rect -160 -116 -156 -84
rect -124 -116 -120 -84
rect -160 -164 -120 -116
rect -160 -196 -156 -164
rect -124 -196 -120 -164
rect -160 -244 -120 -196
rect -160 -276 -156 -244
rect -124 -276 -120 -244
rect -160 -324 -120 -276
rect -160 -356 -156 -324
rect -124 -356 -120 -324
rect -160 -404 -120 -356
rect -160 -436 -156 -404
rect -124 -436 -120 -404
rect -160 -484 -120 -436
rect -160 -516 -156 -484
rect -124 -516 -120 -484
rect -160 -564 -120 -516
rect -160 -596 -156 -564
rect -124 -596 -120 -564
rect -160 -644 -120 -596
rect -160 -676 -156 -644
rect -124 -676 -120 -644
rect -160 -724 -120 -676
rect -160 -756 -156 -724
rect -124 -756 -120 -724
rect -160 -804 -120 -756
rect -160 -836 -156 -804
rect -124 -836 -120 -804
rect -160 -884 -120 -836
rect -160 -916 -156 -884
rect -124 -916 -120 -884
rect -160 -964 -120 -916
rect -160 -996 -156 -964
rect -124 -996 -120 -964
rect -160 -1044 -120 -996
rect -160 -1076 -156 -1044
rect -124 -1076 -120 -1044
rect -160 -1124 -120 -1076
rect -160 -1156 -156 -1124
rect -124 -1156 -120 -1124
rect -160 -1204 -120 -1156
rect -160 -1236 -156 -1204
rect -124 -1236 -120 -1204
rect -160 -1284 -120 -1236
rect -160 -1316 -156 -1284
rect -124 -1316 -120 -1284
rect -160 -1364 -120 -1316
rect -160 -1396 -156 -1364
rect -124 -1396 -120 -1364
rect -160 -1444 -120 -1396
rect -160 -1476 -156 -1444
rect -124 -1476 -120 -1444
rect -160 -1524 -120 -1476
rect -160 -1556 -156 -1524
rect -124 -1556 -120 -1524
rect -160 -1604 -120 -1556
rect -160 -1636 -156 -1604
rect -124 -1636 -120 -1604
rect -160 -1684 -120 -1636
rect -160 -1716 -156 -1684
rect -124 -1716 -120 -1684
rect -160 -1764 -120 -1716
rect -160 -1796 -156 -1764
rect -124 -1796 -120 -1764
rect -160 -1844 -120 -1796
rect -160 -1876 -156 -1844
rect -124 -1876 -120 -1844
rect -160 -1924 -120 -1876
rect -160 -1956 -156 -1924
rect -124 -1956 -120 -1924
rect -160 -2004 -120 -1956
rect -160 -2036 -156 -2004
rect -124 -2036 -120 -2004
rect -160 -2084 -120 -2036
rect -160 -2116 -156 -2084
rect -124 -2116 -120 -2084
rect -160 -2164 -120 -2116
rect -160 -2196 -156 -2164
rect -124 -2196 -120 -2164
rect -160 -2244 -120 -2196
rect -160 -2276 -156 -2244
rect -124 -2276 -120 -2244
rect -160 -2324 -120 -2276
rect -160 -2356 -156 -2324
rect -124 -2356 -120 -2324
rect -160 -2404 -120 -2356
rect -160 -2436 -156 -2404
rect -124 -2436 -120 -2404
rect -160 -2484 -120 -2436
rect -160 -2516 -156 -2484
rect -124 -2516 -120 -2484
rect -160 -2564 -120 -2516
rect -160 -2596 -156 -2564
rect -124 -2596 -120 -2564
rect -160 -2644 -120 -2596
rect -160 -2676 -156 -2644
rect -124 -2676 -120 -2644
rect -160 -2724 -120 -2676
rect -160 -2756 -156 -2724
rect -124 -2756 -120 -2724
rect -160 -2804 -120 -2756
rect -160 -2836 -156 -2804
rect -124 -2836 -120 -2804
rect -160 -2884 -120 -2836
rect -160 -2916 -156 -2884
rect -124 -2916 -120 -2884
rect -160 -2964 -120 -2916
rect -160 -2996 -156 -2964
rect -124 -2996 -120 -2964
rect -160 -3044 -120 -2996
rect -160 -3076 -156 -3044
rect -124 -3076 -120 -3044
rect -160 -3124 -120 -3076
rect -160 -3156 -156 -3124
rect -124 -3156 -120 -3124
rect -160 -3204 -120 -3156
rect -160 -3236 -156 -3204
rect -124 -3236 -120 -3204
rect -160 -3284 -120 -3236
rect -160 -3316 -156 -3284
rect -124 -3316 -120 -3284
rect -160 -3364 -120 -3316
rect -160 -3396 -156 -3364
rect -124 -3396 -120 -3364
rect -160 -3444 -120 -3396
rect -160 -3476 -156 -3444
rect -124 -3476 -120 -3444
rect -160 -3524 -120 -3476
rect -160 -3556 -156 -3524
rect -124 -3556 -120 -3524
rect -160 -3604 -120 -3556
rect -160 -3636 -156 -3604
rect -124 -3636 -120 -3604
rect -160 -3684 -120 -3636
rect -160 -3716 -156 -3684
rect -124 -3716 -120 -3684
rect -160 -3720 -120 -3716
rect -80 1036 -40 1040
rect -80 1004 -76 1036
rect -44 1004 -40 1036
rect -80 956 -40 1004
rect -80 924 -76 956
rect -44 924 -40 956
rect -80 876 -40 924
rect -80 844 -76 876
rect -44 844 -40 876
rect -80 796 -40 844
rect -80 764 -76 796
rect -44 764 -40 796
rect -80 716 -40 764
rect -80 684 -76 716
rect -44 684 -40 716
rect -80 636 -40 684
rect -80 604 -76 636
rect -44 604 -40 636
rect -80 556 -40 604
rect -80 524 -76 556
rect -44 524 -40 556
rect -80 476 -40 524
rect -80 444 -76 476
rect -44 444 -40 476
rect -80 396 -40 444
rect -80 364 -76 396
rect -44 364 -40 396
rect -80 316 -40 364
rect -80 284 -76 316
rect -44 284 -40 316
rect -80 236 -40 284
rect -80 204 -76 236
rect -44 204 -40 236
rect -80 156 -40 204
rect -80 124 -76 156
rect -44 124 -40 156
rect -80 76 -40 124
rect -80 44 -76 76
rect -44 44 -40 76
rect -80 -4 -40 44
rect -80 -36 -76 -4
rect -44 -36 -40 -4
rect -80 -84 -40 -36
rect -80 -116 -76 -84
rect -44 -116 -40 -84
rect -80 -164 -40 -116
rect -80 -196 -76 -164
rect -44 -196 -40 -164
rect -80 -244 -40 -196
rect -80 -276 -76 -244
rect -44 -276 -40 -244
rect -80 -324 -40 -276
rect -80 -356 -76 -324
rect -44 -356 -40 -324
rect -80 -404 -40 -356
rect -80 -436 -76 -404
rect -44 -436 -40 -404
rect -80 -484 -40 -436
rect -80 -516 -76 -484
rect -44 -516 -40 -484
rect -80 -564 -40 -516
rect -80 -596 -76 -564
rect -44 -596 -40 -564
rect -80 -644 -40 -596
rect -80 -676 -76 -644
rect -44 -676 -40 -644
rect -80 -724 -40 -676
rect -80 -756 -76 -724
rect -44 -756 -40 -724
rect -80 -804 -40 -756
rect -80 -836 -76 -804
rect -44 -836 -40 -804
rect -80 -884 -40 -836
rect -80 -916 -76 -884
rect -44 -916 -40 -884
rect -80 -964 -40 -916
rect -80 -996 -76 -964
rect -44 -996 -40 -964
rect -80 -1044 -40 -996
rect -80 -1076 -76 -1044
rect -44 -1076 -40 -1044
rect -80 -1124 -40 -1076
rect -80 -1156 -76 -1124
rect -44 -1156 -40 -1124
rect -80 -1204 -40 -1156
rect -80 -1236 -76 -1204
rect -44 -1236 -40 -1204
rect -80 -1284 -40 -1236
rect -80 -1316 -76 -1284
rect -44 -1316 -40 -1284
rect -80 -1364 -40 -1316
rect -80 -1396 -76 -1364
rect -44 -1396 -40 -1364
rect -80 -1444 -40 -1396
rect -80 -1476 -76 -1444
rect -44 -1476 -40 -1444
rect -80 -1524 -40 -1476
rect -80 -1556 -76 -1524
rect -44 -1556 -40 -1524
rect -80 -1604 -40 -1556
rect -80 -1636 -76 -1604
rect -44 -1636 -40 -1604
rect -80 -1684 -40 -1636
rect -80 -1716 -76 -1684
rect -44 -1716 -40 -1684
rect -80 -1764 -40 -1716
rect -80 -1796 -76 -1764
rect -44 -1796 -40 -1764
rect -80 -1844 -40 -1796
rect -80 -1876 -76 -1844
rect -44 -1876 -40 -1844
rect -80 -1924 -40 -1876
rect -80 -1956 -76 -1924
rect -44 -1956 -40 -1924
rect -80 -2004 -40 -1956
rect -80 -2036 -76 -2004
rect -44 -2036 -40 -2004
rect -80 -2084 -40 -2036
rect -80 -2116 -76 -2084
rect -44 -2116 -40 -2084
rect -80 -2164 -40 -2116
rect -80 -2196 -76 -2164
rect -44 -2196 -40 -2164
rect -80 -2244 -40 -2196
rect -80 -2276 -76 -2244
rect -44 -2276 -40 -2244
rect -80 -2324 -40 -2276
rect -80 -2356 -76 -2324
rect -44 -2356 -40 -2324
rect -80 -2404 -40 -2356
rect -80 -2436 -76 -2404
rect -44 -2436 -40 -2404
rect -80 -2484 -40 -2436
rect -80 -2516 -76 -2484
rect -44 -2516 -40 -2484
rect -80 -2564 -40 -2516
rect -80 -2596 -76 -2564
rect -44 -2596 -40 -2564
rect -80 -2644 -40 -2596
rect -80 -2676 -76 -2644
rect -44 -2676 -40 -2644
rect -80 -2724 -40 -2676
rect -80 -2756 -76 -2724
rect -44 -2756 -40 -2724
rect -80 -2804 -40 -2756
rect -80 -2836 -76 -2804
rect -44 -2836 -40 -2804
rect -80 -2884 -40 -2836
rect -80 -2916 -76 -2884
rect -44 -2916 -40 -2884
rect -80 -2964 -40 -2916
rect -80 -2996 -76 -2964
rect -44 -2996 -40 -2964
rect -80 -3044 -40 -2996
rect -80 -3076 -76 -3044
rect -44 -3076 -40 -3044
rect -80 -3124 -40 -3076
rect -80 -3156 -76 -3124
rect -44 -3156 -40 -3124
rect -80 -3204 -40 -3156
rect -80 -3236 -76 -3204
rect -44 -3236 -40 -3204
rect -80 -3284 -40 -3236
rect -80 -3316 -76 -3284
rect -44 -3316 -40 -3284
rect -80 -3364 -40 -3316
rect -80 -3396 -76 -3364
rect -44 -3396 -40 -3364
rect -80 -3444 -40 -3396
rect -80 -3476 -76 -3444
rect -44 -3476 -40 -3444
rect -80 -3524 -40 -3476
rect -80 -3556 -76 -3524
rect -44 -3556 -40 -3524
rect -80 -3604 -40 -3556
rect -80 -3636 -76 -3604
rect -44 -3636 -40 -3604
rect -80 -3684 -40 -3636
rect -80 -3716 -76 -3684
rect -44 -3716 -40 -3684
rect -80 -3720 -40 -3716
rect 0 1036 40 1040
rect 0 1004 4 1036
rect 36 1004 40 1036
rect 0 956 40 1004
rect 0 924 4 956
rect 36 924 40 956
rect 0 876 40 924
rect 0 844 4 876
rect 36 844 40 876
rect 0 796 40 844
rect 0 764 4 796
rect 36 764 40 796
rect 0 716 40 764
rect 0 684 4 716
rect 36 684 40 716
rect 0 636 40 684
rect 0 604 4 636
rect 36 604 40 636
rect 0 556 40 604
rect 0 524 4 556
rect 36 524 40 556
rect 0 476 40 524
rect 0 444 4 476
rect 36 444 40 476
rect 0 396 40 444
rect 0 364 4 396
rect 36 364 40 396
rect 0 316 40 364
rect 0 284 4 316
rect 36 284 40 316
rect 0 236 40 284
rect 0 204 4 236
rect 36 204 40 236
rect 0 156 40 204
rect 0 124 4 156
rect 36 124 40 156
rect 0 76 40 124
rect 0 44 4 76
rect 36 44 40 76
rect 0 -4 40 44
rect 0 -36 4 -4
rect 36 -36 40 -4
rect 0 -84 40 -36
rect 0 -116 4 -84
rect 36 -116 40 -84
rect 0 -164 40 -116
rect 0 -196 4 -164
rect 36 -196 40 -164
rect 0 -244 40 -196
rect 0 -276 4 -244
rect 36 -276 40 -244
rect 0 -324 40 -276
rect 0 -356 4 -324
rect 36 -356 40 -324
rect 0 -404 40 -356
rect 0 -436 4 -404
rect 36 -436 40 -404
rect 0 -484 40 -436
rect 0 -516 4 -484
rect 36 -516 40 -484
rect 0 -564 40 -516
rect 0 -596 4 -564
rect 36 -596 40 -564
rect 0 -644 40 -596
rect 0 -676 4 -644
rect 36 -676 40 -644
rect 0 -724 40 -676
rect 0 -756 4 -724
rect 36 -756 40 -724
rect 0 -804 40 -756
rect 0 -836 4 -804
rect 36 -836 40 -804
rect 0 -884 40 -836
rect 0 -916 4 -884
rect 36 -916 40 -884
rect 0 -964 40 -916
rect 0 -996 4 -964
rect 36 -996 40 -964
rect 0 -1044 40 -996
rect 0 -1076 4 -1044
rect 36 -1076 40 -1044
rect 0 -1124 40 -1076
rect 0 -1156 4 -1124
rect 36 -1156 40 -1124
rect 0 -1204 40 -1156
rect 0 -1236 4 -1204
rect 36 -1236 40 -1204
rect 0 -1284 40 -1236
rect 0 -1316 4 -1284
rect 36 -1316 40 -1284
rect 0 -1364 40 -1316
rect 0 -1396 4 -1364
rect 36 -1396 40 -1364
rect 0 -1444 40 -1396
rect 0 -1476 4 -1444
rect 36 -1476 40 -1444
rect 0 -1524 40 -1476
rect 0 -1556 4 -1524
rect 36 -1556 40 -1524
rect 0 -1604 40 -1556
rect 0 -1636 4 -1604
rect 36 -1636 40 -1604
rect 0 -1684 40 -1636
rect 0 -1716 4 -1684
rect 36 -1716 40 -1684
rect 0 -1764 40 -1716
rect 0 -1796 4 -1764
rect 36 -1796 40 -1764
rect 0 -1844 40 -1796
rect 0 -1876 4 -1844
rect 36 -1876 40 -1844
rect 0 -1924 40 -1876
rect 0 -1956 4 -1924
rect 36 -1956 40 -1924
rect 0 -2004 40 -1956
rect 0 -2036 4 -2004
rect 36 -2036 40 -2004
rect 0 -2084 40 -2036
rect 0 -2116 4 -2084
rect 36 -2116 40 -2084
rect 0 -2164 40 -2116
rect 0 -2196 4 -2164
rect 36 -2196 40 -2164
rect 0 -2244 40 -2196
rect 0 -2276 4 -2244
rect 36 -2276 40 -2244
rect 0 -2324 40 -2276
rect 0 -2356 4 -2324
rect 36 -2356 40 -2324
rect 0 -2404 40 -2356
rect 0 -2436 4 -2404
rect 36 -2436 40 -2404
rect 0 -2484 40 -2436
rect 0 -2516 4 -2484
rect 36 -2516 40 -2484
rect 0 -2564 40 -2516
rect 0 -2596 4 -2564
rect 36 -2596 40 -2564
rect 0 -2644 40 -2596
rect 0 -2676 4 -2644
rect 36 -2676 40 -2644
rect 0 -2724 40 -2676
rect 0 -2756 4 -2724
rect 36 -2756 40 -2724
rect 0 -2804 40 -2756
rect 0 -2836 4 -2804
rect 36 -2836 40 -2804
rect 0 -2884 40 -2836
rect 0 -2916 4 -2884
rect 36 -2916 40 -2884
rect 0 -2964 40 -2916
rect 0 -2996 4 -2964
rect 36 -2996 40 -2964
rect 0 -3044 40 -2996
rect 0 -3076 4 -3044
rect 36 -3076 40 -3044
rect 0 -3124 40 -3076
rect 0 -3156 4 -3124
rect 36 -3156 40 -3124
rect 0 -3204 40 -3156
rect 0 -3236 4 -3204
rect 36 -3236 40 -3204
rect 0 -3284 40 -3236
rect 0 -3316 4 -3284
rect 36 -3316 40 -3284
rect 0 -3364 40 -3316
rect 0 -3396 4 -3364
rect 36 -3396 40 -3364
rect 0 -3444 40 -3396
rect 0 -3476 4 -3444
rect 36 -3476 40 -3444
rect 0 -3524 40 -3476
rect 0 -3556 4 -3524
rect 36 -3556 40 -3524
rect 0 -3604 40 -3556
rect 0 -3636 4 -3604
rect 36 -3636 40 -3604
rect 0 -3684 40 -3636
rect 0 -3716 4 -3684
rect 36 -3716 40 -3684
rect 0 -3720 40 -3716
rect 80 1036 120 1040
rect 80 1004 84 1036
rect 116 1004 120 1036
rect 80 956 120 1004
rect 80 924 84 956
rect 116 924 120 956
rect 80 876 120 924
rect 80 844 84 876
rect 116 844 120 876
rect 80 796 120 844
rect 80 764 84 796
rect 116 764 120 796
rect 80 716 120 764
rect 80 684 84 716
rect 116 684 120 716
rect 80 636 120 684
rect 80 604 84 636
rect 116 604 120 636
rect 80 556 120 604
rect 80 524 84 556
rect 116 524 120 556
rect 80 476 120 524
rect 80 444 84 476
rect 116 444 120 476
rect 80 396 120 444
rect 80 364 84 396
rect 116 364 120 396
rect 80 316 120 364
rect 80 284 84 316
rect 116 284 120 316
rect 80 236 120 284
rect 80 204 84 236
rect 116 204 120 236
rect 80 156 120 204
rect 80 124 84 156
rect 116 124 120 156
rect 80 76 120 124
rect 80 44 84 76
rect 116 44 120 76
rect 80 -4 120 44
rect 80 -36 84 -4
rect 116 -36 120 -4
rect 80 -84 120 -36
rect 80 -116 84 -84
rect 116 -116 120 -84
rect 80 -164 120 -116
rect 80 -196 84 -164
rect 116 -196 120 -164
rect 80 -244 120 -196
rect 80 -276 84 -244
rect 116 -276 120 -244
rect 80 -324 120 -276
rect 80 -356 84 -324
rect 116 -356 120 -324
rect 80 -404 120 -356
rect 80 -436 84 -404
rect 116 -436 120 -404
rect 80 -484 120 -436
rect 80 -516 84 -484
rect 116 -516 120 -484
rect 80 -564 120 -516
rect 80 -596 84 -564
rect 116 -596 120 -564
rect 80 -644 120 -596
rect 80 -676 84 -644
rect 116 -676 120 -644
rect 80 -724 120 -676
rect 80 -756 84 -724
rect 116 -756 120 -724
rect 80 -804 120 -756
rect 80 -836 84 -804
rect 116 -836 120 -804
rect 80 -884 120 -836
rect 80 -916 84 -884
rect 116 -916 120 -884
rect 80 -964 120 -916
rect 80 -996 84 -964
rect 116 -996 120 -964
rect 80 -1044 120 -996
rect 80 -1076 84 -1044
rect 116 -1076 120 -1044
rect 80 -1124 120 -1076
rect 80 -1156 84 -1124
rect 116 -1156 120 -1124
rect 80 -1204 120 -1156
rect 80 -1236 84 -1204
rect 116 -1236 120 -1204
rect 80 -1284 120 -1236
rect 80 -1316 84 -1284
rect 116 -1316 120 -1284
rect 80 -1364 120 -1316
rect 80 -1396 84 -1364
rect 116 -1396 120 -1364
rect 80 -1444 120 -1396
rect 80 -1476 84 -1444
rect 116 -1476 120 -1444
rect 80 -1524 120 -1476
rect 80 -1556 84 -1524
rect 116 -1556 120 -1524
rect 80 -1604 120 -1556
rect 80 -1636 84 -1604
rect 116 -1636 120 -1604
rect 80 -1684 120 -1636
rect 80 -1716 84 -1684
rect 116 -1716 120 -1684
rect 80 -1764 120 -1716
rect 80 -1796 84 -1764
rect 116 -1796 120 -1764
rect 80 -1844 120 -1796
rect 80 -1876 84 -1844
rect 116 -1876 120 -1844
rect 80 -1924 120 -1876
rect 80 -1956 84 -1924
rect 116 -1956 120 -1924
rect 80 -2004 120 -1956
rect 80 -2036 84 -2004
rect 116 -2036 120 -2004
rect 80 -2084 120 -2036
rect 80 -2116 84 -2084
rect 116 -2116 120 -2084
rect 80 -2164 120 -2116
rect 80 -2196 84 -2164
rect 116 -2196 120 -2164
rect 80 -2244 120 -2196
rect 80 -2276 84 -2244
rect 116 -2276 120 -2244
rect 80 -2324 120 -2276
rect 80 -2356 84 -2324
rect 116 -2356 120 -2324
rect 80 -2404 120 -2356
rect 80 -2436 84 -2404
rect 116 -2436 120 -2404
rect 80 -2484 120 -2436
rect 80 -2516 84 -2484
rect 116 -2516 120 -2484
rect 80 -2564 120 -2516
rect 80 -2596 84 -2564
rect 116 -2596 120 -2564
rect 80 -2644 120 -2596
rect 80 -2676 84 -2644
rect 116 -2676 120 -2644
rect 80 -2724 120 -2676
rect 80 -2756 84 -2724
rect 116 -2756 120 -2724
rect 80 -2804 120 -2756
rect 80 -2836 84 -2804
rect 116 -2836 120 -2804
rect 80 -2884 120 -2836
rect 80 -2916 84 -2884
rect 116 -2916 120 -2884
rect 80 -2964 120 -2916
rect 80 -2996 84 -2964
rect 116 -2996 120 -2964
rect 80 -3044 120 -2996
rect 80 -3076 84 -3044
rect 116 -3076 120 -3044
rect 80 -3124 120 -3076
rect 80 -3156 84 -3124
rect 116 -3156 120 -3124
rect 80 -3204 120 -3156
rect 80 -3236 84 -3204
rect 116 -3236 120 -3204
rect 80 -3284 120 -3236
rect 80 -3316 84 -3284
rect 116 -3316 120 -3284
rect 80 -3364 120 -3316
rect 80 -3396 84 -3364
rect 116 -3396 120 -3364
rect 80 -3444 120 -3396
rect 80 -3476 84 -3444
rect 116 -3476 120 -3444
rect 80 -3524 120 -3476
rect 80 -3556 84 -3524
rect 116 -3556 120 -3524
rect 80 -3604 120 -3556
rect 80 -3636 84 -3604
rect 116 -3636 120 -3604
rect 80 -3684 120 -3636
rect 80 -3716 84 -3684
rect 116 -3716 120 -3684
rect 80 -3720 120 -3716
rect 160 1036 200 1040
rect 160 1004 164 1036
rect 196 1004 200 1036
rect 160 956 200 1004
rect 160 924 164 956
rect 196 924 200 956
rect 160 876 200 924
rect 160 844 164 876
rect 196 844 200 876
rect 160 796 200 844
rect 160 764 164 796
rect 196 764 200 796
rect 160 716 200 764
rect 160 684 164 716
rect 196 684 200 716
rect 160 636 200 684
rect 160 604 164 636
rect 196 604 200 636
rect 160 556 200 604
rect 160 524 164 556
rect 196 524 200 556
rect 160 476 200 524
rect 160 444 164 476
rect 196 444 200 476
rect 160 396 200 444
rect 160 364 164 396
rect 196 364 200 396
rect 160 316 200 364
rect 160 284 164 316
rect 196 284 200 316
rect 160 236 200 284
rect 160 204 164 236
rect 196 204 200 236
rect 160 156 200 204
rect 160 124 164 156
rect 196 124 200 156
rect 160 76 200 124
rect 160 44 164 76
rect 196 44 200 76
rect 160 -4 200 44
rect 160 -36 164 -4
rect 196 -36 200 -4
rect 160 -84 200 -36
rect 160 -116 164 -84
rect 196 -116 200 -84
rect 160 -164 200 -116
rect 160 -196 164 -164
rect 196 -196 200 -164
rect 160 -244 200 -196
rect 160 -276 164 -244
rect 196 -276 200 -244
rect 160 -324 200 -276
rect 160 -356 164 -324
rect 196 -356 200 -324
rect 160 -404 200 -356
rect 160 -436 164 -404
rect 196 -436 200 -404
rect 160 -484 200 -436
rect 160 -516 164 -484
rect 196 -516 200 -484
rect 160 -564 200 -516
rect 160 -596 164 -564
rect 196 -596 200 -564
rect 160 -644 200 -596
rect 160 -676 164 -644
rect 196 -676 200 -644
rect 160 -724 200 -676
rect 160 -756 164 -724
rect 196 -756 200 -724
rect 160 -804 200 -756
rect 160 -836 164 -804
rect 196 -836 200 -804
rect 160 -884 200 -836
rect 160 -916 164 -884
rect 196 -916 200 -884
rect 160 -964 200 -916
rect 160 -996 164 -964
rect 196 -996 200 -964
rect 160 -1044 200 -996
rect 160 -1076 164 -1044
rect 196 -1076 200 -1044
rect 160 -1124 200 -1076
rect 160 -1156 164 -1124
rect 196 -1156 200 -1124
rect 160 -1204 200 -1156
rect 160 -1236 164 -1204
rect 196 -1236 200 -1204
rect 160 -1284 200 -1236
rect 160 -1316 164 -1284
rect 196 -1316 200 -1284
rect 160 -1364 200 -1316
rect 160 -1396 164 -1364
rect 196 -1396 200 -1364
rect 160 -1444 200 -1396
rect 160 -1476 164 -1444
rect 196 -1476 200 -1444
rect 160 -1524 200 -1476
rect 160 -1556 164 -1524
rect 196 -1556 200 -1524
rect 160 -1604 200 -1556
rect 160 -1636 164 -1604
rect 196 -1636 200 -1604
rect 160 -1684 200 -1636
rect 160 -1716 164 -1684
rect 196 -1716 200 -1684
rect 160 -1764 200 -1716
rect 160 -1796 164 -1764
rect 196 -1796 200 -1764
rect 160 -1844 200 -1796
rect 160 -1876 164 -1844
rect 196 -1876 200 -1844
rect 160 -1924 200 -1876
rect 160 -1956 164 -1924
rect 196 -1956 200 -1924
rect 160 -2004 200 -1956
rect 160 -2036 164 -2004
rect 196 -2036 200 -2004
rect 160 -2084 200 -2036
rect 160 -2116 164 -2084
rect 196 -2116 200 -2084
rect 160 -2164 200 -2116
rect 160 -2196 164 -2164
rect 196 -2196 200 -2164
rect 160 -2244 200 -2196
rect 160 -2276 164 -2244
rect 196 -2276 200 -2244
rect 160 -2324 200 -2276
rect 160 -2356 164 -2324
rect 196 -2356 200 -2324
rect 160 -2404 200 -2356
rect 160 -2436 164 -2404
rect 196 -2436 200 -2404
rect 160 -2484 200 -2436
rect 160 -2516 164 -2484
rect 196 -2516 200 -2484
rect 160 -2564 200 -2516
rect 160 -2596 164 -2564
rect 196 -2596 200 -2564
rect 160 -2644 200 -2596
rect 160 -2676 164 -2644
rect 196 -2676 200 -2644
rect 160 -2724 200 -2676
rect 160 -2756 164 -2724
rect 196 -2756 200 -2724
rect 160 -2804 200 -2756
rect 160 -2836 164 -2804
rect 196 -2836 200 -2804
rect 160 -2884 200 -2836
rect 160 -2916 164 -2884
rect 196 -2916 200 -2884
rect 160 -2964 200 -2916
rect 160 -2996 164 -2964
rect 196 -2996 200 -2964
rect 160 -3044 200 -2996
rect 160 -3076 164 -3044
rect 196 -3076 200 -3044
rect 160 -3124 200 -3076
rect 160 -3156 164 -3124
rect 196 -3156 200 -3124
rect 160 -3204 200 -3156
rect 160 -3236 164 -3204
rect 196 -3236 200 -3204
rect 160 -3284 200 -3236
rect 160 -3316 164 -3284
rect 196 -3316 200 -3284
rect 160 -3364 200 -3316
rect 160 -3396 164 -3364
rect 196 -3396 200 -3364
rect 160 -3444 200 -3396
rect 160 -3476 164 -3444
rect 196 -3476 200 -3444
rect 160 -3524 200 -3476
rect 160 -3556 164 -3524
rect 196 -3556 200 -3524
rect 160 -3604 200 -3556
rect 160 -3636 164 -3604
rect 196 -3636 200 -3604
rect 160 -3684 200 -3636
rect 160 -3716 164 -3684
rect 196 -3716 200 -3684
rect 160 -3720 200 -3716
rect 240 1036 280 1040
rect 240 1004 244 1036
rect 276 1004 280 1036
rect 240 956 280 1004
rect 240 924 244 956
rect 276 924 280 956
rect 240 876 280 924
rect 240 844 244 876
rect 276 844 280 876
rect 240 796 280 844
rect 240 764 244 796
rect 276 764 280 796
rect 240 716 280 764
rect 240 684 244 716
rect 276 684 280 716
rect 240 636 280 684
rect 240 604 244 636
rect 276 604 280 636
rect 240 556 280 604
rect 240 524 244 556
rect 276 524 280 556
rect 240 476 280 524
rect 240 444 244 476
rect 276 444 280 476
rect 240 396 280 444
rect 240 364 244 396
rect 276 364 280 396
rect 240 316 280 364
rect 240 284 244 316
rect 276 284 280 316
rect 240 236 280 284
rect 240 204 244 236
rect 276 204 280 236
rect 240 156 280 204
rect 240 124 244 156
rect 276 124 280 156
rect 240 76 280 124
rect 240 44 244 76
rect 276 44 280 76
rect 240 -4 280 44
rect 240 -36 244 -4
rect 276 -36 280 -4
rect 240 -84 280 -36
rect 240 -116 244 -84
rect 276 -116 280 -84
rect 240 -164 280 -116
rect 240 -196 244 -164
rect 276 -196 280 -164
rect 240 -244 280 -196
rect 240 -276 244 -244
rect 276 -276 280 -244
rect 240 -324 280 -276
rect 240 -356 244 -324
rect 276 -356 280 -324
rect 240 -404 280 -356
rect 240 -436 244 -404
rect 276 -436 280 -404
rect 240 -484 280 -436
rect 240 -516 244 -484
rect 276 -516 280 -484
rect 240 -564 280 -516
rect 240 -596 244 -564
rect 276 -596 280 -564
rect 240 -644 280 -596
rect 240 -676 244 -644
rect 276 -676 280 -644
rect 240 -724 280 -676
rect 240 -756 244 -724
rect 276 -756 280 -724
rect 240 -804 280 -756
rect 240 -836 244 -804
rect 276 -836 280 -804
rect 240 -884 280 -836
rect 240 -916 244 -884
rect 276 -916 280 -884
rect 240 -964 280 -916
rect 240 -996 244 -964
rect 276 -996 280 -964
rect 240 -1044 280 -996
rect 240 -1076 244 -1044
rect 276 -1076 280 -1044
rect 240 -1124 280 -1076
rect 240 -1156 244 -1124
rect 276 -1156 280 -1124
rect 240 -1204 280 -1156
rect 240 -1236 244 -1204
rect 276 -1236 280 -1204
rect 240 -1284 280 -1236
rect 240 -1316 244 -1284
rect 276 -1316 280 -1284
rect 240 -1364 280 -1316
rect 240 -1396 244 -1364
rect 276 -1396 280 -1364
rect 240 -1444 280 -1396
rect 240 -1476 244 -1444
rect 276 -1476 280 -1444
rect 240 -1524 280 -1476
rect 240 -1556 244 -1524
rect 276 -1556 280 -1524
rect 240 -1604 280 -1556
rect 240 -1636 244 -1604
rect 276 -1636 280 -1604
rect 240 -1684 280 -1636
rect 240 -1716 244 -1684
rect 276 -1716 280 -1684
rect 240 -1764 280 -1716
rect 240 -1796 244 -1764
rect 276 -1796 280 -1764
rect 240 -1844 280 -1796
rect 240 -1876 244 -1844
rect 276 -1876 280 -1844
rect 240 -1924 280 -1876
rect 240 -1956 244 -1924
rect 276 -1956 280 -1924
rect 240 -2004 280 -1956
rect 240 -2036 244 -2004
rect 276 -2036 280 -2004
rect 240 -2084 280 -2036
rect 240 -2116 244 -2084
rect 276 -2116 280 -2084
rect 240 -2164 280 -2116
rect 240 -2196 244 -2164
rect 276 -2196 280 -2164
rect 240 -2244 280 -2196
rect 240 -2276 244 -2244
rect 276 -2276 280 -2244
rect 240 -2324 280 -2276
rect 240 -2356 244 -2324
rect 276 -2356 280 -2324
rect 240 -2404 280 -2356
rect 240 -2436 244 -2404
rect 276 -2436 280 -2404
rect 240 -2484 280 -2436
rect 240 -2516 244 -2484
rect 276 -2516 280 -2484
rect 240 -2564 280 -2516
rect 240 -2596 244 -2564
rect 276 -2596 280 -2564
rect 240 -2644 280 -2596
rect 240 -2676 244 -2644
rect 276 -2676 280 -2644
rect 240 -2724 280 -2676
rect 240 -2756 244 -2724
rect 276 -2756 280 -2724
rect 240 -2804 280 -2756
rect 240 -2836 244 -2804
rect 276 -2836 280 -2804
rect 240 -2884 280 -2836
rect 240 -2916 244 -2884
rect 276 -2916 280 -2884
rect 240 -2964 280 -2916
rect 240 -2996 244 -2964
rect 276 -2996 280 -2964
rect 240 -3044 280 -2996
rect 240 -3076 244 -3044
rect 276 -3076 280 -3044
rect 240 -3124 280 -3076
rect 240 -3156 244 -3124
rect 276 -3156 280 -3124
rect 240 -3204 280 -3156
rect 240 -3236 244 -3204
rect 276 -3236 280 -3204
rect 240 -3284 280 -3236
rect 240 -3316 244 -3284
rect 276 -3316 280 -3284
rect 240 -3364 280 -3316
rect 240 -3396 244 -3364
rect 276 -3396 280 -3364
rect 240 -3444 280 -3396
rect 240 -3476 244 -3444
rect 276 -3476 280 -3444
rect 240 -3524 280 -3476
rect 240 -3556 244 -3524
rect 276 -3556 280 -3524
rect 240 -3604 280 -3556
rect 240 -3636 244 -3604
rect 276 -3636 280 -3604
rect 240 -3684 280 -3636
rect 240 -3716 244 -3684
rect 276 -3716 280 -3684
rect 240 -3720 280 -3716
rect 320 1036 360 1040
rect 320 1004 324 1036
rect 356 1004 360 1036
rect 320 956 360 1004
rect 320 924 324 956
rect 356 924 360 956
rect 320 876 360 924
rect 320 844 324 876
rect 356 844 360 876
rect 320 796 360 844
rect 320 764 324 796
rect 356 764 360 796
rect 320 716 360 764
rect 320 684 324 716
rect 356 684 360 716
rect 320 636 360 684
rect 320 604 324 636
rect 356 604 360 636
rect 320 556 360 604
rect 320 524 324 556
rect 356 524 360 556
rect 320 476 360 524
rect 320 444 324 476
rect 356 444 360 476
rect 320 396 360 444
rect 320 364 324 396
rect 356 364 360 396
rect 320 316 360 364
rect 320 284 324 316
rect 356 284 360 316
rect 320 236 360 284
rect 320 204 324 236
rect 356 204 360 236
rect 320 156 360 204
rect 320 124 324 156
rect 356 124 360 156
rect 320 76 360 124
rect 320 44 324 76
rect 356 44 360 76
rect 320 -4 360 44
rect 320 -36 324 -4
rect 356 -36 360 -4
rect 320 -84 360 -36
rect 320 -116 324 -84
rect 356 -116 360 -84
rect 320 -164 360 -116
rect 320 -196 324 -164
rect 356 -196 360 -164
rect 320 -244 360 -196
rect 320 -276 324 -244
rect 356 -276 360 -244
rect 320 -324 360 -276
rect 320 -356 324 -324
rect 356 -356 360 -324
rect 320 -404 360 -356
rect 320 -436 324 -404
rect 356 -436 360 -404
rect 320 -484 360 -436
rect 320 -516 324 -484
rect 356 -516 360 -484
rect 320 -564 360 -516
rect 320 -596 324 -564
rect 356 -596 360 -564
rect 320 -644 360 -596
rect 320 -676 324 -644
rect 356 -676 360 -644
rect 320 -724 360 -676
rect 320 -756 324 -724
rect 356 -756 360 -724
rect 320 -804 360 -756
rect 320 -836 324 -804
rect 356 -836 360 -804
rect 320 -884 360 -836
rect 320 -916 324 -884
rect 356 -916 360 -884
rect 320 -964 360 -916
rect 320 -996 324 -964
rect 356 -996 360 -964
rect 320 -1044 360 -996
rect 320 -1076 324 -1044
rect 356 -1076 360 -1044
rect 320 -1124 360 -1076
rect 320 -1156 324 -1124
rect 356 -1156 360 -1124
rect 320 -1204 360 -1156
rect 320 -1236 324 -1204
rect 356 -1236 360 -1204
rect 320 -1284 360 -1236
rect 320 -1316 324 -1284
rect 356 -1316 360 -1284
rect 320 -1364 360 -1316
rect 320 -1396 324 -1364
rect 356 -1396 360 -1364
rect 320 -1444 360 -1396
rect 320 -1476 324 -1444
rect 356 -1476 360 -1444
rect 320 -1524 360 -1476
rect 320 -1556 324 -1524
rect 356 -1556 360 -1524
rect 320 -1604 360 -1556
rect 320 -1636 324 -1604
rect 356 -1636 360 -1604
rect 320 -1684 360 -1636
rect 320 -1716 324 -1684
rect 356 -1716 360 -1684
rect 320 -1764 360 -1716
rect 320 -1796 324 -1764
rect 356 -1796 360 -1764
rect 320 -1844 360 -1796
rect 320 -1876 324 -1844
rect 356 -1876 360 -1844
rect 320 -1924 360 -1876
rect 320 -1956 324 -1924
rect 356 -1956 360 -1924
rect 320 -2004 360 -1956
rect 320 -2036 324 -2004
rect 356 -2036 360 -2004
rect 320 -2084 360 -2036
rect 320 -2116 324 -2084
rect 356 -2116 360 -2084
rect 320 -2164 360 -2116
rect 320 -2196 324 -2164
rect 356 -2196 360 -2164
rect 320 -2244 360 -2196
rect 320 -2276 324 -2244
rect 356 -2276 360 -2244
rect 320 -2324 360 -2276
rect 320 -2356 324 -2324
rect 356 -2356 360 -2324
rect 320 -2404 360 -2356
rect 320 -2436 324 -2404
rect 356 -2436 360 -2404
rect 320 -2484 360 -2436
rect 320 -2516 324 -2484
rect 356 -2516 360 -2484
rect 320 -2564 360 -2516
rect 320 -2596 324 -2564
rect 356 -2596 360 -2564
rect 320 -2644 360 -2596
rect 320 -2676 324 -2644
rect 356 -2676 360 -2644
rect 320 -2724 360 -2676
rect 320 -2756 324 -2724
rect 356 -2756 360 -2724
rect 320 -2804 360 -2756
rect 320 -2836 324 -2804
rect 356 -2836 360 -2804
rect 320 -2884 360 -2836
rect 320 -2916 324 -2884
rect 356 -2916 360 -2884
rect 320 -2964 360 -2916
rect 320 -2996 324 -2964
rect 356 -2996 360 -2964
rect 320 -3044 360 -2996
rect 320 -3076 324 -3044
rect 356 -3076 360 -3044
rect 320 -3124 360 -3076
rect 320 -3156 324 -3124
rect 356 -3156 360 -3124
rect 320 -3204 360 -3156
rect 320 -3236 324 -3204
rect 356 -3236 360 -3204
rect 320 -3284 360 -3236
rect 320 -3316 324 -3284
rect 356 -3316 360 -3284
rect 320 -3364 360 -3316
rect 320 -3396 324 -3364
rect 356 -3396 360 -3364
rect 320 -3444 360 -3396
rect 320 -3476 324 -3444
rect 356 -3476 360 -3444
rect 320 -3524 360 -3476
rect 320 -3556 324 -3524
rect 356 -3556 360 -3524
rect 320 -3604 360 -3556
rect 320 -3636 324 -3604
rect 356 -3636 360 -3604
rect 320 -3684 360 -3636
rect 320 -3716 324 -3684
rect 356 -3716 360 -3684
rect 320 -3720 360 -3716
rect 400 1036 440 1040
rect 400 1004 404 1036
rect 436 1004 440 1036
rect 400 956 440 1004
rect 400 924 404 956
rect 436 924 440 956
rect 400 876 440 924
rect 400 844 404 876
rect 436 844 440 876
rect 400 796 440 844
rect 400 764 404 796
rect 436 764 440 796
rect 400 716 440 764
rect 400 684 404 716
rect 436 684 440 716
rect 400 636 440 684
rect 400 604 404 636
rect 436 604 440 636
rect 400 556 440 604
rect 400 524 404 556
rect 436 524 440 556
rect 400 476 440 524
rect 400 444 404 476
rect 436 444 440 476
rect 400 396 440 444
rect 400 364 404 396
rect 436 364 440 396
rect 400 316 440 364
rect 400 284 404 316
rect 436 284 440 316
rect 400 236 440 284
rect 400 204 404 236
rect 436 204 440 236
rect 400 156 440 204
rect 400 124 404 156
rect 436 124 440 156
rect 400 76 440 124
rect 400 44 404 76
rect 436 44 440 76
rect 400 -4 440 44
rect 400 -36 404 -4
rect 436 -36 440 -4
rect 400 -84 440 -36
rect 400 -116 404 -84
rect 436 -116 440 -84
rect 400 -164 440 -116
rect 400 -196 404 -164
rect 436 -196 440 -164
rect 400 -244 440 -196
rect 400 -276 404 -244
rect 436 -276 440 -244
rect 400 -324 440 -276
rect 400 -356 404 -324
rect 436 -356 440 -324
rect 400 -404 440 -356
rect 400 -436 404 -404
rect 436 -436 440 -404
rect 400 -484 440 -436
rect 400 -516 404 -484
rect 436 -516 440 -484
rect 400 -564 440 -516
rect 400 -596 404 -564
rect 436 -596 440 -564
rect 400 -644 440 -596
rect 400 -676 404 -644
rect 436 -676 440 -644
rect 400 -724 440 -676
rect 400 -756 404 -724
rect 436 -756 440 -724
rect 400 -804 440 -756
rect 400 -836 404 -804
rect 436 -836 440 -804
rect 400 -884 440 -836
rect 400 -916 404 -884
rect 436 -916 440 -884
rect 400 -964 440 -916
rect 400 -996 404 -964
rect 436 -996 440 -964
rect 400 -1044 440 -996
rect 400 -1076 404 -1044
rect 436 -1076 440 -1044
rect 400 -1124 440 -1076
rect 400 -1156 404 -1124
rect 436 -1156 440 -1124
rect 400 -1204 440 -1156
rect 400 -1236 404 -1204
rect 436 -1236 440 -1204
rect 400 -1284 440 -1236
rect 400 -1316 404 -1284
rect 436 -1316 440 -1284
rect 400 -1364 440 -1316
rect 400 -1396 404 -1364
rect 436 -1396 440 -1364
rect 400 -1444 440 -1396
rect 400 -1476 404 -1444
rect 436 -1476 440 -1444
rect 400 -1524 440 -1476
rect 400 -1556 404 -1524
rect 436 -1556 440 -1524
rect 400 -1604 440 -1556
rect 400 -1636 404 -1604
rect 436 -1636 440 -1604
rect 400 -1684 440 -1636
rect 400 -1716 404 -1684
rect 436 -1716 440 -1684
rect 400 -1764 440 -1716
rect 400 -1796 404 -1764
rect 436 -1796 440 -1764
rect 400 -1844 440 -1796
rect 400 -1876 404 -1844
rect 436 -1876 440 -1844
rect 400 -1924 440 -1876
rect 400 -1956 404 -1924
rect 436 -1956 440 -1924
rect 400 -2004 440 -1956
rect 400 -2036 404 -2004
rect 436 -2036 440 -2004
rect 400 -2084 440 -2036
rect 400 -2116 404 -2084
rect 436 -2116 440 -2084
rect 400 -2164 440 -2116
rect 400 -2196 404 -2164
rect 436 -2196 440 -2164
rect 400 -2244 440 -2196
rect 400 -2276 404 -2244
rect 436 -2276 440 -2244
rect 400 -2324 440 -2276
rect 400 -2356 404 -2324
rect 436 -2356 440 -2324
rect 400 -2404 440 -2356
rect 400 -2436 404 -2404
rect 436 -2436 440 -2404
rect 400 -2484 440 -2436
rect 400 -2516 404 -2484
rect 436 -2516 440 -2484
rect 400 -2564 440 -2516
rect 400 -2596 404 -2564
rect 436 -2596 440 -2564
rect 400 -2644 440 -2596
rect 400 -2676 404 -2644
rect 436 -2676 440 -2644
rect 400 -2724 440 -2676
rect 400 -2756 404 -2724
rect 436 -2756 440 -2724
rect 400 -2804 440 -2756
rect 400 -2836 404 -2804
rect 436 -2836 440 -2804
rect 400 -2884 440 -2836
rect 400 -2916 404 -2884
rect 436 -2916 440 -2884
rect 400 -2964 440 -2916
rect 400 -2996 404 -2964
rect 436 -2996 440 -2964
rect 400 -3044 440 -2996
rect 400 -3076 404 -3044
rect 436 -3076 440 -3044
rect 400 -3124 440 -3076
rect 400 -3156 404 -3124
rect 436 -3156 440 -3124
rect 400 -3204 440 -3156
rect 400 -3236 404 -3204
rect 436 -3236 440 -3204
rect 400 -3284 440 -3236
rect 400 -3316 404 -3284
rect 436 -3316 440 -3284
rect 400 -3364 440 -3316
rect 400 -3396 404 -3364
rect 436 -3396 440 -3364
rect 400 -3444 440 -3396
rect 400 -3476 404 -3444
rect 436 -3476 440 -3444
rect 400 -3524 440 -3476
rect 400 -3556 404 -3524
rect 436 -3556 440 -3524
rect 400 -3604 440 -3556
rect 400 -3636 404 -3604
rect 436 -3636 440 -3604
rect 400 -3684 440 -3636
rect 400 -3716 404 -3684
rect 436 -3716 440 -3684
rect 400 -3720 440 -3716
rect 480 1036 520 1040
rect 480 1004 484 1036
rect 516 1004 520 1036
rect 480 956 520 1004
rect 480 924 484 956
rect 516 924 520 956
rect 480 876 520 924
rect 480 844 484 876
rect 516 844 520 876
rect 480 796 520 844
rect 480 764 484 796
rect 516 764 520 796
rect 480 716 520 764
rect 480 684 484 716
rect 516 684 520 716
rect 480 636 520 684
rect 480 604 484 636
rect 516 604 520 636
rect 480 556 520 604
rect 480 524 484 556
rect 516 524 520 556
rect 480 476 520 524
rect 480 444 484 476
rect 516 444 520 476
rect 480 396 520 444
rect 480 364 484 396
rect 516 364 520 396
rect 480 316 520 364
rect 480 284 484 316
rect 516 284 520 316
rect 480 236 520 284
rect 480 204 484 236
rect 516 204 520 236
rect 480 156 520 204
rect 480 124 484 156
rect 516 124 520 156
rect 480 76 520 124
rect 480 44 484 76
rect 516 44 520 76
rect 480 -4 520 44
rect 480 -36 484 -4
rect 516 -36 520 -4
rect 480 -84 520 -36
rect 480 -116 484 -84
rect 516 -116 520 -84
rect 480 -164 520 -116
rect 480 -196 484 -164
rect 516 -196 520 -164
rect 480 -244 520 -196
rect 480 -276 484 -244
rect 516 -276 520 -244
rect 480 -324 520 -276
rect 480 -356 484 -324
rect 516 -356 520 -324
rect 480 -404 520 -356
rect 480 -436 484 -404
rect 516 -436 520 -404
rect 480 -484 520 -436
rect 480 -516 484 -484
rect 516 -516 520 -484
rect 480 -564 520 -516
rect 480 -596 484 -564
rect 516 -596 520 -564
rect 480 -644 520 -596
rect 480 -676 484 -644
rect 516 -676 520 -644
rect 480 -724 520 -676
rect 480 -756 484 -724
rect 516 -756 520 -724
rect 480 -804 520 -756
rect 480 -836 484 -804
rect 516 -836 520 -804
rect 480 -884 520 -836
rect 480 -916 484 -884
rect 516 -916 520 -884
rect 480 -964 520 -916
rect 480 -996 484 -964
rect 516 -996 520 -964
rect 480 -1044 520 -996
rect 480 -1076 484 -1044
rect 516 -1076 520 -1044
rect 480 -1124 520 -1076
rect 480 -1156 484 -1124
rect 516 -1156 520 -1124
rect 480 -1204 520 -1156
rect 480 -1236 484 -1204
rect 516 -1236 520 -1204
rect 480 -1284 520 -1236
rect 480 -1316 484 -1284
rect 516 -1316 520 -1284
rect 480 -1364 520 -1316
rect 480 -1396 484 -1364
rect 516 -1396 520 -1364
rect 480 -1444 520 -1396
rect 480 -1476 484 -1444
rect 516 -1476 520 -1444
rect 480 -1524 520 -1476
rect 480 -1556 484 -1524
rect 516 -1556 520 -1524
rect 480 -1604 520 -1556
rect 480 -1636 484 -1604
rect 516 -1636 520 -1604
rect 480 -1684 520 -1636
rect 480 -1716 484 -1684
rect 516 -1716 520 -1684
rect 480 -1764 520 -1716
rect 480 -1796 484 -1764
rect 516 -1796 520 -1764
rect 480 -1844 520 -1796
rect 480 -1876 484 -1844
rect 516 -1876 520 -1844
rect 480 -1924 520 -1876
rect 480 -1956 484 -1924
rect 516 -1956 520 -1924
rect 480 -2004 520 -1956
rect 480 -2036 484 -2004
rect 516 -2036 520 -2004
rect 480 -2084 520 -2036
rect 480 -2116 484 -2084
rect 516 -2116 520 -2084
rect 480 -2164 520 -2116
rect 480 -2196 484 -2164
rect 516 -2196 520 -2164
rect 480 -2244 520 -2196
rect 480 -2276 484 -2244
rect 516 -2276 520 -2244
rect 480 -2324 520 -2276
rect 480 -2356 484 -2324
rect 516 -2356 520 -2324
rect 480 -2404 520 -2356
rect 480 -2436 484 -2404
rect 516 -2436 520 -2404
rect 480 -2484 520 -2436
rect 480 -2516 484 -2484
rect 516 -2516 520 -2484
rect 480 -2564 520 -2516
rect 480 -2596 484 -2564
rect 516 -2596 520 -2564
rect 480 -2644 520 -2596
rect 480 -2676 484 -2644
rect 516 -2676 520 -2644
rect 480 -2724 520 -2676
rect 480 -2756 484 -2724
rect 516 -2756 520 -2724
rect 480 -2804 520 -2756
rect 480 -2836 484 -2804
rect 516 -2836 520 -2804
rect 480 -2884 520 -2836
rect 480 -2916 484 -2884
rect 516 -2916 520 -2884
rect 480 -2964 520 -2916
rect 480 -2996 484 -2964
rect 516 -2996 520 -2964
rect 480 -3044 520 -2996
rect 480 -3076 484 -3044
rect 516 -3076 520 -3044
rect 480 -3124 520 -3076
rect 480 -3156 484 -3124
rect 516 -3156 520 -3124
rect 480 -3204 520 -3156
rect 480 -3236 484 -3204
rect 516 -3236 520 -3204
rect 480 -3284 520 -3236
rect 480 -3316 484 -3284
rect 516 -3316 520 -3284
rect 480 -3364 520 -3316
rect 480 -3396 484 -3364
rect 516 -3396 520 -3364
rect 480 -3444 520 -3396
rect 480 -3476 484 -3444
rect 516 -3476 520 -3444
rect 480 -3524 520 -3476
rect 480 -3556 484 -3524
rect 516 -3556 520 -3524
rect 480 -3604 520 -3556
rect 480 -3636 484 -3604
rect 516 -3636 520 -3604
rect 480 -3684 520 -3636
rect 480 -3716 484 -3684
rect 516 -3716 520 -3684
rect 480 -3720 520 -3716
rect 560 1036 600 1040
rect 560 1004 564 1036
rect 596 1004 600 1036
rect 560 956 600 1004
rect 560 924 564 956
rect 596 924 600 956
rect 560 876 600 924
rect 560 844 564 876
rect 596 844 600 876
rect 560 796 600 844
rect 560 764 564 796
rect 596 764 600 796
rect 560 716 600 764
rect 560 684 564 716
rect 596 684 600 716
rect 560 636 600 684
rect 560 604 564 636
rect 596 604 600 636
rect 560 556 600 604
rect 560 524 564 556
rect 596 524 600 556
rect 560 476 600 524
rect 560 444 564 476
rect 596 444 600 476
rect 560 396 600 444
rect 560 364 564 396
rect 596 364 600 396
rect 560 316 600 364
rect 560 284 564 316
rect 596 284 600 316
rect 560 236 600 284
rect 560 204 564 236
rect 596 204 600 236
rect 560 156 600 204
rect 560 124 564 156
rect 596 124 600 156
rect 560 76 600 124
rect 560 44 564 76
rect 596 44 600 76
rect 560 -4 600 44
rect 560 -36 564 -4
rect 596 -36 600 -4
rect 560 -84 600 -36
rect 560 -116 564 -84
rect 596 -116 600 -84
rect 560 -164 600 -116
rect 560 -196 564 -164
rect 596 -196 600 -164
rect 560 -244 600 -196
rect 560 -276 564 -244
rect 596 -276 600 -244
rect 560 -324 600 -276
rect 560 -356 564 -324
rect 596 -356 600 -324
rect 560 -404 600 -356
rect 560 -436 564 -404
rect 596 -436 600 -404
rect 560 -484 600 -436
rect 560 -516 564 -484
rect 596 -516 600 -484
rect 560 -564 600 -516
rect 560 -596 564 -564
rect 596 -596 600 -564
rect 560 -644 600 -596
rect 560 -676 564 -644
rect 596 -676 600 -644
rect 560 -724 600 -676
rect 560 -756 564 -724
rect 596 -756 600 -724
rect 560 -804 600 -756
rect 560 -836 564 -804
rect 596 -836 600 -804
rect 560 -884 600 -836
rect 560 -916 564 -884
rect 596 -916 600 -884
rect 560 -964 600 -916
rect 560 -996 564 -964
rect 596 -996 600 -964
rect 560 -1044 600 -996
rect 560 -1076 564 -1044
rect 596 -1076 600 -1044
rect 560 -1124 600 -1076
rect 560 -1156 564 -1124
rect 596 -1156 600 -1124
rect 560 -1204 600 -1156
rect 560 -1236 564 -1204
rect 596 -1236 600 -1204
rect 560 -1284 600 -1236
rect 560 -1316 564 -1284
rect 596 -1316 600 -1284
rect 560 -1364 600 -1316
rect 560 -1396 564 -1364
rect 596 -1396 600 -1364
rect 560 -1444 600 -1396
rect 560 -1476 564 -1444
rect 596 -1476 600 -1444
rect 560 -1524 600 -1476
rect 560 -1556 564 -1524
rect 596 -1556 600 -1524
rect 560 -1604 600 -1556
rect 560 -1636 564 -1604
rect 596 -1636 600 -1604
rect 560 -1684 600 -1636
rect 560 -1716 564 -1684
rect 596 -1716 600 -1684
rect 560 -1764 600 -1716
rect 560 -1796 564 -1764
rect 596 -1796 600 -1764
rect 560 -1844 600 -1796
rect 560 -1876 564 -1844
rect 596 -1876 600 -1844
rect 560 -1924 600 -1876
rect 560 -1956 564 -1924
rect 596 -1956 600 -1924
rect 560 -2004 600 -1956
rect 560 -2036 564 -2004
rect 596 -2036 600 -2004
rect 560 -2084 600 -2036
rect 560 -2116 564 -2084
rect 596 -2116 600 -2084
rect 560 -2164 600 -2116
rect 560 -2196 564 -2164
rect 596 -2196 600 -2164
rect 560 -2244 600 -2196
rect 560 -2276 564 -2244
rect 596 -2276 600 -2244
rect 560 -2324 600 -2276
rect 560 -2356 564 -2324
rect 596 -2356 600 -2324
rect 560 -2404 600 -2356
rect 560 -2436 564 -2404
rect 596 -2436 600 -2404
rect 560 -2484 600 -2436
rect 560 -2516 564 -2484
rect 596 -2516 600 -2484
rect 560 -2564 600 -2516
rect 560 -2596 564 -2564
rect 596 -2596 600 -2564
rect 560 -2644 600 -2596
rect 560 -2676 564 -2644
rect 596 -2676 600 -2644
rect 560 -2724 600 -2676
rect 560 -2756 564 -2724
rect 596 -2756 600 -2724
rect 560 -2804 600 -2756
rect 560 -2836 564 -2804
rect 596 -2836 600 -2804
rect 560 -2884 600 -2836
rect 560 -2916 564 -2884
rect 596 -2916 600 -2884
rect 560 -2964 600 -2916
rect 560 -2996 564 -2964
rect 596 -2996 600 -2964
rect 560 -3044 600 -2996
rect 560 -3076 564 -3044
rect 596 -3076 600 -3044
rect 560 -3124 600 -3076
rect 560 -3156 564 -3124
rect 596 -3156 600 -3124
rect 560 -3204 600 -3156
rect 560 -3236 564 -3204
rect 596 -3236 600 -3204
rect 560 -3284 600 -3236
rect 560 -3316 564 -3284
rect 596 -3316 600 -3284
rect 560 -3364 600 -3316
rect 560 -3396 564 -3364
rect 596 -3396 600 -3364
rect 560 -3444 600 -3396
rect 560 -3476 564 -3444
rect 596 -3476 600 -3444
rect 560 -3524 600 -3476
rect 560 -3556 564 -3524
rect 596 -3556 600 -3524
rect 560 -3604 600 -3556
rect 560 -3636 564 -3604
rect 596 -3636 600 -3604
rect 560 -3684 600 -3636
rect 560 -3716 564 -3684
rect 596 -3716 600 -3684
rect 560 -3720 600 -3716
rect 640 1036 680 1040
rect 640 1004 644 1036
rect 676 1004 680 1036
rect 640 956 680 1004
rect 640 924 644 956
rect 676 924 680 956
rect 640 876 680 924
rect 640 844 644 876
rect 676 844 680 876
rect 640 796 680 844
rect 640 764 644 796
rect 676 764 680 796
rect 640 716 680 764
rect 640 684 644 716
rect 676 684 680 716
rect 640 636 680 684
rect 640 604 644 636
rect 676 604 680 636
rect 640 556 680 604
rect 640 524 644 556
rect 676 524 680 556
rect 640 476 680 524
rect 640 444 644 476
rect 676 444 680 476
rect 640 396 680 444
rect 640 364 644 396
rect 676 364 680 396
rect 640 316 680 364
rect 640 284 644 316
rect 676 284 680 316
rect 640 236 680 284
rect 640 204 644 236
rect 676 204 680 236
rect 640 156 680 204
rect 640 124 644 156
rect 676 124 680 156
rect 640 76 680 124
rect 640 44 644 76
rect 676 44 680 76
rect 640 -4 680 44
rect 640 -36 644 -4
rect 676 -36 680 -4
rect 640 -84 680 -36
rect 640 -116 644 -84
rect 676 -116 680 -84
rect 640 -164 680 -116
rect 640 -196 644 -164
rect 676 -196 680 -164
rect 640 -244 680 -196
rect 640 -276 644 -244
rect 676 -276 680 -244
rect 640 -324 680 -276
rect 640 -356 644 -324
rect 676 -356 680 -324
rect 640 -404 680 -356
rect 640 -436 644 -404
rect 676 -436 680 -404
rect 640 -484 680 -436
rect 640 -516 644 -484
rect 676 -516 680 -484
rect 640 -564 680 -516
rect 640 -596 644 -564
rect 676 -596 680 -564
rect 640 -644 680 -596
rect 640 -676 644 -644
rect 676 -676 680 -644
rect 640 -724 680 -676
rect 640 -756 644 -724
rect 676 -756 680 -724
rect 640 -804 680 -756
rect 640 -836 644 -804
rect 676 -836 680 -804
rect 640 -884 680 -836
rect 640 -916 644 -884
rect 676 -916 680 -884
rect 640 -964 680 -916
rect 640 -996 644 -964
rect 676 -996 680 -964
rect 640 -1044 680 -996
rect 640 -1076 644 -1044
rect 676 -1076 680 -1044
rect 640 -1124 680 -1076
rect 640 -1156 644 -1124
rect 676 -1156 680 -1124
rect 640 -1204 680 -1156
rect 640 -1236 644 -1204
rect 676 -1236 680 -1204
rect 640 -1284 680 -1236
rect 640 -1316 644 -1284
rect 676 -1316 680 -1284
rect 640 -1364 680 -1316
rect 640 -1396 644 -1364
rect 676 -1396 680 -1364
rect 640 -1444 680 -1396
rect 640 -1476 644 -1444
rect 676 -1476 680 -1444
rect 640 -1524 680 -1476
rect 640 -1556 644 -1524
rect 676 -1556 680 -1524
rect 640 -1604 680 -1556
rect 640 -1636 644 -1604
rect 676 -1636 680 -1604
rect 640 -1684 680 -1636
rect 640 -1716 644 -1684
rect 676 -1716 680 -1684
rect 640 -1764 680 -1716
rect 640 -1796 644 -1764
rect 676 -1796 680 -1764
rect 640 -1844 680 -1796
rect 640 -1876 644 -1844
rect 676 -1876 680 -1844
rect 640 -1924 680 -1876
rect 640 -1956 644 -1924
rect 676 -1956 680 -1924
rect 640 -2004 680 -1956
rect 640 -2036 644 -2004
rect 676 -2036 680 -2004
rect 640 -2084 680 -2036
rect 640 -2116 644 -2084
rect 676 -2116 680 -2084
rect 640 -2164 680 -2116
rect 640 -2196 644 -2164
rect 676 -2196 680 -2164
rect 640 -2244 680 -2196
rect 640 -2276 644 -2244
rect 676 -2276 680 -2244
rect 640 -2324 680 -2276
rect 640 -2356 644 -2324
rect 676 -2356 680 -2324
rect 640 -2404 680 -2356
rect 640 -2436 644 -2404
rect 676 -2436 680 -2404
rect 640 -2484 680 -2436
rect 640 -2516 644 -2484
rect 676 -2516 680 -2484
rect 640 -2564 680 -2516
rect 640 -2596 644 -2564
rect 676 -2596 680 -2564
rect 640 -2644 680 -2596
rect 640 -2676 644 -2644
rect 676 -2676 680 -2644
rect 640 -2724 680 -2676
rect 640 -2756 644 -2724
rect 676 -2756 680 -2724
rect 640 -2804 680 -2756
rect 640 -2836 644 -2804
rect 676 -2836 680 -2804
rect 640 -2884 680 -2836
rect 640 -2916 644 -2884
rect 676 -2916 680 -2884
rect 640 -2964 680 -2916
rect 640 -2996 644 -2964
rect 676 -2996 680 -2964
rect 640 -3044 680 -2996
rect 640 -3076 644 -3044
rect 676 -3076 680 -3044
rect 640 -3124 680 -3076
rect 640 -3156 644 -3124
rect 676 -3156 680 -3124
rect 640 -3204 680 -3156
rect 640 -3236 644 -3204
rect 676 -3236 680 -3204
rect 640 -3284 680 -3236
rect 640 -3316 644 -3284
rect 676 -3316 680 -3284
rect 640 -3364 680 -3316
rect 640 -3396 644 -3364
rect 676 -3396 680 -3364
rect 640 -3444 680 -3396
rect 640 -3476 644 -3444
rect 676 -3476 680 -3444
rect 640 -3524 680 -3476
rect 640 -3556 644 -3524
rect 676 -3556 680 -3524
rect 640 -3604 680 -3556
rect 640 -3636 644 -3604
rect 676 -3636 680 -3604
rect 640 -3684 680 -3636
rect 640 -3716 644 -3684
rect 676 -3716 680 -3684
rect 640 -3720 680 -3716
rect 720 1036 760 1040
rect 720 1004 724 1036
rect 756 1004 760 1036
rect 720 956 760 1004
rect 720 924 724 956
rect 756 924 760 956
rect 720 876 760 924
rect 720 844 724 876
rect 756 844 760 876
rect 720 796 760 844
rect 720 764 724 796
rect 756 764 760 796
rect 720 716 760 764
rect 720 684 724 716
rect 756 684 760 716
rect 720 636 760 684
rect 720 604 724 636
rect 756 604 760 636
rect 720 556 760 604
rect 720 524 724 556
rect 756 524 760 556
rect 720 476 760 524
rect 720 444 724 476
rect 756 444 760 476
rect 720 396 760 444
rect 720 364 724 396
rect 756 364 760 396
rect 720 316 760 364
rect 720 284 724 316
rect 756 284 760 316
rect 720 236 760 284
rect 720 204 724 236
rect 756 204 760 236
rect 720 156 760 204
rect 720 124 724 156
rect 756 124 760 156
rect 720 76 760 124
rect 720 44 724 76
rect 756 44 760 76
rect 720 -4 760 44
rect 720 -36 724 -4
rect 756 -36 760 -4
rect 720 -84 760 -36
rect 720 -116 724 -84
rect 756 -116 760 -84
rect 720 -164 760 -116
rect 720 -196 724 -164
rect 756 -196 760 -164
rect 720 -244 760 -196
rect 720 -276 724 -244
rect 756 -276 760 -244
rect 720 -324 760 -276
rect 720 -356 724 -324
rect 756 -356 760 -324
rect 720 -404 760 -356
rect 720 -436 724 -404
rect 756 -436 760 -404
rect 720 -484 760 -436
rect 720 -516 724 -484
rect 756 -516 760 -484
rect 720 -564 760 -516
rect 720 -596 724 -564
rect 756 -596 760 -564
rect 720 -644 760 -596
rect 720 -676 724 -644
rect 756 -676 760 -644
rect 720 -724 760 -676
rect 720 -756 724 -724
rect 756 -756 760 -724
rect 720 -804 760 -756
rect 720 -836 724 -804
rect 756 -836 760 -804
rect 720 -884 760 -836
rect 720 -916 724 -884
rect 756 -916 760 -884
rect 720 -964 760 -916
rect 720 -996 724 -964
rect 756 -996 760 -964
rect 720 -1044 760 -996
rect 720 -1076 724 -1044
rect 756 -1076 760 -1044
rect 720 -1124 760 -1076
rect 720 -1156 724 -1124
rect 756 -1156 760 -1124
rect 720 -1204 760 -1156
rect 720 -1236 724 -1204
rect 756 -1236 760 -1204
rect 720 -1284 760 -1236
rect 720 -1316 724 -1284
rect 756 -1316 760 -1284
rect 720 -1364 760 -1316
rect 720 -1396 724 -1364
rect 756 -1396 760 -1364
rect 720 -1444 760 -1396
rect 720 -1476 724 -1444
rect 756 -1476 760 -1444
rect 720 -1524 760 -1476
rect 720 -1556 724 -1524
rect 756 -1556 760 -1524
rect 720 -1604 760 -1556
rect 720 -1636 724 -1604
rect 756 -1636 760 -1604
rect 720 -1684 760 -1636
rect 720 -1716 724 -1684
rect 756 -1716 760 -1684
rect 720 -1764 760 -1716
rect 720 -1796 724 -1764
rect 756 -1796 760 -1764
rect 720 -1844 760 -1796
rect 720 -1876 724 -1844
rect 756 -1876 760 -1844
rect 720 -1924 760 -1876
rect 720 -1956 724 -1924
rect 756 -1956 760 -1924
rect 720 -2004 760 -1956
rect 720 -2036 724 -2004
rect 756 -2036 760 -2004
rect 720 -2084 760 -2036
rect 720 -2116 724 -2084
rect 756 -2116 760 -2084
rect 720 -2164 760 -2116
rect 720 -2196 724 -2164
rect 756 -2196 760 -2164
rect 720 -2244 760 -2196
rect 720 -2276 724 -2244
rect 756 -2276 760 -2244
rect 720 -2324 760 -2276
rect 720 -2356 724 -2324
rect 756 -2356 760 -2324
rect 720 -2404 760 -2356
rect 720 -2436 724 -2404
rect 756 -2436 760 -2404
rect 720 -2484 760 -2436
rect 720 -2516 724 -2484
rect 756 -2516 760 -2484
rect 720 -2564 760 -2516
rect 720 -2596 724 -2564
rect 756 -2596 760 -2564
rect 720 -2644 760 -2596
rect 720 -2676 724 -2644
rect 756 -2676 760 -2644
rect 720 -2724 760 -2676
rect 720 -2756 724 -2724
rect 756 -2756 760 -2724
rect 720 -2804 760 -2756
rect 720 -2836 724 -2804
rect 756 -2836 760 -2804
rect 720 -2884 760 -2836
rect 720 -2916 724 -2884
rect 756 -2916 760 -2884
rect 720 -2964 760 -2916
rect 720 -2996 724 -2964
rect 756 -2996 760 -2964
rect 720 -3044 760 -2996
rect 720 -3076 724 -3044
rect 756 -3076 760 -3044
rect 720 -3124 760 -3076
rect 720 -3156 724 -3124
rect 756 -3156 760 -3124
rect 720 -3204 760 -3156
rect 720 -3236 724 -3204
rect 756 -3236 760 -3204
rect 720 -3284 760 -3236
rect 720 -3316 724 -3284
rect 756 -3316 760 -3284
rect 720 -3364 760 -3316
rect 720 -3396 724 -3364
rect 756 -3396 760 -3364
rect 720 -3444 760 -3396
rect 720 -3476 724 -3444
rect 756 -3476 760 -3444
rect 720 -3524 760 -3476
rect 720 -3556 724 -3524
rect 756 -3556 760 -3524
rect 720 -3604 760 -3556
rect 720 -3636 724 -3604
rect 756 -3636 760 -3604
rect 720 -3684 760 -3636
rect 720 -3716 724 -3684
rect 756 -3716 760 -3684
rect 720 -3720 760 -3716
rect 800 1036 840 1040
rect 800 1004 804 1036
rect 836 1004 840 1036
rect 800 956 840 1004
rect 800 924 804 956
rect 836 924 840 956
rect 800 876 840 924
rect 800 844 804 876
rect 836 844 840 876
rect 800 796 840 844
rect 800 764 804 796
rect 836 764 840 796
rect 800 716 840 764
rect 800 684 804 716
rect 836 684 840 716
rect 800 636 840 684
rect 800 604 804 636
rect 836 604 840 636
rect 800 556 840 604
rect 800 524 804 556
rect 836 524 840 556
rect 800 476 840 524
rect 800 444 804 476
rect 836 444 840 476
rect 800 396 840 444
rect 800 364 804 396
rect 836 364 840 396
rect 800 316 840 364
rect 800 284 804 316
rect 836 284 840 316
rect 800 236 840 284
rect 800 204 804 236
rect 836 204 840 236
rect 800 156 840 204
rect 800 124 804 156
rect 836 124 840 156
rect 800 76 840 124
rect 800 44 804 76
rect 836 44 840 76
rect 800 -4 840 44
rect 800 -36 804 -4
rect 836 -36 840 -4
rect 800 -84 840 -36
rect 800 -116 804 -84
rect 836 -116 840 -84
rect 800 -164 840 -116
rect 800 -196 804 -164
rect 836 -196 840 -164
rect 800 -244 840 -196
rect 800 -276 804 -244
rect 836 -276 840 -244
rect 800 -324 840 -276
rect 800 -356 804 -324
rect 836 -356 840 -324
rect 800 -404 840 -356
rect 800 -436 804 -404
rect 836 -436 840 -404
rect 800 -484 840 -436
rect 800 -516 804 -484
rect 836 -516 840 -484
rect 800 -564 840 -516
rect 800 -596 804 -564
rect 836 -596 840 -564
rect 800 -644 840 -596
rect 800 -676 804 -644
rect 836 -676 840 -644
rect 800 -724 840 -676
rect 800 -756 804 -724
rect 836 -756 840 -724
rect 800 -804 840 -756
rect 800 -836 804 -804
rect 836 -836 840 -804
rect 800 -884 840 -836
rect 800 -916 804 -884
rect 836 -916 840 -884
rect 800 -964 840 -916
rect 800 -996 804 -964
rect 836 -996 840 -964
rect 800 -1044 840 -996
rect 800 -1076 804 -1044
rect 836 -1076 840 -1044
rect 800 -1124 840 -1076
rect 800 -1156 804 -1124
rect 836 -1156 840 -1124
rect 800 -1204 840 -1156
rect 800 -1236 804 -1204
rect 836 -1236 840 -1204
rect 800 -1284 840 -1236
rect 800 -1316 804 -1284
rect 836 -1316 840 -1284
rect 800 -1364 840 -1316
rect 800 -1396 804 -1364
rect 836 -1396 840 -1364
rect 800 -1444 840 -1396
rect 800 -1476 804 -1444
rect 836 -1476 840 -1444
rect 800 -1524 840 -1476
rect 800 -1556 804 -1524
rect 836 -1556 840 -1524
rect 800 -1604 840 -1556
rect 800 -1636 804 -1604
rect 836 -1636 840 -1604
rect 800 -1684 840 -1636
rect 800 -1716 804 -1684
rect 836 -1716 840 -1684
rect 800 -1764 840 -1716
rect 800 -1796 804 -1764
rect 836 -1796 840 -1764
rect 800 -1844 840 -1796
rect 800 -1876 804 -1844
rect 836 -1876 840 -1844
rect 800 -1924 840 -1876
rect 800 -1956 804 -1924
rect 836 -1956 840 -1924
rect 800 -2004 840 -1956
rect 800 -2036 804 -2004
rect 836 -2036 840 -2004
rect 800 -2084 840 -2036
rect 800 -2116 804 -2084
rect 836 -2116 840 -2084
rect 800 -2164 840 -2116
rect 800 -2196 804 -2164
rect 836 -2196 840 -2164
rect 800 -2244 840 -2196
rect 800 -2276 804 -2244
rect 836 -2276 840 -2244
rect 800 -2324 840 -2276
rect 800 -2356 804 -2324
rect 836 -2356 840 -2324
rect 800 -2404 840 -2356
rect 800 -2436 804 -2404
rect 836 -2436 840 -2404
rect 800 -2484 840 -2436
rect 800 -2516 804 -2484
rect 836 -2516 840 -2484
rect 800 -2564 840 -2516
rect 800 -2596 804 -2564
rect 836 -2596 840 -2564
rect 800 -2644 840 -2596
rect 800 -2676 804 -2644
rect 836 -2676 840 -2644
rect 800 -2724 840 -2676
rect 800 -2756 804 -2724
rect 836 -2756 840 -2724
rect 800 -2804 840 -2756
rect 800 -2836 804 -2804
rect 836 -2836 840 -2804
rect 800 -2884 840 -2836
rect 800 -2916 804 -2884
rect 836 -2916 840 -2884
rect 800 -2964 840 -2916
rect 800 -2996 804 -2964
rect 836 -2996 840 -2964
rect 800 -3044 840 -2996
rect 800 -3076 804 -3044
rect 836 -3076 840 -3044
rect 800 -3124 840 -3076
rect 800 -3156 804 -3124
rect 836 -3156 840 -3124
rect 800 -3204 840 -3156
rect 800 -3236 804 -3204
rect 836 -3236 840 -3204
rect 800 -3284 840 -3236
rect 800 -3316 804 -3284
rect 836 -3316 840 -3284
rect 800 -3364 840 -3316
rect 800 -3396 804 -3364
rect 836 -3396 840 -3364
rect 800 -3444 840 -3396
rect 800 -3476 804 -3444
rect 836 -3476 840 -3444
rect 800 -3524 840 -3476
rect 800 -3556 804 -3524
rect 836 -3556 840 -3524
rect 800 -3604 840 -3556
rect 800 -3636 804 -3604
rect 836 -3636 840 -3604
rect 800 -3684 840 -3636
rect 800 -3716 804 -3684
rect 836 -3716 840 -3684
rect 800 -3720 840 -3716
rect 880 1036 920 1040
rect 880 1004 884 1036
rect 916 1004 920 1036
rect 880 956 920 1004
rect 880 924 884 956
rect 916 924 920 956
rect 880 876 920 924
rect 880 844 884 876
rect 916 844 920 876
rect 880 796 920 844
rect 880 764 884 796
rect 916 764 920 796
rect 880 716 920 764
rect 880 684 884 716
rect 916 684 920 716
rect 880 636 920 684
rect 880 604 884 636
rect 916 604 920 636
rect 880 556 920 604
rect 880 524 884 556
rect 916 524 920 556
rect 880 476 920 524
rect 880 444 884 476
rect 916 444 920 476
rect 880 396 920 444
rect 880 364 884 396
rect 916 364 920 396
rect 880 316 920 364
rect 880 284 884 316
rect 916 284 920 316
rect 880 236 920 284
rect 880 204 884 236
rect 916 204 920 236
rect 880 156 920 204
rect 880 124 884 156
rect 916 124 920 156
rect 880 76 920 124
rect 880 44 884 76
rect 916 44 920 76
rect 880 -4 920 44
rect 880 -36 884 -4
rect 916 -36 920 -4
rect 880 -84 920 -36
rect 880 -116 884 -84
rect 916 -116 920 -84
rect 880 -164 920 -116
rect 880 -196 884 -164
rect 916 -196 920 -164
rect 880 -244 920 -196
rect 880 -276 884 -244
rect 916 -276 920 -244
rect 880 -324 920 -276
rect 880 -356 884 -324
rect 916 -356 920 -324
rect 880 -404 920 -356
rect 880 -436 884 -404
rect 916 -436 920 -404
rect 880 -484 920 -436
rect 880 -516 884 -484
rect 916 -516 920 -484
rect 880 -564 920 -516
rect 880 -596 884 -564
rect 916 -596 920 -564
rect 880 -644 920 -596
rect 880 -676 884 -644
rect 916 -676 920 -644
rect 880 -724 920 -676
rect 880 -756 884 -724
rect 916 -756 920 -724
rect 880 -804 920 -756
rect 880 -836 884 -804
rect 916 -836 920 -804
rect 880 -884 920 -836
rect 880 -916 884 -884
rect 916 -916 920 -884
rect 880 -964 920 -916
rect 880 -996 884 -964
rect 916 -996 920 -964
rect 880 -1044 920 -996
rect 880 -1076 884 -1044
rect 916 -1076 920 -1044
rect 880 -1124 920 -1076
rect 880 -1156 884 -1124
rect 916 -1156 920 -1124
rect 880 -1204 920 -1156
rect 880 -1236 884 -1204
rect 916 -1236 920 -1204
rect 880 -1284 920 -1236
rect 880 -1316 884 -1284
rect 916 -1316 920 -1284
rect 880 -1364 920 -1316
rect 880 -1396 884 -1364
rect 916 -1396 920 -1364
rect 880 -1444 920 -1396
rect 880 -1476 884 -1444
rect 916 -1476 920 -1444
rect 880 -1524 920 -1476
rect 880 -1556 884 -1524
rect 916 -1556 920 -1524
rect 880 -1604 920 -1556
rect 880 -1636 884 -1604
rect 916 -1636 920 -1604
rect 880 -1684 920 -1636
rect 880 -1716 884 -1684
rect 916 -1716 920 -1684
rect 880 -1764 920 -1716
rect 880 -1796 884 -1764
rect 916 -1796 920 -1764
rect 880 -1844 920 -1796
rect 880 -1876 884 -1844
rect 916 -1876 920 -1844
rect 880 -1924 920 -1876
rect 880 -1956 884 -1924
rect 916 -1956 920 -1924
rect 880 -2004 920 -1956
rect 880 -2036 884 -2004
rect 916 -2036 920 -2004
rect 880 -2084 920 -2036
rect 880 -2116 884 -2084
rect 916 -2116 920 -2084
rect 880 -2164 920 -2116
rect 880 -2196 884 -2164
rect 916 -2196 920 -2164
rect 880 -2244 920 -2196
rect 880 -2276 884 -2244
rect 916 -2276 920 -2244
rect 880 -2324 920 -2276
rect 880 -2356 884 -2324
rect 916 -2356 920 -2324
rect 880 -2404 920 -2356
rect 880 -2436 884 -2404
rect 916 -2436 920 -2404
rect 880 -2484 920 -2436
rect 880 -2516 884 -2484
rect 916 -2516 920 -2484
rect 880 -2564 920 -2516
rect 880 -2596 884 -2564
rect 916 -2596 920 -2564
rect 880 -2644 920 -2596
rect 880 -2676 884 -2644
rect 916 -2676 920 -2644
rect 880 -2724 920 -2676
rect 880 -2756 884 -2724
rect 916 -2756 920 -2724
rect 880 -2804 920 -2756
rect 880 -2836 884 -2804
rect 916 -2836 920 -2804
rect 880 -2884 920 -2836
rect 880 -2916 884 -2884
rect 916 -2916 920 -2884
rect 880 -2964 920 -2916
rect 880 -2996 884 -2964
rect 916 -2996 920 -2964
rect 880 -3044 920 -2996
rect 880 -3076 884 -3044
rect 916 -3076 920 -3044
rect 880 -3124 920 -3076
rect 880 -3156 884 -3124
rect 916 -3156 920 -3124
rect 880 -3204 920 -3156
rect 880 -3236 884 -3204
rect 916 -3236 920 -3204
rect 880 -3284 920 -3236
rect 880 -3316 884 -3284
rect 916 -3316 920 -3284
rect 880 -3364 920 -3316
rect 880 -3396 884 -3364
rect 916 -3396 920 -3364
rect 880 -3444 920 -3396
rect 880 -3476 884 -3444
rect 916 -3476 920 -3444
rect 880 -3524 920 -3476
rect 880 -3556 884 -3524
rect 916 -3556 920 -3524
rect 880 -3604 920 -3556
rect 880 -3636 884 -3604
rect 916 -3636 920 -3604
rect 880 -3684 920 -3636
rect 880 -3716 884 -3684
rect 916 -3716 920 -3684
rect 880 -3720 920 -3716
rect 960 1036 1000 1040
rect 960 1004 964 1036
rect 996 1004 1000 1036
rect 960 956 1000 1004
rect 960 924 964 956
rect 996 924 1000 956
rect 960 876 1000 924
rect 960 844 964 876
rect 996 844 1000 876
rect 960 796 1000 844
rect 960 764 964 796
rect 996 764 1000 796
rect 960 716 1000 764
rect 960 684 964 716
rect 996 684 1000 716
rect 960 636 1000 684
rect 960 604 964 636
rect 996 604 1000 636
rect 960 556 1000 604
rect 960 524 964 556
rect 996 524 1000 556
rect 960 476 1000 524
rect 960 444 964 476
rect 996 444 1000 476
rect 960 396 1000 444
rect 960 364 964 396
rect 996 364 1000 396
rect 960 316 1000 364
rect 960 284 964 316
rect 996 284 1000 316
rect 960 236 1000 284
rect 960 204 964 236
rect 996 204 1000 236
rect 960 156 1000 204
rect 960 124 964 156
rect 996 124 1000 156
rect 960 76 1000 124
rect 960 44 964 76
rect 996 44 1000 76
rect 960 -4 1000 44
rect 960 -36 964 -4
rect 996 -36 1000 -4
rect 960 -84 1000 -36
rect 960 -116 964 -84
rect 996 -116 1000 -84
rect 960 -164 1000 -116
rect 960 -196 964 -164
rect 996 -196 1000 -164
rect 960 -244 1000 -196
rect 960 -276 964 -244
rect 996 -276 1000 -244
rect 960 -324 1000 -276
rect 960 -356 964 -324
rect 996 -356 1000 -324
rect 960 -404 1000 -356
rect 960 -436 964 -404
rect 996 -436 1000 -404
rect 960 -484 1000 -436
rect 960 -516 964 -484
rect 996 -516 1000 -484
rect 960 -564 1000 -516
rect 960 -596 964 -564
rect 996 -596 1000 -564
rect 960 -644 1000 -596
rect 960 -676 964 -644
rect 996 -676 1000 -644
rect 960 -724 1000 -676
rect 960 -756 964 -724
rect 996 -756 1000 -724
rect 960 -804 1000 -756
rect 960 -836 964 -804
rect 996 -836 1000 -804
rect 960 -884 1000 -836
rect 960 -916 964 -884
rect 996 -916 1000 -884
rect 960 -964 1000 -916
rect 960 -996 964 -964
rect 996 -996 1000 -964
rect 960 -1044 1000 -996
rect 960 -1076 964 -1044
rect 996 -1076 1000 -1044
rect 960 -1124 1000 -1076
rect 960 -1156 964 -1124
rect 996 -1156 1000 -1124
rect 960 -1204 1000 -1156
rect 960 -1236 964 -1204
rect 996 -1236 1000 -1204
rect 960 -1284 1000 -1236
rect 960 -1316 964 -1284
rect 996 -1316 1000 -1284
rect 960 -1364 1000 -1316
rect 960 -1396 964 -1364
rect 996 -1396 1000 -1364
rect 960 -1444 1000 -1396
rect 960 -1476 964 -1444
rect 996 -1476 1000 -1444
rect 960 -1524 1000 -1476
rect 960 -1556 964 -1524
rect 996 -1556 1000 -1524
rect 960 -1604 1000 -1556
rect 960 -1636 964 -1604
rect 996 -1636 1000 -1604
rect 960 -1684 1000 -1636
rect 960 -1716 964 -1684
rect 996 -1716 1000 -1684
rect 960 -1764 1000 -1716
rect 960 -1796 964 -1764
rect 996 -1796 1000 -1764
rect 960 -1844 1000 -1796
rect 960 -1876 964 -1844
rect 996 -1876 1000 -1844
rect 960 -1924 1000 -1876
rect 960 -1956 964 -1924
rect 996 -1956 1000 -1924
rect 960 -2004 1000 -1956
rect 960 -2036 964 -2004
rect 996 -2036 1000 -2004
rect 960 -2084 1000 -2036
rect 960 -2116 964 -2084
rect 996 -2116 1000 -2084
rect 960 -2164 1000 -2116
rect 960 -2196 964 -2164
rect 996 -2196 1000 -2164
rect 960 -2244 1000 -2196
rect 960 -2276 964 -2244
rect 996 -2276 1000 -2244
rect 960 -2324 1000 -2276
rect 960 -2356 964 -2324
rect 996 -2356 1000 -2324
rect 960 -2404 1000 -2356
rect 960 -2436 964 -2404
rect 996 -2436 1000 -2404
rect 960 -2484 1000 -2436
rect 960 -2516 964 -2484
rect 996 -2516 1000 -2484
rect 960 -2564 1000 -2516
rect 960 -2596 964 -2564
rect 996 -2596 1000 -2564
rect 960 -2644 1000 -2596
rect 960 -2676 964 -2644
rect 996 -2676 1000 -2644
rect 960 -2724 1000 -2676
rect 960 -2756 964 -2724
rect 996 -2756 1000 -2724
rect 960 -2804 1000 -2756
rect 960 -2836 964 -2804
rect 996 -2836 1000 -2804
rect 960 -2884 1000 -2836
rect 960 -2916 964 -2884
rect 996 -2916 1000 -2884
rect 960 -2964 1000 -2916
rect 960 -2996 964 -2964
rect 996 -2996 1000 -2964
rect 960 -3044 1000 -2996
rect 960 -3076 964 -3044
rect 996 -3076 1000 -3044
rect 960 -3124 1000 -3076
rect 960 -3156 964 -3124
rect 996 -3156 1000 -3124
rect 960 -3204 1000 -3156
rect 960 -3236 964 -3204
rect 996 -3236 1000 -3204
rect 960 -3284 1000 -3236
rect 960 -3316 964 -3284
rect 996 -3316 1000 -3284
rect 960 -3364 1000 -3316
rect 960 -3396 964 -3364
rect 996 -3396 1000 -3364
rect 960 -3444 1000 -3396
rect 960 -3476 964 -3444
rect 996 -3476 1000 -3444
rect 960 -3524 1000 -3476
rect 960 -3556 964 -3524
rect 996 -3556 1000 -3524
rect 960 -3604 1000 -3556
rect 960 -3636 964 -3604
rect 996 -3636 1000 -3604
rect 960 -3684 1000 -3636
rect 960 -3716 964 -3684
rect 996 -3716 1000 -3684
rect 960 -3720 1000 -3716
rect 1040 1036 1080 1040
rect 1040 1004 1044 1036
rect 1076 1004 1080 1036
rect 1040 956 1080 1004
rect 1040 924 1044 956
rect 1076 924 1080 956
rect 1040 876 1080 924
rect 1040 844 1044 876
rect 1076 844 1080 876
rect 1040 796 1080 844
rect 1040 764 1044 796
rect 1076 764 1080 796
rect 1040 716 1080 764
rect 1040 684 1044 716
rect 1076 684 1080 716
rect 1040 636 1080 684
rect 1040 604 1044 636
rect 1076 604 1080 636
rect 1040 556 1080 604
rect 1040 524 1044 556
rect 1076 524 1080 556
rect 1040 476 1080 524
rect 1040 444 1044 476
rect 1076 444 1080 476
rect 1040 396 1080 444
rect 1040 364 1044 396
rect 1076 364 1080 396
rect 1040 316 1080 364
rect 1040 284 1044 316
rect 1076 284 1080 316
rect 1040 236 1080 284
rect 1040 204 1044 236
rect 1076 204 1080 236
rect 1040 156 1080 204
rect 1040 124 1044 156
rect 1076 124 1080 156
rect 1040 76 1080 124
rect 1040 44 1044 76
rect 1076 44 1080 76
rect 1040 -4 1080 44
rect 1040 -36 1044 -4
rect 1076 -36 1080 -4
rect 1040 -84 1080 -36
rect 1040 -116 1044 -84
rect 1076 -116 1080 -84
rect 1040 -164 1080 -116
rect 1040 -196 1044 -164
rect 1076 -196 1080 -164
rect 1040 -244 1080 -196
rect 1040 -276 1044 -244
rect 1076 -276 1080 -244
rect 1040 -324 1080 -276
rect 1040 -356 1044 -324
rect 1076 -356 1080 -324
rect 1040 -404 1080 -356
rect 1040 -436 1044 -404
rect 1076 -436 1080 -404
rect 1040 -484 1080 -436
rect 1040 -516 1044 -484
rect 1076 -516 1080 -484
rect 1040 -564 1080 -516
rect 1040 -596 1044 -564
rect 1076 -596 1080 -564
rect 1040 -644 1080 -596
rect 1040 -676 1044 -644
rect 1076 -676 1080 -644
rect 1040 -724 1080 -676
rect 1040 -756 1044 -724
rect 1076 -756 1080 -724
rect 1040 -804 1080 -756
rect 1040 -836 1044 -804
rect 1076 -836 1080 -804
rect 1040 -884 1080 -836
rect 1040 -916 1044 -884
rect 1076 -916 1080 -884
rect 1040 -964 1080 -916
rect 1040 -996 1044 -964
rect 1076 -996 1080 -964
rect 1040 -1044 1080 -996
rect 1040 -1076 1044 -1044
rect 1076 -1076 1080 -1044
rect 1040 -1124 1080 -1076
rect 1040 -1156 1044 -1124
rect 1076 -1156 1080 -1124
rect 1040 -1204 1080 -1156
rect 1040 -1236 1044 -1204
rect 1076 -1236 1080 -1204
rect 1040 -1284 1080 -1236
rect 1040 -1316 1044 -1284
rect 1076 -1316 1080 -1284
rect 1040 -1364 1080 -1316
rect 1040 -1396 1044 -1364
rect 1076 -1396 1080 -1364
rect 1040 -1444 1080 -1396
rect 1040 -1476 1044 -1444
rect 1076 -1476 1080 -1444
rect 1040 -1524 1080 -1476
rect 1040 -1556 1044 -1524
rect 1076 -1556 1080 -1524
rect 1040 -1604 1080 -1556
rect 1040 -1636 1044 -1604
rect 1076 -1636 1080 -1604
rect 1040 -1684 1080 -1636
rect 1040 -1716 1044 -1684
rect 1076 -1716 1080 -1684
rect 1040 -1764 1080 -1716
rect 1040 -1796 1044 -1764
rect 1076 -1796 1080 -1764
rect 1040 -1844 1080 -1796
rect 1040 -1876 1044 -1844
rect 1076 -1876 1080 -1844
rect 1040 -1924 1080 -1876
rect 1040 -1956 1044 -1924
rect 1076 -1956 1080 -1924
rect 1040 -2004 1080 -1956
rect 1040 -2036 1044 -2004
rect 1076 -2036 1080 -2004
rect 1040 -2084 1080 -2036
rect 1040 -2116 1044 -2084
rect 1076 -2116 1080 -2084
rect 1040 -2164 1080 -2116
rect 1040 -2196 1044 -2164
rect 1076 -2196 1080 -2164
rect 1040 -2244 1080 -2196
rect 1040 -2276 1044 -2244
rect 1076 -2276 1080 -2244
rect 1040 -2324 1080 -2276
rect 1040 -2356 1044 -2324
rect 1076 -2356 1080 -2324
rect 1040 -2404 1080 -2356
rect 1040 -2436 1044 -2404
rect 1076 -2436 1080 -2404
rect 1040 -2484 1080 -2436
rect 1040 -2516 1044 -2484
rect 1076 -2516 1080 -2484
rect 1040 -2564 1080 -2516
rect 1040 -2596 1044 -2564
rect 1076 -2596 1080 -2564
rect 1040 -2644 1080 -2596
rect 1040 -2676 1044 -2644
rect 1076 -2676 1080 -2644
rect 1040 -2724 1080 -2676
rect 1040 -2756 1044 -2724
rect 1076 -2756 1080 -2724
rect 1040 -2804 1080 -2756
rect 1040 -2836 1044 -2804
rect 1076 -2836 1080 -2804
rect 1040 -2884 1080 -2836
rect 1040 -2916 1044 -2884
rect 1076 -2916 1080 -2884
rect 1040 -2964 1080 -2916
rect 1040 -2996 1044 -2964
rect 1076 -2996 1080 -2964
rect 1040 -3044 1080 -2996
rect 1040 -3076 1044 -3044
rect 1076 -3076 1080 -3044
rect 1040 -3124 1080 -3076
rect 1040 -3156 1044 -3124
rect 1076 -3156 1080 -3124
rect 1040 -3204 1080 -3156
rect 1040 -3236 1044 -3204
rect 1076 -3236 1080 -3204
rect 1040 -3284 1080 -3236
rect 1040 -3316 1044 -3284
rect 1076 -3316 1080 -3284
rect 1040 -3364 1080 -3316
rect 1040 -3396 1044 -3364
rect 1076 -3396 1080 -3364
rect 1040 -3444 1080 -3396
rect 1040 -3476 1044 -3444
rect 1076 -3476 1080 -3444
rect 1040 -3524 1080 -3476
rect 1040 -3556 1044 -3524
rect 1076 -3556 1080 -3524
rect 1040 -3604 1080 -3556
rect 1040 -3636 1044 -3604
rect 1076 -3636 1080 -3604
rect 1040 -3684 1080 -3636
rect 1040 -3716 1044 -3684
rect 1076 -3716 1080 -3684
rect 1040 -3720 1080 -3716
rect 1120 1036 1160 1040
rect 1120 1004 1124 1036
rect 1156 1004 1160 1036
rect 1120 956 1160 1004
rect 1120 924 1124 956
rect 1156 924 1160 956
rect 1120 876 1160 924
rect 1120 844 1124 876
rect 1156 844 1160 876
rect 1120 796 1160 844
rect 1120 764 1124 796
rect 1156 764 1160 796
rect 1120 716 1160 764
rect 1120 684 1124 716
rect 1156 684 1160 716
rect 1120 636 1160 684
rect 1120 604 1124 636
rect 1156 604 1160 636
rect 1120 556 1160 604
rect 1120 524 1124 556
rect 1156 524 1160 556
rect 1120 476 1160 524
rect 1120 444 1124 476
rect 1156 444 1160 476
rect 1120 396 1160 444
rect 1120 364 1124 396
rect 1156 364 1160 396
rect 1120 316 1160 364
rect 1120 284 1124 316
rect 1156 284 1160 316
rect 1120 236 1160 284
rect 1120 204 1124 236
rect 1156 204 1160 236
rect 1120 156 1160 204
rect 1120 124 1124 156
rect 1156 124 1160 156
rect 1120 76 1160 124
rect 1120 44 1124 76
rect 1156 44 1160 76
rect 1120 -4 1160 44
rect 1120 -36 1124 -4
rect 1156 -36 1160 -4
rect 1120 -84 1160 -36
rect 1120 -116 1124 -84
rect 1156 -116 1160 -84
rect 1120 -164 1160 -116
rect 1120 -196 1124 -164
rect 1156 -196 1160 -164
rect 1120 -244 1160 -196
rect 1120 -276 1124 -244
rect 1156 -276 1160 -244
rect 1120 -324 1160 -276
rect 1120 -356 1124 -324
rect 1156 -356 1160 -324
rect 1120 -404 1160 -356
rect 1120 -436 1124 -404
rect 1156 -436 1160 -404
rect 1120 -484 1160 -436
rect 1120 -516 1124 -484
rect 1156 -516 1160 -484
rect 1120 -564 1160 -516
rect 1120 -596 1124 -564
rect 1156 -596 1160 -564
rect 1120 -644 1160 -596
rect 1120 -676 1124 -644
rect 1156 -676 1160 -644
rect 1120 -724 1160 -676
rect 1120 -756 1124 -724
rect 1156 -756 1160 -724
rect 1120 -804 1160 -756
rect 1120 -836 1124 -804
rect 1156 -836 1160 -804
rect 1120 -884 1160 -836
rect 1120 -916 1124 -884
rect 1156 -916 1160 -884
rect 1120 -964 1160 -916
rect 1120 -996 1124 -964
rect 1156 -996 1160 -964
rect 1120 -1044 1160 -996
rect 1120 -1076 1124 -1044
rect 1156 -1076 1160 -1044
rect 1120 -1124 1160 -1076
rect 1120 -1156 1124 -1124
rect 1156 -1156 1160 -1124
rect 1120 -1204 1160 -1156
rect 1120 -1236 1124 -1204
rect 1156 -1236 1160 -1204
rect 1120 -1284 1160 -1236
rect 1120 -1316 1124 -1284
rect 1156 -1316 1160 -1284
rect 1120 -1364 1160 -1316
rect 1120 -1396 1124 -1364
rect 1156 -1396 1160 -1364
rect 1120 -1444 1160 -1396
rect 1120 -1476 1124 -1444
rect 1156 -1476 1160 -1444
rect 1120 -1524 1160 -1476
rect 1120 -1556 1124 -1524
rect 1156 -1556 1160 -1524
rect 1120 -1604 1160 -1556
rect 1120 -1636 1124 -1604
rect 1156 -1636 1160 -1604
rect 1120 -1684 1160 -1636
rect 1120 -1716 1124 -1684
rect 1156 -1716 1160 -1684
rect 1120 -1764 1160 -1716
rect 1120 -1796 1124 -1764
rect 1156 -1796 1160 -1764
rect 1120 -1844 1160 -1796
rect 1120 -1876 1124 -1844
rect 1156 -1876 1160 -1844
rect 1120 -1924 1160 -1876
rect 1120 -1956 1124 -1924
rect 1156 -1956 1160 -1924
rect 1120 -2004 1160 -1956
rect 1120 -2036 1124 -2004
rect 1156 -2036 1160 -2004
rect 1120 -2084 1160 -2036
rect 1120 -2116 1124 -2084
rect 1156 -2116 1160 -2084
rect 1120 -2164 1160 -2116
rect 1120 -2196 1124 -2164
rect 1156 -2196 1160 -2164
rect 1120 -2244 1160 -2196
rect 1120 -2276 1124 -2244
rect 1156 -2276 1160 -2244
rect 1120 -2324 1160 -2276
rect 1120 -2356 1124 -2324
rect 1156 -2356 1160 -2324
rect 1120 -2404 1160 -2356
rect 1120 -2436 1124 -2404
rect 1156 -2436 1160 -2404
rect 1120 -2484 1160 -2436
rect 1120 -2516 1124 -2484
rect 1156 -2516 1160 -2484
rect 1120 -2564 1160 -2516
rect 1120 -2596 1124 -2564
rect 1156 -2596 1160 -2564
rect 1120 -2644 1160 -2596
rect 1120 -2676 1124 -2644
rect 1156 -2676 1160 -2644
rect 1120 -2724 1160 -2676
rect 1120 -2756 1124 -2724
rect 1156 -2756 1160 -2724
rect 1120 -2804 1160 -2756
rect 1120 -2836 1124 -2804
rect 1156 -2836 1160 -2804
rect 1120 -2884 1160 -2836
rect 1120 -2916 1124 -2884
rect 1156 -2916 1160 -2884
rect 1120 -2964 1160 -2916
rect 1120 -2996 1124 -2964
rect 1156 -2996 1160 -2964
rect 1120 -3044 1160 -2996
rect 1120 -3076 1124 -3044
rect 1156 -3076 1160 -3044
rect 1120 -3124 1160 -3076
rect 1120 -3156 1124 -3124
rect 1156 -3156 1160 -3124
rect 1120 -3204 1160 -3156
rect 1120 -3236 1124 -3204
rect 1156 -3236 1160 -3204
rect 1120 -3284 1160 -3236
rect 1120 -3316 1124 -3284
rect 1156 -3316 1160 -3284
rect 1120 -3364 1160 -3316
rect 1120 -3396 1124 -3364
rect 1156 -3396 1160 -3364
rect 1120 -3444 1160 -3396
rect 1120 -3476 1124 -3444
rect 1156 -3476 1160 -3444
rect 1120 -3524 1160 -3476
rect 1120 -3556 1124 -3524
rect 1156 -3556 1160 -3524
rect 1120 -3604 1160 -3556
rect 1120 -3636 1124 -3604
rect 1156 -3636 1160 -3604
rect 1120 -3684 1160 -3636
rect 1120 -3716 1124 -3684
rect 1156 -3716 1160 -3684
rect 1120 -3720 1160 -3716
rect 1200 1036 1240 1040
rect 1200 1004 1204 1036
rect 1236 1004 1240 1036
rect 1200 956 1240 1004
rect 1200 924 1204 956
rect 1236 924 1240 956
rect 1200 876 1240 924
rect 1200 844 1204 876
rect 1236 844 1240 876
rect 1200 796 1240 844
rect 1200 764 1204 796
rect 1236 764 1240 796
rect 1200 716 1240 764
rect 1200 684 1204 716
rect 1236 684 1240 716
rect 1200 636 1240 684
rect 1200 604 1204 636
rect 1236 604 1240 636
rect 1200 556 1240 604
rect 1200 524 1204 556
rect 1236 524 1240 556
rect 1200 476 1240 524
rect 1200 444 1204 476
rect 1236 444 1240 476
rect 1200 396 1240 444
rect 1200 364 1204 396
rect 1236 364 1240 396
rect 1200 316 1240 364
rect 1200 284 1204 316
rect 1236 284 1240 316
rect 1200 236 1240 284
rect 1200 204 1204 236
rect 1236 204 1240 236
rect 1200 156 1240 204
rect 1200 124 1204 156
rect 1236 124 1240 156
rect 1200 76 1240 124
rect 1200 44 1204 76
rect 1236 44 1240 76
rect 1200 -4 1240 44
rect 1200 -36 1204 -4
rect 1236 -36 1240 -4
rect 1200 -84 1240 -36
rect 1200 -116 1204 -84
rect 1236 -116 1240 -84
rect 1200 -164 1240 -116
rect 1200 -196 1204 -164
rect 1236 -196 1240 -164
rect 1200 -244 1240 -196
rect 1200 -276 1204 -244
rect 1236 -276 1240 -244
rect 1200 -324 1240 -276
rect 1200 -356 1204 -324
rect 1236 -356 1240 -324
rect 1200 -404 1240 -356
rect 1200 -436 1204 -404
rect 1236 -436 1240 -404
rect 1200 -484 1240 -436
rect 1200 -516 1204 -484
rect 1236 -516 1240 -484
rect 1200 -564 1240 -516
rect 1200 -596 1204 -564
rect 1236 -596 1240 -564
rect 1200 -644 1240 -596
rect 1200 -676 1204 -644
rect 1236 -676 1240 -644
rect 1200 -724 1240 -676
rect 1200 -756 1204 -724
rect 1236 -756 1240 -724
rect 1200 -804 1240 -756
rect 1200 -836 1204 -804
rect 1236 -836 1240 -804
rect 1200 -884 1240 -836
rect 1200 -916 1204 -884
rect 1236 -916 1240 -884
rect 1200 -964 1240 -916
rect 1200 -996 1204 -964
rect 1236 -996 1240 -964
rect 1200 -1044 1240 -996
rect 1200 -1076 1204 -1044
rect 1236 -1076 1240 -1044
rect 1200 -1124 1240 -1076
rect 1200 -1156 1204 -1124
rect 1236 -1156 1240 -1124
rect 1200 -1204 1240 -1156
rect 1200 -1236 1204 -1204
rect 1236 -1236 1240 -1204
rect 1200 -1284 1240 -1236
rect 1200 -1316 1204 -1284
rect 1236 -1316 1240 -1284
rect 1200 -1364 1240 -1316
rect 1200 -1396 1204 -1364
rect 1236 -1396 1240 -1364
rect 1200 -1444 1240 -1396
rect 1200 -1476 1204 -1444
rect 1236 -1476 1240 -1444
rect 1200 -1524 1240 -1476
rect 1200 -1556 1204 -1524
rect 1236 -1556 1240 -1524
rect 1200 -1604 1240 -1556
rect 1200 -1636 1204 -1604
rect 1236 -1636 1240 -1604
rect 1200 -1684 1240 -1636
rect 1200 -1716 1204 -1684
rect 1236 -1716 1240 -1684
rect 1200 -1764 1240 -1716
rect 1200 -1796 1204 -1764
rect 1236 -1796 1240 -1764
rect 1200 -1844 1240 -1796
rect 1200 -1876 1204 -1844
rect 1236 -1876 1240 -1844
rect 1200 -1924 1240 -1876
rect 1200 -1956 1204 -1924
rect 1236 -1956 1240 -1924
rect 1200 -2004 1240 -1956
rect 1200 -2036 1204 -2004
rect 1236 -2036 1240 -2004
rect 1200 -2084 1240 -2036
rect 1200 -2116 1204 -2084
rect 1236 -2116 1240 -2084
rect 1200 -2164 1240 -2116
rect 1200 -2196 1204 -2164
rect 1236 -2196 1240 -2164
rect 1200 -2244 1240 -2196
rect 1200 -2276 1204 -2244
rect 1236 -2276 1240 -2244
rect 1200 -2324 1240 -2276
rect 1200 -2356 1204 -2324
rect 1236 -2356 1240 -2324
rect 1200 -2404 1240 -2356
rect 1200 -2436 1204 -2404
rect 1236 -2436 1240 -2404
rect 1200 -2484 1240 -2436
rect 1200 -2516 1204 -2484
rect 1236 -2516 1240 -2484
rect 1200 -2564 1240 -2516
rect 1200 -2596 1204 -2564
rect 1236 -2596 1240 -2564
rect 1200 -2644 1240 -2596
rect 1200 -2676 1204 -2644
rect 1236 -2676 1240 -2644
rect 1200 -2724 1240 -2676
rect 1200 -2756 1204 -2724
rect 1236 -2756 1240 -2724
rect 1200 -2804 1240 -2756
rect 1200 -2836 1204 -2804
rect 1236 -2836 1240 -2804
rect 1200 -2884 1240 -2836
rect 1200 -2916 1204 -2884
rect 1236 -2916 1240 -2884
rect 1200 -2964 1240 -2916
rect 1200 -2996 1204 -2964
rect 1236 -2996 1240 -2964
rect 1200 -3044 1240 -2996
rect 1200 -3076 1204 -3044
rect 1236 -3076 1240 -3044
rect 1200 -3124 1240 -3076
rect 1200 -3156 1204 -3124
rect 1236 -3156 1240 -3124
rect 1200 -3204 1240 -3156
rect 1200 -3236 1204 -3204
rect 1236 -3236 1240 -3204
rect 1200 -3284 1240 -3236
rect 1200 -3316 1204 -3284
rect 1236 -3316 1240 -3284
rect 1200 -3364 1240 -3316
rect 1200 -3396 1204 -3364
rect 1236 -3396 1240 -3364
rect 1200 -3444 1240 -3396
rect 1200 -3476 1204 -3444
rect 1236 -3476 1240 -3444
rect 1200 -3524 1240 -3476
rect 1200 -3556 1204 -3524
rect 1236 -3556 1240 -3524
rect 1200 -3604 1240 -3556
rect 1200 -3636 1204 -3604
rect 1236 -3636 1240 -3604
rect 1200 -3684 1240 -3636
rect 1200 -3716 1204 -3684
rect 1236 -3716 1240 -3684
rect 1200 -3720 1240 -3716
rect 1280 1036 1320 1040
rect 1280 1004 1284 1036
rect 1316 1004 1320 1036
rect 1280 956 1320 1004
rect 1280 924 1284 956
rect 1316 924 1320 956
rect 1280 876 1320 924
rect 1280 844 1284 876
rect 1316 844 1320 876
rect 1280 796 1320 844
rect 1280 764 1284 796
rect 1316 764 1320 796
rect 1280 716 1320 764
rect 1280 684 1284 716
rect 1316 684 1320 716
rect 1280 636 1320 684
rect 1280 604 1284 636
rect 1316 604 1320 636
rect 1280 556 1320 604
rect 1280 524 1284 556
rect 1316 524 1320 556
rect 1280 476 1320 524
rect 1280 444 1284 476
rect 1316 444 1320 476
rect 1280 396 1320 444
rect 1280 364 1284 396
rect 1316 364 1320 396
rect 1280 316 1320 364
rect 1280 284 1284 316
rect 1316 284 1320 316
rect 1280 236 1320 284
rect 1280 204 1284 236
rect 1316 204 1320 236
rect 1280 156 1320 204
rect 1280 124 1284 156
rect 1316 124 1320 156
rect 1280 76 1320 124
rect 1280 44 1284 76
rect 1316 44 1320 76
rect 1280 -4 1320 44
rect 1280 -36 1284 -4
rect 1316 -36 1320 -4
rect 1280 -84 1320 -36
rect 1280 -116 1284 -84
rect 1316 -116 1320 -84
rect 1280 -164 1320 -116
rect 1280 -196 1284 -164
rect 1316 -196 1320 -164
rect 1280 -244 1320 -196
rect 1280 -276 1284 -244
rect 1316 -276 1320 -244
rect 1280 -324 1320 -276
rect 1280 -356 1284 -324
rect 1316 -356 1320 -324
rect 1280 -404 1320 -356
rect 1280 -436 1284 -404
rect 1316 -436 1320 -404
rect 1280 -484 1320 -436
rect 1280 -516 1284 -484
rect 1316 -516 1320 -484
rect 1280 -564 1320 -516
rect 1280 -596 1284 -564
rect 1316 -596 1320 -564
rect 1280 -644 1320 -596
rect 1280 -676 1284 -644
rect 1316 -676 1320 -644
rect 1280 -724 1320 -676
rect 1280 -756 1284 -724
rect 1316 -756 1320 -724
rect 1280 -804 1320 -756
rect 1280 -836 1284 -804
rect 1316 -836 1320 -804
rect 1280 -884 1320 -836
rect 1280 -916 1284 -884
rect 1316 -916 1320 -884
rect 1280 -964 1320 -916
rect 1280 -996 1284 -964
rect 1316 -996 1320 -964
rect 1280 -1044 1320 -996
rect 1280 -1076 1284 -1044
rect 1316 -1076 1320 -1044
rect 1280 -1124 1320 -1076
rect 1280 -1156 1284 -1124
rect 1316 -1156 1320 -1124
rect 1280 -1204 1320 -1156
rect 1280 -1236 1284 -1204
rect 1316 -1236 1320 -1204
rect 1280 -1284 1320 -1236
rect 1280 -1316 1284 -1284
rect 1316 -1316 1320 -1284
rect 1280 -1364 1320 -1316
rect 1280 -1396 1284 -1364
rect 1316 -1396 1320 -1364
rect 1280 -1444 1320 -1396
rect 1280 -1476 1284 -1444
rect 1316 -1476 1320 -1444
rect 1280 -1524 1320 -1476
rect 1280 -1556 1284 -1524
rect 1316 -1556 1320 -1524
rect 1280 -1604 1320 -1556
rect 1280 -1636 1284 -1604
rect 1316 -1636 1320 -1604
rect 1280 -1684 1320 -1636
rect 1280 -1716 1284 -1684
rect 1316 -1716 1320 -1684
rect 1280 -1764 1320 -1716
rect 1280 -1796 1284 -1764
rect 1316 -1796 1320 -1764
rect 1280 -1844 1320 -1796
rect 1280 -1876 1284 -1844
rect 1316 -1876 1320 -1844
rect 1280 -1924 1320 -1876
rect 1280 -1956 1284 -1924
rect 1316 -1956 1320 -1924
rect 1280 -2004 1320 -1956
rect 1280 -2036 1284 -2004
rect 1316 -2036 1320 -2004
rect 1280 -2084 1320 -2036
rect 1280 -2116 1284 -2084
rect 1316 -2116 1320 -2084
rect 1280 -2164 1320 -2116
rect 1280 -2196 1284 -2164
rect 1316 -2196 1320 -2164
rect 1280 -2244 1320 -2196
rect 1280 -2276 1284 -2244
rect 1316 -2276 1320 -2244
rect 1280 -2324 1320 -2276
rect 1280 -2356 1284 -2324
rect 1316 -2356 1320 -2324
rect 1280 -2404 1320 -2356
rect 1280 -2436 1284 -2404
rect 1316 -2436 1320 -2404
rect 1280 -2484 1320 -2436
rect 1280 -2516 1284 -2484
rect 1316 -2516 1320 -2484
rect 1280 -2564 1320 -2516
rect 1280 -2596 1284 -2564
rect 1316 -2596 1320 -2564
rect 1280 -2644 1320 -2596
rect 1280 -2676 1284 -2644
rect 1316 -2676 1320 -2644
rect 1280 -2724 1320 -2676
rect 1280 -2756 1284 -2724
rect 1316 -2756 1320 -2724
rect 1280 -2804 1320 -2756
rect 1280 -2836 1284 -2804
rect 1316 -2836 1320 -2804
rect 1280 -2884 1320 -2836
rect 1280 -2916 1284 -2884
rect 1316 -2916 1320 -2884
rect 1280 -2964 1320 -2916
rect 1280 -2996 1284 -2964
rect 1316 -2996 1320 -2964
rect 1280 -3044 1320 -2996
rect 1280 -3076 1284 -3044
rect 1316 -3076 1320 -3044
rect 1280 -3124 1320 -3076
rect 1280 -3156 1284 -3124
rect 1316 -3156 1320 -3124
rect 1280 -3204 1320 -3156
rect 1280 -3236 1284 -3204
rect 1316 -3236 1320 -3204
rect 1280 -3284 1320 -3236
rect 1280 -3316 1284 -3284
rect 1316 -3316 1320 -3284
rect 1280 -3364 1320 -3316
rect 1280 -3396 1284 -3364
rect 1316 -3396 1320 -3364
rect 1280 -3444 1320 -3396
rect 1280 -3476 1284 -3444
rect 1316 -3476 1320 -3444
rect 1280 -3524 1320 -3476
rect 1280 -3556 1284 -3524
rect 1316 -3556 1320 -3524
rect 1280 -3604 1320 -3556
rect 1280 -3636 1284 -3604
rect 1316 -3636 1320 -3604
rect 1280 -3684 1320 -3636
rect 1280 -3716 1284 -3684
rect 1316 -3716 1320 -3684
rect 1280 -3720 1320 -3716
rect 1360 1036 1400 1040
rect 1360 1004 1364 1036
rect 1396 1004 1400 1036
rect 1360 956 1400 1004
rect 1360 924 1364 956
rect 1396 924 1400 956
rect 1360 876 1400 924
rect 1360 844 1364 876
rect 1396 844 1400 876
rect 1360 796 1400 844
rect 1360 764 1364 796
rect 1396 764 1400 796
rect 1360 716 1400 764
rect 1360 684 1364 716
rect 1396 684 1400 716
rect 1360 636 1400 684
rect 1360 604 1364 636
rect 1396 604 1400 636
rect 1360 556 1400 604
rect 1360 524 1364 556
rect 1396 524 1400 556
rect 1360 476 1400 524
rect 1360 444 1364 476
rect 1396 444 1400 476
rect 1360 396 1400 444
rect 1360 364 1364 396
rect 1396 364 1400 396
rect 1360 316 1400 364
rect 1360 284 1364 316
rect 1396 284 1400 316
rect 1360 236 1400 284
rect 1360 204 1364 236
rect 1396 204 1400 236
rect 1360 156 1400 204
rect 1360 124 1364 156
rect 1396 124 1400 156
rect 1360 76 1400 124
rect 1360 44 1364 76
rect 1396 44 1400 76
rect 1360 -4 1400 44
rect 1360 -36 1364 -4
rect 1396 -36 1400 -4
rect 1360 -84 1400 -36
rect 1360 -116 1364 -84
rect 1396 -116 1400 -84
rect 1360 -164 1400 -116
rect 1360 -196 1364 -164
rect 1396 -196 1400 -164
rect 1360 -244 1400 -196
rect 1360 -276 1364 -244
rect 1396 -276 1400 -244
rect 1360 -324 1400 -276
rect 1360 -356 1364 -324
rect 1396 -356 1400 -324
rect 1360 -404 1400 -356
rect 1360 -436 1364 -404
rect 1396 -436 1400 -404
rect 1360 -484 1400 -436
rect 1360 -516 1364 -484
rect 1396 -516 1400 -484
rect 1360 -564 1400 -516
rect 1360 -596 1364 -564
rect 1396 -596 1400 -564
rect 1360 -644 1400 -596
rect 1360 -676 1364 -644
rect 1396 -676 1400 -644
rect 1360 -724 1400 -676
rect 1360 -756 1364 -724
rect 1396 -756 1400 -724
rect 1360 -804 1400 -756
rect 1360 -836 1364 -804
rect 1396 -836 1400 -804
rect 1360 -884 1400 -836
rect 1360 -916 1364 -884
rect 1396 -916 1400 -884
rect 1360 -964 1400 -916
rect 1360 -996 1364 -964
rect 1396 -996 1400 -964
rect 1360 -1044 1400 -996
rect 1360 -1076 1364 -1044
rect 1396 -1076 1400 -1044
rect 1360 -1124 1400 -1076
rect 1360 -1156 1364 -1124
rect 1396 -1156 1400 -1124
rect 1360 -1204 1400 -1156
rect 1360 -1236 1364 -1204
rect 1396 -1236 1400 -1204
rect 1360 -1284 1400 -1236
rect 1360 -1316 1364 -1284
rect 1396 -1316 1400 -1284
rect 1360 -1364 1400 -1316
rect 1360 -1396 1364 -1364
rect 1396 -1396 1400 -1364
rect 1360 -1444 1400 -1396
rect 1360 -1476 1364 -1444
rect 1396 -1476 1400 -1444
rect 1360 -1524 1400 -1476
rect 1360 -1556 1364 -1524
rect 1396 -1556 1400 -1524
rect 1360 -1604 1400 -1556
rect 1360 -1636 1364 -1604
rect 1396 -1636 1400 -1604
rect 1360 -1684 1400 -1636
rect 1360 -1716 1364 -1684
rect 1396 -1716 1400 -1684
rect 1360 -1764 1400 -1716
rect 1360 -1796 1364 -1764
rect 1396 -1796 1400 -1764
rect 1360 -1844 1400 -1796
rect 1360 -1876 1364 -1844
rect 1396 -1876 1400 -1844
rect 1360 -1924 1400 -1876
rect 1360 -1956 1364 -1924
rect 1396 -1956 1400 -1924
rect 1360 -2004 1400 -1956
rect 1360 -2036 1364 -2004
rect 1396 -2036 1400 -2004
rect 1360 -2084 1400 -2036
rect 1360 -2116 1364 -2084
rect 1396 -2116 1400 -2084
rect 1360 -2164 1400 -2116
rect 1360 -2196 1364 -2164
rect 1396 -2196 1400 -2164
rect 1360 -2244 1400 -2196
rect 1360 -2276 1364 -2244
rect 1396 -2276 1400 -2244
rect 1360 -2324 1400 -2276
rect 1360 -2356 1364 -2324
rect 1396 -2356 1400 -2324
rect 1360 -2404 1400 -2356
rect 1360 -2436 1364 -2404
rect 1396 -2436 1400 -2404
rect 1360 -2484 1400 -2436
rect 1360 -2516 1364 -2484
rect 1396 -2516 1400 -2484
rect 1360 -2564 1400 -2516
rect 1360 -2596 1364 -2564
rect 1396 -2596 1400 -2564
rect 1360 -2644 1400 -2596
rect 1360 -2676 1364 -2644
rect 1396 -2676 1400 -2644
rect 1360 -2724 1400 -2676
rect 1360 -2756 1364 -2724
rect 1396 -2756 1400 -2724
rect 1360 -2804 1400 -2756
rect 1360 -2836 1364 -2804
rect 1396 -2836 1400 -2804
rect 1360 -2884 1400 -2836
rect 1360 -2916 1364 -2884
rect 1396 -2916 1400 -2884
rect 1360 -2964 1400 -2916
rect 1360 -2996 1364 -2964
rect 1396 -2996 1400 -2964
rect 1360 -3044 1400 -2996
rect 1360 -3076 1364 -3044
rect 1396 -3076 1400 -3044
rect 1360 -3124 1400 -3076
rect 1360 -3156 1364 -3124
rect 1396 -3156 1400 -3124
rect 1360 -3204 1400 -3156
rect 1360 -3236 1364 -3204
rect 1396 -3236 1400 -3204
rect 1360 -3284 1400 -3236
rect 1360 -3316 1364 -3284
rect 1396 -3316 1400 -3284
rect 1360 -3364 1400 -3316
rect 1360 -3396 1364 -3364
rect 1396 -3396 1400 -3364
rect 1360 -3444 1400 -3396
rect 1360 -3476 1364 -3444
rect 1396 -3476 1400 -3444
rect 1360 -3524 1400 -3476
rect 1360 -3556 1364 -3524
rect 1396 -3556 1400 -3524
rect 1360 -3604 1400 -3556
rect 1360 -3636 1364 -3604
rect 1396 -3636 1400 -3604
rect 1360 -3684 1400 -3636
rect 1360 -3716 1364 -3684
rect 1396 -3716 1400 -3684
rect 1360 -3720 1400 -3716
rect 1440 1036 1480 1040
rect 1440 1004 1444 1036
rect 1476 1004 1480 1036
rect 1440 956 1480 1004
rect 1440 924 1444 956
rect 1476 924 1480 956
rect 1440 876 1480 924
rect 1440 844 1444 876
rect 1476 844 1480 876
rect 1440 796 1480 844
rect 1440 764 1444 796
rect 1476 764 1480 796
rect 1440 716 1480 764
rect 1440 684 1444 716
rect 1476 684 1480 716
rect 1440 636 1480 684
rect 1440 604 1444 636
rect 1476 604 1480 636
rect 1440 556 1480 604
rect 1440 524 1444 556
rect 1476 524 1480 556
rect 1440 476 1480 524
rect 1440 444 1444 476
rect 1476 444 1480 476
rect 1440 396 1480 444
rect 1440 364 1444 396
rect 1476 364 1480 396
rect 1440 316 1480 364
rect 1440 284 1444 316
rect 1476 284 1480 316
rect 1440 236 1480 284
rect 1440 204 1444 236
rect 1476 204 1480 236
rect 1440 156 1480 204
rect 1440 124 1444 156
rect 1476 124 1480 156
rect 1440 76 1480 124
rect 1440 44 1444 76
rect 1476 44 1480 76
rect 1440 -4 1480 44
rect 1440 -36 1444 -4
rect 1476 -36 1480 -4
rect 1440 -84 1480 -36
rect 1440 -116 1444 -84
rect 1476 -116 1480 -84
rect 1440 -164 1480 -116
rect 1440 -196 1444 -164
rect 1476 -196 1480 -164
rect 1440 -244 1480 -196
rect 1440 -276 1444 -244
rect 1476 -276 1480 -244
rect 1440 -324 1480 -276
rect 1440 -356 1444 -324
rect 1476 -356 1480 -324
rect 1440 -404 1480 -356
rect 1440 -436 1444 -404
rect 1476 -436 1480 -404
rect 1440 -484 1480 -436
rect 1440 -516 1444 -484
rect 1476 -516 1480 -484
rect 1440 -564 1480 -516
rect 1440 -596 1444 -564
rect 1476 -596 1480 -564
rect 1440 -644 1480 -596
rect 1440 -676 1444 -644
rect 1476 -676 1480 -644
rect 1440 -724 1480 -676
rect 1440 -756 1444 -724
rect 1476 -756 1480 -724
rect 1440 -804 1480 -756
rect 1440 -836 1444 -804
rect 1476 -836 1480 -804
rect 1440 -884 1480 -836
rect 1440 -916 1444 -884
rect 1476 -916 1480 -884
rect 1440 -964 1480 -916
rect 1440 -996 1444 -964
rect 1476 -996 1480 -964
rect 1440 -1044 1480 -996
rect 1440 -1076 1444 -1044
rect 1476 -1076 1480 -1044
rect 1440 -1124 1480 -1076
rect 1440 -1156 1444 -1124
rect 1476 -1156 1480 -1124
rect 1440 -1204 1480 -1156
rect 1440 -1236 1444 -1204
rect 1476 -1236 1480 -1204
rect 1440 -1284 1480 -1236
rect 1440 -1316 1444 -1284
rect 1476 -1316 1480 -1284
rect 1440 -1364 1480 -1316
rect 1440 -1396 1444 -1364
rect 1476 -1396 1480 -1364
rect 1440 -1444 1480 -1396
rect 1440 -1476 1444 -1444
rect 1476 -1476 1480 -1444
rect 1440 -1524 1480 -1476
rect 1440 -1556 1444 -1524
rect 1476 -1556 1480 -1524
rect 1440 -1604 1480 -1556
rect 1440 -1636 1444 -1604
rect 1476 -1636 1480 -1604
rect 1440 -1684 1480 -1636
rect 1440 -1716 1444 -1684
rect 1476 -1716 1480 -1684
rect 1440 -1764 1480 -1716
rect 1440 -1796 1444 -1764
rect 1476 -1796 1480 -1764
rect 1440 -1844 1480 -1796
rect 1440 -1876 1444 -1844
rect 1476 -1876 1480 -1844
rect 1440 -1924 1480 -1876
rect 1440 -1956 1444 -1924
rect 1476 -1956 1480 -1924
rect 1440 -2004 1480 -1956
rect 1440 -2036 1444 -2004
rect 1476 -2036 1480 -2004
rect 1440 -2084 1480 -2036
rect 1440 -2116 1444 -2084
rect 1476 -2116 1480 -2084
rect 1440 -2164 1480 -2116
rect 1440 -2196 1444 -2164
rect 1476 -2196 1480 -2164
rect 1440 -2244 1480 -2196
rect 1440 -2276 1444 -2244
rect 1476 -2276 1480 -2244
rect 1440 -2324 1480 -2276
rect 1440 -2356 1444 -2324
rect 1476 -2356 1480 -2324
rect 1440 -2404 1480 -2356
rect 1440 -2436 1444 -2404
rect 1476 -2436 1480 -2404
rect 1440 -2484 1480 -2436
rect 1440 -2516 1444 -2484
rect 1476 -2516 1480 -2484
rect 1440 -2564 1480 -2516
rect 1440 -2596 1444 -2564
rect 1476 -2596 1480 -2564
rect 1440 -2644 1480 -2596
rect 1440 -2676 1444 -2644
rect 1476 -2676 1480 -2644
rect 1440 -2724 1480 -2676
rect 1440 -2756 1444 -2724
rect 1476 -2756 1480 -2724
rect 1440 -2804 1480 -2756
rect 1440 -2836 1444 -2804
rect 1476 -2836 1480 -2804
rect 1440 -2884 1480 -2836
rect 1440 -2916 1444 -2884
rect 1476 -2916 1480 -2884
rect 1440 -2964 1480 -2916
rect 1440 -2996 1444 -2964
rect 1476 -2996 1480 -2964
rect 1440 -3044 1480 -2996
rect 1440 -3076 1444 -3044
rect 1476 -3076 1480 -3044
rect 1440 -3124 1480 -3076
rect 1440 -3156 1444 -3124
rect 1476 -3156 1480 -3124
rect 1440 -3204 1480 -3156
rect 1440 -3236 1444 -3204
rect 1476 -3236 1480 -3204
rect 1440 -3284 1480 -3236
rect 1440 -3316 1444 -3284
rect 1476 -3316 1480 -3284
rect 1440 -3364 1480 -3316
rect 1440 -3396 1444 -3364
rect 1476 -3396 1480 -3364
rect 1440 -3444 1480 -3396
rect 1440 -3476 1444 -3444
rect 1476 -3476 1480 -3444
rect 1440 -3524 1480 -3476
rect 1440 -3556 1444 -3524
rect 1476 -3556 1480 -3524
rect 1440 -3604 1480 -3556
rect 1440 -3636 1444 -3604
rect 1476 -3636 1480 -3604
rect 1440 -3684 1480 -3636
rect 1440 -3716 1444 -3684
rect 1476 -3716 1480 -3684
rect 1440 -3720 1480 -3716
rect 1520 1036 1560 1040
rect 1520 1004 1524 1036
rect 1556 1004 1560 1036
rect 1520 956 1560 1004
rect 1520 924 1524 956
rect 1556 924 1560 956
rect 1520 876 1560 924
rect 1520 844 1524 876
rect 1556 844 1560 876
rect 1520 796 1560 844
rect 1520 764 1524 796
rect 1556 764 1560 796
rect 1520 716 1560 764
rect 1520 684 1524 716
rect 1556 684 1560 716
rect 1520 636 1560 684
rect 1520 604 1524 636
rect 1556 604 1560 636
rect 1520 556 1560 604
rect 1520 524 1524 556
rect 1556 524 1560 556
rect 1520 476 1560 524
rect 1520 444 1524 476
rect 1556 444 1560 476
rect 1520 396 1560 444
rect 1520 364 1524 396
rect 1556 364 1560 396
rect 1520 316 1560 364
rect 1520 284 1524 316
rect 1556 284 1560 316
rect 1520 236 1560 284
rect 1520 204 1524 236
rect 1556 204 1560 236
rect 1520 156 1560 204
rect 1520 124 1524 156
rect 1556 124 1560 156
rect 1520 76 1560 124
rect 1520 44 1524 76
rect 1556 44 1560 76
rect 1520 -4 1560 44
rect 1520 -36 1524 -4
rect 1556 -36 1560 -4
rect 1520 -84 1560 -36
rect 1520 -116 1524 -84
rect 1556 -116 1560 -84
rect 1520 -164 1560 -116
rect 1520 -196 1524 -164
rect 1556 -196 1560 -164
rect 1520 -244 1560 -196
rect 1520 -276 1524 -244
rect 1556 -276 1560 -244
rect 1520 -324 1560 -276
rect 1520 -356 1524 -324
rect 1556 -356 1560 -324
rect 1520 -404 1560 -356
rect 1520 -436 1524 -404
rect 1556 -436 1560 -404
rect 1520 -484 1560 -436
rect 1520 -516 1524 -484
rect 1556 -516 1560 -484
rect 1520 -564 1560 -516
rect 1520 -596 1524 -564
rect 1556 -596 1560 -564
rect 1520 -644 1560 -596
rect 1520 -676 1524 -644
rect 1556 -676 1560 -644
rect 1520 -724 1560 -676
rect 1520 -756 1524 -724
rect 1556 -756 1560 -724
rect 1520 -804 1560 -756
rect 1520 -836 1524 -804
rect 1556 -836 1560 -804
rect 1520 -884 1560 -836
rect 1520 -916 1524 -884
rect 1556 -916 1560 -884
rect 1520 -964 1560 -916
rect 1520 -996 1524 -964
rect 1556 -996 1560 -964
rect 1520 -1044 1560 -996
rect 1520 -1076 1524 -1044
rect 1556 -1076 1560 -1044
rect 1520 -1124 1560 -1076
rect 1520 -1156 1524 -1124
rect 1556 -1156 1560 -1124
rect 1520 -1204 1560 -1156
rect 1520 -1236 1524 -1204
rect 1556 -1236 1560 -1204
rect 1520 -1284 1560 -1236
rect 1520 -1316 1524 -1284
rect 1556 -1316 1560 -1284
rect 1520 -1364 1560 -1316
rect 1520 -1396 1524 -1364
rect 1556 -1396 1560 -1364
rect 1520 -1444 1560 -1396
rect 1520 -1476 1524 -1444
rect 1556 -1476 1560 -1444
rect 1520 -1524 1560 -1476
rect 1520 -1556 1524 -1524
rect 1556 -1556 1560 -1524
rect 1520 -1604 1560 -1556
rect 1520 -1636 1524 -1604
rect 1556 -1636 1560 -1604
rect 1520 -1684 1560 -1636
rect 1520 -1716 1524 -1684
rect 1556 -1716 1560 -1684
rect 1520 -1764 1560 -1716
rect 1520 -1796 1524 -1764
rect 1556 -1796 1560 -1764
rect 1520 -1844 1560 -1796
rect 1520 -1876 1524 -1844
rect 1556 -1876 1560 -1844
rect 1520 -1924 1560 -1876
rect 1520 -1956 1524 -1924
rect 1556 -1956 1560 -1924
rect 1520 -2004 1560 -1956
rect 1520 -2036 1524 -2004
rect 1556 -2036 1560 -2004
rect 1520 -2084 1560 -2036
rect 1520 -2116 1524 -2084
rect 1556 -2116 1560 -2084
rect 1520 -2164 1560 -2116
rect 1520 -2196 1524 -2164
rect 1556 -2196 1560 -2164
rect 1520 -2244 1560 -2196
rect 1520 -2276 1524 -2244
rect 1556 -2276 1560 -2244
rect 1520 -2324 1560 -2276
rect 1520 -2356 1524 -2324
rect 1556 -2356 1560 -2324
rect 1520 -2404 1560 -2356
rect 1520 -2436 1524 -2404
rect 1556 -2436 1560 -2404
rect 1520 -2484 1560 -2436
rect 1520 -2516 1524 -2484
rect 1556 -2516 1560 -2484
rect 1520 -2564 1560 -2516
rect 1520 -2596 1524 -2564
rect 1556 -2596 1560 -2564
rect 1520 -2644 1560 -2596
rect 1520 -2676 1524 -2644
rect 1556 -2676 1560 -2644
rect 1520 -2724 1560 -2676
rect 1520 -2756 1524 -2724
rect 1556 -2756 1560 -2724
rect 1520 -2804 1560 -2756
rect 1520 -2836 1524 -2804
rect 1556 -2836 1560 -2804
rect 1520 -2884 1560 -2836
rect 1520 -2916 1524 -2884
rect 1556 -2916 1560 -2884
rect 1520 -2964 1560 -2916
rect 1520 -2996 1524 -2964
rect 1556 -2996 1560 -2964
rect 1520 -3044 1560 -2996
rect 1520 -3076 1524 -3044
rect 1556 -3076 1560 -3044
rect 1520 -3124 1560 -3076
rect 1520 -3156 1524 -3124
rect 1556 -3156 1560 -3124
rect 1520 -3204 1560 -3156
rect 1520 -3236 1524 -3204
rect 1556 -3236 1560 -3204
rect 1520 -3284 1560 -3236
rect 1520 -3316 1524 -3284
rect 1556 -3316 1560 -3284
rect 1520 -3364 1560 -3316
rect 1520 -3396 1524 -3364
rect 1556 -3396 1560 -3364
rect 1520 -3444 1560 -3396
rect 1520 -3476 1524 -3444
rect 1556 -3476 1560 -3444
rect 1520 -3524 1560 -3476
rect 1520 -3556 1524 -3524
rect 1556 -3556 1560 -3524
rect 1520 -3604 1560 -3556
rect 1520 -3636 1524 -3604
rect 1556 -3636 1560 -3604
rect 1520 -3684 1560 -3636
rect 1520 -3716 1524 -3684
rect 1556 -3716 1560 -3684
rect 1520 -3720 1560 -3716
rect 1600 1036 1640 1040
rect 1600 1004 1604 1036
rect 1636 1004 1640 1036
rect 1600 956 1640 1004
rect 1600 924 1604 956
rect 1636 924 1640 956
rect 1600 876 1640 924
rect 1600 844 1604 876
rect 1636 844 1640 876
rect 1600 796 1640 844
rect 1600 764 1604 796
rect 1636 764 1640 796
rect 1600 716 1640 764
rect 1600 684 1604 716
rect 1636 684 1640 716
rect 1600 636 1640 684
rect 1600 604 1604 636
rect 1636 604 1640 636
rect 1600 556 1640 604
rect 1600 524 1604 556
rect 1636 524 1640 556
rect 1600 476 1640 524
rect 1600 444 1604 476
rect 1636 444 1640 476
rect 1600 396 1640 444
rect 1600 364 1604 396
rect 1636 364 1640 396
rect 1600 316 1640 364
rect 1600 284 1604 316
rect 1636 284 1640 316
rect 1600 236 1640 284
rect 1600 204 1604 236
rect 1636 204 1640 236
rect 1600 156 1640 204
rect 1600 124 1604 156
rect 1636 124 1640 156
rect 1600 76 1640 124
rect 1600 44 1604 76
rect 1636 44 1640 76
rect 1600 -4 1640 44
rect 1600 -36 1604 -4
rect 1636 -36 1640 -4
rect 1600 -84 1640 -36
rect 1600 -116 1604 -84
rect 1636 -116 1640 -84
rect 1600 -164 1640 -116
rect 1600 -196 1604 -164
rect 1636 -196 1640 -164
rect 1600 -244 1640 -196
rect 1600 -276 1604 -244
rect 1636 -276 1640 -244
rect 1600 -324 1640 -276
rect 1600 -356 1604 -324
rect 1636 -356 1640 -324
rect 1600 -404 1640 -356
rect 1600 -436 1604 -404
rect 1636 -436 1640 -404
rect 1600 -484 1640 -436
rect 1600 -516 1604 -484
rect 1636 -516 1640 -484
rect 1600 -564 1640 -516
rect 1600 -596 1604 -564
rect 1636 -596 1640 -564
rect 1600 -644 1640 -596
rect 1600 -676 1604 -644
rect 1636 -676 1640 -644
rect 1600 -724 1640 -676
rect 1600 -756 1604 -724
rect 1636 -756 1640 -724
rect 1600 -804 1640 -756
rect 1600 -836 1604 -804
rect 1636 -836 1640 -804
rect 1600 -884 1640 -836
rect 1600 -916 1604 -884
rect 1636 -916 1640 -884
rect 1600 -964 1640 -916
rect 1600 -996 1604 -964
rect 1636 -996 1640 -964
rect 1600 -1044 1640 -996
rect 1600 -1076 1604 -1044
rect 1636 -1076 1640 -1044
rect 1600 -1124 1640 -1076
rect 1600 -1156 1604 -1124
rect 1636 -1156 1640 -1124
rect 1600 -1204 1640 -1156
rect 1600 -1236 1604 -1204
rect 1636 -1236 1640 -1204
rect 1600 -1284 1640 -1236
rect 1600 -1316 1604 -1284
rect 1636 -1316 1640 -1284
rect 1600 -1364 1640 -1316
rect 1600 -1396 1604 -1364
rect 1636 -1396 1640 -1364
rect 1600 -1444 1640 -1396
rect 1600 -1476 1604 -1444
rect 1636 -1476 1640 -1444
rect 1600 -1524 1640 -1476
rect 1600 -1556 1604 -1524
rect 1636 -1556 1640 -1524
rect 1600 -1604 1640 -1556
rect 1600 -1636 1604 -1604
rect 1636 -1636 1640 -1604
rect 1600 -1684 1640 -1636
rect 1600 -1716 1604 -1684
rect 1636 -1716 1640 -1684
rect 1600 -1764 1640 -1716
rect 1600 -1796 1604 -1764
rect 1636 -1796 1640 -1764
rect 1600 -1844 1640 -1796
rect 1600 -1876 1604 -1844
rect 1636 -1876 1640 -1844
rect 1600 -1924 1640 -1876
rect 1600 -1956 1604 -1924
rect 1636 -1956 1640 -1924
rect 1600 -2004 1640 -1956
rect 1600 -2036 1604 -2004
rect 1636 -2036 1640 -2004
rect 1600 -2084 1640 -2036
rect 1600 -2116 1604 -2084
rect 1636 -2116 1640 -2084
rect 1600 -2164 1640 -2116
rect 1600 -2196 1604 -2164
rect 1636 -2196 1640 -2164
rect 1600 -2244 1640 -2196
rect 1600 -2276 1604 -2244
rect 1636 -2276 1640 -2244
rect 1600 -2324 1640 -2276
rect 1600 -2356 1604 -2324
rect 1636 -2356 1640 -2324
rect 1600 -2404 1640 -2356
rect 1600 -2436 1604 -2404
rect 1636 -2436 1640 -2404
rect 1600 -2484 1640 -2436
rect 1600 -2516 1604 -2484
rect 1636 -2516 1640 -2484
rect 1600 -2564 1640 -2516
rect 1600 -2596 1604 -2564
rect 1636 -2596 1640 -2564
rect 1600 -2644 1640 -2596
rect 1600 -2676 1604 -2644
rect 1636 -2676 1640 -2644
rect 1600 -2724 1640 -2676
rect 1600 -2756 1604 -2724
rect 1636 -2756 1640 -2724
rect 1600 -2804 1640 -2756
rect 1600 -2836 1604 -2804
rect 1636 -2836 1640 -2804
rect 1600 -2884 1640 -2836
rect 1600 -2916 1604 -2884
rect 1636 -2916 1640 -2884
rect 1600 -2964 1640 -2916
rect 1600 -2996 1604 -2964
rect 1636 -2996 1640 -2964
rect 1600 -3044 1640 -2996
rect 1600 -3076 1604 -3044
rect 1636 -3076 1640 -3044
rect 1600 -3124 1640 -3076
rect 1600 -3156 1604 -3124
rect 1636 -3156 1640 -3124
rect 1600 -3204 1640 -3156
rect 1600 -3236 1604 -3204
rect 1636 -3236 1640 -3204
rect 1600 -3284 1640 -3236
rect 1600 -3316 1604 -3284
rect 1636 -3316 1640 -3284
rect 1600 -3364 1640 -3316
rect 1600 -3396 1604 -3364
rect 1636 -3396 1640 -3364
rect 1600 -3444 1640 -3396
rect 1600 -3476 1604 -3444
rect 1636 -3476 1640 -3444
rect 1600 -3524 1640 -3476
rect 1600 -3556 1604 -3524
rect 1636 -3556 1640 -3524
rect 1600 -3604 1640 -3556
rect 1600 -3636 1604 -3604
rect 1636 -3636 1640 -3604
rect 1600 -3684 1640 -3636
rect 1600 -3716 1604 -3684
rect 1636 -3716 1640 -3684
rect 1600 -3720 1640 -3716
rect 1680 1036 1720 1040
rect 1680 1004 1684 1036
rect 1716 1004 1720 1036
rect 1680 956 1720 1004
rect 1680 924 1684 956
rect 1716 924 1720 956
rect 1680 876 1720 924
rect 1680 844 1684 876
rect 1716 844 1720 876
rect 1680 796 1720 844
rect 1680 764 1684 796
rect 1716 764 1720 796
rect 1680 716 1720 764
rect 1680 684 1684 716
rect 1716 684 1720 716
rect 1680 636 1720 684
rect 1680 604 1684 636
rect 1716 604 1720 636
rect 1680 556 1720 604
rect 1680 524 1684 556
rect 1716 524 1720 556
rect 1680 476 1720 524
rect 1680 444 1684 476
rect 1716 444 1720 476
rect 1680 396 1720 444
rect 1680 364 1684 396
rect 1716 364 1720 396
rect 1680 316 1720 364
rect 1680 284 1684 316
rect 1716 284 1720 316
rect 1680 236 1720 284
rect 1680 204 1684 236
rect 1716 204 1720 236
rect 1680 156 1720 204
rect 1680 124 1684 156
rect 1716 124 1720 156
rect 1680 76 1720 124
rect 1680 44 1684 76
rect 1716 44 1720 76
rect 1680 -4 1720 44
rect 1680 -36 1684 -4
rect 1716 -36 1720 -4
rect 1680 -84 1720 -36
rect 1680 -116 1684 -84
rect 1716 -116 1720 -84
rect 1680 -164 1720 -116
rect 1680 -196 1684 -164
rect 1716 -196 1720 -164
rect 1680 -244 1720 -196
rect 1680 -276 1684 -244
rect 1716 -276 1720 -244
rect 1680 -324 1720 -276
rect 1680 -356 1684 -324
rect 1716 -356 1720 -324
rect 1680 -404 1720 -356
rect 1680 -436 1684 -404
rect 1716 -436 1720 -404
rect 1680 -484 1720 -436
rect 1680 -516 1684 -484
rect 1716 -516 1720 -484
rect 1680 -564 1720 -516
rect 1680 -596 1684 -564
rect 1716 -596 1720 -564
rect 1680 -644 1720 -596
rect 1680 -676 1684 -644
rect 1716 -676 1720 -644
rect 1680 -724 1720 -676
rect 1680 -756 1684 -724
rect 1716 -756 1720 -724
rect 1680 -804 1720 -756
rect 1680 -836 1684 -804
rect 1716 -836 1720 -804
rect 1680 -884 1720 -836
rect 1680 -916 1684 -884
rect 1716 -916 1720 -884
rect 1680 -964 1720 -916
rect 1680 -996 1684 -964
rect 1716 -996 1720 -964
rect 1680 -1044 1720 -996
rect 1680 -1076 1684 -1044
rect 1716 -1076 1720 -1044
rect 1680 -1124 1720 -1076
rect 1680 -1156 1684 -1124
rect 1716 -1156 1720 -1124
rect 1680 -1204 1720 -1156
rect 1680 -1236 1684 -1204
rect 1716 -1236 1720 -1204
rect 1680 -1284 1720 -1236
rect 1680 -1316 1684 -1284
rect 1716 -1316 1720 -1284
rect 1680 -1364 1720 -1316
rect 1680 -1396 1684 -1364
rect 1716 -1396 1720 -1364
rect 1680 -1444 1720 -1396
rect 1680 -1476 1684 -1444
rect 1716 -1476 1720 -1444
rect 1680 -1524 1720 -1476
rect 1680 -1556 1684 -1524
rect 1716 -1556 1720 -1524
rect 1680 -1604 1720 -1556
rect 1680 -1636 1684 -1604
rect 1716 -1636 1720 -1604
rect 1680 -1684 1720 -1636
rect 1680 -1716 1684 -1684
rect 1716 -1716 1720 -1684
rect 1680 -1764 1720 -1716
rect 1680 -1796 1684 -1764
rect 1716 -1796 1720 -1764
rect 1680 -1844 1720 -1796
rect 1680 -1876 1684 -1844
rect 1716 -1876 1720 -1844
rect 1680 -1924 1720 -1876
rect 1680 -1956 1684 -1924
rect 1716 -1956 1720 -1924
rect 1680 -2004 1720 -1956
rect 1680 -2036 1684 -2004
rect 1716 -2036 1720 -2004
rect 1680 -2084 1720 -2036
rect 1680 -2116 1684 -2084
rect 1716 -2116 1720 -2084
rect 1680 -2164 1720 -2116
rect 1680 -2196 1684 -2164
rect 1716 -2196 1720 -2164
rect 1680 -2244 1720 -2196
rect 1680 -2276 1684 -2244
rect 1716 -2276 1720 -2244
rect 1680 -2324 1720 -2276
rect 1680 -2356 1684 -2324
rect 1716 -2356 1720 -2324
rect 1680 -2404 1720 -2356
rect 1680 -2436 1684 -2404
rect 1716 -2436 1720 -2404
rect 1680 -2484 1720 -2436
rect 1680 -2516 1684 -2484
rect 1716 -2516 1720 -2484
rect 1680 -2564 1720 -2516
rect 1680 -2596 1684 -2564
rect 1716 -2596 1720 -2564
rect 1680 -2644 1720 -2596
rect 1680 -2676 1684 -2644
rect 1716 -2676 1720 -2644
rect 1680 -2724 1720 -2676
rect 1680 -2756 1684 -2724
rect 1716 -2756 1720 -2724
rect 1680 -2804 1720 -2756
rect 1680 -2836 1684 -2804
rect 1716 -2836 1720 -2804
rect 1680 -2884 1720 -2836
rect 1680 -2916 1684 -2884
rect 1716 -2916 1720 -2884
rect 1680 -2964 1720 -2916
rect 1680 -2996 1684 -2964
rect 1716 -2996 1720 -2964
rect 1680 -3044 1720 -2996
rect 1680 -3076 1684 -3044
rect 1716 -3076 1720 -3044
rect 1680 -3124 1720 -3076
rect 1680 -3156 1684 -3124
rect 1716 -3156 1720 -3124
rect 1680 -3204 1720 -3156
rect 1680 -3236 1684 -3204
rect 1716 -3236 1720 -3204
rect 1680 -3284 1720 -3236
rect 1680 -3316 1684 -3284
rect 1716 -3316 1720 -3284
rect 1680 -3364 1720 -3316
rect 1680 -3396 1684 -3364
rect 1716 -3396 1720 -3364
rect 1680 -3444 1720 -3396
rect 1680 -3476 1684 -3444
rect 1716 -3476 1720 -3444
rect 1680 -3524 1720 -3476
rect 1680 -3556 1684 -3524
rect 1716 -3556 1720 -3524
rect 1680 -3604 1720 -3556
rect 1680 -3636 1684 -3604
rect 1716 -3636 1720 -3604
rect 1680 -3684 1720 -3636
rect 1680 -3716 1684 -3684
rect 1716 -3716 1720 -3684
rect 1680 -3720 1720 -3716
rect 1760 1036 1800 1040
rect 1760 1004 1764 1036
rect 1796 1004 1800 1036
rect 1760 956 1800 1004
rect 1760 924 1764 956
rect 1796 924 1800 956
rect 1760 876 1800 924
rect 1760 844 1764 876
rect 1796 844 1800 876
rect 1760 796 1800 844
rect 1760 764 1764 796
rect 1796 764 1800 796
rect 1760 716 1800 764
rect 1760 684 1764 716
rect 1796 684 1800 716
rect 1760 636 1800 684
rect 1760 604 1764 636
rect 1796 604 1800 636
rect 1760 556 1800 604
rect 1760 524 1764 556
rect 1796 524 1800 556
rect 1760 476 1800 524
rect 1760 444 1764 476
rect 1796 444 1800 476
rect 1760 396 1800 444
rect 1760 364 1764 396
rect 1796 364 1800 396
rect 1760 316 1800 364
rect 1760 284 1764 316
rect 1796 284 1800 316
rect 1760 236 1800 284
rect 1760 204 1764 236
rect 1796 204 1800 236
rect 1760 156 1800 204
rect 1760 124 1764 156
rect 1796 124 1800 156
rect 1760 76 1800 124
rect 1760 44 1764 76
rect 1796 44 1800 76
rect 1760 -4 1800 44
rect 1760 -36 1764 -4
rect 1796 -36 1800 -4
rect 1760 -84 1800 -36
rect 1760 -116 1764 -84
rect 1796 -116 1800 -84
rect 1760 -164 1800 -116
rect 1760 -196 1764 -164
rect 1796 -196 1800 -164
rect 1760 -244 1800 -196
rect 1760 -276 1764 -244
rect 1796 -276 1800 -244
rect 1760 -324 1800 -276
rect 1760 -356 1764 -324
rect 1796 -356 1800 -324
rect 1760 -404 1800 -356
rect 1760 -436 1764 -404
rect 1796 -436 1800 -404
rect 1760 -484 1800 -436
rect 1760 -516 1764 -484
rect 1796 -516 1800 -484
rect 1760 -564 1800 -516
rect 1760 -596 1764 -564
rect 1796 -596 1800 -564
rect 1760 -644 1800 -596
rect 1760 -676 1764 -644
rect 1796 -676 1800 -644
rect 1760 -724 1800 -676
rect 1760 -756 1764 -724
rect 1796 -756 1800 -724
rect 1760 -804 1800 -756
rect 1760 -836 1764 -804
rect 1796 -836 1800 -804
rect 1760 -884 1800 -836
rect 1760 -916 1764 -884
rect 1796 -916 1800 -884
rect 1760 -964 1800 -916
rect 1760 -996 1764 -964
rect 1796 -996 1800 -964
rect 1760 -1044 1800 -996
rect 1760 -1076 1764 -1044
rect 1796 -1076 1800 -1044
rect 1760 -1124 1800 -1076
rect 1760 -1156 1764 -1124
rect 1796 -1156 1800 -1124
rect 1760 -1204 1800 -1156
rect 1760 -1236 1764 -1204
rect 1796 -1236 1800 -1204
rect 1760 -1284 1800 -1236
rect 1760 -1316 1764 -1284
rect 1796 -1316 1800 -1284
rect 1760 -1364 1800 -1316
rect 1760 -1396 1764 -1364
rect 1796 -1396 1800 -1364
rect 1760 -1444 1800 -1396
rect 1760 -1476 1764 -1444
rect 1796 -1476 1800 -1444
rect 1760 -1524 1800 -1476
rect 1760 -1556 1764 -1524
rect 1796 -1556 1800 -1524
rect 1760 -1604 1800 -1556
rect 1760 -1636 1764 -1604
rect 1796 -1636 1800 -1604
rect 1760 -1684 1800 -1636
rect 1760 -1716 1764 -1684
rect 1796 -1716 1800 -1684
rect 1760 -1764 1800 -1716
rect 1760 -1796 1764 -1764
rect 1796 -1796 1800 -1764
rect 1760 -1844 1800 -1796
rect 1760 -1876 1764 -1844
rect 1796 -1876 1800 -1844
rect 1760 -1924 1800 -1876
rect 1760 -1956 1764 -1924
rect 1796 -1956 1800 -1924
rect 1760 -2004 1800 -1956
rect 1760 -2036 1764 -2004
rect 1796 -2036 1800 -2004
rect 1760 -2084 1800 -2036
rect 1760 -2116 1764 -2084
rect 1796 -2116 1800 -2084
rect 1760 -2164 1800 -2116
rect 1760 -2196 1764 -2164
rect 1796 -2196 1800 -2164
rect 1760 -2244 1800 -2196
rect 1760 -2276 1764 -2244
rect 1796 -2276 1800 -2244
rect 1760 -2324 1800 -2276
rect 1760 -2356 1764 -2324
rect 1796 -2356 1800 -2324
rect 1760 -2404 1800 -2356
rect 1760 -2436 1764 -2404
rect 1796 -2436 1800 -2404
rect 1760 -2484 1800 -2436
rect 1760 -2516 1764 -2484
rect 1796 -2516 1800 -2484
rect 1760 -2564 1800 -2516
rect 1760 -2596 1764 -2564
rect 1796 -2596 1800 -2564
rect 1760 -2644 1800 -2596
rect 1760 -2676 1764 -2644
rect 1796 -2676 1800 -2644
rect 1760 -2724 1800 -2676
rect 1760 -2756 1764 -2724
rect 1796 -2756 1800 -2724
rect 1760 -2804 1800 -2756
rect 1760 -2836 1764 -2804
rect 1796 -2836 1800 -2804
rect 1760 -2884 1800 -2836
rect 1760 -2916 1764 -2884
rect 1796 -2916 1800 -2884
rect 1760 -2964 1800 -2916
rect 1760 -2996 1764 -2964
rect 1796 -2996 1800 -2964
rect 1760 -3044 1800 -2996
rect 1760 -3076 1764 -3044
rect 1796 -3076 1800 -3044
rect 1760 -3124 1800 -3076
rect 1760 -3156 1764 -3124
rect 1796 -3156 1800 -3124
rect 1760 -3204 1800 -3156
rect 1760 -3236 1764 -3204
rect 1796 -3236 1800 -3204
rect 1760 -3284 1800 -3236
rect 1760 -3316 1764 -3284
rect 1796 -3316 1800 -3284
rect 1760 -3364 1800 -3316
rect 1760 -3396 1764 -3364
rect 1796 -3396 1800 -3364
rect 1760 -3444 1800 -3396
rect 1760 -3476 1764 -3444
rect 1796 -3476 1800 -3444
rect 1760 -3524 1800 -3476
rect 1760 -3556 1764 -3524
rect 1796 -3556 1800 -3524
rect 1760 -3604 1800 -3556
rect 1760 -3636 1764 -3604
rect 1796 -3636 1800 -3604
rect 1760 -3684 1800 -3636
rect 1760 -3716 1764 -3684
rect 1796 -3716 1800 -3684
rect 1760 -3720 1800 -3716
rect 1840 1036 1880 1040
rect 1840 1004 1844 1036
rect 1876 1004 1880 1036
rect 1840 956 1880 1004
rect 1840 924 1844 956
rect 1876 924 1880 956
rect 1840 876 1880 924
rect 1840 844 1844 876
rect 1876 844 1880 876
rect 1840 796 1880 844
rect 1840 764 1844 796
rect 1876 764 1880 796
rect 1840 716 1880 764
rect 1840 684 1844 716
rect 1876 684 1880 716
rect 1840 636 1880 684
rect 1840 604 1844 636
rect 1876 604 1880 636
rect 1840 556 1880 604
rect 1840 524 1844 556
rect 1876 524 1880 556
rect 1840 476 1880 524
rect 1840 444 1844 476
rect 1876 444 1880 476
rect 1840 396 1880 444
rect 1840 364 1844 396
rect 1876 364 1880 396
rect 1840 316 1880 364
rect 1840 284 1844 316
rect 1876 284 1880 316
rect 1840 236 1880 284
rect 1840 204 1844 236
rect 1876 204 1880 236
rect 1840 156 1880 204
rect 1840 124 1844 156
rect 1876 124 1880 156
rect 1840 76 1880 124
rect 1840 44 1844 76
rect 1876 44 1880 76
rect 1840 -4 1880 44
rect 1840 -36 1844 -4
rect 1876 -36 1880 -4
rect 1840 -84 1880 -36
rect 1840 -116 1844 -84
rect 1876 -116 1880 -84
rect 1840 -164 1880 -116
rect 1840 -196 1844 -164
rect 1876 -196 1880 -164
rect 1840 -244 1880 -196
rect 1840 -276 1844 -244
rect 1876 -276 1880 -244
rect 1840 -324 1880 -276
rect 1840 -356 1844 -324
rect 1876 -356 1880 -324
rect 1840 -404 1880 -356
rect 1840 -436 1844 -404
rect 1876 -436 1880 -404
rect 1840 -484 1880 -436
rect 1840 -516 1844 -484
rect 1876 -516 1880 -484
rect 1840 -564 1880 -516
rect 1840 -596 1844 -564
rect 1876 -596 1880 -564
rect 1840 -644 1880 -596
rect 1840 -676 1844 -644
rect 1876 -676 1880 -644
rect 1840 -724 1880 -676
rect 1840 -756 1844 -724
rect 1876 -756 1880 -724
rect 1840 -804 1880 -756
rect 1840 -836 1844 -804
rect 1876 -836 1880 -804
rect 1840 -884 1880 -836
rect 1840 -916 1844 -884
rect 1876 -916 1880 -884
rect 1840 -964 1880 -916
rect 1840 -996 1844 -964
rect 1876 -996 1880 -964
rect 1840 -1044 1880 -996
rect 1840 -1076 1844 -1044
rect 1876 -1076 1880 -1044
rect 1840 -1124 1880 -1076
rect 1840 -1156 1844 -1124
rect 1876 -1156 1880 -1124
rect 1840 -1204 1880 -1156
rect 1840 -1236 1844 -1204
rect 1876 -1236 1880 -1204
rect 1840 -1284 1880 -1236
rect 1840 -1316 1844 -1284
rect 1876 -1316 1880 -1284
rect 1840 -1364 1880 -1316
rect 1840 -1396 1844 -1364
rect 1876 -1396 1880 -1364
rect 1840 -1444 1880 -1396
rect 1840 -1476 1844 -1444
rect 1876 -1476 1880 -1444
rect 1840 -1524 1880 -1476
rect 1840 -1556 1844 -1524
rect 1876 -1556 1880 -1524
rect 1840 -1604 1880 -1556
rect 1840 -1636 1844 -1604
rect 1876 -1636 1880 -1604
rect 1840 -1684 1880 -1636
rect 1840 -1716 1844 -1684
rect 1876 -1716 1880 -1684
rect 1840 -1764 1880 -1716
rect 1840 -1796 1844 -1764
rect 1876 -1796 1880 -1764
rect 1840 -1844 1880 -1796
rect 1840 -1876 1844 -1844
rect 1876 -1876 1880 -1844
rect 1840 -1924 1880 -1876
rect 1840 -1956 1844 -1924
rect 1876 -1956 1880 -1924
rect 1840 -2004 1880 -1956
rect 1840 -2036 1844 -2004
rect 1876 -2036 1880 -2004
rect 1840 -2084 1880 -2036
rect 1840 -2116 1844 -2084
rect 1876 -2116 1880 -2084
rect 1840 -2164 1880 -2116
rect 1840 -2196 1844 -2164
rect 1876 -2196 1880 -2164
rect 1840 -2244 1880 -2196
rect 1840 -2276 1844 -2244
rect 1876 -2276 1880 -2244
rect 1840 -2324 1880 -2276
rect 1840 -2356 1844 -2324
rect 1876 -2356 1880 -2324
rect 1840 -2404 1880 -2356
rect 1840 -2436 1844 -2404
rect 1876 -2436 1880 -2404
rect 1840 -2484 1880 -2436
rect 1840 -2516 1844 -2484
rect 1876 -2516 1880 -2484
rect 1840 -2564 1880 -2516
rect 1840 -2596 1844 -2564
rect 1876 -2596 1880 -2564
rect 1840 -2644 1880 -2596
rect 1840 -2676 1844 -2644
rect 1876 -2676 1880 -2644
rect 1840 -2724 1880 -2676
rect 1840 -2756 1844 -2724
rect 1876 -2756 1880 -2724
rect 1840 -2804 1880 -2756
rect 1840 -2836 1844 -2804
rect 1876 -2836 1880 -2804
rect 1840 -2884 1880 -2836
rect 1840 -2916 1844 -2884
rect 1876 -2916 1880 -2884
rect 1840 -2964 1880 -2916
rect 1840 -2996 1844 -2964
rect 1876 -2996 1880 -2964
rect 1840 -3044 1880 -2996
rect 1840 -3076 1844 -3044
rect 1876 -3076 1880 -3044
rect 1840 -3124 1880 -3076
rect 1840 -3156 1844 -3124
rect 1876 -3156 1880 -3124
rect 1840 -3204 1880 -3156
rect 1840 -3236 1844 -3204
rect 1876 -3236 1880 -3204
rect 1840 -3284 1880 -3236
rect 1840 -3316 1844 -3284
rect 1876 -3316 1880 -3284
rect 1840 -3364 1880 -3316
rect 1840 -3396 1844 -3364
rect 1876 -3396 1880 -3364
rect 1840 -3444 1880 -3396
rect 1840 -3476 1844 -3444
rect 1876 -3476 1880 -3444
rect 1840 -3524 1880 -3476
rect 1840 -3556 1844 -3524
rect 1876 -3556 1880 -3524
rect 1840 -3604 1880 -3556
rect 1840 -3636 1844 -3604
rect 1876 -3636 1880 -3604
rect 1840 -3684 1880 -3636
rect 1840 -3716 1844 -3684
rect 1876 -3716 1880 -3684
rect 1840 -3720 1880 -3716
rect 1920 1036 1960 1040
rect 1920 1004 1924 1036
rect 1956 1004 1960 1036
rect 1920 956 1960 1004
rect 1920 924 1924 956
rect 1956 924 1960 956
rect 1920 876 1960 924
rect 1920 844 1924 876
rect 1956 844 1960 876
rect 1920 796 1960 844
rect 1920 764 1924 796
rect 1956 764 1960 796
rect 1920 716 1960 764
rect 1920 684 1924 716
rect 1956 684 1960 716
rect 1920 636 1960 684
rect 1920 604 1924 636
rect 1956 604 1960 636
rect 1920 556 1960 604
rect 1920 524 1924 556
rect 1956 524 1960 556
rect 1920 476 1960 524
rect 1920 444 1924 476
rect 1956 444 1960 476
rect 1920 396 1960 444
rect 1920 364 1924 396
rect 1956 364 1960 396
rect 1920 316 1960 364
rect 1920 284 1924 316
rect 1956 284 1960 316
rect 1920 236 1960 284
rect 1920 204 1924 236
rect 1956 204 1960 236
rect 1920 156 1960 204
rect 1920 124 1924 156
rect 1956 124 1960 156
rect 1920 76 1960 124
rect 1920 44 1924 76
rect 1956 44 1960 76
rect 1920 -4 1960 44
rect 1920 -36 1924 -4
rect 1956 -36 1960 -4
rect 1920 -84 1960 -36
rect 1920 -116 1924 -84
rect 1956 -116 1960 -84
rect 1920 -164 1960 -116
rect 1920 -196 1924 -164
rect 1956 -196 1960 -164
rect 1920 -244 1960 -196
rect 1920 -276 1924 -244
rect 1956 -276 1960 -244
rect 1920 -324 1960 -276
rect 1920 -356 1924 -324
rect 1956 -356 1960 -324
rect 1920 -404 1960 -356
rect 1920 -436 1924 -404
rect 1956 -436 1960 -404
rect 1920 -484 1960 -436
rect 1920 -516 1924 -484
rect 1956 -516 1960 -484
rect 1920 -564 1960 -516
rect 1920 -596 1924 -564
rect 1956 -596 1960 -564
rect 1920 -644 1960 -596
rect 1920 -676 1924 -644
rect 1956 -676 1960 -644
rect 1920 -724 1960 -676
rect 1920 -756 1924 -724
rect 1956 -756 1960 -724
rect 1920 -804 1960 -756
rect 1920 -836 1924 -804
rect 1956 -836 1960 -804
rect 1920 -884 1960 -836
rect 1920 -916 1924 -884
rect 1956 -916 1960 -884
rect 1920 -964 1960 -916
rect 1920 -996 1924 -964
rect 1956 -996 1960 -964
rect 1920 -1044 1960 -996
rect 1920 -1076 1924 -1044
rect 1956 -1076 1960 -1044
rect 1920 -1124 1960 -1076
rect 1920 -1156 1924 -1124
rect 1956 -1156 1960 -1124
rect 1920 -1204 1960 -1156
rect 1920 -1236 1924 -1204
rect 1956 -1236 1960 -1204
rect 1920 -1284 1960 -1236
rect 1920 -1316 1924 -1284
rect 1956 -1316 1960 -1284
rect 1920 -1364 1960 -1316
rect 1920 -1396 1924 -1364
rect 1956 -1396 1960 -1364
rect 1920 -1444 1960 -1396
rect 1920 -1476 1924 -1444
rect 1956 -1476 1960 -1444
rect 1920 -1524 1960 -1476
rect 1920 -1556 1924 -1524
rect 1956 -1556 1960 -1524
rect 1920 -1604 1960 -1556
rect 1920 -1636 1924 -1604
rect 1956 -1636 1960 -1604
rect 1920 -1684 1960 -1636
rect 1920 -1716 1924 -1684
rect 1956 -1716 1960 -1684
rect 1920 -1764 1960 -1716
rect 1920 -1796 1924 -1764
rect 1956 -1796 1960 -1764
rect 1920 -1844 1960 -1796
rect 1920 -1876 1924 -1844
rect 1956 -1876 1960 -1844
rect 1920 -1924 1960 -1876
rect 1920 -1956 1924 -1924
rect 1956 -1956 1960 -1924
rect 1920 -2004 1960 -1956
rect 1920 -2036 1924 -2004
rect 1956 -2036 1960 -2004
rect 1920 -2084 1960 -2036
rect 1920 -2116 1924 -2084
rect 1956 -2116 1960 -2084
rect 1920 -2164 1960 -2116
rect 1920 -2196 1924 -2164
rect 1956 -2196 1960 -2164
rect 1920 -2244 1960 -2196
rect 1920 -2276 1924 -2244
rect 1956 -2276 1960 -2244
rect 1920 -2324 1960 -2276
rect 1920 -2356 1924 -2324
rect 1956 -2356 1960 -2324
rect 1920 -2404 1960 -2356
rect 1920 -2436 1924 -2404
rect 1956 -2436 1960 -2404
rect 1920 -2484 1960 -2436
rect 1920 -2516 1924 -2484
rect 1956 -2516 1960 -2484
rect 1920 -2564 1960 -2516
rect 1920 -2596 1924 -2564
rect 1956 -2596 1960 -2564
rect 1920 -2644 1960 -2596
rect 1920 -2676 1924 -2644
rect 1956 -2676 1960 -2644
rect 1920 -2724 1960 -2676
rect 1920 -2756 1924 -2724
rect 1956 -2756 1960 -2724
rect 1920 -2804 1960 -2756
rect 1920 -2836 1924 -2804
rect 1956 -2836 1960 -2804
rect 1920 -2884 1960 -2836
rect 1920 -2916 1924 -2884
rect 1956 -2916 1960 -2884
rect 1920 -2964 1960 -2916
rect 1920 -2996 1924 -2964
rect 1956 -2996 1960 -2964
rect 1920 -3044 1960 -2996
rect 1920 -3076 1924 -3044
rect 1956 -3076 1960 -3044
rect 1920 -3124 1960 -3076
rect 1920 -3156 1924 -3124
rect 1956 -3156 1960 -3124
rect 1920 -3204 1960 -3156
rect 1920 -3236 1924 -3204
rect 1956 -3236 1960 -3204
rect 1920 -3284 1960 -3236
rect 1920 -3316 1924 -3284
rect 1956 -3316 1960 -3284
rect 1920 -3364 1960 -3316
rect 1920 -3396 1924 -3364
rect 1956 -3396 1960 -3364
rect 1920 -3444 1960 -3396
rect 1920 -3476 1924 -3444
rect 1956 -3476 1960 -3444
rect 1920 -3524 1960 -3476
rect 1920 -3556 1924 -3524
rect 1956 -3556 1960 -3524
rect 1920 -3604 1960 -3556
rect 1920 -3636 1924 -3604
rect 1956 -3636 1960 -3604
rect 1920 -3684 1960 -3636
rect 1920 -3716 1924 -3684
rect 1956 -3716 1960 -3684
rect 1920 -3720 1960 -3716
rect 2000 1036 2040 1040
rect 2000 1004 2004 1036
rect 2036 1004 2040 1036
rect 2000 956 2040 1004
rect 2000 924 2004 956
rect 2036 924 2040 956
rect 2000 876 2040 924
rect 2000 844 2004 876
rect 2036 844 2040 876
rect 2000 796 2040 844
rect 2000 764 2004 796
rect 2036 764 2040 796
rect 2000 716 2040 764
rect 2000 684 2004 716
rect 2036 684 2040 716
rect 2000 636 2040 684
rect 2000 604 2004 636
rect 2036 604 2040 636
rect 2000 556 2040 604
rect 2000 524 2004 556
rect 2036 524 2040 556
rect 2000 476 2040 524
rect 2000 444 2004 476
rect 2036 444 2040 476
rect 2000 396 2040 444
rect 2000 364 2004 396
rect 2036 364 2040 396
rect 2000 316 2040 364
rect 2000 284 2004 316
rect 2036 284 2040 316
rect 2000 236 2040 284
rect 2000 204 2004 236
rect 2036 204 2040 236
rect 2000 156 2040 204
rect 2000 124 2004 156
rect 2036 124 2040 156
rect 2000 76 2040 124
rect 2000 44 2004 76
rect 2036 44 2040 76
rect 2000 -4 2040 44
rect 2000 -36 2004 -4
rect 2036 -36 2040 -4
rect 2000 -84 2040 -36
rect 2000 -116 2004 -84
rect 2036 -116 2040 -84
rect 2000 -164 2040 -116
rect 2000 -196 2004 -164
rect 2036 -196 2040 -164
rect 2000 -244 2040 -196
rect 2000 -276 2004 -244
rect 2036 -276 2040 -244
rect 2000 -324 2040 -276
rect 2000 -356 2004 -324
rect 2036 -356 2040 -324
rect 2000 -404 2040 -356
rect 2000 -436 2004 -404
rect 2036 -436 2040 -404
rect 2000 -484 2040 -436
rect 2000 -516 2004 -484
rect 2036 -516 2040 -484
rect 2000 -564 2040 -516
rect 2000 -596 2004 -564
rect 2036 -596 2040 -564
rect 2000 -644 2040 -596
rect 2000 -676 2004 -644
rect 2036 -676 2040 -644
rect 2000 -724 2040 -676
rect 2000 -756 2004 -724
rect 2036 -756 2040 -724
rect 2000 -804 2040 -756
rect 2000 -836 2004 -804
rect 2036 -836 2040 -804
rect 2000 -884 2040 -836
rect 2000 -916 2004 -884
rect 2036 -916 2040 -884
rect 2000 -964 2040 -916
rect 2000 -996 2004 -964
rect 2036 -996 2040 -964
rect 2000 -1044 2040 -996
rect 2000 -1076 2004 -1044
rect 2036 -1076 2040 -1044
rect 2000 -1124 2040 -1076
rect 2000 -1156 2004 -1124
rect 2036 -1156 2040 -1124
rect 2000 -1204 2040 -1156
rect 2000 -1236 2004 -1204
rect 2036 -1236 2040 -1204
rect 2000 -1284 2040 -1236
rect 2000 -1316 2004 -1284
rect 2036 -1316 2040 -1284
rect 2000 -1364 2040 -1316
rect 2000 -1396 2004 -1364
rect 2036 -1396 2040 -1364
rect 2000 -1444 2040 -1396
rect 2000 -1476 2004 -1444
rect 2036 -1476 2040 -1444
rect 2000 -1524 2040 -1476
rect 2000 -1556 2004 -1524
rect 2036 -1556 2040 -1524
rect 2000 -1604 2040 -1556
rect 2000 -1636 2004 -1604
rect 2036 -1636 2040 -1604
rect 2000 -1684 2040 -1636
rect 2000 -1716 2004 -1684
rect 2036 -1716 2040 -1684
rect 2000 -1764 2040 -1716
rect 2000 -1796 2004 -1764
rect 2036 -1796 2040 -1764
rect 2000 -1844 2040 -1796
rect 2000 -1876 2004 -1844
rect 2036 -1876 2040 -1844
rect 2000 -1924 2040 -1876
rect 2000 -1956 2004 -1924
rect 2036 -1956 2040 -1924
rect 2000 -2004 2040 -1956
rect 2000 -2036 2004 -2004
rect 2036 -2036 2040 -2004
rect 2000 -2084 2040 -2036
rect 2000 -2116 2004 -2084
rect 2036 -2116 2040 -2084
rect 2000 -2164 2040 -2116
rect 2000 -2196 2004 -2164
rect 2036 -2196 2040 -2164
rect 2000 -2244 2040 -2196
rect 2000 -2276 2004 -2244
rect 2036 -2276 2040 -2244
rect 2000 -2324 2040 -2276
rect 2000 -2356 2004 -2324
rect 2036 -2356 2040 -2324
rect 2000 -2404 2040 -2356
rect 2000 -2436 2004 -2404
rect 2036 -2436 2040 -2404
rect 2000 -2484 2040 -2436
rect 2000 -2516 2004 -2484
rect 2036 -2516 2040 -2484
rect 2000 -2564 2040 -2516
rect 2000 -2596 2004 -2564
rect 2036 -2596 2040 -2564
rect 2000 -2644 2040 -2596
rect 2000 -2676 2004 -2644
rect 2036 -2676 2040 -2644
rect 2000 -2724 2040 -2676
rect 2000 -2756 2004 -2724
rect 2036 -2756 2040 -2724
rect 2000 -2804 2040 -2756
rect 2000 -2836 2004 -2804
rect 2036 -2836 2040 -2804
rect 2000 -2884 2040 -2836
rect 2000 -2916 2004 -2884
rect 2036 -2916 2040 -2884
rect 2000 -2964 2040 -2916
rect 2000 -2996 2004 -2964
rect 2036 -2996 2040 -2964
rect 2000 -3044 2040 -2996
rect 2000 -3076 2004 -3044
rect 2036 -3076 2040 -3044
rect 2000 -3124 2040 -3076
rect 2000 -3156 2004 -3124
rect 2036 -3156 2040 -3124
rect 2000 -3204 2040 -3156
rect 2000 -3236 2004 -3204
rect 2036 -3236 2040 -3204
rect 2000 -3284 2040 -3236
rect 2000 -3316 2004 -3284
rect 2036 -3316 2040 -3284
rect 2000 -3364 2040 -3316
rect 2000 -3396 2004 -3364
rect 2036 -3396 2040 -3364
rect 2000 -3444 2040 -3396
rect 2000 -3476 2004 -3444
rect 2036 -3476 2040 -3444
rect 2000 -3524 2040 -3476
rect 2000 -3556 2004 -3524
rect 2036 -3556 2040 -3524
rect 2000 -3604 2040 -3556
rect 2000 -3636 2004 -3604
rect 2036 -3636 2040 -3604
rect 2000 -3684 2040 -3636
rect 2000 -3716 2004 -3684
rect 2036 -3716 2040 -3684
rect 2000 -3720 2040 -3716
rect 2080 1036 2120 1040
rect 2080 1004 2084 1036
rect 2116 1004 2120 1036
rect 2080 956 2120 1004
rect 2080 924 2084 956
rect 2116 924 2120 956
rect 2080 876 2120 924
rect 2080 844 2084 876
rect 2116 844 2120 876
rect 2080 796 2120 844
rect 2080 764 2084 796
rect 2116 764 2120 796
rect 2080 716 2120 764
rect 2080 684 2084 716
rect 2116 684 2120 716
rect 2080 636 2120 684
rect 2080 604 2084 636
rect 2116 604 2120 636
rect 2080 556 2120 604
rect 2080 524 2084 556
rect 2116 524 2120 556
rect 2080 476 2120 524
rect 2080 444 2084 476
rect 2116 444 2120 476
rect 2080 396 2120 444
rect 2080 364 2084 396
rect 2116 364 2120 396
rect 2080 316 2120 364
rect 2080 284 2084 316
rect 2116 284 2120 316
rect 2080 236 2120 284
rect 2080 204 2084 236
rect 2116 204 2120 236
rect 2080 156 2120 204
rect 2080 124 2084 156
rect 2116 124 2120 156
rect 2080 76 2120 124
rect 2080 44 2084 76
rect 2116 44 2120 76
rect 2080 -4 2120 44
rect 2080 -36 2084 -4
rect 2116 -36 2120 -4
rect 2080 -84 2120 -36
rect 2080 -116 2084 -84
rect 2116 -116 2120 -84
rect 2080 -164 2120 -116
rect 2080 -196 2084 -164
rect 2116 -196 2120 -164
rect 2080 -244 2120 -196
rect 2080 -276 2084 -244
rect 2116 -276 2120 -244
rect 2080 -324 2120 -276
rect 2080 -356 2084 -324
rect 2116 -356 2120 -324
rect 2080 -404 2120 -356
rect 2080 -436 2084 -404
rect 2116 -436 2120 -404
rect 2080 -484 2120 -436
rect 2080 -516 2084 -484
rect 2116 -516 2120 -484
rect 2080 -564 2120 -516
rect 2080 -596 2084 -564
rect 2116 -596 2120 -564
rect 2080 -644 2120 -596
rect 2080 -676 2084 -644
rect 2116 -676 2120 -644
rect 2080 -724 2120 -676
rect 2080 -756 2084 -724
rect 2116 -756 2120 -724
rect 2080 -804 2120 -756
rect 2080 -836 2084 -804
rect 2116 -836 2120 -804
rect 2080 -884 2120 -836
rect 2080 -916 2084 -884
rect 2116 -916 2120 -884
rect 2080 -964 2120 -916
rect 2080 -996 2084 -964
rect 2116 -996 2120 -964
rect 2080 -1044 2120 -996
rect 2080 -1076 2084 -1044
rect 2116 -1076 2120 -1044
rect 2080 -1124 2120 -1076
rect 2080 -1156 2084 -1124
rect 2116 -1156 2120 -1124
rect 2080 -1204 2120 -1156
rect 2080 -1236 2084 -1204
rect 2116 -1236 2120 -1204
rect 2080 -1284 2120 -1236
rect 2080 -1316 2084 -1284
rect 2116 -1316 2120 -1284
rect 2080 -1364 2120 -1316
rect 2080 -1396 2084 -1364
rect 2116 -1396 2120 -1364
rect 2080 -1444 2120 -1396
rect 2080 -1476 2084 -1444
rect 2116 -1476 2120 -1444
rect 2080 -1524 2120 -1476
rect 2080 -1556 2084 -1524
rect 2116 -1556 2120 -1524
rect 2080 -1604 2120 -1556
rect 2080 -1636 2084 -1604
rect 2116 -1636 2120 -1604
rect 2080 -1684 2120 -1636
rect 2080 -1716 2084 -1684
rect 2116 -1716 2120 -1684
rect 2080 -1764 2120 -1716
rect 2080 -1796 2084 -1764
rect 2116 -1796 2120 -1764
rect 2080 -1844 2120 -1796
rect 2080 -1876 2084 -1844
rect 2116 -1876 2120 -1844
rect 2080 -1924 2120 -1876
rect 2080 -1956 2084 -1924
rect 2116 -1956 2120 -1924
rect 2080 -2004 2120 -1956
rect 2080 -2036 2084 -2004
rect 2116 -2036 2120 -2004
rect 2080 -2084 2120 -2036
rect 2080 -2116 2084 -2084
rect 2116 -2116 2120 -2084
rect 2080 -2164 2120 -2116
rect 2080 -2196 2084 -2164
rect 2116 -2196 2120 -2164
rect 2080 -2244 2120 -2196
rect 2080 -2276 2084 -2244
rect 2116 -2276 2120 -2244
rect 2080 -2324 2120 -2276
rect 2080 -2356 2084 -2324
rect 2116 -2356 2120 -2324
rect 2080 -2404 2120 -2356
rect 2080 -2436 2084 -2404
rect 2116 -2436 2120 -2404
rect 2080 -2484 2120 -2436
rect 2080 -2516 2084 -2484
rect 2116 -2516 2120 -2484
rect 2080 -2564 2120 -2516
rect 2080 -2596 2084 -2564
rect 2116 -2596 2120 -2564
rect 2080 -2644 2120 -2596
rect 2080 -2676 2084 -2644
rect 2116 -2676 2120 -2644
rect 2080 -2724 2120 -2676
rect 2080 -2756 2084 -2724
rect 2116 -2756 2120 -2724
rect 2080 -2804 2120 -2756
rect 2080 -2836 2084 -2804
rect 2116 -2836 2120 -2804
rect 2080 -2884 2120 -2836
rect 2080 -2916 2084 -2884
rect 2116 -2916 2120 -2884
rect 2080 -2964 2120 -2916
rect 2080 -2996 2084 -2964
rect 2116 -2996 2120 -2964
rect 2080 -3044 2120 -2996
rect 2080 -3076 2084 -3044
rect 2116 -3076 2120 -3044
rect 2080 -3124 2120 -3076
rect 2080 -3156 2084 -3124
rect 2116 -3156 2120 -3124
rect 2080 -3204 2120 -3156
rect 2080 -3236 2084 -3204
rect 2116 -3236 2120 -3204
rect 2080 -3284 2120 -3236
rect 2080 -3316 2084 -3284
rect 2116 -3316 2120 -3284
rect 2080 -3364 2120 -3316
rect 2080 -3396 2084 -3364
rect 2116 -3396 2120 -3364
rect 2080 -3444 2120 -3396
rect 2080 -3476 2084 -3444
rect 2116 -3476 2120 -3444
rect 2080 -3524 2120 -3476
rect 2080 -3556 2084 -3524
rect 2116 -3556 2120 -3524
rect 2080 -3604 2120 -3556
rect 2080 -3636 2084 -3604
rect 2116 -3636 2120 -3604
rect 2080 -3684 2120 -3636
rect 2080 -3716 2084 -3684
rect 2116 -3716 2120 -3684
rect 2080 -3720 2120 -3716
rect 2160 1036 2200 1040
rect 2160 1004 2164 1036
rect 2196 1004 2200 1036
rect 2160 956 2200 1004
rect 2160 924 2164 956
rect 2196 924 2200 956
rect 2160 876 2200 924
rect 2160 844 2164 876
rect 2196 844 2200 876
rect 2160 796 2200 844
rect 2160 764 2164 796
rect 2196 764 2200 796
rect 2160 716 2200 764
rect 2160 684 2164 716
rect 2196 684 2200 716
rect 2160 636 2200 684
rect 2160 604 2164 636
rect 2196 604 2200 636
rect 2160 556 2200 604
rect 2160 524 2164 556
rect 2196 524 2200 556
rect 2160 476 2200 524
rect 2160 444 2164 476
rect 2196 444 2200 476
rect 2160 396 2200 444
rect 2160 364 2164 396
rect 2196 364 2200 396
rect 2160 316 2200 364
rect 2160 284 2164 316
rect 2196 284 2200 316
rect 2160 236 2200 284
rect 2160 204 2164 236
rect 2196 204 2200 236
rect 2160 156 2200 204
rect 2160 124 2164 156
rect 2196 124 2200 156
rect 2160 76 2200 124
rect 2160 44 2164 76
rect 2196 44 2200 76
rect 2160 -4 2200 44
rect 2160 -36 2164 -4
rect 2196 -36 2200 -4
rect 2160 -84 2200 -36
rect 2160 -116 2164 -84
rect 2196 -116 2200 -84
rect 2160 -164 2200 -116
rect 2160 -196 2164 -164
rect 2196 -196 2200 -164
rect 2160 -244 2200 -196
rect 2160 -276 2164 -244
rect 2196 -276 2200 -244
rect 2160 -324 2200 -276
rect 2160 -356 2164 -324
rect 2196 -356 2200 -324
rect 2160 -404 2200 -356
rect 2160 -436 2164 -404
rect 2196 -436 2200 -404
rect 2160 -484 2200 -436
rect 2160 -516 2164 -484
rect 2196 -516 2200 -484
rect 2160 -564 2200 -516
rect 2160 -596 2164 -564
rect 2196 -596 2200 -564
rect 2160 -644 2200 -596
rect 2160 -676 2164 -644
rect 2196 -676 2200 -644
rect 2160 -724 2200 -676
rect 2160 -756 2164 -724
rect 2196 -756 2200 -724
rect 2160 -804 2200 -756
rect 2160 -836 2164 -804
rect 2196 -836 2200 -804
rect 2160 -884 2200 -836
rect 2160 -916 2164 -884
rect 2196 -916 2200 -884
rect 2160 -964 2200 -916
rect 2160 -996 2164 -964
rect 2196 -996 2200 -964
rect 2160 -1044 2200 -996
rect 2160 -1076 2164 -1044
rect 2196 -1076 2200 -1044
rect 2160 -1124 2200 -1076
rect 2160 -1156 2164 -1124
rect 2196 -1156 2200 -1124
rect 2160 -1204 2200 -1156
rect 2160 -1236 2164 -1204
rect 2196 -1236 2200 -1204
rect 2160 -1284 2200 -1236
rect 2160 -1316 2164 -1284
rect 2196 -1316 2200 -1284
rect 2160 -1364 2200 -1316
rect 2160 -1396 2164 -1364
rect 2196 -1396 2200 -1364
rect 2160 -1444 2200 -1396
rect 2160 -1476 2164 -1444
rect 2196 -1476 2200 -1444
rect 2160 -1524 2200 -1476
rect 2160 -1556 2164 -1524
rect 2196 -1556 2200 -1524
rect 2160 -1604 2200 -1556
rect 2160 -1636 2164 -1604
rect 2196 -1636 2200 -1604
rect 2160 -1684 2200 -1636
rect 2160 -1716 2164 -1684
rect 2196 -1716 2200 -1684
rect 2160 -1764 2200 -1716
rect 2160 -1796 2164 -1764
rect 2196 -1796 2200 -1764
rect 2160 -1844 2200 -1796
rect 2160 -1876 2164 -1844
rect 2196 -1876 2200 -1844
rect 2160 -1924 2200 -1876
rect 2160 -1956 2164 -1924
rect 2196 -1956 2200 -1924
rect 2160 -2004 2200 -1956
rect 2160 -2036 2164 -2004
rect 2196 -2036 2200 -2004
rect 2160 -2084 2200 -2036
rect 2160 -2116 2164 -2084
rect 2196 -2116 2200 -2084
rect 2160 -2164 2200 -2116
rect 2160 -2196 2164 -2164
rect 2196 -2196 2200 -2164
rect 2160 -2244 2200 -2196
rect 2160 -2276 2164 -2244
rect 2196 -2276 2200 -2244
rect 2160 -2324 2200 -2276
rect 2160 -2356 2164 -2324
rect 2196 -2356 2200 -2324
rect 2160 -2404 2200 -2356
rect 2160 -2436 2164 -2404
rect 2196 -2436 2200 -2404
rect 2160 -2484 2200 -2436
rect 2160 -2516 2164 -2484
rect 2196 -2516 2200 -2484
rect 2160 -2564 2200 -2516
rect 2160 -2596 2164 -2564
rect 2196 -2596 2200 -2564
rect 2160 -2644 2200 -2596
rect 2160 -2676 2164 -2644
rect 2196 -2676 2200 -2644
rect 2160 -2724 2200 -2676
rect 2160 -2756 2164 -2724
rect 2196 -2756 2200 -2724
rect 2160 -2804 2200 -2756
rect 2160 -2836 2164 -2804
rect 2196 -2836 2200 -2804
rect 2160 -2884 2200 -2836
rect 2160 -2916 2164 -2884
rect 2196 -2916 2200 -2884
rect 2160 -2964 2200 -2916
rect 2160 -2996 2164 -2964
rect 2196 -2996 2200 -2964
rect 2160 -3044 2200 -2996
rect 2160 -3076 2164 -3044
rect 2196 -3076 2200 -3044
rect 2160 -3124 2200 -3076
rect 2160 -3156 2164 -3124
rect 2196 -3156 2200 -3124
rect 2160 -3204 2200 -3156
rect 2160 -3236 2164 -3204
rect 2196 -3236 2200 -3204
rect 2160 -3284 2200 -3236
rect 2160 -3316 2164 -3284
rect 2196 -3316 2200 -3284
rect 2160 -3364 2200 -3316
rect 2160 -3396 2164 -3364
rect 2196 -3396 2200 -3364
rect 2160 -3444 2200 -3396
rect 2160 -3476 2164 -3444
rect 2196 -3476 2200 -3444
rect 2160 -3524 2200 -3476
rect 2160 -3556 2164 -3524
rect 2196 -3556 2200 -3524
rect 2160 -3604 2200 -3556
rect 2160 -3636 2164 -3604
rect 2196 -3636 2200 -3604
rect 2160 -3684 2200 -3636
rect 2160 -3716 2164 -3684
rect 2196 -3716 2200 -3684
rect 2160 -3720 2200 -3716
rect 2240 1036 2280 1040
rect 2240 1004 2244 1036
rect 2276 1004 2280 1036
rect 2240 956 2280 1004
rect 2240 924 2244 956
rect 2276 924 2280 956
rect 2240 876 2280 924
rect 2240 844 2244 876
rect 2276 844 2280 876
rect 2240 796 2280 844
rect 2240 764 2244 796
rect 2276 764 2280 796
rect 2240 716 2280 764
rect 2240 684 2244 716
rect 2276 684 2280 716
rect 2240 636 2280 684
rect 2240 604 2244 636
rect 2276 604 2280 636
rect 2240 556 2280 604
rect 2240 524 2244 556
rect 2276 524 2280 556
rect 2240 476 2280 524
rect 2240 444 2244 476
rect 2276 444 2280 476
rect 2240 396 2280 444
rect 2240 364 2244 396
rect 2276 364 2280 396
rect 2240 316 2280 364
rect 2240 284 2244 316
rect 2276 284 2280 316
rect 2240 236 2280 284
rect 2240 204 2244 236
rect 2276 204 2280 236
rect 2240 156 2280 204
rect 2240 124 2244 156
rect 2276 124 2280 156
rect 2240 76 2280 124
rect 2240 44 2244 76
rect 2276 44 2280 76
rect 2240 -4 2280 44
rect 2240 -36 2244 -4
rect 2276 -36 2280 -4
rect 2240 -84 2280 -36
rect 2240 -116 2244 -84
rect 2276 -116 2280 -84
rect 2240 -164 2280 -116
rect 2240 -196 2244 -164
rect 2276 -196 2280 -164
rect 2240 -244 2280 -196
rect 2240 -276 2244 -244
rect 2276 -276 2280 -244
rect 2240 -324 2280 -276
rect 2240 -356 2244 -324
rect 2276 -356 2280 -324
rect 2240 -404 2280 -356
rect 2240 -436 2244 -404
rect 2276 -436 2280 -404
rect 2240 -484 2280 -436
rect 2240 -516 2244 -484
rect 2276 -516 2280 -484
rect 2240 -564 2280 -516
rect 2240 -596 2244 -564
rect 2276 -596 2280 -564
rect 2240 -644 2280 -596
rect 2240 -676 2244 -644
rect 2276 -676 2280 -644
rect 2240 -724 2280 -676
rect 2240 -756 2244 -724
rect 2276 -756 2280 -724
rect 2240 -804 2280 -756
rect 2240 -836 2244 -804
rect 2276 -836 2280 -804
rect 2240 -884 2280 -836
rect 2240 -916 2244 -884
rect 2276 -916 2280 -884
rect 2240 -964 2280 -916
rect 2240 -996 2244 -964
rect 2276 -996 2280 -964
rect 2240 -1044 2280 -996
rect 2240 -1076 2244 -1044
rect 2276 -1076 2280 -1044
rect 2240 -1124 2280 -1076
rect 2240 -1156 2244 -1124
rect 2276 -1156 2280 -1124
rect 2240 -1204 2280 -1156
rect 2240 -1236 2244 -1204
rect 2276 -1236 2280 -1204
rect 2240 -1284 2280 -1236
rect 2240 -1316 2244 -1284
rect 2276 -1316 2280 -1284
rect 2240 -1364 2280 -1316
rect 2240 -1396 2244 -1364
rect 2276 -1396 2280 -1364
rect 2240 -1444 2280 -1396
rect 2240 -1476 2244 -1444
rect 2276 -1476 2280 -1444
rect 2240 -1524 2280 -1476
rect 2240 -1556 2244 -1524
rect 2276 -1556 2280 -1524
rect 2240 -1604 2280 -1556
rect 2240 -1636 2244 -1604
rect 2276 -1636 2280 -1604
rect 2240 -1684 2280 -1636
rect 2240 -1716 2244 -1684
rect 2276 -1716 2280 -1684
rect 2240 -1764 2280 -1716
rect 2240 -1796 2244 -1764
rect 2276 -1796 2280 -1764
rect 2240 -1844 2280 -1796
rect 2240 -1876 2244 -1844
rect 2276 -1876 2280 -1844
rect 2240 -1924 2280 -1876
rect 2240 -1956 2244 -1924
rect 2276 -1956 2280 -1924
rect 2240 -2004 2280 -1956
rect 2240 -2036 2244 -2004
rect 2276 -2036 2280 -2004
rect 2240 -2084 2280 -2036
rect 2240 -2116 2244 -2084
rect 2276 -2116 2280 -2084
rect 2240 -2164 2280 -2116
rect 2240 -2196 2244 -2164
rect 2276 -2196 2280 -2164
rect 2240 -2244 2280 -2196
rect 2240 -2276 2244 -2244
rect 2276 -2276 2280 -2244
rect 2240 -2324 2280 -2276
rect 2240 -2356 2244 -2324
rect 2276 -2356 2280 -2324
rect 2240 -2404 2280 -2356
rect 2240 -2436 2244 -2404
rect 2276 -2436 2280 -2404
rect 2240 -2484 2280 -2436
rect 2240 -2516 2244 -2484
rect 2276 -2516 2280 -2484
rect 2240 -2564 2280 -2516
rect 2240 -2596 2244 -2564
rect 2276 -2596 2280 -2564
rect 2240 -2644 2280 -2596
rect 2240 -2676 2244 -2644
rect 2276 -2676 2280 -2644
rect 2240 -2724 2280 -2676
rect 2240 -2756 2244 -2724
rect 2276 -2756 2280 -2724
rect 2240 -2804 2280 -2756
rect 2240 -2836 2244 -2804
rect 2276 -2836 2280 -2804
rect 2240 -2884 2280 -2836
rect 2240 -2916 2244 -2884
rect 2276 -2916 2280 -2884
rect 2240 -2964 2280 -2916
rect 2240 -2996 2244 -2964
rect 2276 -2996 2280 -2964
rect 2240 -3044 2280 -2996
rect 2240 -3076 2244 -3044
rect 2276 -3076 2280 -3044
rect 2240 -3124 2280 -3076
rect 2240 -3156 2244 -3124
rect 2276 -3156 2280 -3124
rect 2240 -3204 2280 -3156
rect 2240 -3236 2244 -3204
rect 2276 -3236 2280 -3204
rect 2240 -3284 2280 -3236
rect 2240 -3316 2244 -3284
rect 2276 -3316 2280 -3284
rect 2240 -3364 2280 -3316
rect 2240 -3396 2244 -3364
rect 2276 -3396 2280 -3364
rect 2240 -3444 2280 -3396
rect 2240 -3476 2244 -3444
rect 2276 -3476 2280 -3444
rect 2240 -3524 2280 -3476
rect 2240 -3556 2244 -3524
rect 2276 -3556 2280 -3524
rect 2240 -3604 2280 -3556
rect 2240 -3636 2244 -3604
rect 2276 -3636 2280 -3604
rect 2240 -3684 2280 -3636
rect 2240 -3716 2244 -3684
rect 2276 -3716 2280 -3684
rect 2240 -3720 2280 -3716
rect 2320 1036 2360 1040
rect 2320 1004 2324 1036
rect 2356 1004 2360 1036
rect 2320 956 2360 1004
rect 2320 924 2324 956
rect 2356 924 2360 956
rect 2320 876 2360 924
rect 2320 844 2324 876
rect 2356 844 2360 876
rect 2320 796 2360 844
rect 2320 764 2324 796
rect 2356 764 2360 796
rect 2320 716 2360 764
rect 2320 684 2324 716
rect 2356 684 2360 716
rect 2320 636 2360 684
rect 2320 604 2324 636
rect 2356 604 2360 636
rect 2320 556 2360 604
rect 2320 524 2324 556
rect 2356 524 2360 556
rect 2320 476 2360 524
rect 2320 444 2324 476
rect 2356 444 2360 476
rect 2320 396 2360 444
rect 2320 364 2324 396
rect 2356 364 2360 396
rect 2320 316 2360 364
rect 2320 284 2324 316
rect 2356 284 2360 316
rect 2320 236 2360 284
rect 2320 204 2324 236
rect 2356 204 2360 236
rect 2320 156 2360 204
rect 2320 124 2324 156
rect 2356 124 2360 156
rect 2320 76 2360 124
rect 2320 44 2324 76
rect 2356 44 2360 76
rect 2320 -4 2360 44
rect 2320 -36 2324 -4
rect 2356 -36 2360 -4
rect 2320 -84 2360 -36
rect 2320 -116 2324 -84
rect 2356 -116 2360 -84
rect 2320 -164 2360 -116
rect 2320 -196 2324 -164
rect 2356 -196 2360 -164
rect 2320 -244 2360 -196
rect 2320 -276 2324 -244
rect 2356 -276 2360 -244
rect 2320 -324 2360 -276
rect 2320 -356 2324 -324
rect 2356 -356 2360 -324
rect 2320 -404 2360 -356
rect 2320 -436 2324 -404
rect 2356 -436 2360 -404
rect 2320 -484 2360 -436
rect 2320 -516 2324 -484
rect 2356 -516 2360 -484
rect 2320 -564 2360 -516
rect 2320 -596 2324 -564
rect 2356 -596 2360 -564
rect 2320 -644 2360 -596
rect 2320 -676 2324 -644
rect 2356 -676 2360 -644
rect 2320 -724 2360 -676
rect 2320 -756 2324 -724
rect 2356 -756 2360 -724
rect 2320 -804 2360 -756
rect 2320 -836 2324 -804
rect 2356 -836 2360 -804
rect 2320 -884 2360 -836
rect 2320 -916 2324 -884
rect 2356 -916 2360 -884
rect 2320 -964 2360 -916
rect 2320 -996 2324 -964
rect 2356 -996 2360 -964
rect 2320 -1044 2360 -996
rect 2320 -1076 2324 -1044
rect 2356 -1076 2360 -1044
rect 2320 -1124 2360 -1076
rect 2320 -1156 2324 -1124
rect 2356 -1156 2360 -1124
rect 2320 -1204 2360 -1156
rect 2320 -1236 2324 -1204
rect 2356 -1236 2360 -1204
rect 2320 -1284 2360 -1236
rect 2320 -1316 2324 -1284
rect 2356 -1316 2360 -1284
rect 2320 -1364 2360 -1316
rect 2320 -1396 2324 -1364
rect 2356 -1396 2360 -1364
rect 2320 -1444 2360 -1396
rect 2320 -1476 2324 -1444
rect 2356 -1476 2360 -1444
rect 2320 -1524 2360 -1476
rect 2320 -1556 2324 -1524
rect 2356 -1556 2360 -1524
rect 2320 -1604 2360 -1556
rect 2320 -1636 2324 -1604
rect 2356 -1636 2360 -1604
rect 2320 -1684 2360 -1636
rect 2320 -1716 2324 -1684
rect 2356 -1716 2360 -1684
rect 2320 -1764 2360 -1716
rect 2320 -1796 2324 -1764
rect 2356 -1796 2360 -1764
rect 2320 -1844 2360 -1796
rect 2320 -1876 2324 -1844
rect 2356 -1876 2360 -1844
rect 2320 -1924 2360 -1876
rect 2320 -1956 2324 -1924
rect 2356 -1956 2360 -1924
rect 2320 -2004 2360 -1956
rect 2320 -2036 2324 -2004
rect 2356 -2036 2360 -2004
rect 2320 -2084 2360 -2036
rect 2320 -2116 2324 -2084
rect 2356 -2116 2360 -2084
rect 2320 -2164 2360 -2116
rect 2320 -2196 2324 -2164
rect 2356 -2196 2360 -2164
rect 2320 -2244 2360 -2196
rect 2320 -2276 2324 -2244
rect 2356 -2276 2360 -2244
rect 2320 -2324 2360 -2276
rect 2320 -2356 2324 -2324
rect 2356 -2356 2360 -2324
rect 2320 -2404 2360 -2356
rect 2320 -2436 2324 -2404
rect 2356 -2436 2360 -2404
rect 2320 -2484 2360 -2436
rect 2320 -2516 2324 -2484
rect 2356 -2516 2360 -2484
rect 2320 -2564 2360 -2516
rect 2320 -2596 2324 -2564
rect 2356 -2596 2360 -2564
rect 2320 -2644 2360 -2596
rect 2320 -2676 2324 -2644
rect 2356 -2676 2360 -2644
rect 2320 -2724 2360 -2676
rect 2320 -2756 2324 -2724
rect 2356 -2756 2360 -2724
rect 2320 -2804 2360 -2756
rect 2320 -2836 2324 -2804
rect 2356 -2836 2360 -2804
rect 2320 -2884 2360 -2836
rect 2320 -2916 2324 -2884
rect 2356 -2916 2360 -2884
rect 2320 -2964 2360 -2916
rect 2320 -2996 2324 -2964
rect 2356 -2996 2360 -2964
rect 2320 -3044 2360 -2996
rect 2320 -3076 2324 -3044
rect 2356 -3076 2360 -3044
rect 2320 -3124 2360 -3076
rect 2320 -3156 2324 -3124
rect 2356 -3156 2360 -3124
rect 2320 -3204 2360 -3156
rect 2320 -3236 2324 -3204
rect 2356 -3236 2360 -3204
rect 2320 -3284 2360 -3236
rect 2320 -3316 2324 -3284
rect 2356 -3316 2360 -3284
rect 2320 -3364 2360 -3316
rect 2320 -3396 2324 -3364
rect 2356 -3396 2360 -3364
rect 2320 -3444 2360 -3396
rect 2320 -3476 2324 -3444
rect 2356 -3476 2360 -3444
rect 2320 -3524 2360 -3476
rect 2320 -3556 2324 -3524
rect 2356 -3556 2360 -3524
rect 2320 -3604 2360 -3556
rect 2320 -3636 2324 -3604
rect 2356 -3636 2360 -3604
rect 2320 -3684 2360 -3636
rect 2320 -3716 2324 -3684
rect 2356 -3716 2360 -3684
rect 2320 -3720 2360 -3716
rect 2400 1036 2440 1040
rect 2400 1004 2404 1036
rect 2436 1004 2440 1036
rect 2400 956 2440 1004
rect 2400 924 2404 956
rect 2436 924 2440 956
rect 2400 876 2440 924
rect 2400 844 2404 876
rect 2436 844 2440 876
rect 2400 796 2440 844
rect 2400 764 2404 796
rect 2436 764 2440 796
rect 2400 716 2440 764
rect 2400 684 2404 716
rect 2436 684 2440 716
rect 2400 636 2440 684
rect 2400 604 2404 636
rect 2436 604 2440 636
rect 2400 556 2440 604
rect 2400 524 2404 556
rect 2436 524 2440 556
rect 2400 476 2440 524
rect 2400 444 2404 476
rect 2436 444 2440 476
rect 2400 396 2440 444
rect 2400 364 2404 396
rect 2436 364 2440 396
rect 2400 316 2440 364
rect 2400 284 2404 316
rect 2436 284 2440 316
rect 2400 236 2440 284
rect 2400 204 2404 236
rect 2436 204 2440 236
rect 2400 156 2440 204
rect 2400 124 2404 156
rect 2436 124 2440 156
rect 2400 76 2440 124
rect 2400 44 2404 76
rect 2436 44 2440 76
rect 2400 -4 2440 44
rect 2400 -36 2404 -4
rect 2436 -36 2440 -4
rect 2400 -84 2440 -36
rect 2400 -116 2404 -84
rect 2436 -116 2440 -84
rect 2400 -164 2440 -116
rect 2400 -196 2404 -164
rect 2436 -196 2440 -164
rect 2400 -244 2440 -196
rect 2400 -276 2404 -244
rect 2436 -276 2440 -244
rect 2400 -324 2440 -276
rect 2400 -356 2404 -324
rect 2436 -356 2440 -324
rect 2400 -404 2440 -356
rect 2400 -436 2404 -404
rect 2436 -436 2440 -404
rect 2400 -484 2440 -436
rect 2400 -516 2404 -484
rect 2436 -516 2440 -484
rect 2400 -564 2440 -516
rect 2400 -596 2404 -564
rect 2436 -596 2440 -564
rect 2400 -644 2440 -596
rect 2400 -676 2404 -644
rect 2436 -676 2440 -644
rect 2400 -724 2440 -676
rect 2400 -756 2404 -724
rect 2436 -756 2440 -724
rect 2400 -804 2440 -756
rect 2400 -836 2404 -804
rect 2436 -836 2440 -804
rect 2400 -884 2440 -836
rect 2400 -916 2404 -884
rect 2436 -916 2440 -884
rect 2400 -964 2440 -916
rect 2400 -996 2404 -964
rect 2436 -996 2440 -964
rect 2400 -1044 2440 -996
rect 2400 -1076 2404 -1044
rect 2436 -1076 2440 -1044
rect 2400 -1124 2440 -1076
rect 2400 -1156 2404 -1124
rect 2436 -1156 2440 -1124
rect 2400 -1204 2440 -1156
rect 2400 -1236 2404 -1204
rect 2436 -1236 2440 -1204
rect 2400 -1284 2440 -1236
rect 2400 -1316 2404 -1284
rect 2436 -1316 2440 -1284
rect 2400 -1364 2440 -1316
rect 2400 -1396 2404 -1364
rect 2436 -1396 2440 -1364
rect 2400 -1444 2440 -1396
rect 2400 -1476 2404 -1444
rect 2436 -1476 2440 -1444
rect 2400 -1524 2440 -1476
rect 2400 -1556 2404 -1524
rect 2436 -1556 2440 -1524
rect 2400 -1604 2440 -1556
rect 2400 -1636 2404 -1604
rect 2436 -1636 2440 -1604
rect 2400 -1684 2440 -1636
rect 2400 -1716 2404 -1684
rect 2436 -1716 2440 -1684
rect 2400 -1764 2440 -1716
rect 2400 -1796 2404 -1764
rect 2436 -1796 2440 -1764
rect 2400 -1844 2440 -1796
rect 2400 -1876 2404 -1844
rect 2436 -1876 2440 -1844
rect 2400 -1924 2440 -1876
rect 2400 -1956 2404 -1924
rect 2436 -1956 2440 -1924
rect 2400 -2004 2440 -1956
rect 2400 -2036 2404 -2004
rect 2436 -2036 2440 -2004
rect 2400 -2084 2440 -2036
rect 2400 -2116 2404 -2084
rect 2436 -2116 2440 -2084
rect 2400 -2164 2440 -2116
rect 2400 -2196 2404 -2164
rect 2436 -2196 2440 -2164
rect 2400 -2244 2440 -2196
rect 2400 -2276 2404 -2244
rect 2436 -2276 2440 -2244
rect 2400 -2324 2440 -2276
rect 2400 -2356 2404 -2324
rect 2436 -2356 2440 -2324
rect 2400 -2404 2440 -2356
rect 2400 -2436 2404 -2404
rect 2436 -2436 2440 -2404
rect 2400 -2484 2440 -2436
rect 2400 -2516 2404 -2484
rect 2436 -2516 2440 -2484
rect 2400 -2564 2440 -2516
rect 2400 -2596 2404 -2564
rect 2436 -2596 2440 -2564
rect 2400 -2644 2440 -2596
rect 2400 -2676 2404 -2644
rect 2436 -2676 2440 -2644
rect 2400 -2724 2440 -2676
rect 2400 -2756 2404 -2724
rect 2436 -2756 2440 -2724
rect 2400 -2804 2440 -2756
rect 2400 -2836 2404 -2804
rect 2436 -2836 2440 -2804
rect 2400 -2884 2440 -2836
rect 2400 -2916 2404 -2884
rect 2436 -2916 2440 -2884
rect 2400 -2964 2440 -2916
rect 2400 -2996 2404 -2964
rect 2436 -2996 2440 -2964
rect 2400 -3044 2440 -2996
rect 2400 -3076 2404 -3044
rect 2436 -3076 2440 -3044
rect 2400 -3124 2440 -3076
rect 2400 -3156 2404 -3124
rect 2436 -3156 2440 -3124
rect 2400 -3204 2440 -3156
rect 2400 -3236 2404 -3204
rect 2436 -3236 2440 -3204
rect 2400 -3284 2440 -3236
rect 2400 -3316 2404 -3284
rect 2436 -3316 2440 -3284
rect 2400 -3364 2440 -3316
rect 2400 -3396 2404 -3364
rect 2436 -3396 2440 -3364
rect 2400 -3444 2440 -3396
rect 2400 -3476 2404 -3444
rect 2436 -3476 2440 -3444
rect 2400 -3524 2440 -3476
rect 2400 -3556 2404 -3524
rect 2436 -3556 2440 -3524
rect 2400 -3604 2440 -3556
rect 2400 -3636 2404 -3604
rect 2436 -3636 2440 -3604
rect 2400 -3684 2440 -3636
rect 2400 -3716 2404 -3684
rect 2436 -3716 2440 -3684
rect 2400 -3720 2440 -3716
rect 2480 1036 2520 1040
rect 2480 1004 2484 1036
rect 2516 1004 2520 1036
rect 2480 956 2520 1004
rect 2480 924 2484 956
rect 2516 924 2520 956
rect 2480 876 2520 924
rect 2480 844 2484 876
rect 2516 844 2520 876
rect 2480 796 2520 844
rect 2480 764 2484 796
rect 2516 764 2520 796
rect 2480 716 2520 764
rect 2480 684 2484 716
rect 2516 684 2520 716
rect 2480 636 2520 684
rect 2480 604 2484 636
rect 2516 604 2520 636
rect 2480 556 2520 604
rect 2480 524 2484 556
rect 2516 524 2520 556
rect 2480 476 2520 524
rect 2480 444 2484 476
rect 2516 444 2520 476
rect 2480 396 2520 444
rect 2480 364 2484 396
rect 2516 364 2520 396
rect 2480 316 2520 364
rect 2480 284 2484 316
rect 2516 284 2520 316
rect 2480 236 2520 284
rect 2480 204 2484 236
rect 2516 204 2520 236
rect 2480 156 2520 204
rect 2480 124 2484 156
rect 2516 124 2520 156
rect 2480 76 2520 124
rect 2480 44 2484 76
rect 2516 44 2520 76
rect 2480 -4 2520 44
rect 2480 -36 2484 -4
rect 2516 -36 2520 -4
rect 2480 -84 2520 -36
rect 2480 -116 2484 -84
rect 2516 -116 2520 -84
rect 2480 -164 2520 -116
rect 2480 -196 2484 -164
rect 2516 -196 2520 -164
rect 2480 -244 2520 -196
rect 2480 -276 2484 -244
rect 2516 -276 2520 -244
rect 2480 -324 2520 -276
rect 2480 -356 2484 -324
rect 2516 -356 2520 -324
rect 2480 -404 2520 -356
rect 2480 -436 2484 -404
rect 2516 -436 2520 -404
rect 2480 -484 2520 -436
rect 2480 -516 2484 -484
rect 2516 -516 2520 -484
rect 2480 -564 2520 -516
rect 2480 -596 2484 -564
rect 2516 -596 2520 -564
rect 2480 -644 2520 -596
rect 2480 -676 2484 -644
rect 2516 -676 2520 -644
rect 2480 -724 2520 -676
rect 2480 -756 2484 -724
rect 2516 -756 2520 -724
rect 2480 -804 2520 -756
rect 2480 -836 2484 -804
rect 2516 -836 2520 -804
rect 2480 -884 2520 -836
rect 2480 -916 2484 -884
rect 2516 -916 2520 -884
rect 2480 -964 2520 -916
rect 2480 -996 2484 -964
rect 2516 -996 2520 -964
rect 2480 -1044 2520 -996
rect 2480 -1076 2484 -1044
rect 2516 -1076 2520 -1044
rect 2480 -1124 2520 -1076
rect 2480 -1156 2484 -1124
rect 2516 -1156 2520 -1124
rect 2480 -1204 2520 -1156
rect 2480 -1236 2484 -1204
rect 2516 -1236 2520 -1204
rect 2480 -1284 2520 -1236
rect 2480 -1316 2484 -1284
rect 2516 -1316 2520 -1284
rect 2480 -1364 2520 -1316
rect 2480 -1396 2484 -1364
rect 2516 -1396 2520 -1364
rect 2480 -1444 2520 -1396
rect 2480 -1476 2484 -1444
rect 2516 -1476 2520 -1444
rect 2480 -1524 2520 -1476
rect 2480 -1556 2484 -1524
rect 2516 -1556 2520 -1524
rect 2480 -1604 2520 -1556
rect 2480 -1636 2484 -1604
rect 2516 -1636 2520 -1604
rect 2480 -1684 2520 -1636
rect 2480 -1716 2484 -1684
rect 2516 -1716 2520 -1684
rect 2480 -1764 2520 -1716
rect 2480 -1796 2484 -1764
rect 2516 -1796 2520 -1764
rect 2480 -1844 2520 -1796
rect 2480 -1876 2484 -1844
rect 2516 -1876 2520 -1844
rect 2480 -1924 2520 -1876
rect 2480 -1956 2484 -1924
rect 2516 -1956 2520 -1924
rect 2480 -2004 2520 -1956
rect 2480 -2036 2484 -2004
rect 2516 -2036 2520 -2004
rect 2480 -2084 2520 -2036
rect 2480 -2116 2484 -2084
rect 2516 -2116 2520 -2084
rect 2480 -2164 2520 -2116
rect 2480 -2196 2484 -2164
rect 2516 -2196 2520 -2164
rect 2480 -2244 2520 -2196
rect 2480 -2276 2484 -2244
rect 2516 -2276 2520 -2244
rect 2480 -2324 2520 -2276
rect 2480 -2356 2484 -2324
rect 2516 -2356 2520 -2324
rect 2480 -2404 2520 -2356
rect 2480 -2436 2484 -2404
rect 2516 -2436 2520 -2404
rect 2480 -2484 2520 -2436
rect 2480 -2516 2484 -2484
rect 2516 -2516 2520 -2484
rect 2480 -2564 2520 -2516
rect 2480 -2596 2484 -2564
rect 2516 -2596 2520 -2564
rect 2480 -2644 2520 -2596
rect 2480 -2676 2484 -2644
rect 2516 -2676 2520 -2644
rect 2480 -2724 2520 -2676
rect 2480 -2756 2484 -2724
rect 2516 -2756 2520 -2724
rect 2480 -2804 2520 -2756
rect 2480 -2836 2484 -2804
rect 2516 -2836 2520 -2804
rect 2480 -2884 2520 -2836
rect 2480 -2916 2484 -2884
rect 2516 -2916 2520 -2884
rect 2480 -2964 2520 -2916
rect 2480 -2996 2484 -2964
rect 2516 -2996 2520 -2964
rect 2480 -3044 2520 -2996
rect 2480 -3076 2484 -3044
rect 2516 -3076 2520 -3044
rect 2480 -3124 2520 -3076
rect 2480 -3156 2484 -3124
rect 2516 -3156 2520 -3124
rect 2480 -3204 2520 -3156
rect 2480 -3236 2484 -3204
rect 2516 -3236 2520 -3204
rect 2480 -3284 2520 -3236
rect 2480 -3316 2484 -3284
rect 2516 -3316 2520 -3284
rect 2480 -3364 2520 -3316
rect 2480 -3396 2484 -3364
rect 2516 -3396 2520 -3364
rect 2480 -3444 2520 -3396
rect 2480 -3476 2484 -3444
rect 2516 -3476 2520 -3444
rect 2480 -3524 2520 -3476
rect 2480 -3556 2484 -3524
rect 2516 -3556 2520 -3524
rect 2480 -3604 2520 -3556
rect 2480 -3636 2484 -3604
rect 2516 -3636 2520 -3604
rect 2480 -3684 2520 -3636
rect 2480 -3716 2484 -3684
rect 2516 -3716 2520 -3684
rect 2480 -3720 2520 -3716
rect 2560 1036 2600 1040
rect 2560 1004 2564 1036
rect 2596 1004 2600 1036
rect 2560 956 2600 1004
rect 2560 924 2564 956
rect 2596 924 2600 956
rect 2560 876 2600 924
rect 2560 844 2564 876
rect 2596 844 2600 876
rect 2560 796 2600 844
rect 2560 764 2564 796
rect 2596 764 2600 796
rect 2560 716 2600 764
rect 2560 684 2564 716
rect 2596 684 2600 716
rect 2560 636 2600 684
rect 2560 604 2564 636
rect 2596 604 2600 636
rect 2560 556 2600 604
rect 2560 524 2564 556
rect 2596 524 2600 556
rect 2560 476 2600 524
rect 2560 444 2564 476
rect 2596 444 2600 476
rect 2560 396 2600 444
rect 2560 364 2564 396
rect 2596 364 2600 396
rect 2560 316 2600 364
rect 2560 284 2564 316
rect 2596 284 2600 316
rect 2560 236 2600 284
rect 2560 204 2564 236
rect 2596 204 2600 236
rect 2560 156 2600 204
rect 2560 124 2564 156
rect 2596 124 2600 156
rect 2560 76 2600 124
rect 2560 44 2564 76
rect 2596 44 2600 76
rect 2560 -4 2600 44
rect 2560 -36 2564 -4
rect 2596 -36 2600 -4
rect 2560 -84 2600 -36
rect 2560 -116 2564 -84
rect 2596 -116 2600 -84
rect 2560 -164 2600 -116
rect 2560 -196 2564 -164
rect 2596 -196 2600 -164
rect 2560 -244 2600 -196
rect 2560 -276 2564 -244
rect 2596 -276 2600 -244
rect 2560 -324 2600 -276
rect 2560 -356 2564 -324
rect 2596 -356 2600 -324
rect 2560 -404 2600 -356
rect 2560 -436 2564 -404
rect 2596 -436 2600 -404
rect 2560 -484 2600 -436
rect 2560 -516 2564 -484
rect 2596 -516 2600 -484
rect 2560 -564 2600 -516
rect 2560 -596 2564 -564
rect 2596 -596 2600 -564
rect 2560 -644 2600 -596
rect 2560 -676 2564 -644
rect 2596 -676 2600 -644
rect 2560 -724 2600 -676
rect 2560 -756 2564 -724
rect 2596 -756 2600 -724
rect 2560 -804 2600 -756
rect 2560 -836 2564 -804
rect 2596 -836 2600 -804
rect 2560 -884 2600 -836
rect 2560 -916 2564 -884
rect 2596 -916 2600 -884
rect 2560 -964 2600 -916
rect 2560 -996 2564 -964
rect 2596 -996 2600 -964
rect 2560 -1044 2600 -996
rect 2560 -1076 2564 -1044
rect 2596 -1076 2600 -1044
rect 2560 -1124 2600 -1076
rect 2560 -1156 2564 -1124
rect 2596 -1156 2600 -1124
rect 2560 -1204 2600 -1156
rect 2560 -1236 2564 -1204
rect 2596 -1236 2600 -1204
rect 2560 -1284 2600 -1236
rect 2560 -1316 2564 -1284
rect 2596 -1316 2600 -1284
rect 2560 -1364 2600 -1316
rect 2560 -1396 2564 -1364
rect 2596 -1396 2600 -1364
rect 2560 -1444 2600 -1396
rect 2560 -1476 2564 -1444
rect 2596 -1476 2600 -1444
rect 2560 -1524 2600 -1476
rect 2560 -1556 2564 -1524
rect 2596 -1556 2600 -1524
rect 2560 -1604 2600 -1556
rect 2560 -1636 2564 -1604
rect 2596 -1636 2600 -1604
rect 2560 -1684 2600 -1636
rect 2560 -1716 2564 -1684
rect 2596 -1716 2600 -1684
rect 2560 -1764 2600 -1716
rect 2560 -1796 2564 -1764
rect 2596 -1796 2600 -1764
rect 2560 -1844 2600 -1796
rect 2560 -1876 2564 -1844
rect 2596 -1876 2600 -1844
rect 2560 -1924 2600 -1876
rect 2560 -1956 2564 -1924
rect 2596 -1956 2600 -1924
rect 2560 -2004 2600 -1956
rect 2560 -2036 2564 -2004
rect 2596 -2036 2600 -2004
rect 2560 -2084 2600 -2036
rect 2560 -2116 2564 -2084
rect 2596 -2116 2600 -2084
rect 2560 -2164 2600 -2116
rect 2560 -2196 2564 -2164
rect 2596 -2196 2600 -2164
rect 2560 -2244 2600 -2196
rect 2560 -2276 2564 -2244
rect 2596 -2276 2600 -2244
rect 2560 -2324 2600 -2276
rect 2560 -2356 2564 -2324
rect 2596 -2356 2600 -2324
rect 2560 -2404 2600 -2356
rect 2560 -2436 2564 -2404
rect 2596 -2436 2600 -2404
rect 2560 -2484 2600 -2436
rect 2560 -2516 2564 -2484
rect 2596 -2516 2600 -2484
rect 2560 -2564 2600 -2516
rect 2560 -2596 2564 -2564
rect 2596 -2596 2600 -2564
rect 2560 -2644 2600 -2596
rect 2560 -2676 2564 -2644
rect 2596 -2676 2600 -2644
rect 2560 -2724 2600 -2676
rect 2560 -2756 2564 -2724
rect 2596 -2756 2600 -2724
rect 2560 -2804 2600 -2756
rect 2560 -2836 2564 -2804
rect 2596 -2836 2600 -2804
rect 2560 -2884 2600 -2836
rect 2560 -2916 2564 -2884
rect 2596 -2916 2600 -2884
rect 2560 -2964 2600 -2916
rect 2560 -2996 2564 -2964
rect 2596 -2996 2600 -2964
rect 2560 -3044 2600 -2996
rect 2560 -3076 2564 -3044
rect 2596 -3076 2600 -3044
rect 2560 -3124 2600 -3076
rect 2560 -3156 2564 -3124
rect 2596 -3156 2600 -3124
rect 2560 -3204 2600 -3156
rect 2560 -3236 2564 -3204
rect 2596 -3236 2600 -3204
rect 2560 -3284 2600 -3236
rect 2560 -3316 2564 -3284
rect 2596 -3316 2600 -3284
rect 2560 -3364 2600 -3316
rect 2560 -3396 2564 -3364
rect 2596 -3396 2600 -3364
rect 2560 -3444 2600 -3396
rect 2560 -3476 2564 -3444
rect 2596 -3476 2600 -3444
rect 2560 -3524 2600 -3476
rect 2560 -3556 2564 -3524
rect 2596 -3556 2600 -3524
rect 2560 -3604 2600 -3556
rect 2560 -3636 2564 -3604
rect 2596 -3636 2600 -3604
rect 2560 -3684 2600 -3636
rect 2560 -3716 2564 -3684
rect 2596 -3716 2600 -3684
rect 2560 -3720 2600 -3716
rect 2640 1036 2680 1040
rect 2640 1004 2644 1036
rect 2676 1004 2680 1036
rect 2640 956 2680 1004
rect 2640 924 2644 956
rect 2676 924 2680 956
rect 2640 876 2680 924
rect 2640 844 2644 876
rect 2676 844 2680 876
rect 2640 796 2680 844
rect 2640 764 2644 796
rect 2676 764 2680 796
rect 2640 716 2680 764
rect 2640 684 2644 716
rect 2676 684 2680 716
rect 2640 636 2680 684
rect 2640 604 2644 636
rect 2676 604 2680 636
rect 2640 556 2680 604
rect 2640 524 2644 556
rect 2676 524 2680 556
rect 2640 476 2680 524
rect 2640 444 2644 476
rect 2676 444 2680 476
rect 2640 396 2680 444
rect 2640 364 2644 396
rect 2676 364 2680 396
rect 2640 316 2680 364
rect 2640 284 2644 316
rect 2676 284 2680 316
rect 2640 236 2680 284
rect 2640 204 2644 236
rect 2676 204 2680 236
rect 2640 156 2680 204
rect 2640 124 2644 156
rect 2676 124 2680 156
rect 2640 76 2680 124
rect 2640 44 2644 76
rect 2676 44 2680 76
rect 2640 -4 2680 44
rect 2640 -36 2644 -4
rect 2676 -36 2680 -4
rect 2640 -84 2680 -36
rect 2640 -116 2644 -84
rect 2676 -116 2680 -84
rect 2640 -164 2680 -116
rect 2640 -196 2644 -164
rect 2676 -196 2680 -164
rect 2640 -244 2680 -196
rect 2640 -276 2644 -244
rect 2676 -276 2680 -244
rect 2640 -324 2680 -276
rect 2640 -356 2644 -324
rect 2676 -356 2680 -324
rect 2640 -404 2680 -356
rect 2640 -436 2644 -404
rect 2676 -436 2680 -404
rect 2640 -484 2680 -436
rect 2640 -516 2644 -484
rect 2676 -516 2680 -484
rect 2640 -564 2680 -516
rect 2640 -596 2644 -564
rect 2676 -596 2680 -564
rect 2640 -644 2680 -596
rect 2640 -676 2644 -644
rect 2676 -676 2680 -644
rect 2640 -724 2680 -676
rect 2640 -756 2644 -724
rect 2676 -756 2680 -724
rect 2640 -804 2680 -756
rect 2640 -836 2644 -804
rect 2676 -836 2680 -804
rect 2640 -884 2680 -836
rect 2640 -916 2644 -884
rect 2676 -916 2680 -884
rect 2640 -964 2680 -916
rect 2640 -996 2644 -964
rect 2676 -996 2680 -964
rect 2640 -1044 2680 -996
rect 2640 -1076 2644 -1044
rect 2676 -1076 2680 -1044
rect 2640 -1124 2680 -1076
rect 2640 -1156 2644 -1124
rect 2676 -1156 2680 -1124
rect 2640 -1204 2680 -1156
rect 2640 -1236 2644 -1204
rect 2676 -1236 2680 -1204
rect 2640 -1284 2680 -1236
rect 2640 -1316 2644 -1284
rect 2676 -1316 2680 -1284
rect 2640 -1364 2680 -1316
rect 2640 -1396 2644 -1364
rect 2676 -1396 2680 -1364
rect 2640 -1444 2680 -1396
rect 2640 -1476 2644 -1444
rect 2676 -1476 2680 -1444
rect 2640 -1524 2680 -1476
rect 2640 -1556 2644 -1524
rect 2676 -1556 2680 -1524
rect 2640 -1604 2680 -1556
rect 2640 -1636 2644 -1604
rect 2676 -1636 2680 -1604
rect 2640 -1684 2680 -1636
rect 2640 -1716 2644 -1684
rect 2676 -1716 2680 -1684
rect 2640 -1764 2680 -1716
rect 2640 -1796 2644 -1764
rect 2676 -1796 2680 -1764
rect 2640 -1844 2680 -1796
rect 2640 -1876 2644 -1844
rect 2676 -1876 2680 -1844
rect 2640 -1924 2680 -1876
rect 2640 -1956 2644 -1924
rect 2676 -1956 2680 -1924
rect 2640 -2004 2680 -1956
rect 2640 -2036 2644 -2004
rect 2676 -2036 2680 -2004
rect 2640 -2084 2680 -2036
rect 2640 -2116 2644 -2084
rect 2676 -2116 2680 -2084
rect 2640 -2164 2680 -2116
rect 2640 -2196 2644 -2164
rect 2676 -2196 2680 -2164
rect 2640 -2244 2680 -2196
rect 2640 -2276 2644 -2244
rect 2676 -2276 2680 -2244
rect 2640 -2324 2680 -2276
rect 2640 -2356 2644 -2324
rect 2676 -2356 2680 -2324
rect 2640 -2404 2680 -2356
rect 2640 -2436 2644 -2404
rect 2676 -2436 2680 -2404
rect 2640 -2484 2680 -2436
rect 2640 -2516 2644 -2484
rect 2676 -2516 2680 -2484
rect 2640 -2564 2680 -2516
rect 2640 -2596 2644 -2564
rect 2676 -2596 2680 -2564
rect 2640 -2644 2680 -2596
rect 2640 -2676 2644 -2644
rect 2676 -2676 2680 -2644
rect 2640 -2724 2680 -2676
rect 2640 -2756 2644 -2724
rect 2676 -2756 2680 -2724
rect 2640 -2804 2680 -2756
rect 2640 -2836 2644 -2804
rect 2676 -2836 2680 -2804
rect 2640 -2884 2680 -2836
rect 2640 -2916 2644 -2884
rect 2676 -2916 2680 -2884
rect 2640 -2964 2680 -2916
rect 2640 -2996 2644 -2964
rect 2676 -2996 2680 -2964
rect 2640 -3044 2680 -2996
rect 2640 -3076 2644 -3044
rect 2676 -3076 2680 -3044
rect 2640 -3124 2680 -3076
rect 2640 -3156 2644 -3124
rect 2676 -3156 2680 -3124
rect 2640 -3204 2680 -3156
rect 2640 -3236 2644 -3204
rect 2676 -3236 2680 -3204
rect 2640 -3284 2680 -3236
rect 2640 -3316 2644 -3284
rect 2676 -3316 2680 -3284
rect 2640 -3364 2680 -3316
rect 2640 -3396 2644 -3364
rect 2676 -3396 2680 -3364
rect 2640 -3444 2680 -3396
rect 2640 -3476 2644 -3444
rect 2676 -3476 2680 -3444
rect 2640 -3524 2680 -3476
rect 2640 -3556 2644 -3524
rect 2676 -3556 2680 -3524
rect 2640 -3604 2680 -3556
rect 2640 -3636 2644 -3604
rect 2676 -3636 2680 -3604
rect 2640 -3684 2680 -3636
rect 2640 -3716 2644 -3684
rect 2676 -3716 2680 -3684
rect 2640 -3720 2680 -3716
rect 2720 1036 2760 1040
rect 2720 1004 2724 1036
rect 2756 1004 2760 1036
rect 2720 956 2760 1004
rect 2720 924 2724 956
rect 2756 924 2760 956
rect 2720 876 2760 924
rect 2720 844 2724 876
rect 2756 844 2760 876
rect 2720 796 2760 844
rect 2720 764 2724 796
rect 2756 764 2760 796
rect 2720 716 2760 764
rect 2720 684 2724 716
rect 2756 684 2760 716
rect 2720 636 2760 684
rect 2720 604 2724 636
rect 2756 604 2760 636
rect 2720 556 2760 604
rect 2720 524 2724 556
rect 2756 524 2760 556
rect 2720 476 2760 524
rect 2720 444 2724 476
rect 2756 444 2760 476
rect 2720 396 2760 444
rect 2720 364 2724 396
rect 2756 364 2760 396
rect 2720 316 2760 364
rect 2720 284 2724 316
rect 2756 284 2760 316
rect 2720 236 2760 284
rect 2720 204 2724 236
rect 2756 204 2760 236
rect 2720 156 2760 204
rect 2720 124 2724 156
rect 2756 124 2760 156
rect 2720 76 2760 124
rect 2720 44 2724 76
rect 2756 44 2760 76
rect 2720 -4 2760 44
rect 2720 -36 2724 -4
rect 2756 -36 2760 -4
rect 2720 -84 2760 -36
rect 2720 -116 2724 -84
rect 2756 -116 2760 -84
rect 2720 -164 2760 -116
rect 2720 -196 2724 -164
rect 2756 -196 2760 -164
rect 2720 -244 2760 -196
rect 2720 -276 2724 -244
rect 2756 -276 2760 -244
rect 2720 -324 2760 -276
rect 2720 -356 2724 -324
rect 2756 -356 2760 -324
rect 2720 -404 2760 -356
rect 2720 -436 2724 -404
rect 2756 -436 2760 -404
rect 2720 -484 2760 -436
rect 2720 -516 2724 -484
rect 2756 -516 2760 -484
rect 2720 -564 2760 -516
rect 2720 -596 2724 -564
rect 2756 -596 2760 -564
rect 2720 -644 2760 -596
rect 2720 -676 2724 -644
rect 2756 -676 2760 -644
rect 2720 -724 2760 -676
rect 2720 -756 2724 -724
rect 2756 -756 2760 -724
rect 2720 -804 2760 -756
rect 2720 -836 2724 -804
rect 2756 -836 2760 -804
rect 2720 -884 2760 -836
rect 2720 -916 2724 -884
rect 2756 -916 2760 -884
rect 2720 -964 2760 -916
rect 2720 -996 2724 -964
rect 2756 -996 2760 -964
rect 2720 -1044 2760 -996
rect 2720 -1076 2724 -1044
rect 2756 -1076 2760 -1044
rect 2720 -1124 2760 -1076
rect 2720 -1156 2724 -1124
rect 2756 -1156 2760 -1124
rect 2720 -1204 2760 -1156
rect 2720 -1236 2724 -1204
rect 2756 -1236 2760 -1204
rect 2720 -1284 2760 -1236
rect 2720 -1316 2724 -1284
rect 2756 -1316 2760 -1284
rect 2720 -1364 2760 -1316
rect 2720 -1396 2724 -1364
rect 2756 -1396 2760 -1364
rect 2720 -1444 2760 -1396
rect 2720 -1476 2724 -1444
rect 2756 -1476 2760 -1444
rect 2720 -1524 2760 -1476
rect 2720 -1556 2724 -1524
rect 2756 -1556 2760 -1524
rect 2720 -1604 2760 -1556
rect 2720 -1636 2724 -1604
rect 2756 -1636 2760 -1604
rect 2720 -1684 2760 -1636
rect 2720 -1716 2724 -1684
rect 2756 -1716 2760 -1684
rect 2720 -1764 2760 -1716
rect 2720 -1796 2724 -1764
rect 2756 -1796 2760 -1764
rect 2720 -1844 2760 -1796
rect 2720 -1876 2724 -1844
rect 2756 -1876 2760 -1844
rect 2720 -1924 2760 -1876
rect 2720 -1956 2724 -1924
rect 2756 -1956 2760 -1924
rect 2720 -2004 2760 -1956
rect 2720 -2036 2724 -2004
rect 2756 -2036 2760 -2004
rect 2720 -2084 2760 -2036
rect 2720 -2116 2724 -2084
rect 2756 -2116 2760 -2084
rect 2720 -2164 2760 -2116
rect 2720 -2196 2724 -2164
rect 2756 -2196 2760 -2164
rect 2720 -2244 2760 -2196
rect 2720 -2276 2724 -2244
rect 2756 -2276 2760 -2244
rect 2720 -2324 2760 -2276
rect 2720 -2356 2724 -2324
rect 2756 -2356 2760 -2324
rect 2720 -2404 2760 -2356
rect 2720 -2436 2724 -2404
rect 2756 -2436 2760 -2404
rect 2720 -2484 2760 -2436
rect 2720 -2516 2724 -2484
rect 2756 -2516 2760 -2484
rect 2720 -2564 2760 -2516
rect 2720 -2596 2724 -2564
rect 2756 -2596 2760 -2564
rect 2720 -2644 2760 -2596
rect 2720 -2676 2724 -2644
rect 2756 -2676 2760 -2644
rect 2720 -2724 2760 -2676
rect 2720 -2756 2724 -2724
rect 2756 -2756 2760 -2724
rect 2720 -2804 2760 -2756
rect 2720 -2836 2724 -2804
rect 2756 -2836 2760 -2804
rect 2720 -2884 2760 -2836
rect 2720 -2916 2724 -2884
rect 2756 -2916 2760 -2884
rect 2720 -2964 2760 -2916
rect 2720 -2996 2724 -2964
rect 2756 -2996 2760 -2964
rect 2720 -3044 2760 -2996
rect 2720 -3076 2724 -3044
rect 2756 -3076 2760 -3044
rect 2720 -3124 2760 -3076
rect 2720 -3156 2724 -3124
rect 2756 -3156 2760 -3124
rect 2720 -3204 2760 -3156
rect 2720 -3236 2724 -3204
rect 2756 -3236 2760 -3204
rect 2720 -3284 2760 -3236
rect 2720 -3316 2724 -3284
rect 2756 -3316 2760 -3284
rect 2720 -3364 2760 -3316
rect 2720 -3396 2724 -3364
rect 2756 -3396 2760 -3364
rect 2720 -3444 2760 -3396
rect 2720 -3476 2724 -3444
rect 2756 -3476 2760 -3444
rect 2720 -3524 2760 -3476
rect 2720 -3556 2724 -3524
rect 2756 -3556 2760 -3524
rect 2720 -3604 2760 -3556
rect 2720 -3636 2724 -3604
rect 2756 -3636 2760 -3604
rect 2720 -3684 2760 -3636
rect 2720 -3716 2724 -3684
rect 2756 -3716 2760 -3684
rect 2720 -3720 2760 -3716
rect 2800 1036 2840 1040
rect 2800 1004 2804 1036
rect 2836 1004 2840 1036
rect 2800 956 2840 1004
rect 2800 924 2804 956
rect 2836 924 2840 956
rect 2800 876 2840 924
rect 2800 844 2804 876
rect 2836 844 2840 876
rect 2800 796 2840 844
rect 2800 764 2804 796
rect 2836 764 2840 796
rect 2800 716 2840 764
rect 2800 684 2804 716
rect 2836 684 2840 716
rect 2800 636 2840 684
rect 2800 604 2804 636
rect 2836 604 2840 636
rect 2800 556 2840 604
rect 2800 524 2804 556
rect 2836 524 2840 556
rect 2800 476 2840 524
rect 2800 444 2804 476
rect 2836 444 2840 476
rect 2800 396 2840 444
rect 2800 364 2804 396
rect 2836 364 2840 396
rect 2800 316 2840 364
rect 2800 284 2804 316
rect 2836 284 2840 316
rect 2800 236 2840 284
rect 2800 204 2804 236
rect 2836 204 2840 236
rect 2800 156 2840 204
rect 2800 124 2804 156
rect 2836 124 2840 156
rect 2800 76 2840 124
rect 2800 44 2804 76
rect 2836 44 2840 76
rect 2800 -4 2840 44
rect 2800 -36 2804 -4
rect 2836 -36 2840 -4
rect 2800 -84 2840 -36
rect 2800 -116 2804 -84
rect 2836 -116 2840 -84
rect 2800 -164 2840 -116
rect 2800 -196 2804 -164
rect 2836 -196 2840 -164
rect 2800 -244 2840 -196
rect 2800 -276 2804 -244
rect 2836 -276 2840 -244
rect 2800 -324 2840 -276
rect 2800 -356 2804 -324
rect 2836 -356 2840 -324
rect 2800 -404 2840 -356
rect 2800 -436 2804 -404
rect 2836 -436 2840 -404
rect 2800 -484 2840 -436
rect 2800 -516 2804 -484
rect 2836 -516 2840 -484
rect 2800 -564 2840 -516
rect 2800 -596 2804 -564
rect 2836 -596 2840 -564
rect 2800 -644 2840 -596
rect 2800 -676 2804 -644
rect 2836 -676 2840 -644
rect 2800 -724 2840 -676
rect 2800 -756 2804 -724
rect 2836 -756 2840 -724
rect 2800 -804 2840 -756
rect 2800 -836 2804 -804
rect 2836 -836 2840 -804
rect 2800 -884 2840 -836
rect 2800 -916 2804 -884
rect 2836 -916 2840 -884
rect 2800 -964 2840 -916
rect 2800 -996 2804 -964
rect 2836 -996 2840 -964
rect 2800 -1044 2840 -996
rect 2800 -1076 2804 -1044
rect 2836 -1076 2840 -1044
rect 2800 -1124 2840 -1076
rect 2800 -1156 2804 -1124
rect 2836 -1156 2840 -1124
rect 2800 -1204 2840 -1156
rect 2800 -1236 2804 -1204
rect 2836 -1236 2840 -1204
rect 2800 -1284 2840 -1236
rect 2800 -1316 2804 -1284
rect 2836 -1316 2840 -1284
rect 2800 -1364 2840 -1316
rect 2800 -1396 2804 -1364
rect 2836 -1396 2840 -1364
rect 2800 -1444 2840 -1396
rect 2800 -1476 2804 -1444
rect 2836 -1476 2840 -1444
rect 2800 -1524 2840 -1476
rect 2800 -1556 2804 -1524
rect 2836 -1556 2840 -1524
rect 2800 -1604 2840 -1556
rect 2800 -1636 2804 -1604
rect 2836 -1636 2840 -1604
rect 2800 -1684 2840 -1636
rect 2800 -1716 2804 -1684
rect 2836 -1716 2840 -1684
rect 2800 -1764 2840 -1716
rect 2800 -1796 2804 -1764
rect 2836 -1796 2840 -1764
rect 2800 -1844 2840 -1796
rect 2800 -1876 2804 -1844
rect 2836 -1876 2840 -1844
rect 2800 -1924 2840 -1876
rect 2800 -1956 2804 -1924
rect 2836 -1956 2840 -1924
rect 2800 -2004 2840 -1956
rect 2800 -2036 2804 -2004
rect 2836 -2036 2840 -2004
rect 2800 -2084 2840 -2036
rect 2800 -2116 2804 -2084
rect 2836 -2116 2840 -2084
rect 2800 -2164 2840 -2116
rect 2800 -2196 2804 -2164
rect 2836 -2196 2840 -2164
rect 2800 -2244 2840 -2196
rect 2800 -2276 2804 -2244
rect 2836 -2276 2840 -2244
rect 2800 -2324 2840 -2276
rect 2800 -2356 2804 -2324
rect 2836 -2356 2840 -2324
rect 2800 -2404 2840 -2356
rect 2800 -2436 2804 -2404
rect 2836 -2436 2840 -2404
rect 2800 -2484 2840 -2436
rect 2800 -2516 2804 -2484
rect 2836 -2516 2840 -2484
rect 2800 -2564 2840 -2516
rect 2800 -2596 2804 -2564
rect 2836 -2596 2840 -2564
rect 2800 -2644 2840 -2596
rect 2800 -2676 2804 -2644
rect 2836 -2676 2840 -2644
rect 2800 -2724 2840 -2676
rect 2800 -2756 2804 -2724
rect 2836 -2756 2840 -2724
rect 2800 -2804 2840 -2756
rect 2800 -2836 2804 -2804
rect 2836 -2836 2840 -2804
rect 2800 -2884 2840 -2836
rect 2800 -2916 2804 -2884
rect 2836 -2916 2840 -2884
rect 2800 -2964 2840 -2916
rect 2800 -2996 2804 -2964
rect 2836 -2996 2840 -2964
rect 2800 -3044 2840 -2996
rect 2800 -3076 2804 -3044
rect 2836 -3076 2840 -3044
rect 2800 -3124 2840 -3076
rect 2800 -3156 2804 -3124
rect 2836 -3156 2840 -3124
rect 2800 -3204 2840 -3156
rect 2800 -3236 2804 -3204
rect 2836 -3236 2840 -3204
rect 2800 -3284 2840 -3236
rect 2800 -3316 2804 -3284
rect 2836 -3316 2840 -3284
rect 2800 -3364 2840 -3316
rect 2800 -3396 2804 -3364
rect 2836 -3396 2840 -3364
rect 2800 -3444 2840 -3396
rect 2800 -3476 2804 -3444
rect 2836 -3476 2840 -3444
rect 2800 -3524 2840 -3476
rect 2800 -3556 2804 -3524
rect 2836 -3556 2840 -3524
rect 2800 -3604 2840 -3556
rect 2800 -3636 2804 -3604
rect 2836 -3636 2840 -3604
rect 2800 -3684 2840 -3636
rect 2800 -3716 2804 -3684
rect 2836 -3716 2840 -3684
rect 2800 -3720 2840 -3716
rect 2880 1036 2920 1040
rect 2880 1004 2884 1036
rect 2916 1004 2920 1036
rect 2880 956 2920 1004
rect 2880 924 2884 956
rect 2916 924 2920 956
rect 2880 876 2920 924
rect 2880 844 2884 876
rect 2916 844 2920 876
rect 2880 796 2920 844
rect 2880 764 2884 796
rect 2916 764 2920 796
rect 2880 716 2920 764
rect 2880 684 2884 716
rect 2916 684 2920 716
rect 2880 636 2920 684
rect 2880 604 2884 636
rect 2916 604 2920 636
rect 2880 556 2920 604
rect 2880 524 2884 556
rect 2916 524 2920 556
rect 2880 476 2920 524
rect 2880 444 2884 476
rect 2916 444 2920 476
rect 2880 396 2920 444
rect 2880 364 2884 396
rect 2916 364 2920 396
rect 2880 316 2920 364
rect 2880 284 2884 316
rect 2916 284 2920 316
rect 2880 236 2920 284
rect 2880 204 2884 236
rect 2916 204 2920 236
rect 2880 156 2920 204
rect 2880 124 2884 156
rect 2916 124 2920 156
rect 2880 76 2920 124
rect 2880 44 2884 76
rect 2916 44 2920 76
rect 2880 -4 2920 44
rect 2880 -36 2884 -4
rect 2916 -36 2920 -4
rect 2880 -84 2920 -36
rect 2880 -116 2884 -84
rect 2916 -116 2920 -84
rect 2880 -164 2920 -116
rect 2880 -196 2884 -164
rect 2916 -196 2920 -164
rect 2880 -244 2920 -196
rect 2880 -276 2884 -244
rect 2916 -276 2920 -244
rect 2880 -324 2920 -276
rect 2880 -356 2884 -324
rect 2916 -356 2920 -324
rect 2880 -404 2920 -356
rect 2880 -436 2884 -404
rect 2916 -436 2920 -404
rect 2880 -484 2920 -436
rect 2880 -516 2884 -484
rect 2916 -516 2920 -484
rect 2880 -564 2920 -516
rect 2880 -596 2884 -564
rect 2916 -596 2920 -564
rect 2880 -644 2920 -596
rect 2880 -676 2884 -644
rect 2916 -676 2920 -644
rect 2880 -724 2920 -676
rect 2880 -756 2884 -724
rect 2916 -756 2920 -724
rect 2880 -804 2920 -756
rect 2880 -836 2884 -804
rect 2916 -836 2920 -804
rect 2880 -884 2920 -836
rect 2880 -916 2884 -884
rect 2916 -916 2920 -884
rect 2880 -964 2920 -916
rect 2880 -996 2884 -964
rect 2916 -996 2920 -964
rect 2880 -1044 2920 -996
rect 2880 -1076 2884 -1044
rect 2916 -1076 2920 -1044
rect 2880 -1124 2920 -1076
rect 2880 -1156 2884 -1124
rect 2916 -1156 2920 -1124
rect 2880 -1204 2920 -1156
rect 2880 -1236 2884 -1204
rect 2916 -1236 2920 -1204
rect 2880 -1284 2920 -1236
rect 2880 -1316 2884 -1284
rect 2916 -1316 2920 -1284
rect 2880 -1364 2920 -1316
rect 2880 -1396 2884 -1364
rect 2916 -1396 2920 -1364
rect 2880 -1444 2920 -1396
rect 2880 -1476 2884 -1444
rect 2916 -1476 2920 -1444
rect 2880 -1524 2920 -1476
rect 2880 -1556 2884 -1524
rect 2916 -1556 2920 -1524
rect 2880 -1604 2920 -1556
rect 2880 -1636 2884 -1604
rect 2916 -1636 2920 -1604
rect 2880 -1684 2920 -1636
rect 2880 -1716 2884 -1684
rect 2916 -1716 2920 -1684
rect 2880 -1764 2920 -1716
rect 2880 -1796 2884 -1764
rect 2916 -1796 2920 -1764
rect 2880 -1844 2920 -1796
rect 2880 -1876 2884 -1844
rect 2916 -1876 2920 -1844
rect 2880 -1924 2920 -1876
rect 2880 -1956 2884 -1924
rect 2916 -1956 2920 -1924
rect 2880 -2004 2920 -1956
rect 2880 -2036 2884 -2004
rect 2916 -2036 2920 -2004
rect 2880 -2084 2920 -2036
rect 2880 -2116 2884 -2084
rect 2916 -2116 2920 -2084
rect 2880 -2164 2920 -2116
rect 2880 -2196 2884 -2164
rect 2916 -2196 2920 -2164
rect 2880 -2244 2920 -2196
rect 2880 -2276 2884 -2244
rect 2916 -2276 2920 -2244
rect 2880 -2324 2920 -2276
rect 2880 -2356 2884 -2324
rect 2916 -2356 2920 -2324
rect 2880 -2404 2920 -2356
rect 2880 -2436 2884 -2404
rect 2916 -2436 2920 -2404
rect 2880 -2484 2920 -2436
rect 2880 -2516 2884 -2484
rect 2916 -2516 2920 -2484
rect 2880 -2564 2920 -2516
rect 2880 -2596 2884 -2564
rect 2916 -2596 2920 -2564
rect 2880 -2644 2920 -2596
rect 2880 -2676 2884 -2644
rect 2916 -2676 2920 -2644
rect 2880 -2724 2920 -2676
rect 2880 -2756 2884 -2724
rect 2916 -2756 2920 -2724
rect 2880 -2804 2920 -2756
rect 2880 -2836 2884 -2804
rect 2916 -2836 2920 -2804
rect 2880 -2884 2920 -2836
rect 2880 -2916 2884 -2884
rect 2916 -2916 2920 -2884
rect 2880 -2964 2920 -2916
rect 2880 -2996 2884 -2964
rect 2916 -2996 2920 -2964
rect 2880 -3044 2920 -2996
rect 2880 -3076 2884 -3044
rect 2916 -3076 2920 -3044
rect 2880 -3124 2920 -3076
rect 2880 -3156 2884 -3124
rect 2916 -3156 2920 -3124
rect 2880 -3204 2920 -3156
rect 2880 -3236 2884 -3204
rect 2916 -3236 2920 -3204
rect 2880 -3284 2920 -3236
rect 2880 -3316 2884 -3284
rect 2916 -3316 2920 -3284
rect 2880 -3364 2920 -3316
rect 2880 -3396 2884 -3364
rect 2916 -3396 2920 -3364
rect 2880 -3444 2920 -3396
rect 2880 -3476 2884 -3444
rect 2916 -3476 2920 -3444
rect 2880 -3524 2920 -3476
rect 2880 -3556 2884 -3524
rect 2916 -3556 2920 -3524
rect 2880 -3604 2920 -3556
rect 2880 -3636 2884 -3604
rect 2916 -3636 2920 -3604
rect 2880 -3684 2920 -3636
rect 2880 -3716 2884 -3684
rect 2916 -3716 2920 -3684
rect 2880 -3720 2920 -3716
rect 2960 1036 3000 1040
rect 2960 1004 2964 1036
rect 2996 1004 3000 1036
rect 2960 956 3000 1004
rect 2960 924 2964 956
rect 2996 924 3000 956
rect 2960 876 3000 924
rect 2960 844 2964 876
rect 2996 844 3000 876
rect 2960 796 3000 844
rect 2960 764 2964 796
rect 2996 764 3000 796
rect 2960 716 3000 764
rect 2960 684 2964 716
rect 2996 684 3000 716
rect 2960 636 3000 684
rect 2960 604 2964 636
rect 2996 604 3000 636
rect 2960 556 3000 604
rect 2960 524 2964 556
rect 2996 524 3000 556
rect 2960 476 3000 524
rect 2960 444 2964 476
rect 2996 444 3000 476
rect 2960 396 3000 444
rect 2960 364 2964 396
rect 2996 364 3000 396
rect 2960 316 3000 364
rect 2960 284 2964 316
rect 2996 284 3000 316
rect 2960 236 3000 284
rect 2960 204 2964 236
rect 2996 204 3000 236
rect 2960 156 3000 204
rect 2960 124 2964 156
rect 2996 124 3000 156
rect 2960 76 3000 124
rect 2960 44 2964 76
rect 2996 44 3000 76
rect 2960 -4 3000 44
rect 2960 -36 2964 -4
rect 2996 -36 3000 -4
rect 2960 -84 3000 -36
rect 2960 -116 2964 -84
rect 2996 -116 3000 -84
rect 2960 -164 3000 -116
rect 2960 -196 2964 -164
rect 2996 -196 3000 -164
rect 2960 -244 3000 -196
rect 2960 -276 2964 -244
rect 2996 -276 3000 -244
rect 2960 -324 3000 -276
rect 2960 -356 2964 -324
rect 2996 -356 3000 -324
rect 2960 -404 3000 -356
rect 2960 -436 2964 -404
rect 2996 -436 3000 -404
rect 2960 -484 3000 -436
rect 2960 -516 2964 -484
rect 2996 -516 3000 -484
rect 2960 -564 3000 -516
rect 2960 -596 2964 -564
rect 2996 -596 3000 -564
rect 2960 -644 3000 -596
rect 2960 -676 2964 -644
rect 2996 -676 3000 -644
rect 2960 -724 3000 -676
rect 2960 -756 2964 -724
rect 2996 -756 3000 -724
rect 2960 -804 3000 -756
rect 2960 -836 2964 -804
rect 2996 -836 3000 -804
rect 2960 -884 3000 -836
rect 2960 -916 2964 -884
rect 2996 -916 3000 -884
rect 2960 -964 3000 -916
rect 2960 -996 2964 -964
rect 2996 -996 3000 -964
rect 2960 -1044 3000 -996
rect 2960 -1076 2964 -1044
rect 2996 -1076 3000 -1044
rect 2960 -1124 3000 -1076
rect 2960 -1156 2964 -1124
rect 2996 -1156 3000 -1124
rect 2960 -1204 3000 -1156
rect 2960 -1236 2964 -1204
rect 2996 -1236 3000 -1204
rect 2960 -1284 3000 -1236
rect 2960 -1316 2964 -1284
rect 2996 -1316 3000 -1284
rect 2960 -1364 3000 -1316
rect 2960 -1396 2964 -1364
rect 2996 -1396 3000 -1364
rect 2960 -1444 3000 -1396
rect 2960 -1476 2964 -1444
rect 2996 -1476 3000 -1444
rect 2960 -1524 3000 -1476
rect 2960 -1556 2964 -1524
rect 2996 -1556 3000 -1524
rect 2960 -1604 3000 -1556
rect 2960 -1636 2964 -1604
rect 2996 -1636 3000 -1604
rect 2960 -1684 3000 -1636
rect 2960 -1716 2964 -1684
rect 2996 -1716 3000 -1684
rect 2960 -1764 3000 -1716
rect 2960 -1796 2964 -1764
rect 2996 -1796 3000 -1764
rect 2960 -1844 3000 -1796
rect 2960 -1876 2964 -1844
rect 2996 -1876 3000 -1844
rect 2960 -1924 3000 -1876
rect 2960 -1956 2964 -1924
rect 2996 -1956 3000 -1924
rect 2960 -2004 3000 -1956
rect 2960 -2036 2964 -2004
rect 2996 -2036 3000 -2004
rect 2960 -2084 3000 -2036
rect 2960 -2116 2964 -2084
rect 2996 -2116 3000 -2084
rect 2960 -2164 3000 -2116
rect 2960 -2196 2964 -2164
rect 2996 -2196 3000 -2164
rect 2960 -2244 3000 -2196
rect 2960 -2276 2964 -2244
rect 2996 -2276 3000 -2244
rect 2960 -2324 3000 -2276
rect 2960 -2356 2964 -2324
rect 2996 -2356 3000 -2324
rect 2960 -2404 3000 -2356
rect 2960 -2436 2964 -2404
rect 2996 -2436 3000 -2404
rect 2960 -2484 3000 -2436
rect 2960 -2516 2964 -2484
rect 2996 -2516 3000 -2484
rect 2960 -2564 3000 -2516
rect 2960 -2596 2964 -2564
rect 2996 -2596 3000 -2564
rect 2960 -2644 3000 -2596
rect 2960 -2676 2964 -2644
rect 2996 -2676 3000 -2644
rect 2960 -2724 3000 -2676
rect 2960 -2756 2964 -2724
rect 2996 -2756 3000 -2724
rect 2960 -2804 3000 -2756
rect 2960 -2836 2964 -2804
rect 2996 -2836 3000 -2804
rect 2960 -2884 3000 -2836
rect 2960 -2916 2964 -2884
rect 2996 -2916 3000 -2884
rect 2960 -2964 3000 -2916
rect 2960 -2996 2964 -2964
rect 2996 -2996 3000 -2964
rect 2960 -3044 3000 -2996
rect 2960 -3076 2964 -3044
rect 2996 -3076 3000 -3044
rect 2960 -3124 3000 -3076
rect 2960 -3156 2964 -3124
rect 2996 -3156 3000 -3124
rect 2960 -3204 3000 -3156
rect 2960 -3236 2964 -3204
rect 2996 -3236 3000 -3204
rect 2960 -3284 3000 -3236
rect 2960 -3316 2964 -3284
rect 2996 -3316 3000 -3284
rect 2960 -3364 3000 -3316
rect 2960 -3396 2964 -3364
rect 2996 -3396 3000 -3364
rect 2960 -3444 3000 -3396
rect 2960 -3476 2964 -3444
rect 2996 -3476 3000 -3444
rect 2960 -3524 3000 -3476
rect 2960 -3556 2964 -3524
rect 2996 -3556 3000 -3524
rect 2960 -3604 3000 -3556
rect 2960 -3636 2964 -3604
rect 2996 -3636 3000 -3604
rect 2960 -3684 3000 -3636
rect 2960 -3716 2964 -3684
rect 2996 -3716 3000 -3684
rect 2960 -3720 3000 -3716
rect 3040 1036 3080 1040
rect 3040 1004 3044 1036
rect 3076 1004 3080 1036
rect 3040 956 3080 1004
rect 3040 924 3044 956
rect 3076 924 3080 956
rect 3040 876 3080 924
rect 3040 844 3044 876
rect 3076 844 3080 876
rect 3040 796 3080 844
rect 3040 764 3044 796
rect 3076 764 3080 796
rect 3040 716 3080 764
rect 3040 684 3044 716
rect 3076 684 3080 716
rect 3040 636 3080 684
rect 3040 604 3044 636
rect 3076 604 3080 636
rect 3040 556 3080 604
rect 3040 524 3044 556
rect 3076 524 3080 556
rect 3040 476 3080 524
rect 3040 444 3044 476
rect 3076 444 3080 476
rect 3040 396 3080 444
rect 3040 364 3044 396
rect 3076 364 3080 396
rect 3040 316 3080 364
rect 3040 284 3044 316
rect 3076 284 3080 316
rect 3040 236 3080 284
rect 3040 204 3044 236
rect 3076 204 3080 236
rect 3040 156 3080 204
rect 3040 124 3044 156
rect 3076 124 3080 156
rect 3040 76 3080 124
rect 3040 44 3044 76
rect 3076 44 3080 76
rect 3040 -4 3080 44
rect 3040 -36 3044 -4
rect 3076 -36 3080 -4
rect 3040 -84 3080 -36
rect 3040 -116 3044 -84
rect 3076 -116 3080 -84
rect 3040 -164 3080 -116
rect 3040 -196 3044 -164
rect 3076 -196 3080 -164
rect 3040 -244 3080 -196
rect 3040 -276 3044 -244
rect 3076 -276 3080 -244
rect 3040 -324 3080 -276
rect 3040 -356 3044 -324
rect 3076 -356 3080 -324
rect 3040 -404 3080 -356
rect 3040 -436 3044 -404
rect 3076 -436 3080 -404
rect 3040 -484 3080 -436
rect 3040 -516 3044 -484
rect 3076 -516 3080 -484
rect 3040 -564 3080 -516
rect 3040 -596 3044 -564
rect 3076 -596 3080 -564
rect 3040 -644 3080 -596
rect 3040 -676 3044 -644
rect 3076 -676 3080 -644
rect 3040 -724 3080 -676
rect 3040 -756 3044 -724
rect 3076 -756 3080 -724
rect 3040 -804 3080 -756
rect 3040 -836 3044 -804
rect 3076 -836 3080 -804
rect 3040 -884 3080 -836
rect 3040 -916 3044 -884
rect 3076 -916 3080 -884
rect 3040 -964 3080 -916
rect 3040 -996 3044 -964
rect 3076 -996 3080 -964
rect 3040 -1044 3080 -996
rect 3040 -1076 3044 -1044
rect 3076 -1076 3080 -1044
rect 3040 -1124 3080 -1076
rect 3040 -1156 3044 -1124
rect 3076 -1156 3080 -1124
rect 3040 -1204 3080 -1156
rect 3040 -1236 3044 -1204
rect 3076 -1236 3080 -1204
rect 3040 -1284 3080 -1236
rect 3040 -1316 3044 -1284
rect 3076 -1316 3080 -1284
rect 3040 -1364 3080 -1316
rect 3040 -1396 3044 -1364
rect 3076 -1396 3080 -1364
rect 3040 -1444 3080 -1396
rect 3040 -1476 3044 -1444
rect 3076 -1476 3080 -1444
rect 3040 -1524 3080 -1476
rect 3040 -1556 3044 -1524
rect 3076 -1556 3080 -1524
rect 3040 -1604 3080 -1556
rect 3040 -1636 3044 -1604
rect 3076 -1636 3080 -1604
rect 3040 -1684 3080 -1636
rect 3040 -1716 3044 -1684
rect 3076 -1716 3080 -1684
rect 3040 -1764 3080 -1716
rect 3040 -1796 3044 -1764
rect 3076 -1796 3080 -1764
rect 3040 -1844 3080 -1796
rect 3040 -1876 3044 -1844
rect 3076 -1876 3080 -1844
rect 3040 -1924 3080 -1876
rect 3040 -1956 3044 -1924
rect 3076 -1956 3080 -1924
rect 3040 -2004 3080 -1956
rect 3040 -2036 3044 -2004
rect 3076 -2036 3080 -2004
rect 3040 -2084 3080 -2036
rect 3040 -2116 3044 -2084
rect 3076 -2116 3080 -2084
rect 3040 -2164 3080 -2116
rect 3040 -2196 3044 -2164
rect 3076 -2196 3080 -2164
rect 3040 -2244 3080 -2196
rect 3040 -2276 3044 -2244
rect 3076 -2276 3080 -2244
rect 3040 -2324 3080 -2276
rect 3040 -2356 3044 -2324
rect 3076 -2356 3080 -2324
rect 3040 -2404 3080 -2356
rect 3040 -2436 3044 -2404
rect 3076 -2436 3080 -2404
rect 3040 -2484 3080 -2436
rect 3040 -2516 3044 -2484
rect 3076 -2516 3080 -2484
rect 3040 -2564 3080 -2516
rect 3040 -2596 3044 -2564
rect 3076 -2596 3080 -2564
rect 3040 -2644 3080 -2596
rect 3040 -2676 3044 -2644
rect 3076 -2676 3080 -2644
rect 3040 -2724 3080 -2676
rect 3040 -2756 3044 -2724
rect 3076 -2756 3080 -2724
rect 3040 -2804 3080 -2756
rect 3040 -2836 3044 -2804
rect 3076 -2836 3080 -2804
rect 3040 -2884 3080 -2836
rect 3040 -2916 3044 -2884
rect 3076 -2916 3080 -2884
rect 3040 -2964 3080 -2916
rect 3040 -2996 3044 -2964
rect 3076 -2996 3080 -2964
rect 3040 -3044 3080 -2996
rect 3040 -3076 3044 -3044
rect 3076 -3076 3080 -3044
rect 3040 -3124 3080 -3076
rect 3040 -3156 3044 -3124
rect 3076 -3156 3080 -3124
rect 3040 -3204 3080 -3156
rect 3040 -3236 3044 -3204
rect 3076 -3236 3080 -3204
rect 3040 -3284 3080 -3236
rect 3040 -3316 3044 -3284
rect 3076 -3316 3080 -3284
rect 3040 -3364 3080 -3316
rect 3040 -3396 3044 -3364
rect 3076 -3396 3080 -3364
rect 3040 -3444 3080 -3396
rect 3040 -3476 3044 -3444
rect 3076 -3476 3080 -3444
rect 3040 -3524 3080 -3476
rect 3040 -3556 3044 -3524
rect 3076 -3556 3080 -3524
rect 3040 -3604 3080 -3556
rect 3040 -3636 3044 -3604
rect 3076 -3636 3080 -3604
rect 3040 -3684 3080 -3636
rect 3040 -3716 3044 -3684
rect 3076 -3716 3080 -3684
rect 3040 -3720 3080 -3716
rect 3120 1036 3160 1040
rect 3120 1004 3124 1036
rect 3156 1004 3160 1036
rect 3120 956 3160 1004
rect 3120 924 3124 956
rect 3156 924 3160 956
rect 3120 876 3160 924
rect 3120 844 3124 876
rect 3156 844 3160 876
rect 3120 796 3160 844
rect 3120 764 3124 796
rect 3156 764 3160 796
rect 3120 716 3160 764
rect 3120 684 3124 716
rect 3156 684 3160 716
rect 3120 636 3160 684
rect 3120 604 3124 636
rect 3156 604 3160 636
rect 3120 556 3160 604
rect 3120 524 3124 556
rect 3156 524 3160 556
rect 3120 476 3160 524
rect 3120 444 3124 476
rect 3156 444 3160 476
rect 3120 396 3160 444
rect 3120 364 3124 396
rect 3156 364 3160 396
rect 3120 316 3160 364
rect 3120 284 3124 316
rect 3156 284 3160 316
rect 3120 236 3160 284
rect 3120 204 3124 236
rect 3156 204 3160 236
rect 3120 156 3160 204
rect 3120 124 3124 156
rect 3156 124 3160 156
rect 3120 76 3160 124
rect 3120 44 3124 76
rect 3156 44 3160 76
rect 3120 -4 3160 44
rect 3120 -36 3124 -4
rect 3156 -36 3160 -4
rect 3120 -84 3160 -36
rect 3120 -116 3124 -84
rect 3156 -116 3160 -84
rect 3120 -164 3160 -116
rect 3120 -196 3124 -164
rect 3156 -196 3160 -164
rect 3120 -244 3160 -196
rect 3120 -276 3124 -244
rect 3156 -276 3160 -244
rect 3120 -324 3160 -276
rect 3120 -356 3124 -324
rect 3156 -356 3160 -324
rect 3120 -404 3160 -356
rect 3120 -436 3124 -404
rect 3156 -436 3160 -404
rect 3120 -484 3160 -436
rect 3120 -516 3124 -484
rect 3156 -516 3160 -484
rect 3120 -564 3160 -516
rect 3120 -596 3124 -564
rect 3156 -596 3160 -564
rect 3120 -644 3160 -596
rect 3120 -676 3124 -644
rect 3156 -676 3160 -644
rect 3120 -724 3160 -676
rect 3120 -756 3124 -724
rect 3156 -756 3160 -724
rect 3120 -804 3160 -756
rect 3120 -836 3124 -804
rect 3156 -836 3160 -804
rect 3120 -884 3160 -836
rect 3120 -916 3124 -884
rect 3156 -916 3160 -884
rect 3120 -964 3160 -916
rect 3120 -996 3124 -964
rect 3156 -996 3160 -964
rect 3120 -1044 3160 -996
rect 3120 -1076 3124 -1044
rect 3156 -1076 3160 -1044
rect 3120 -1124 3160 -1076
rect 3120 -1156 3124 -1124
rect 3156 -1156 3160 -1124
rect 3120 -1204 3160 -1156
rect 3120 -1236 3124 -1204
rect 3156 -1236 3160 -1204
rect 3120 -1284 3160 -1236
rect 3120 -1316 3124 -1284
rect 3156 -1316 3160 -1284
rect 3120 -1364 3160 -1316
rect 3120 -1396 3124 -1364
rect 3156 -1396 3160 -1364
rect 3120 -1444 3160 -1396
rect 3120 -1476 3124 -1444
rect 3156 -1476 3160 -1444
rect 3120 -1524 3160 -1476
rect 3120 -1556 3124 -1524
rect 3156 -1556 3160 -1524
rect 3120 -1604 3160 -1556
rect 3120 -1636 3124 -1604
rect 3156 -1636 3160 -1604
rect 3120 -1684 3160 -1636
rect 3120 -1716 3124 -1684
rect 3156 -1716 3160 -1684
rect 3120 -1764 3160 -1716
rect 3120 -1796 3124 -1764
rect 3156 -1796 3160 -1764
rect 3120 -1844 3160 -1796
rect 3120 -1876 3124 -1844
rect 3156 -1876 3160 -1844
rect 3120 -1924 3160 -1876
rect 3120 -1956 3124 -1924
rect 3156 -1956 3160 -1924
rect 3120 -2004 3160 -1956
rect 3120 -2036 3124 -2004
rect 3156 -2036 3160 -2004
rect 3120 -2084 3160 -2036
rect 3120 -2116 3124 -2084
rect 3156 -2116 3160 -2084
rect 3120 -2164 3160 -2116
rect 3120 -2196 3124 -2164
rect 3156 -2196 3160 -2164
rect 3120 -2244 3160 -2196
rect 3120 -2276 3124 -2244
rect 3156 -2276 3160 -2244
rect 3120 -2324 3160 -2276
rect 3120 -2356 3124 -2324
rect 3156 -2356 3160 -2324
rect 3120 -2404 3160 -2356
rect 3120 -2436 3124 -2404
rect 3156 -2436 3160 -2404
rect 3120 -2484 3160 -2436
rect 3120 -2516 3124 -2484
rect 3156 -2516 3160 -2484
rect 3120 -2564 3160 -2516
rect 3120 -2596 3124 -2564
rect 3156 -2596 3160 -2564
rect 3120 -2644 3160 -2596
rect 3120 -2676 3124 -2644
rect 3156 -2676 3160 -2644
rect 3120 -2724 3160 -2676
rect 3120 -2756 3124 -2724
rect 3156 -2756 3160 -2724
rect 3120 -2804 3160 -2756
rect 3120 -2836 3124 -2804
rect 3156 -2836 3160 -2804
rect 3120 -2884 3160 -2836
rect 3120 -2916 3124 -2884
rect 3156 -2916 3160 -2884
rect 3120 -2964 3160 -2916
rect 3120 -2996 3124 -2964
rect 3156 -2996 3160 -2964
rect 3120 -3044 3160 -2996
rect 3120 -3076 3124 -3044
rect 3156 -3076 3160 -3044
rect 3120 -3124 3160 -3076
rect 3120 -3156 3124 -3124
rect 3156 -3156 3160 -3124
rect 3120 -3204 3160 -3156
rect 3120 -3236 3124 -3204
rect 3156 -3236 3160 -3204
rect 3120 -3284 3160 -3236
rect 3120 -3316 3124 -3284
rect 3156 -3316 3160 -3284
rect 3120 -3364 3160 -3316
rect 3120 -3396 3124 -3364
rect 3156 -3396 3160 -3364
rect 3120 -3444 3160 -3396
rect 3120 -3476 3124 -3444
rect 3156 -3476 3160 -3444
rect 3120 -3524 3160 -3476
rect 3120 -3556 3124 -3524
rect 3156 -3556 3160 -3524
rect 3120 -3604 3160 -3556
rect 3120 -3636 3124 -3604
rect 3156 -3636 3160 -3604
rect 3120 -3684 3160 -3636
rect 3120 -3716 3124 -3684
rect 3156 -3716 3160 -3684
rect 3120 -3720 3160 -3716
rect 3200 1036 3240 1040
rect 3200 1004 3204 1036
rect 3236 1004 3240 1036
rect 3200 956 3240 1004
rect 3200 924 3204 956
rect 3236 924 3240 956
rect 3200 876 3240 924
rect 3200 844 3204 876
rect 3236 844 3240 876
rect 3200 796 3240 844
rect 3200 764 3204 796
rect 3236 764 3240 796
rect 3200 716 3240 764
rect 3200 684 3204 716
rect 3236 684 3240 716
rect 3200 636 3240 684
rect 3200 604 3204 636
rect 3236 604 3240 636
rect 3200 556 3240 604
rect 3200 524 3204 556
rect 3236 524 3240 556
rect 3200 476 3240 524
rect 3200 444 3204 476
rect 3236 444 3240 476
rect 3200 396 3240 444
rect 3200 364 3204 396
rect 3236 364 3240 396
rect 3200 316 3240 364
rect 3200 284 3204 316
rect 3236 284 3240 316
rect 3200 236 3240 284
rect 3200 204 3204 236
rect 3236 204 3240 236
rect 3200 156 3240 204
rect 3200 124 3204 156
rect 3236 124 3240 156
rect 3200 76 3240 124
rect 3200 44 3204 76
rect 3236 44 3240 76
rect 3200 -4 3240 44
rect 3200 -36 3204 -4
rect 3236 -36 3240 -4
rect 3200 -84 3240 -36
rect 3200 -116 3204 -84
rect 3236 -116 3240 -84
rect 3200 -164 3240 -116
rect 3200 -196 3204 -164
rect 3236 -196 3240 -164
rect 3200 -244 3240 -196
rect 3200 -276 3204 -244
rect 3236 -276 3240 -244
rect 3200 -324 3240 -276
rect 3200 -356 3204 -324
rect 3236 -356 3240 -324
rect 3200 -404 3240 -356
rect 3200 -436 3204 -404
rect 3236 -436 3240 -404
rect 3200 -484 3240 -436
rect 3200 -516 3204 -484
rect 3236 -516 3240 -484
rect 3200 -564 3240 -516
rect 3200 -596 3204 -564
rect 3236 -596 3240 -564
rect 3200 -644 3240 -596
rect 3200 -676 3204 -644
rect 3236 -676 3240 -644
rect 3200 -724 3240 -676
rect 3200 -756 3204 -724
rect 3236 -756 3240 -724
rect 3200 -804 3240 -756
rect 3200 -836 3204 -804
rect 3236 -836 3240 -804
rect 3200 -884 3240 -836
rect 3200 -916 3204 -884
rect 3236 -916 3240 -884
rect 3200 -964 3240 -916
rect 3200 -996 3204 -964
rect 3236 -996 3240 -964
rect 3200 -1044 3240 -996
rect 3200 -1076 3204 -1044
rect 3236 -1076 3240 -1044
rect 3200 -1124 3240 -1076
rect 3200 -1156 3204 -1124
rect 3236 -1156 3240 -1124
rect 3200 -1204 3240 -1156
rect 3200 -1236 3204 -1204
rect 3236 -1236 3240 -1204
rect 3200 -1284 3240 -1236
rect 3200 -1316 3204 -1284
rect 3236 -1316 3240 -1284
rect 3200 -1364 3240 -1316
rect 3200 -1396 3204 -1364
rect 3236 -1396 3240 -1364
rect 3200 -1444 3240 -1396
rect 3200 -1476 3204 -1444
rect 3236 -1476 3240 -1444
rect 3200 -1524 3240 -1476
rect 3200 -1556 3204 -1524
rect 3236 -1556 3240 -1524
rect 3200 -1604 3240 -1556
rect 3200 -1636 3204 -1604
rect 3236 -1636 3240 -1604
rect 3200 -1684 3240 -1636
rect 3200 -1716 3204 -1684
rect 3236 -1716 3240 -1684
rect 3200 -1764 3240 -1716
rect 3200 -1796 3204 -1764
rect 3236 -1796 3240 -1764
rect 3200 -1844 3240 -1796
rect 3200 -1876 3204 -1844
rect 3236 -1876 3240 -1844
rect 3200 -1924 3240 -1876
rect 3200 -1956 3204 -1924
rect 3236 -1956 3240 -1924
rect 3200 -2004 3240 -1956
rect 3200 -2036 3204 -2004
rect 3236 -2036 3240 -2004
rect 3200 -2084 3240 -2036
rect 3200 -2116 3204 -2084
rect 3236 -2116 3240 -2084
rect 3200 -2164 3240 -2116
rect 3200 -2196 3204 -2164
rect 3236 -2196 3240 -2164
rect 3200 -2244 3240 -2196
rect 3200 -2276 3204 -2244
rect 3236 -2276 3240 -2244
rect 3200 -2324 3240 -2276
rect 3200 -2356 3204 -2324
rect 3236 -2356 3240 -2324
rect 3200 -2404 3240 -2356
rect 3200 -2436 3204 -2404
rect 3236 -2436 3240 -2404
rect 3200 -2484 3240 -2436
rect 3200 -2516 3204 -2484
rect 3236 -2516 3240 -2484
rect 3200 -2564 3240 -2516
rect 3200 -2596 3204 -2564
rect 3236 -2596 3240 -2564
rect 3200 -2644 3240 -2596
rect 3200 -2676 3204 -2644
rect 3236 -2676 3240 -2644
rect 3200 -2724 3240 -2676
rect 3200 -2756 3204 -2724
rect 3236 -2756 3240 -2724
rect 3200 -2804 3240 -2756
rect 3200 -2836 3204 -2804
rect 3236 -2836 3240 -2804
rect 3200 -2884 3240 -2836
rect 3200 -2916 3204 -2884
rect 3236 -2916 3240 -2884
rect 3200 -2964 3240 -2916
rect 3200 -2996 3204 -2964
rect 3236 -2996 3240 -2964
rect 3200 -3044 3240 -2996
rect 3200 -3076 3204 -3044
rect 3236 -3076 3240 -3044
rect 3200 -3124 3240 -3076
rect 3200 -3156 3204 -3124
rect 3236 -3156 3240 -3124
rect 3200 -3204 3240 -3156
rect 3200 -3236 3204 -3204
rect 3236 -3236 3240 -3204
rect 3200 -3284 3240 -3236
rect 3200 -3316 3204 -3284
rect 3236 -3316 3240 -3284
rect 3200 -3364 3240 -3316
rect 3200 -3396 3204 -3364
rect 3236 -3396 3240 -3364
rect 3200 -3444 3240 -3396
rect 3200 -3476 3204 -3444
rect 3236 -3476 3240 -3444
rect 3200 -3524 3240 -3476
rect 3200 -3556 3204 -3524
rect 3236 -3556 3240 -3524
rect 3200 -3604 3240 -3556
rect 3200 -3636 3204 -3604
rect 3236 -3636 3240 -3604
rect 3200 -3684 3240 -3636
rect 3200 -3716 3204 -3684
rect 3236 -3716 3240 -3684
rect 3200 -3720 3240 -3716
rect 3280 1036 3320 1040
rect 3280 1004 3284 1036
rect 3316 1004 3320 1036
rect 3280 956 3320 1004
rect 3280 924 3284 956
rect 3316 924 3320 956
rect 3280 876 3320 924
rect 3280 844 3284 876
rect 3316 844 3320 876
rect 3280 796 3320 844
rect 3280 764 3284 796
rect 3316 764 3320 796
rect 3280 716 3320 764
rect 3280 684 3284 716
rect 3316 684 3320 716
rect 3280 636 3320 684
rect 3280 604 3284 636
rect 3316 604 3320 636
rect 3280 556 3320 604
rect 3280 524 3284 556
rect 3316 524 3320 556
rect 3280 476 3320 524
rect 3280 444 3284 476
rect 3316 444 3320 476
rect 3280 396 3320 444
rect 3280 364 3284 396
rect 3316 364 3320 396
rect 3280 316 3320 364
rect 3280 284 3284 316
rect 3316 284 3320 316
rect 3280 236 3320 284
rect 3280 204 3284 236
rect 3316 204 3320 236
rect 3280 156 3320 204
rect 3280 124 3284 156
rect 3316 124 3320 156
rect 3280 76 3320 124
rect 3280 44 3284 76
rect 3316 44 3320 76
rect 3280 -4 3320 44
rect 3280 -36 3284 -4
rect 3316 -36 3320 -4
rect 3280 -84 3320 -36
rect 3280 -116 3284 -84
rect 3316 -116 3320 -84
rect 3280 -164 3320 -116
rect 3280 -196 3284 -164
rect 3316 -196 3320 -164
rect 3280 -244 3320 -196
rect 3280 -276 3284 -244
rect 3316 -276 3320 -244
rect 3280 -324 3320 -276
rect 3280 -356 3284 -324
rect 3316 -356 3320 -324
rect 3280 -404 3320 -356
rect 3280 -436 3284 -404
rect 3316 -436 3320 -404
rect 3280 -484 3320 -436
rect 3280 -516 3284 -484
rect 3316 -516 3320 -484
rect 3280 -564 3320 -516
rect 3280 -596 3284 -564
rect 3316 -596 3320 -564
rect 3280 -644 3320 -596
rect 3280 -676 3284 -644
rect 3316 -676 3320 -644
rect 3280 -724 3320 -676
rect 3280 -756 3284 -724
rect 3316 -756 3320 -724
rect 3280 -804 3320 -756
rect 3280 -836 3284 -804
rect 3316 -836 3320 -804
rect 3280 -884 3320 -836
rect 3280 -916 3284 -884
rect 3316 -916 3320 -884
rect 3280 -964 3320 -916
rect 3280 -996 3284 -964
rect 3316 -996 3320 -964
rect 3280 -1044 3320 -996
rect 3280 -1076 3284 -1044
rect 3316 -1076 3320 -1044
rect 3280 -1124 3320 -1076
rect 3280 -1156 3284 -1124
rect 3316 -1156 3320 -1124
rect 3280 -1204 3320 -1156
rect 3280 -1236 3284 -1204
rect 3316 -1236 3320 -1204
rect 3280 -1284 3320 -1236
rect 3280 -1316 3284 -1284
rect 3316 -1316 3320 -1284
rect 3280 -1364 3320 -1316
rect 3280 -1396 3284 -1364
rect 3316 -1396 3320 -1364
rect 3280 -1444 3320 -1396
rect 3280 -1476 3284 -1444
rect 3316 -1476 3320 -1444
rect 3280 -1524 3320 -1476
rect 3280 -1556 3284 -1524
rect 3316 -1556 3320 -1524
rect 3280 -1604 3320 -1556
rect 3280 -1636 3284 -1604
rect 3316 -1636 3320 -1604
rect 3280 -1684 3320 -1636
rect 3280 -1716 3284 -1684
rect 3316 -1716 3320 -1684
rect 3280 -1764 3320 -1716
rect 3280 -1796 3284 -1764
rect 3316 -1796 3320 -1764
rect 3280 -1844 3320 -1796
rect 3280 -1876 3284 -1844
rect 3316 -1876 3320 -1844
rect 3280 -1924 3320 -1876
rect 3280 -1956 3284 -1924
rect 3316 -1956 3320 -1924
rect 3280 -2004 3320 -1956
rect 3280 -2036 3284 -2004
rect 3316 -2036 3320 -2004
rect 3280 -2084 3320 -2036
rect 3280 -2116 3284 -2084
rect 3316 -2116 3320 -2084
rect 3280 -2164 3320 -2116
rect 3280 -2196 3284 -2164
rect 3316 -2196 3320 -2164
rect 3280 -2244 3320 -2196
rect 3280 -2276 3284 -2244
rect 3316 -2276 3320 -2244
rect 3280 -2324 3320 -2276
rect 3280 -2356 3284 -2324
rect 3316 -2356 3320 -2324
rect 3280 -2404 3320 -2356
rect 3280 -2436 3284 -2404
rect 3316 -2436 3320 -2404
rect 3280 -2484 3320 -2436
rect 3280 -2516 3284 -2484
rect 3316 -2516 3320 -2484
rect 3280 -2564 3320 -2516
rect 3280 -2596 3284 -2564
rect 3316 -2596 3320 -2564
rect 3280 -2644 3320 -2596
rect 3280 -2676 3284 -2644
rect 3316 -2676 3320 -2644
rect 3280 -2724 3320 -2676
rect 3280 -2756 3284 -2724
rect 3316 -2756 3320 -2724
rect 3280 -2804 3320 -2756
rect 3280 -2836 3284 -2804
rect 3316 -2836 3320 -2804
rect 3280 -2884 3320 -2836
rect 3280 -2916 3284 -2884
rect 3316 -2916 3320 -2884
rect 3280 -2964 3320 -2916
rect 3280 -2996 3284 -2964
rect 3316 -2996 3320 -2964
rect 3280 -3044 3320 -2996
rect 3280 -3076 3284 -3044
rect 3316 -3076 3320 -3044
rect 3280 -3124 3320 -3076
rect 3280 -3156 3284 -3124
rect 3316 -3156 3320 -3124
rect 3280 -3204 3320 -3156
rect 3280 -3236 3284 -3204
rect 3316 -3236 3320 -3204
rect 3280 -3284 3320 -3236
rect 3280 -3316 3284 -3284
rect 3316 -3316 3320 -3284
rect 3280 -3364 3320 -3316
rect 3280 -3396 3284 -3364
rect 3316 -3396 3320 -3364
rect 3280 -3444 3320 -3396
rect 3280 -3476 3284 -3444
rect 3316 -3476 3320 -3444
rect 3280 -3524 3320 -3476
rect 3280 -3556 3284 -3524
rect 3316 -3556 3320 -3524
rect 3280 -3604 3320 -3556
rect 3280 -3636 3284 -3604
rect 3316 -3636 3320 -3604
rect 3280 -3684 3320 -3636
rect 3280 -3716 3284 -3684
rect 3316 -3716 3320 -3684
rect 3280 -3720 3320 -3716
rect 3360 1036 3400 1040
rect 3360 1004 3364 1036
rect 3396 1004 3400 1036
rect 3360 956 3400 1004
rect 3360 924 3364 956
rect 3396 924 3400 956
rect 3360 876 3400 924
rect 3360 844 3364 876
rect 3396 844 3400 876
rect 3360 796 3400 844
rect 3360 764 3364 796
rect 3396 764 3400 796
rect 3360 716 3400 764
rect 3360 684 3364 716
rect 3396 684 3400 716
rect 3360 636 3400 684
rect 3360 604 3364 636
rect 3396 604 3400 636
rect 3360 556 3400 604
rect 3360 524 3364 556
rect 3396 524 3400 556
rect 3360 476 3400 524
rect 3360 444 3364 476
rect 3396 444 3400 476
rect 3360 396 3400 444
rect 3360 364 3364 396
rect 3396 364 3400 396
rect 3360 316 3400 364
rect 3360 284 3364 316
rect 3396 284 3400 316
rect 3360 236 3400 284
rect 3360 204 3364 236
rect 3396 204 3400 236
rect 3360 156 3400 204
rect 3360 124 3364 156
rect 3396 124 3400 156
rect 3360 76 3400 124
rect 3360 44 3364 76
rect 3396 44 3400 76
rect 3360 -4 3400 44
rect 3360 -36 3364 -4
rect 3396 -36 3400 -4
rect 3360 -84 3400 -36
rect 3360 -116 3364 -84
rect 3396 -116 3400 -84
rect 3360 -164 3400 -116
rect 3360 -196 3364 -164
rect 3396 -196 3400 -164
rect 3360 -244 3400 -196
rect 3360 -276 3364 -244
rect 3396 -276 3400 -244
rect 3360 -324 3400 -276
rect 3360 -356 3364 -324
rect 3396 -356 3400 -324
rect 3360 -404 3400 -356
rect 3360 -436 3364 -404
rect 3396 -436 3400 -404
rect 3360 -484 3400 -436
rect 3360 -516 3364 -484
rect 3396 -516 3400 -484
rect 3360 -564 3400 -516
rect 3360 -596 3364 -564
rect 3396 -596 3400 -564
rect 3360 -644 3400 -596
rect 3360 -676 3364 -644
rect 3396 -676 3400 -644
rect 3360 -724 3400 -676
rect 3360 -756 3364 -724
rect 3396 -756 3400 -724
rect 3360 -804 3400 -756
rect 3360 -836 3364 -804
rect 3396 -836 3400 -804
rect 3360 -884 3400 -836
rect 3360 -916 3364 -884
rect 3396 -916 3400 -884
rect 3360 -964 3400 -916
rect 3360 -996 3364 -964
rect 3396 -996 3400 -964
rect 3360 -1044 3400 -996
rect 3360 -1076 3364 -1044
rect 3396 -1076 3400 -1044
rect 3360 -1124 3400 -1076
rect 3360 -1156 3364 -1124
rect 3396 -1156 3400 -1124
rect 3360 -1204 3400 -1156
rect 3360 -1236 3364 -1204
rect 3396 -1236 3400 -1204
rect 3360 -1284 3400 -1236
rect 3360 -1316 3364 -1284
rect 3396 -1316 3400 -1284
rect 3360 -1364 3400 -1316
rect 3360 -1396 3364 -1364
rect 3396 -1396 3400 -1364
rect 3360 -1444 3400 -1396
rect 3360 -1476 3364 -1444
rect 3396 -1476 3400 -1444
rect 3360 -1524 3400 -1476
rect 3360 -1556 3364 -1524
rect 3396 -1556 3400 -1524
rect 3360 -1604 3400 -1556
rect 3360 -1636 3364 -1604
rect 3396 -1636 3400 -1604
rect 3360 -1684 3400 -1636
rect 3360 -1716 3364 -1684
rect 3396 -1716 3400 -1684
rect 3360 -1764 3400 -1716
rect 3360 -1796 3364 -1764
rect 3396 -1796 3400 -1764
rect 3360 -1844 3400 -1796
rect 3360 -1876 3364 -1844
rect 3396 -1876 3400 -1844
rect 3360 -1924 3400 -1876
rect 3360 -1956 3364 -1924
rect 3396 -1956 3400 -1924
rect 3360 -2004 3400 -1956
rect 3360 -2036 3364 -2004
rect 3396 -2036 3400 -2004
rect 3360 -2084 3400 -2036
rect 3360 -2116 3364 -2084
rect 3396 -2116 3400 -2084
rect 3360 -2164 3400 -2116
rect 3360 -2196 3364 -2164
rect 3396 -2196 3400 -2164
rect 3360 -2244 3400 -2196
rect 3360 -2276 3364 -2244
rect 3396 -2276 3400 -2244
rect 3360 -2324 3400 -2276
rect 3360 -2356 3364 -2324
rect 3396 -2356 3400 -2324
rect 3360 -2404 3400 -2356
rect 3360 -2436 3364 -2404
rect 3396 -2436 3400 -2404
rect 3360 -2484 3400 -2436
rect 3360 -2516 3364 -2484
rect 3396 -2516 3400 -2484
rect 3360 -2564 3400 -2516
rect 3360 -2596 3364 -2564
rect 3396 -2596 3400 -2564
rect 3360 -2644 3400 -2596
rect 3360 -2676 3364 -2644
rect 3396 -2676 3400 -2644
rect 3360 -2724 3400 -2676
rect 3360 -2756 3364 -2724
rect 3396 -2756 3400 -2724
rect 3360 -2804 3400 -2756
rect 3360 -2836 3364 -2804
rect 3396 -2836 3400 -2804
rect 3360 -2884 3400 -2836
rect 3360 -2916 3364 -2884
rect 3396 -2916 3400 -2884
rect 3360 -2964 3400 -2916
rect 3360 -2996 3364 -2964
rect 3396 -2996 3400 -2964
rect 3360 -3044 3400 -2996
rect 3360 -3076 3364 -3044
rect 3396 -3076 3400 -3044
rect 3360 -3124 3400 -3076
rect 3360 -3156 3364 -3124
rect 3396 -3156 3400 -3124
rect 3360 -3204 3400 -3156
rect 3360 -3236 3364 -3204
rect 3396 -3236 3400 -3204
rect 3360 -3284 3400 -3236
rect 3360 -3316 3364 -3284
rect 3396 -3316 3400 -3284
rect 3360 -3364 3400 -3316
rect 3360 -3396 3364 -3364
rect 3396 -3396 3400 -3364
rect 3360 -3444 3400 -3396
rect 3360 -3476 3364 -3444
rect 3396 -3476 3400 -3444
rect 3360 -3524 3400 -3476
rect 3360 -3556 3364 -3524
rect 3396 -3556 3400 -3524
rect 3360 -3604 3400 -3556
rect 3360 -3636 3364 -3604
rect 3396 -3636 3400 -3604
rect 3360 -3684 3400 -3636
rect 3360 -3716 3364 -3684
rect 3396 -3716 3400 -3684
rect 3360 -3720 3400 -3716
rect 3440 1036 3480 1040
rect 3440 1004 3444 1036
rect 3476 1004 3480 1036
rect 3440 956 3480 1004
rect 3440 924 3444 956
rect 3476 924 3480 956
rect 3440 876 3480 924
rect 3440 844 3444 876
rect 3476 844 3480 876
rect 3440 796 3480 844
rect 3440 764 3444 796
rect 3476 764 3480 796
rect 3440 716 3480 764
rect 3440 684 3444 716
rect 3476 684 3480 716
rect 3440 636 3480 684
rect 3440 604 3444 636
rect 3476 604 3480 636
rect 3440 556 3480 604
rect 3440 524 3444 556
rect 3476 524 3480 556
rect 3440 476 3480 524
rect 3440 444 3444 476
rect 3476 444 3480 476
rect 3440 396 3480 444
rect 3440 364 3444 396
rect 3476 364 3480 396
rect 3440 316 3480 364
rect 3440 284 3444 316
rect 3476 284 3480 316
rect 3440 236 3480 284
rect 3440 204 3444 236
rect 3476 204 3480 236
rect 3440 156 3480 204
rect 3440 124 3444 156
rect 3476 124 3480 156
rect 3440 76 3480 124
rect 3440 44 3444 76
rect 3476 44 3480 76
rect 3440 -4 3480 44
rect 3440 -36 3444 -4
rect 3476 -36 3480 -4
rect 3440 -84 3480 -36
rect 3440 -116 3444 -84
rect 3476 -116 3480 -84
rect 3440 -164 3480 -116
rect 3440 -196 3444 -164
rect 3476 -196 3480 -164
rect 3440 -244 3480 -196
rect 3440 -276 3444 -244
rect 3476 -276 3480 -244
rect 3440 -324 3480 -276
rect 3440 -356 3444 -324
rect 3476 -356 3480 -324
rect 3440 -404 3480 -356
rect 3440 -436 3444 -404
rect 3476 -436 3480 -404
rect 3440 -484 3480 -436
rect 3440 -516 3444 -484
rect 3476 -516 3480 -484
rect 3440 -564 3480 -516
rect 3440 -596 3444 -564
rect 3476 -596 3480 -564
rect 3440 -644 3480 -596
rect 3440 -676 3444 -644
rect 3476 -676 3480 -644
rect 3440 -724 3480 -676
rect 3440 -756 3444 -724
rect 3476 -756 3480 -724
rect 3440 -804 3480 -756
rect 3440 -836 3444 -804
rect 3476 -836 3480 -804
rect 3440 -884 3480 -836
rect 3440 -916 3444 -884
rect 3476 -916 3480 -884
rect 3440 -964 3480 -916
rect 3440 -996 3444 -964
rect 3476 -996 3480 -964
rect 3440 -1044 3480 -996
rect 3440 -1076 3444 -1044
rect 3476 -1076 3480 -1044
rect 3440 -1124 3480 -1076
rect 3440 -1156 3444 -1124
rect 3476 -1156 3480 -1124
rect 3440 -1204 3480 -1156
rect 3440 -1236 3444 -1204
rect 3476 -1236 3480 -1204
rect 3440 -1284 3480 -1236
rect 3440 -1316 3444 -1284
rect 3476 -1316 3480 -1284
rect 3440 -1364 3480 -1316
rect 3440 -1396 3444 -1364
rect 3476 -1396 3480 -1364
rect 3440 -1444 3480 -1396
rect 3440 -1476 3444 -1444
rect 3476 -1476 3480 -1444
rect 3440 -1524 3480 -1476
rect 3440 -1556 3444 -1524
rect 3476 -1556 3480 -1524
rect 3440 -1604 3480 -1556
rect 3440 -1636 3444 -1604
rect 3476 -1636 3480 -1604
rect 3440 -1684 3480 -1636
rect 3440 -1716 3444 -1684
rect 3476 -1716 3480 -1684
rect 3440 -1764 3480 -1716
rect 3440 -1796 3444 -1764
rect 3476 -1796 3480 -1764
rect 3440 -1844 3480 -1796
rect 3440 -1876 3444 -1844
rect 3476 -1876 3480 -1844
rect 3440 -1924 3480 -1876
rect 3440 -1956 3444 -1924
rect 3476 -1956 3480 -1924
rect 3440 -2004 3480 -1956
rect 3440 -2036 3444 -2004
rect 3476 -2036 3480 -2004
rect 3440 -2084 3480 -2036
rect 3440 -2116 3444 -2084
rect 3476 -2116 3480 -2084
rect 3440 -2164 3480 -2116
rect 3440 -2196 3444 -2164
rect 3476 -2196 3480 -2164
rect 3440 -2244 3480 -2196
rect 3440 -2276 3444 -2244
rect 3476 -2276 3480 -2244
rect 3440 -2324 3480 -2276
rect 3440 -2356 3444 -2324
rect 3476 -2356 3480 -2324
rect 3440 -2404 3480 -2356
rect 3440 -2436 3444 -2404
rect 3476 -2436 3480 -2404
rect 3440 -2484 3480 -2436
rect 3440 -2516 3444 -2484
rect 3476 -2516 3480 -2484
rect 3440 -2564 3480 -2516
rect 3440 -2596 3444 -2564
rect 3476 -2596 3480 -2564
rect 3440 -2644 3480 -2596
rect 3440 -2676 3444 -2644
rect 3476 -2676 3480 -2644
rect 3440 -2724 3480 -2676
rect 3440 -2756 3444 -2724
rect 3476 -2756 3480 -2724
rect 3440 -2804 3480 -2756
rect 3440 -2836 3444 -2804
rect 3476 -2836 3480 -2804
rect 3440 -2884 3480 -2836
rect 3440 -2916 3444 -2884
rect 3476 -2916 3480 -2884
rect 3440 -2964 3480 -2916
rect 3440 -2996 3444 -2964
rect 3476 -2996 3480 -2964
rect 3440 -3044 3480 -2996
rect 3440 -3076 3444 -3044
rect 3476 -3076 3480 -3044
rect 3440 -3124 3480 -3076
rect 3440 -3156 3444 -3124
rect 3476 -3156 3480 -3124
rect 3440 -3204 3480 -3156
rect 3440 -3236 3444 -3204
rect 3476 -3236 3480 -3204
rect 3440 -3284 3480 -3236
rect 3440 -3316 3444 -3284
rect 3476 -3316 3480 -3284
rect 3440 -3364 3480 -3316
rect 3440 -3396 3444 -3364
rect 3476 -3396 3480 -3364
rect 3440 -3444 3480 -3396
rect 3440 -3476 3444 -3444
rect 3476 -3476 3480 -3444
rect 3440 -3524 3480 -3476
rect 3440 -3556 3444 -3524
rect 3476 -3556 3480 -3524
rect 3440 -3604 3480 -3556
rect 3440 -3636 3444 -3604
rect 3476 -3636 3480 -3604
rect 3440 -3684 3480 -3636
rect 3440 -3716 3444 -3684
rect 3476 -3716 3480 -3684
rect 3440 -3720 3480 -3716
rect 3520 1036 3560 1040
rect 3520 1004 3524 1036
rect 3556 1004 3560 1036
rect 3520 956 3560 1004
rect 3520 924 3524 956
rect 3556 924 3560 956
rect 3520 876 3560 924
rect 3520 844 3524 876
rect 3556 844 3560 876
rect 3520 796 3560 844
rect 3520 764 3524 796
rect 3556 764 3560 796
rect 3520 716 3560 764
rect 3520 684 3524 716
rect 3556 684 3560 716
rect 3520 636 3560 684
rect 3520 604 3524 636
rect 3556 604 3560 636
rect 3520 556 3560 604
rect 3520 524 3524 556
rect 3556 524 3560 556
rect 3520 476 3560 524
rect 3520 444 3524 476
rect 3556 444 3560 476
rect 3520 396 3560 444
rect 3520 364 3524 396
rect 3556 364 3560 396
rect 3520 316 3560 364
rect 3520 284 3524 316
rect 3556 284 3560 316
rect 3520 236 3560 284
rect 3520 204 3524 236
rect 3556 204 3560 236
rect 3520 156 3560 204
rect 3520 124 3524 156
rect 3556 124 3560 156
rect 3520 76 3560 124
rect 3520 44 3524 76
rect 3556 44 3560 76
rect 3520 -4 3560 44
rect 3520 -36 3524 -4
rect 3556 -36 3560 -4
rect 3520 -84 3560 -36
rect 3520 -116 3524 -84
rect 3556 -116 3560 -84
rect 3520 -164 3560 -116
rect 3520 -196 3524 -164
rect 3556 -196 3560 -164
rect 3520 -244 3560 -196
rect 3520 -276 3524 -244
rect 3556 -276 3560 -244
rect 3520 -324 3560 -276
rect 3520 -356 3524 -324
rect 3556 -356 3560 -324
rect 3520 -404 3560 -356
rect 3520 -436 3524 -404
rect 3556 -436 3560 -404
rect 3520 -484 3560 -436
rect 3520 -516 3524 -484
rect 3556 -516 3560 -484
rect 3520 -564 3560 -516
rect 3520 -596 3524 -564
rect 3556 -596 3560 -564
rect 3520 -644 3560 -596
rect 3520 -676 3524 -644
rect 3556 -676 3560 -644
rect 3520 -724 3560 -676
rect 3520 -756 3524 -724
rect 3556 -756 3560 -724
rect 3520 -804 3560 -756
rect 3520 -836 3524 -804
rect 3556 -836 3560 -804
rect 3520 -884 3560 -836
rect 3520 -916 3524 -884
rect 3556 -916 3560 -884
rect 3520 -964 3560 -916
rect 3520 -996 3524 -964
rect 3556 -996 3560 -964
rect 3520 -1044 3560 -996
rect 3520 -1076 3524 -1044
rect 3556 -1076 3560 -1044
rect 3520 -1124 3560 -1076
rect 3520 -1156 3524 -1124
rect 3556 -1156 3560 -1124
rect 3520 -1204 3560 -1156
rect 3520 -1236 3524 -1204
rect 3556 -1236 3560 -1204
rect 3520 -1284 3560 -1236
rect 3520 -1316 3524 -1284
rect 3556 -1316 3560 -1284
rect 3520 -1364 3560 -1316
rect 3520 -1396 3524 -1364
rect 3556 -1396 3560 -1364
rect 3520 -1444 3560 -1396
rect 3520 -1476 3524 -1444
rect 3556 -1476 3560 -1444
rect 3520 -1524 3560 -1476
rect 3520 -1556 3524 -1524
rect 3556 -1556 3560 -1524
rect 3520 -1604 3560 -1556
rect 3520 -1636 3524 -1604
rect 3556 -1636 3560 -1604
rect 3520 -1684 3560 -1636
rect 3520 -1716 3524 -1684
rect 3556 -1716 3560 -1684
rect 3520 -1764 3560 -1716
rect 3520 -1796 3524 -1764
rect 3556 -1796 3560 -1764
rect 3520 -1844 3560 -1796
rect 3520 -1876 3524 -1844
rect 3556 -1876 3560 -1844
rect 3520 -1924 3560 -1876
rect 3520 -1956 3524 -1924
rect 3556 -1956 3560 -1924
rect 3520 -2004 3560 -1956
rect 3520 -2036 3524 -2004
rect 3556 -2036 3560 -2004
rect 3520 -2084 3560 -2036
rect 3520 -2116 3524 -2084
rect 3556 -2116 3560 -2084
rect 3520 -2164 3560 -2116
rect 3520 -2196 3524 -2164
rect 3556 -2196 3560 -2164
rect 3520 -2244 3560 -2196
rect 3520 -2276 3524 -2244
rect 3556 -2276 3560 -2244
rect 3520 -2324 3560 -2276
rect 3520 -2356 3524 -2324
rect 3556 -2356 3560 -2324
rect 3520 -2404 3560 -2356
rect 3520 -2436 3524 -2404
rect 3556 -2436 3560 -2404
rect 3520 -2484 3560 -2436
rect 3520 -2516 3524 -2484
rect 3556 -2516 3560 -2484
rect 3520 -2564 3560 -2516
rect 3520 -2596 3524 -2564
rect 3556 -2596 3560 -2564
rect 3520 -2644 3560 -2596
rect 3520 -2676 3524 -2644
rect 3556 -2676 3560 -2644
rect 3520 -2724 3560 -2676
rect 3520 -2756 3524 -2724
rect 3556 -2756 3560 -2724
rect 3520 -2804 3560 -2756
rect 3520 -2836 3524 -2804
rect 3556 -2836 3560 -2804
rect 3520 -2884 3560 -2836
rect 3520 -2916 3524 -2884
rect 3556 -2916 3560 -2884
rect 3520 -2964 3560 -2916
rect 3520 -2996 3524 -2964
rect 3556 -2996 3560 -2964
rect 3520 -3044 3560 -2996
rect 3520 -3076 3524 -3044
rect 3556 -3076 3560 -3044
rect 3520 -3124 3560 -3076
rect 3520 -3156 3524 -3124
rect 3556 -3156 3560 -3124
rect 3520 -3204 3560 -3156
rect 3520 -3236 3524 -3204
rect 3556 -3236 3560 -3204
rect 3520 -3284 3560 -3236
rect 3520 -3316 3524 -3284
rect 3556 -3316 3560 -3284
rect 3520 -3364 3560 -3316
rect 3520 -3396 3524 -3364
rect 3556 -3396 3560 -3364
rect 3520 -3444 3560 -3396
rect 3520 -3476 3524 -3444
rect 3556 -3476 3560 -3444
rect 3520 -3524 3560 -3476
rect 3520 -3556 3524 -3524
rect 3556 -3556 3560 -3524
rect 3520 -3604 3560 -3556
rect 3520 -3636 3524 -3604
rect 3556 -3636 3560 -3604
rect 3520 -3684 3560 -3636
rect 3520 -3716 3524 -3684
rect 3556 -3716 3560 -3684
rect 3520 -3720 3560 -3716
rect 3600 1036 3640 1040
rect 3600 1004 3604 1036
rect 3636 1004 3640 1036
rect 3600 956 3640 1004
rect 3600 924 3604 956
rect 3636 924 3640 956
rect 3600 876 3640 924
rect 3600 844 3604 876
rect 3636 844 3640 876
rect 3600 796 3640 844
rect 3600 764 3604 796
rect 3636 764 3640 796
rect 3600 716 3640 764
rect 3600 684 3604 716
rect 3636 684 3640 716
rect 3600 636 3640 684
rect 3600 604 3604 636
rect 3636 604 3640 636
rect 3600 556 3640 604
rect 3600 524 3604 556
rect 3636 524 3640 556
rect 3600 476 3640 524
rect 3600 444 3604 476
rect 3636 444 3640 476
rect 3600 396 3640 444
rect 3600 364 3604 396
rect 3636 364 3640 396
rect 3600 316 3640 364
rect 3600 284 3604 316
rect 3636 284 3640 316
rect 3600 236 3640 284
rect 3600 204 3604 236
rect 3636 204 3640 236
rect 3600 156 3640 204
rect 3600 124 3604 156
rect 3636 124 3640 156
rect 3600 76 3640 124
rect 3600 44 3604 76
rect 3636 44 3640 76
rect 3600 -4 3640 44
rect 3600 -36 3604 -4
rect 3636 -36 3640 -4
rect 3600 -84 3640 -36
rect 3600 -116 3604 -84
rect 3636 -116 3640 -84
rect 3600 -164 3640 -116
rect 3600 -196 3604 -164
rect 3636 -196 3640 -164
rect 3600 -244 3640 -196
rect 3600 -276 3604 -244
rect 3636 -276 3640 -244
rect 3600 -324 3640 -276
rect 3600 -356 3604 -324
rect 3636 -356 3640 -324
rect 3600 -404 3640 -356
rect 3600 -436 3604 -404
rect 3636 -436 3640 -404
rect 3600 -484 3640 -436
rect 3600 -516 3604 -484
rect 3636 -516 3640 -484
rect 3600 -564 3640 -516
rect 3600 -596 3604 -564
rect 3636 -596 3640 -564
rect 3600 -644 3640 -596
rect 3600 -676 3604 -644
rect 3636 -676 3640 -644
rect 3600 -724 3640 -676
rect 3600 -756 3604 -724
rect 3636 -756 3640 -724
rect 3600 -804 3640 -756
rect 3600 -836 3604 -804
rect 3636 -836 3640 -804
rect 3600 -884 3640 -836
rect 3600 -916 3604 -884
rect 3636 -916 3640 -884
rect 3600 -964 3640 -916
rect 3600 -996 3604 -964
rect 3636 -996 3640 -964
rect 3600 -1044 3640 -996
rect 3600 -1076 3604 -1044
rect 3636 -1076 3640 -1044
rect 3600 -1124 3640 -1076
rect 3600 -1156 3604 -1124
rect 3636 -1156 3640 -1124
rect 3600 -1204 3640 -1156
rect 3600 -1236 3604 -1204
rect 3636 -1236 3640 -1204
rect 3600 -1284 3640 -1236
rect 3600 -1316 3604 -1284
rect 3636 -1316 3640 -1284
rect 3600 -1364 3640 -1316
rect 3600 -1396 3604 -1364
rect 3636 -1396 3640 -1364
rect 3600 -1444 3640 -1396
rect 3600 -1476 3604 -1444
rect 3636 -1476 3640 -1444
rect 3600 -1524 3640 -1476
rect 3600 -1556 3604 -1524
rect 3636 -1556 3640 -1524
rect 3600 -1604 3640 -1556
rect 3600 -1636 3604 -1604
rect 3636 -1636 3640 -1604
rect 3600 -1684 3640 -1636
rect 3600 -1716 3604 -1684
rect 3636 -1716 3640 -1684
rect 3600 -1764 3640 -1716
rect 3600 -1796 3604 -1764
rect 3636 -1796 3640 -1764
rect 3600 -1844 3640 -1796
rect 3600 -1876 3604 -1844
rect 3636 -1876 3640 -1844
rect 3600 -1924 3640 -1876
rect 3600 -1956 3604 -1924
rect 3636 -1956 3640 -1924
rect 3600 -2004 3640 -1956
rect 3600 -2036 3604 -2004
rect 3636 -2036 3640 -2004
rect 3600 -2084 3640 -2036
rect 3600 -2116 3604 -2084
rect 3636 -2116 3640 -2084
rect 3600 -2164 3640 -2116
rect 3600 -2196 3604 -2164
rect 3636 -2196 3640 -2164
rect 3600 -2244 3640 -2196
rect 3600 -2276 3604 -2244
rect 3636 -2276 3640 -2244
rect 3600 -2324 3640 -2276
rect 3600 -2356 3604 -2324
rect 3636 -2356 3640 -2324
rect 3600 -2404 3640 -2356
rect 3600 -2436 3604 -2404
rect 3636 -2436 3640 -2404
rect 3600 -2484 3640 -2436
rect 3600 -2516 3604 -2484
rect 3636 -2516 3640 -2484
rect 3600 -2564 3640 -2516
rect 3600 -2596 3604 -2564
rect 3636 -2596 3640 -2564
rect 3600 -2644 3640 -2596
rect 3600 -2676 3604 -2644
rect 3636 -2676 3640 -2644
rect 3600 -2724 3640 -2676
rect 3600 -2756 3604 -2724
rect 3636 -2756 3640 -2724
rect 3600 -2804 3640 -2756
rect 3600 -2836 3604 -2804
rect 3636 -2836 3640 -2804
rect 3600 -2884 3640 -2836
rect 3600 -2916 3604 -2884
rect 3636 -2916 3640 -2884
rect 3600 -2964 3640 -2916
rect 3600 -2996 3604 -2964
rect 3636 -2996 3640 -2964
rect 3600 -3044 3640 -2996
rect 3600 -3076 3604 -3044
rect 3636 -3076 3640 -3044
rect 3600 -3124 3640 -3076
rect 3600 -3156 3604 -3124
rect 3636 -3156 3640 -3124
rect 3600 -3204 3640 -3156
rect 3600 -3236 3604 -3204
rect 3636 -3236 3640 -3204
rect 3600 -3284 3640 -3236
rect 3600 -3316 3604 -3284
rect 3636 -3316 3640 -3284
rect 3600 -3364 3640 -3316
rect 3600 -3396 3604 -3364
rect 3636 -3396 3640 -3364
rect 3600 -3444 3640 -3396
rect 3600 -3476 3604 -3444
rect 3636 -3476 3640 -3444
rect 3600 -3524 3640 -3476
rect 3600 -3556 3604 -3524
rect 3636 -3556 3640 -3524
rect 3600 -3604 3640 -3556
rect 3600 -3636 3604 -3604
rect 3636 -3636 3640 -3604
rect 3600 -3684 3640 -3636
rect 3600 -3716 3604 -3684
rect 3636 -3716 3640 -3684
rect 3600 -3720 3640 -3716
rect 3680 1036 3720 1040
rect 3680 1004 3684 1036
rect 3716 1004 3720 1036
rect 3680 956 3720 1004
rect 3680 924 3684 956
rect 3716 924 3720 956
rect 3680 876 3720 924
rect 3680 844 3684 876
rect 3716 844 3720 876
rect 3680 796 3720 844
rect 3680 764 3684 796
rect 3716 764 3720 796
rect 3680 716 3720 764
rect 3680 684 3684 716
rect 3716 684 3720 716
rect 3680 636 3720 684
rect 3680 604 3684 636
rect 3716 604 3720 636
rect 3680 556 3720 604
rect 3680 524 3684 556
rect 3716 524 3720 556
rect 3680 476 3720 524
rect 3680 444 3684 476
rect 3716 444 3720 476
rect 3680 396 3720 444
rect 3680 364 3684 396
rect 3716 364 3720 396
rect 3680 316 3720 364
rect 3680 284 3684 316
rect 3716 284 3720 316
rect 3680 236 3720 284
rect 3680 204 3684 236
rect 3716 204 3720 236
rect 3680 156 3720 204
rect 3680 124 3684 156
rect 3716 124 3720 156
rect 3680 76 3720 124
rect 3680 44 3684 76
rect 3716 44 3720 76
rect 3680 -4 3720 44
rect 3680 -36 3684 -4
rect 3716 -36 3720 -4
rect 3680 -84 3720 -36
rect 3680 -116 3684 -84
rect 3716 -116 3720 -84
rect 3680 -164 3720 -116
rect 3680 -196 3684 -164
rect 3716 -196 3720 -164
rect 3680 -244 3720 -196
rect 3680 -276 3684 -244
rect 3716 -276 3720 -244
rect 3680 -324 3720 -276
rect 3680 -356 3684 -324
rect 3716 -356 3720 -324
rect 3680 -404 3720 -356
rect 3680 -436 3684 -404
rect 3716 -436 3720 -404
rect 3680 -484 3720 -436
rect 3680 -516 3684 -484
rect 3716 -516 3720 -484
rect 3680 -564 3720 -516
rect 3680 -596 3684 -564
rect 3716 -596 3720 -564
rect 3680 -644 3720 -596
rect 3680 -676 3684 -644
rect 3716 -676 3720 -644
rect 3680 -724 3720 -676
rect 3680 -756 3684 -724
rect 3716 -756 3720 -724
rect 3680 -804 3720 -756
rect 3680 -836 3684 -804
rect 3716 -836 3720 -804
rect 3680 -884 3720 -836
rect 3680 -916 3684 -884
rect 3716 -916 3720 -884
rect 3680 -964 3720 -916
rect 3680 -996 3684 -964
rect 3716 -996 3720 -964
rect 3680 -1044 3720 -996
rect 3680 -1076 3684 -1044
rect 3716 -1076 3720 -1044
rect 3680 -1124 3720 -1076
rect 3680 -1156 3684 -1124
rect 3716 -1156 3720 -1124
rect 3680 -1204 3720 -1156
rect 3680 -1236 3684 -1204
rect 3716 -1236 3720 -1204
rect 3680 -1284 3720 -1236
rect 3680 -1316 3684 -1284
rect 3716 -1316 3720 -1284
rect 3680 -1364 3720 -1316
rect 3680 -1396 3684 -1364
rect 3716 -1396 3720 -1364
rect 3680 -1444 3720 -1396
rect 3680 -1476 3684 -1444
rect 3716 -1476 3720 -1444
rect 3680 -1524 3720 -1476
rect 3680 -1556 3684 -1524
rect 3716 -1556 3720 -1524
rect 3680 -1604 3720 -1556
rect 3680 -1636 3684 -1604
rect 3716 -1636 3720 -1604
rect 3680 -1684 3720 -1636
rect 3680 -1716 3684 -1684
rect 3716 -1716 3720 -1684
rect 3680 -1764 3720 -1716
rect 3680 -1796 3684 -1764
rect 3716 -1796 3720 -1764
rect 3680 -1844 3720 -1796
rect 3680 -1876 3684 -1844
rect 3716 -1876 3720 -1844
rect 3680 -1924 3720 -1876
rect 3680 -1956 3684 -1924
rect 3716 -1956 3720 -1924
rect 3680 -2004 3720 -1956
rect 3680 -2036 3684 -2004
rect 3716 -2036 3720 -2004
rect 3680 -2084 3720 -2036
rect 3680 -2116 3684 -2084
rect 3716 -2116 3720 -2084
rect 3680 -2164 3720 -2116
rect 3680 -2196 3684 -2164
rect 3716 -2196 3720 -2164
rect 3680 -2244 3720 -2196
rect 3680 -2276 3684 -2244
rect 3716 -2276 3720 -2244
rect 3680 -2324 3720 -2276
rect 3680 -2356 3684 -2324
rect 3716 -2356 3720 -2324
rect 3680 -2404 3720 -2356
rect 3680 -2436 3684 -2404
rect 3716 -2436 3720 -2404
rect 3680 -2484 3720 -2436
rect 3680 -2516 3684 -2484
rect 3716 -2516 3720 -2484
rect 3680 -2564 3720 -2516
rect 3680 -2596 3684 -2564
rect 3716 -2596 3720 -2564
rect 3680 -2644 3720 -2596
rect 3680 -2676 3684 -2644
rect 3716 -2676 3720 -2644
rect 3680 -2724 3720 -2676
rect 3680 -2756 3684 -2724
rect 3716 -2756 3720 -2724
rect 3680 -2804 3720 -2756
rect 3680 -2836 3684 -2804
rect 3716 -2836 3720 -2804
rect 3680 -2884 3720 -2836
rect 3680 -2916 3684 -2884
rect 3716 -2916 3720 -2884
rect 3680 -2964 3720 -2916
rect 3680 -2996 3684 -2964
rect 3716 -2996 3720 -2964
rect 3680 -3044 3720 -2996
rect 3680 -3076 3684 -3044
rect 3716 -3076 3720 -3044
rect 3680 -3124 3720 -3076
rect 3680 -3156 3684 -3124
rect 3716 -3156 3720 -3124
rect 3680 -3204 3720 -3156
rect 3680 -3236 3684 -3204
rect 3716 -3236 3720 -3204
rect 3680 -3284 3720 -3236
rect 3680 -3316 3684 -3284
rect 3716 -3316 3720 -3284
rect 3680 -3364 3720 -3316
rect 3680 -3396 3684 -3364
rect 3716 -3396 3720 -3364
rect 3680 -3444 3720 -3396
rect 3680 -3476 3684 -3444
rect 3716 -3476 3720 -3444
rect 3680 -3524 3720 -3476
rect 3680 -3556 3684 -3524
rect 3716 -3556 3720 -3524
rect 3680 -3604 3720 -3556
rect 3680 -3636 3684 -3604
rect 3716 -3636 3720 -3604
rect 3680 -3684 3720 -3636
rect 3680 -3716 3684 -3684
rect 3716 -3716 3720 -3684
rect 3680 -3720 3720 -3716
rect 3760 1036 3800 1040
rect 3760 1004 3764 1036
rect 3796 1004 3800 1036
rect 3760 956 3800 1004
rect 3760 924 3764 956
rect 3796 924 3800 956
rect 3760 876 3800 924
rect 3760 844 3764 876
rect 3796 844 3800 876
rect 3760 796 3800 844
rect 3760 764 3764 796
rect 3796 764 3800 796
rect 3760 716 3800 764
rect 3760 684 3764 716
rect 3796 684 3800 716
rect 3760 636 3800 684
rect 3760 604 3764 636
rect 3796 604 3800 636
rect 3760 556 3800 604
rect 3760 524 3764 556
rect 3796 524 3800 556
rect 3760 476 3800 524
rect 3760 444 3764 476
rect 3796 444 3800 476
rect 3760 396 3800 444
rect 3760 364 3764 396
rect 3796 364 3800 396
rect 3760 316 3800 364
rect 3760 284 3764 316
rect 3796 284 3800 316
rect 3760 236 3800 284
rect 3760 204 3764 236
rect 3796 204 3800 236
rect 3760 156 3800 204
rect 3760 124 3764 156
rect 3796 124 3800 156
rect 3760 76 3800 124
rect 3760 44 3764 76
rect 3796 44 3800 76
rect 3760 -4 3800 44
rect 3760 -36 3764 -4
rect 3796 -36 3800 -4
rect 3760 -84 3800 -36
rect 3760 -116 3764 -84
rect 3796 -116 3800 -84
rect 3760 -164 3800 -116
rect 3760 -196 3764 -164
rect 3796 -196 3800 -164
rect 3760 -244 3800 -196
rect 3760 -276 3764 -244
rect 3796 -276 3800 -244
rect 3760 -324 3800 -276
rect 3760 -356 3764 -324
rect 3796 -356 3800 -324
rect 3760 -404 3800 -356
rect 3760 -436 3764 -404
rect 3796 -436 3800 -404
rect 3760 -484 3800 -436
rect 3760 -516 3764 -484
rect 3796 -516 3800 -484
rect 3760 -564 3800 -516
rect 3760 -596 3764 -564
rect 3796 -596 3800 -564
rect 3760 -644 3800 -596
rect 3760 -676 3764 -644
rect 3796 -676 3800 -644
rect 3760 -724 3800 -676
rect 3760 -756 3764 -724
rect 3796 -756 3800 -724
rect 3760 -804 3800 -756
rect 3760 -836 3764 -804
rect 3796 -836 3800 -804
rect 3760 -884 3800 -836
rect 3760 -916 3764 -884
rect 3796 -916 3800 -884
rect 3760 -964 3800 -916
rect 3760 -996 3764 -964
rect 3796 -996 3800 -964
rect 3760 -1044 3800 -996
rect 3760 -1076 3764 -1044
rect 3796 -1076 3800 -1044
rect 3760 -1124 3800 -1076
rect 3760 -1156 3764 -1124
rect 3796 -1156 3800 -1124
rect 3760 -1204 3800 -1156
rect 3760 -1236 3764 -1204
rect 3796 -1236 3800 -1204
rect 3760 -1284 3800 -1236
rect 3760 -1316 3764 -1284
rect 3796 -1316 3800 -1284
rect 3760 -1364 3800 -1316
rect 3760 -1396 3764 -1364
rect 3796 -1396 3800 -1364
rect 3760 -1444 3800 -1396
rect 3760 -1476 3764 -1444
rect 3796 -1476 3800 -1444
rect 3760 -1524 3800 -1476
rect 3760 -1556 3764 -1524
rect 3796 -1556 3800 -1524
rect 3760 -1604 3800 -1556
rect 3760 -1636 3764 -1604
rect 3796 -1636 3800 -1604
rect 3760 -1684 3800 -1636
rect 3760 -1716 3764 -1684
rect 3796 -1716 3800 -1684
rect 3760 -1764 3800 -1716
rect 3760 -1796 3764 -1764
rect 3796 -1796 3800 -1764
rect 3760 -1844 3800 -1796
rect 3760 -1876 3764 -1844
rect 3796 -1876 3800 -1844
rect 3760 -1924 3800 -1876
rect 3760 -1956 3764 -1924
rect 3796 -1956 3800 -1924
rect 3760 -2004 3800 -1956
rect 3760 -2036 3764 -2004
rect 3796 -2036 3800 -2004
rect 3760 -2084 3800 -2036
rect 3760 -2116 3764 -2084
rect 3796 -2116 3800 -2084
rect 3760 -2164 3800 -2116
rect 3760 -2196 3764 -2164
rect 3796 -2196 3800 -2164
rect 3760 -2244 3800 -2196
rect 3760 -2276 3764 -2244
rect 3796 -2276 3800 -2244
rect 3760 -2324 3800 -2276
rect 3760 -2356 3764 -2324
rect 3796 -2356 3800 -2324
rect 3760 -2404 3800 -2356
rect 3760 -2436 3764 -2404
rect 3796 -2436 3800 -2404
rect 3760 -2484 3800 -2436
rect 3760 -2516 3764 -2484
rect 3796 -2516 3800 -2484
rect 3760 -2564 3800 -2516
rect 3760 -2596 3764 -2564
rect 3796 -2596 3800 -2564
rect 3760 -2644 3800 -2596
rect 3760 -2676 3764 -2644
rect 3796 -2676 3800 -2644
rect 3760 -2724 3800 -2676
rect 3760 -2756 3764 -2724
rect 3796 -2756 3800 -2724
rect 3760 -2804 3800 -2756
rect 3760 -2836 3764 -2804
rect 3796 -2836 3800 -2804
rect 3760 -2884 3800 -2836
rect 3760 -2916 3764 -2884
rect 3796 -2916 3800 -2884
rect 3760 -2964 3800 -2916
rect 3760 -2996 3764 -2964
rect 3796 -2996 3800 -2964
rect 3760 -3044 3800 -2996
rect 3760 -3076 3764 -3044
rect 3796 -3076 3800 -3044
rect 3760 -3124 3800 -3076
rect 3760 -3156 3764 -3124
rect 3796 -3156 3800 -3124
rect 3760 -3204 3800 -3156
rect 3760 -3236 3764 -3204
rect 3796 -3236 3800 -3204
rect 3760 -3284 3800 -3236
rect 3760 -3316 3764 -3284
rect 3796 -3316 3800 -3284
rect 3760 -3364 3800 -3316
rect 3760 -3396 3764 -3364
rect 3796 -3396 3800 -3364
rect 3760 -3444 3800 -3396
rect 3760 -3476 3764 -3444
rect 3796 -3476 3800 -3444
rect 3760 -3524 3800 -3476
rect 3760 -3556 3764 -3524
rect 3796 -3556 3800 -3524
rect 3760 -3604 3800 -3556
rect 3760 -3636 3764 -3604
rect 3796 -3636 3800 -3604
rect 3760 -3684 3800 -3636
rect 3760 -3716 3764 -3684
rect 3796 -3716 3800 -3684
rect 3760 -3720 3800 -3716
rect 3840 1036 3880 1040
rect 3840 1004 3844 1036
rect 3876 1004 3880 1036
rect 3840 956 3880 1004
rect 3840 924 3844 956
rect 3876 924 3880 956
rect 3840 876 3880 924
rect 3840 844 3844 876
rect 3876 844 3880 876
rect 3840 796 3880 844
rect 3840 764 3844 796
rect 3876 764 3880 796
rect 3840 716 3880 764
rect 3840 684 3844 716
rect 3876 684 3880 716
rect 3840 636 3880 684
rect 3840 604 3844 636
rect 3876 604 3880 636
rect 3840 556 3880 604
rect 3840 524 3844 556
rect 3876 524 3880 556
rect 3840 476 3880 524
rect 3840 444 3844 476
rect 3876 444 3880 476
rect 3840 396 3880 444
rect 3840 364 3844 396
rect 3876 364 3880 396
rect 3840 316 3880 364
rect 3840 284 3844 316
rect 3876 284 3880 316
rect 3840 236 3880 284
rect 3840 204 3844 236
rect 3876 204 3880 236
rect 3840 156 3880 204
rect 3840 124 3844 156
rect 3876 124 3880 156
rect 3840 76 3880 124
rect 3840 44 3844 76
rect 3876 44 3880 76
rect 3840 -4 3880 44
rect 3840 -36 3844 -4
rect 3876 -36 3880 -4
rect 3840 -84 3880 -36
rect 3840 -116 3844 -84
rect 3876 -116 3880 -84
rect 3840 -164 3880 -116
rect 3840 -196 3844 -164
rect 3876 -196 3880 -164
rect 3840 -244 3880 -196
rect 3840 -276 3844 -244
rect 3876 -276 3880 -244
rect 3840 -324 3880 -276
rect 3840 -356 3844 -324
rect 3876 -356 3880 -324
rect 3840 -404 3880 -356
rect 3840 -436 3844 -404
rect 3876 -436 3880 -404
rect 3840 -484 3880 -436
rect 3840 -516 3844 -484
rect 3876 -516 3880 -484
rect 3840 -564 3880 -516
rect 3840 -596 3844 -564
rect 3876 -596 3880 -564
rect 3840 -644 3880 -596
rect 3840 -676 3844 -644
rect 3876 -676 3880 -644
rect 3840 -724 3880 -676
rect 3840 -756 3844 -724
rect 3876 -756 3880 -724
rect 3840 -804 3880 -756
rect 3840 -836 3844 -804
rect 3876 -836 3880 -804
rect 3840 -884 3880 -836
rect 3840 -916 3844 -884
rect 3876 -916 3880 -884
rect 3840 -964 3880 -916
rect 3840 -996 3844 -964
rect 3876 -996 3880 -964
rect 3840 -1044 3880 -996
rect 3840 -1076 3844 -1044
rect 3876 -1076 3880 -1044
rect 3840 -1124 3880 -1076
rect 3840 -1156 3844 -1124
rect 3876 -1156 3880 -1124
rect 3840 -1204 3880 -1156
rect 3840 -1236 3844 -1204
rect 3876 -1236 3880 -1204
rect 3840 -1284 3880 -1236
rect 3840 -1316 3844 -1284
rect 3876 -1316 3880 -1284
rect 3840 -1364 3880 -1316
rect 3840 -1396 3844 -1364
rect 3876 -1396 3880 -1364
rect 3840 -1444 3880 -1396
rect 3840 -1476 3844 -1444
rect 3876 -1476 3880 -1444
rect 3840 -1524 3880 -1476
rect 3840 -1556 3844 -1524
rect 3876 -1556 3880 -1524
rect 3840 -1604 3880 -1556
rect 3840 -1636 3844 -1604
rect 3876 -1636 3880 -1604
rect 3840 -1684 3880 -1636
rect 3840 -1716 3844 -1684
rect 3876 -1716 3880 -1684
rect 3840 -1764 3880 -1716
rect 3840 -1796 3844 -1764
rect 3876 -1796 3880 -1764
rect 3840 -1844 3880 -1796
rect 3840 -1876 3844 -1844
rect 3876 -1876 3880 -1844
rect 3840 -1924 3880 -1876
rect 3840 -1956 3844 -1924
rect 3876 -1956 3880 -1924
rect 3840 -2004 3880 -1956
rect 3840 -2036 3844 -2004
rect 3876 -2036 3880 -2004
rect 3840 -2084 3880 -2036
rect 3840 -2116 3844 -2084
rect 3876 -2116 3880 -2084
rect 3840 -2164 3880 -2116
rect 3840 -2196 3844 -2164
rect 3876 -2196 3880 -2164
rect 3840 -2244 3880 -2196
rect 3840 -2276 3844 -2244
rect 3876 -2276 3880 -2244
rect 3840 -2324 3880 -2276
rect 3840 -2356 3844 -2324
rect 3876 -2356 3880 -2324
rect 3840 -2404 3880 -2356
rect 3840 -2436 3844 -2404
rect 3876 -2436 3880 -2404
rect 3840 -2484 3880 -2436
rect 3840 -2516 3844 -2484
rect 3876 -2516 3880 -2484
rect 3840 -2564 3880 -2516
rect 3840 -2596 3844 -2564
rect 3876 -2596 3880 -2564
rect 3840 -2644 3880 -2596
rect 3840 -2676 3844 -2644
rect 3876 -2676 3880 -2644
rect 3840 -2724 3880 -2676
rect 3840 -2756 3844 -2724
rect 3876 -2756 3880 -2724
rect 3840 -2804 3880 -2756
rect 3840 -2836 3844 -2804
rect 3876 -2836 3880 -2804
rect 3840 -2884 3880 -2836
rect 3840 -2916 3844 -2884
rect 3876 -2916 3880 -2884
rect 3840 -2964 3880 -2916
rect 3840 -2996 3844 -2964
rect 3876 -2996 3880 -2964
rect 3840 -3044 3880 -2996
rect 3840 -3076 3844 -3044
rect 3876 -3076 3880 -3044
rect 3840 -3124 3880 -3076
rect 3840 -3156 3844 -3124
rect 3876 -3156 3880 -3124
rect 3840 -3204 3880 -3156
rect 3840 -3236 3844 -3204
rect 3876 -3236 3880 -3204
rect 3840 -3284 3880 -3236
rect 3840 -3316 3844 -3284
rect 3876 -3316 3880 -3284
rect 3840 -3364 3880 -3316
rect 3840 -3396 3844 -3364
rect 3876 -3396 3880 -3364
rect 3840 -3444 3880 -3396
rect 3840 -3476 3844 -3444
rect 3876 -3476 3880 -3444
rect 3840 -3524 3880 -3476
rect 3840 -3556 3844 -3524
rect 3876 -3556 3880 -3524
rect 3840 -3604 3880 -3556
rect 3840 -3636 3844 -3604
rect 3876 -3636 3880 -3604
rect 3840 -3684 3880 -3636
rect 3840 -3716 3844 -3684
rect 3876 -3716 3880 -3684
rect 3840 -3720 3880 -3716
rect 3920 1036 3960 1040
rect 3920 1004 3924 1036
rect 3956 1004 3960 1036
rect 3920 956 3960 1004
rect 3920 924 3924 956
rect 3956 924 3960 956
rect 3920 876 3960 924
rect 3920 844 3924 876
rect 3956 844 3960 876
rect 3920 796 3960 844
rect 3920 764 3924 796
rect 3956 764 3960 796
rect 3920 716 3960 764
rect 3920 684 3924 716
rect 3956 684 3960 716
rect 3920 636 3960 684
rect 3920 604 3924 636
rect 3956 604 3960 636
rect 3920 556 3960 604
rect 3920 524 3924 556
rect 3956 524 3960 556
rect 3920 476 3960 524
rect 3920 444 3924 476
rect 3956 444 3960 476
rect 3920 396 3960 444
rect 3920 364 3924 396
rect 3956 364 3960 396
rect 3920 316 3960 364
rect 3920 284 3924 316
rect 3956 284 3960 316
rect 3920 236 3960 284
rect 3920 204 3924 236
rect 3956 204 3960 236
rect 3920 156 3960 204
rect 3920 124 3924 156
rect 3956 124 3960 156
rect 3920 76 3960 124
rect 3920 44 3924 76
rect 3956 44 3960 76
rect 3920 -4 3960 44
rect 3920 -36 3924 -4
rect 3956 -36 3960 -4
rect 3920 -84 3960 -36
rect 3920 -116 3924 -84
rect 3956 -116 3960 -84
rect 3920 -164 3960 -116
rect 3920 -196 3924 -164
rect 3956 -196 3960 -164
rect 3920 -244 3960 -196
rect 3920 -276 3924 -244
rect 3956 -276 3960 -244
rect 3920 -324 3960 -276
rect 3920 -356 3924 -324
rect 3956 -356 3960 -324
rect 3920 -404 3960 -356
rect 3920 -436 3924 -404
rect 3956 -436 3960 -404
rect 3920 -484 3960 -436
rect 3920 -516 3924 -484
rect 3956 -516 3960 -484
rect 3920 -564 3960 -516
rect 3920 -596 3924 -564
rect 3956 -596 3960 -564
rect 3920 -644 3960 -596
rect 3920 -676 3924 -644
rect 3956 -676 3960 -644
rect 3920 -724 3960 -676
rect 3920 -756 3924 -724
rect 3956 -756 3960 -724
rect 3920 -804 3960 -756
rect 3920 -836 3924 -804
rect 3956 -836 3960 -804
rect 3920 -884 3960 -836
rect 3920 -916 3924 -884
rect 3956 -916 3960 -884
rect 3920 -964 3960 -916
rect 3920 -996 3924 -964
rect 3956 -996 3960 -964
rect 3920 -1044 3960 -996
rect 3920 -1076 3924 -1044
rect 3956 -1076 3960 -1044
rect 3920 -1124 3960 -1076
rect 3920 -1156 3924 -1124
rect 3956 -1156 3960 -1124
rect 3920 -1204 3960 -1156
rect 3920 -1236 3924 -1204
rect 3956 -1236 3960 -1204
rect 3920 -1284 3960 -1236
rect 3920 -1316 3924 -1284
rect 3956 -1316 3960 -1284
rect 3920 -1364 3960 -1316
rect 3920 -1396 3924 -1364
rect 3956 -1396 3960 -1364
rect 3920 -1444 3960 -1396
rect 3920 -1476 3924 -1444
rect 3956 -1476 3960 -1444
rect 3920 -1524 3960 -1476
rect 3920 -1556 3924 -1524
rect 3956 -1556 3960 -1524
rect 3920 -1604 3960 -1556
rect 3920 -1636 3924 -1604
rect 3956 -1636 3960 -1604
rect 3920 -1684 3960 -1636
rect 3920 -1716 3924 -1684
rect 3956 -1716 3960 -1684
rect 3920 -1764 3960 -1716
rect 3920 -1796 3924 -1764
rect 3956 -1796 3960 -1764
rect 3920 -1844 3960 -1796
rect 3920 -1876 3924 -1844
rect 3956 -1876 3960 -1844
rect 3920 -1924 3960 -1876
rect 3920 -1956 3924 -1924
rect 3956 -1956 3960 -1924
rect 3920 -2004 3960 -1956
rect 3920 -2036 3924 -2004
rect 3956 -2036 3960 -2004
rect 3920 -2084 3960 -2036
rect 3920 -2116 3924 -2084
rect 3956 -2116 3960 -2084
rect 3920 -2164 3960 -2116
rect 3920 -2196 3924 -2164
rect 3956 -2196 3960 -2164
rect 3920 -2244 3960 -2196
rect 3920 -2276 3924 -2244
rect 3956 -2276 3960 -2244
rect 3920 -2324 3960 -2276
rect 3920 -2356 3924 -2324
rect 3956 -2356 3960 -2324
rect 3920 -2404 3960 -2356
rect 3920 -2436 3924 -2404
rect 3956 -2436 3960 -2404
rect 3920 -2484 3960 -2436
rect 3920 -2516 3924 -2484
rect 3956 -2516 3960 -2484
rect 3920 -2564 3960 -2516
rect 3920 -2596 3924 -2564
rect 3956 -2596 3960 -2564
rect 3920 -2644 3960 -2596
rect 3920 -2676 3924 -2644
rect 3956 -2676 3960 -2644
rect 3920 -2724 3960 -2676
rect 3920 -2756 3924 -2724
rect 3956 -2756 3960 -2724
rect 3920 -2804 3960 -2756
rect 3920 -2836 3924 -2804
rect 3956 -2836 3960 -2804
rect 3920 -2884 3960 -2836
rect 3920 -2916 3924 -2884
rect 3956 -2916 3960 -2884
rect 3920 -2964 3960 -2916
rect 3920 -2996 3924 -2964
rect 3956 -2996 3960 -2964
rect 3920 -3044 3960 -2996
rect 3920 -3076 3924 -3044
rect 3956 -3076 3960 -3044
rect 3920 -3124 3960 -3076
rect 3920 -3156 3924 -3124
rect 3956 -3156 3960 -3124
rect 3920 -3204 3960 -3156
rect 3920 -3236 3924 -3204
rect 3956 -3236 3960 -3204
rect 3920 -3284 3960 -3236
rect 3920 -3316 3924 -3284
rect 3956 -3316 3960 -3284
rect 3920 -3364 3960 -3316
rect 3920 -3396 3924 -3364
rect 3956 -3396 3960 -3364
rect 3920 -3444 3960 -3396
rect 3920 -3476 3924 -3444
rect 3956 -3476 3960 -3444
rect 3920 -3524 3960 -3476
rect 3920 -3556 3924 -3524
rect 3956 -3556 3960 -3524
rect 3920 -3604 3960 -3556
rect 3920 -3636 3924 -3604
rect 3956 -3636 3960 -3604
rect 3920 -3684 3960 -3636
rect 3920 -3716 3924 -3684
rect 3956 -3716 3960 -3684
rect 3920 -3720 3960 -3716
rect 4000 1036 4040 1040
rect 4000 1004 4004 1036
rect 4036 1004 4040 1036
rect 4000 956 4040 1004
rect 4000 924 4004 956
rect 4036 924 4040 956
rect 4000 876 4040 924
rect 4000 844 4004 876
rect 4036 844 4040 876
rect 4000 796 4040 844
rect 4000 764 4004 796
rect 4036 764 4040 796
rect 4000 716 4040 764
rect 4000 684 4004 716
rect 4036 684 4040 716
rect 4000 636 4040 684
rect 4000 604 4004 636
rect 4036 604 4040 636
rect 4000 556 4040 604
rect 4000 524 4004 556
rect 4036 524 4040 556
rect 4000 476 4040 524
rect 4000 444 4004 476
rect 4036 444 4040 476
rect 4000 396 4040 444
rect 4000 364 4004 396
rect 4036 364 4040 396
rect 4000 316 4040 364
rect 4000 284 4004 316
rect 4036 284 4040 316
rect 4000 236 4040 284
rect 4000 204 4004 236
rect 4036 204 4040 236
rect 4000 156 4040 204
rect 4000 124 4004 156
rect 4036 124 4040 156
rect 4000 76 4040 124
rect 4000 44 4004 76
rect 4036 44 4040 76
rect 4000 -4 4040 44
rect 4000 -36 4004 -4
rect 4036 -36 4040 -4
rect 4000 -84 4040 -36
rect 4000 -116 4004 -84
rect 4036 -116 4040 -84
rect 4000 -164 4040 -116
rect 4000 -196 4004 -164
rect 4036 -196 4040 -164
rect 4000 -244 4040 -196
rect 4000 -276 4004 -244
rect 4036 -276 4040 -244
rect 4000 -324 4040 -276
rect 4000 -356 4004 -324
rect 4036 -356 4040 -324
rect 4000 -404 4040 -356
rect 4000 -436 4004 -404
rect 4036 -436 4040 -404
rect 4000 -484 4040 -436
rect 4000 -516 4004 -484
rect 4036 -516 4040 -484
rect 4000 -564 4040 -516
rect 4000 -596 4004 -564
rect 4036 -596 4040 -564
rect 4000 -644 4040 -596
rect 4000 -676 4004 -644
rect 4036 -676 4040 -644
rect 4000 -724 4040 -676
rect 4000 -756 4004 -724
rect 4036 -756 4040 -724
rect 4000 -804 4040 -756
rect 4000 -836 4004 -804
rect 4036 -836 4040 -804
rect 4000 -884 4040 -836
rect 4000 -916 4004 -884
rect 4036 -916 4040 -884
rect 4000 -964 4040 -916
rect 4000 -996 4004 -964
rect 4036 -996 4040 -964
rect 4000 -1044 4040 -996
rect 4000 -1076 4004 -1044
rect 4036 -1076 4040 -1044
rect 4000 -1124 4040 -1076
rect 4000 -1156 4004 -1124
rect 4036 -1156 4040 -1124
rect 4000 -1204 4040 -1156
rect 4000 -1236 4004 -1204
rect 4036 -1236 4040 -1204
rect 4000 -1284 4040 -1236
rect 4000 -1316 4004 -1284
rect 4036 -1316 4040 -1284
rect 4000 -1364 4040 -1316
rect 4000 -1396 4004 -1364
rect 4036 -1396 4040 -1364
rect 4000 -1444 4040 -1396
rect 4000 -1476 4004 -1444
rect 4036 -1476 4040 -1444
rect 4000 -1524 4040 -1476
rect 4000 -1556 4004 -1524
rect 4036 -1556 4040 -1524
rect 4000 -1604 4040 -1556
rect 4000 -1636 4004 -1604
rect 4036 -1636 4040 -1604
rect 4000 -1684 4040 -1636
rect 4000 -1716 4004 -1684
rect 4036 -1716 4040 -1684
rect 4000 -1764 4040 -1716
rect 4000 -1796 4004 -1764
rect 4036 -1796 4040 -1764
rect 4000 -1844 4040 -1796
rect 4000 -1876 4004 -1844
rect 4036 -1876 4040 -1844
rect 4000 -1924 4040 -1876
rect 4000 -1956 4004 -1924
rect 4036 -1956 4040 -1924
rect 4000 -2004 4040 -1956
rect 4000 -2036 4004 -2004
rect 4036 -2036 4040 -2004
rect 4000 -2084 4040 -2036
rect 4000 -2116 4004 -2084
rect 4036 -2116 4040 -2084
rect 4000 -2164 4040 -2116
rect 4000 -2196 4004 -2164
rect 4036 -2196 4040 -2164
rect 4000 -2244 4040 -2196
rect 4000 -2276 4004 -2244
rect 4036 -2276 4040 -2244
rect 4000 -2324 4040 -2276
rect 4000 -2356 4004 -2324
rect 4036 -2356 4040 -2324
rect 4000 -2404 4040 -2356
rect 4000 -2436 4004 -2404
rect 4036 -2436 4040 -2404
rect 4000 -2484 4040 -2436
rect 4000 -2516 4004 -2484
rect 4036 -2516 4040 -2484
rect 4000 -2564 4040 -2516
rect 4000 -2596 4004 -2564
rect 4036 -2596 4040 -2564
rect 4000 -2644 4040 -2596
rect 4000 -2676 4004 -2644
rect 4036 -2676 4040 -2644
rect 4000 -2724 4040 -2676
rect 4000 -2756 4004 -2724
rect 4036 -2756 4040 -2724
rect 4000 -2804 4040 -2756
rect 4000 -2836 4004 -2804
rect 4036 -2836 4040 -2804
rect 4000 -2884 4040 -2836
rect 4000 -2916 4004 -2884
rect 4036 -2916 4040 -2884
rect 4000 -2964 4040 -2916
rect 4000 -2996 4004 -2964
rect 4036 -2996 4040 -2964
rect 4000 -3044 4040 -2996
rect 4000 -3076 4004 -3044
rect 4036 -3076 4040 -3044
rect 4000 -3124 4040 -3076
rect 4000 -3156 4004 -3124
rect 4036 -3156 4040 -3124
rect 4000 -3204 4040 -3156
rect 4000 -3236 4004 -3204
rect 4036 -3236 4040 -3204
rect 4000 -3284 4040 -3236
rect 4000 -3316 4004 -3284
rect 4036 -3316 4040 -3284
rect 4000 -3364 4040 -3316
rect 4000 -3396 4004 -3364
rect 4036 -3396 4040 -3364
rect 4000 -3444 4040 -3396
rect 4000 -3476 4004 -3444
rect 4036 -3476 4040 -3444
rect 4000 -3524 4040 -3476
rect 4000 -3556 4004 -3524
rect 4036 -3556 4040 -3524
rect 4000 -3604 4040 -3556
rect 4000 -3636 4004 -3604
rect 4036 -3636 4040 -3604
rect 4000 -3684 4040 -3636
rect 4000 -3716 4004 -3684
rect 4036 -3716 4040 -3684
rect 4000 -3720 4040 -3716
rect 4080 1036 4120 1040
rect 4080 1004 4084 1036
rect 4116 1004 4120 1036
rect 4080 956 4120 1004
rect 4080 924 4084 956
rect 4116 924 4120 956
rect 4080 876 4120 924
rect 4080 844 4084 876
rect 4116 844 4120 876
rect 4080 796 4120 844
rect 4080 764 4084 796
rect 4116 764 4120 796
rect 4080 716 4120 764
rect 4080 684 4084 716
rect 4116 684 4120 716
rect 4080 636 4120 684
rect 4080 604 4084 636
rect 4116 604 4120 636
rect 4080 556 4120 604
rect 4080 524 4084 556
rect 4116 524 4120 556
rect 4080 476 4120 524
rect 4080 444 4084 476
rect 4116 444 4120 476
rect 4080 396 4120 444
rect 4080 364 4084 396
rect 4116 364 4120 396
rect 4080 316 4120 364
rect 4080 284 4084 316
rect 4116 284 4120 316
rect 4080 236 4120 284
rect 4080 204 4084 236
rect 4116 204 4120 236
rect 4080 156 4120 204
rect 4080 124 4084 156
rect 4116 124 4120 156
rect 4080 76 4120 124
rect 4080 44 4084 76
rect 4116 44 4120 76
rect 4080 -4 4120 44
rect 4080 -36 4084 -4
rect 4116 -36 4120 -4
rect 4080 -84 4120 -36
rect 4080 -116 4084 -84
rect 4116 -116 4120 -84
rect 4080 -164 4120 -116
rect 4080 -196 4084 -164
rect 4116 -196 4120 -164
rect 4080 -244 4120 -196
rect 4080 -276 4084 -244
rect 4116 -276 4120 -244
rect 4080 -324 4120 -276
rect 4080 -356 4084 -324
rect 4116 -356 4120 -324
rect 4080 -404 4120 -356
rect 4080 -436 4084 -404
rect 4116 -436 4120 -404
rect 4080 -484 4120 -436
rect 4080 -516 4084 -484
rect 4116 -516 4120 -484
rect 4080 -564 4120 -516
rect 4080 -596 4084 -564
rect 4116 -596 4120 -564
rect 4080 -644 4120 -596
rect 4080 -676 4084 -644
rect 4116 -676 4120 -644
rect 4080 -724 4120 -676
rect 4080 -756 4084 -724
rect 4116 -756 4120 -724
rect 4080 -804 4120 -756
rect 4080 -836 4084 -804
rect 4116 -836 4120 -804
rect 4080 -884 4120 -836
rect 4080 -916 4084 -884
rect 4116 -916 4120 -884
rect 4080 -964 4120 -916
rect 4080 -996 4084 -964
rect 4116 -996 4120 -964
rect 4080 -1044 4120 -996
rect 4080 -1076 4084 -1044
rect 4116 -1076 4120 -1044
rect 4080 -1124 4120 -1076
rect 4080 -1156 4084 -1124
rect 4116 -1156 4120 -1124
rect 4080 -1204 4120 -1156
rect 4080 -1236 4084 -1204
rect 4116 -1236 4120 -1204
rect 4080 -1284 4120 -1236
rect 4080 -1316 4084 -1284
rect 4116 -1316 4120 -1284
rect 4080 -1364 4120 -1316
rect 4080 -1396 4084 -1364
rect 4116 -1396 4120 -1364
rect 4080 -1444 4120 -1396
rect 4080 -1476 4084 -1444
rect 4116 -1476 4120 -1444
rect 4080 -1524 4120 -1476
rect 4080 -1556 4084 -1524
rect 4116 -1556 4120 -1524
rect 4080 -1604 4120 -1556
rect 4080 -1636 4084 -1604
rect 4116 -1636 4120 -1604
rect 4080 -1684 4120 -1636
rect 4080 -1716 4084 -1684
rect 4116 -1716 4120 -1684
rect 4080 -1764 4120 -1716
rect 4080 -1796 4084 -1764
rect 4116 -1796 4120 -1764
rect 4080 -1844 4120 -1796
rect 4080 -1876 4084 -1844
rect 4116 -1876 4120 -1844
rect 4080 -1924 4120 -1876
rect 4080 -1956 4084 -1924
rect 4116 -1956 4120 -1924
rect 4080 -2004 4120 -1956
rect 4080 -2036 4084 -2004
rect 4116 -2036 4120 -2004
rect 4080 -2084 4120 -2036
rect 4080 -2116 4084 -2084
rect 4116 -2116 4120 -2084
rect 4080 -2164 4120 -2116
rect 4080 -2196 4084 -2164
rect 4116 -2196 4120 -2164
rect 4080 -2244 4120 -2196
rect 4080 -2276 4084 -2244
rect 4116 -2276 4120 -2244
rect 4080 -2324 4120 -2276
rect 4080 -2356 4084 -2324
rect 4116 -2356 4120 -2324
rect 4080 -2404 4120 -2356
rect 4080 -2436 4084 -2404
rect 4116 -2436 4120 -2404
rect 4080 -2484 4120 -2436
rect 4080 -2516 4084 -2484
rect 4116 -2516 4120 -2484
rect 4080 -2564 4120 -2516
rect 4080 -2596 4084 -2564
rect 4116 -2596 4120 -2564
rect 4080 -2644 4120 -2596
rect 4080 -2676 4084 -2644
rect 4116 -2676 4120 -2644
rect 4080 -2724 4120 -2676
rect 4080 -2756 4084 -2724
rect 4116 -2756 4120 -2724
rect 4080 -2804 4120 -2756
rect 4080 -2836 4084 -2804
rect 4116 -2836 4120 -2804
rect 4080 -2884 4120 -2836
rect 4080 -2916 4084 -2884
rect 4116 -2916 4120 -2884
rect 4080 -2964 4120 -2916
rect 4080 -2996 4084 -2964
rect 4116 -2996 4120 -2964
rect 4080 -3044 4120 -2996
rect 4080 -3076 4084 -3044
rect 4116 -3076 4120 -3044
rect 4080 -3124 4120 -3076
rect 4080 -3156 4084 -3124
rect 4116 -3156 4120 -3124
rect 4080 -3204 4120 -3156
rect 4080 -3236 4084 -3204
rect 4116 -3236 4120 -3204
rect 4080 -3284 4120 -3236
rect 4080 -3316 4084 -3284
rect 4116 -3316 4120 -3284
rect 4080 -3364 4120 -3316
rect 4080 -3396 4084 -3364
rect 4116 -3396 4120 -3364
rect 4080 -3444 4120 -3396
rect 4080 -3476 4084 -3444
rect 4116 -3476 4120 -3444
rect 4080 -3524 4120 -3476
rect 4080 -3556 4084 -3524
rect 4116 -3556 4120 -3524
rect 4080 -3604 4120 -3556
rect 4080 -3636 4084 -3604
rect 4116 -3636 4120 -3604
rect 4080 -3684 4120 -3636
rect 4080 -3716 4084 -3684
rect 4116 -3716 4120 -3684
rect 4080 -3720 4120 -3716
rect 4160 1036 4200 1040
rect 4160 1004 4164 1036
rect 4196 1004 4200 1036
rect 4160 956 4200 1004
rect 4160 924 4164 956
rect 4196 924 4200 956
rect 4160 876 4200 924
rect 4160 844 4164 876
rect 4196 844 4200 876
rect 4160 796 4200 844
rect 4160 764 4164 796
rect 4196 764 4200 796
rect 4160 716 4200 764
rect 4160 684 4164 716
rect 4196 684 4200 716
rect 4160 636 4200 684
rect 4160 604 4164 636
rect 4196 604 4200 636
rect 4160 556 4200 604
rect 4160 524 4164 556
rect 4196 524 4200 556
rect 4160 476 4200 524
rect 4160 444 4164 476
rect 4196 444 4200 476
rect 4160 396 4200 444
rect 4160 364 4164 396
rect 4196 364 4200 396
rect 4160 316 4200 364
rect 4160 284 4164 316
rect 4196 284 4200 316
rect 4160 236 4200 284
rect 4160 204 4164 236
rect 4196 204 4200 236
rect 4160 156 4200 204
rect 4160 124 4164 156
rect 4196 124 4200 156
rect 4160 76 4200 124
rect 4160 44 4164 76
rect 4196 44 4200 76
rect 4160 -4 4200 44
rect 4160 -36 4164 -4
rect 4196 -36 4200 -4
rect 4160 -84 4200 -36
rect 4160 -116 4164 -84
rect 4196 -116 4200 -84
rect 4160 -164 4200 -116
rect 4160 -196 4164 -164
rect 4196 -196 4200 -164
rect 4160 -244 4200 -196
rect 4160 -276 4164 -244
rect 4196 -276 4200 -244
rect 4160 -324 4200 -276
rect 4160 -356 4164 -324
rect 4196 -356 4200 -324
rect 4160 -404 4200 -356
rect 4160 -436 4164 -404
rect 4196 -436 4200 -404
rect 4160 -484 4200 -436
rect 4160 -516 4164 -484
rect 4196 -516 4200 -484
rect 4160 -564 4200 -516
rect 4160 -596 4164 -564
rect 4196 -596 4200 -564
rect 4160 -644 4200 -596
rect 4160 -676 4164 -644
rect 4196 -676 4200 -644
rect 4160 -724 4200 -676
rect 4160 -756 4164 -724
rect 4196 -756 4200 -724
rect 4160 -804 4200 -756
rect 4160 -836 4164 -804
rect 4196 -836 4200 -804
rect 4160 -884 4200 -836
rect 4160 -916 4164 -884
rect 4196 -916 4200 -884
rect 4160 -964 4200 -916
rect 4160 -996 4164 -964
rect 4196 -996 4200 -964
rect 4160 -1044 4200 -996
rect 4160 -1076 4164 -1044
rect 4196 -1076 4200 -1044
rect 4160 -1124 4200 -1076
rect 4160 -1156 4164 -1124
rect 4196 -1156 4200 -1124
rect 4160 -1204 4200 -1156
rect 4160 -1236 4164 -1204
rect 4196 -1236 4200 -1204
rect 4160 -1284 4200 -1236
rect 4160 -1316 4164 -1284
rect 4196 -1316 4200 -1284
rect 4160 -1364 4200 -1316
rect 4160 -1396 4164 -1364
rect 4196 -1396 4200 -1364
rect 4160 -1444 4200 -1396
rect 4160 -1476 4164 -1444
rect 4196 -1476 4200 -1444
rect 4160 -1524 4200 -1476
rect 4160 -1556 4164 -1524
rect 4196 -1556 4200 -1524
rect 4160 -1604 4200 -1556
rect 4160 -1636 4164 -1604
rect 4196 -1636 4200 -1604
rect 4160 -1684 4200 -1636
rect 4160 -1716 4164 -1684
rect 4196 -1716 4200 -1684
rect 4160 -1764 4200 -1716
rect 4160 -1796 4164 -1764
rect 4196 -1796 4200 -1764
rect 4160 -1844 4200 -1796
rect 4160 -1876 4164 -1844
rect 4196 -1876 4200 -1844
rect 4160 -1924 4200 -1876
rect 4160 -1956 4164 -1924
rect 4196 -1956 4200 -1924
rect 4160 -2004 4200 -1956
rect 4160 -2036 4164 -2004
rect 4196 -2036 4200 -2004
rect 4160 -2084 4200 -2036
rect 4160 -2116 4164 -2084
rect 4196 -2116 4200 -2084
rect 4160 -2164 4200 -2116
rect 4160 -2196 4164 -2164
rect 4196 -2196 4200 -2164
rect 4160 -2244 4200 -2196
rect 4160 -2276 4164 -2244
rect 4196 -2276 4200 -2244
rect 4160 -2324 4200 -2276
rect 4160 -2356 4164 -2324
rect 4196 -2356 4200 -2324
rect 4160 -2404 4200 -2356
rect 4160 -2436 4164 -2404
rect 4196 -2436 4200 -2404
rect 4160 -2484 4200 -2436
rect 4160 -2516 4164 -2484
rect 4196 -2516 4200 -2484
rect 4160 -2564 4200 -2516
rect 4160 -2596 4164 -2564
rect 4196 -2596 4200 -2564
rect 4160 -2644 4200 -2596
rect 4160 -2676 4164 -2644
rect 4196 -2676 4200 -2644
rect 4160 -2724 4200 -2676
rect 4160 -2756 4164 -2724
rect 4196 -2756 4200 -2724
rect 4160 -2804 4200 -2756
rect 4160 -2836 4164 -2804
rect 4196 -2836 4200 -2804
rect 4160 -2884 4200 -2836
rect 4160 -2916 4164 -2884
rect 4196 -2916 4200 -2884
rect 4160 -2964 4200 -2916
rect 4160 -2996 4164 -2964
rect 4196 -2996 4200 -2964
rect 4160 -3044 4200 -2996
rect 4160 -3076 4164 -3044
rect 4196 -3076 4200 -3044
rect 4160 -3124 4200 -3076
rect 4160 -3156 4164 -3124
rect 4196 -3156 4200 -3124
rect 4160 -3204 4200 -3156
rect 4160 -3236 4164 -3204
rect 4196 -3236 4200 -3204
rect 4160 -3284 4200 -3236
rect 4160 -3316 4164 -3284
rect 4196 -3316 4200 -3284
rect 4160 -3364 4200 -3316
rect 4160 -3396 4164 -3364
rect 4196 -3396 4200 -3364
rect 4160 -3444 4200 -3396
rect 4160 -3476 4164 -3444
rect 4196 -3476 4200 -3444
rect 4160 -3524 4200 -3476
rect 4160 -3556 4164 -3524
rect 4196 -3556 4200 -3524
rect 4160 -3604 4200 -3556
rect 4160 -3636 4164 -3604
rect 4196 -3636 4200 -3604
rect 4160 -3684 4200 -3636
rect 4160 -3716 4164 -3684
rect 4196 -3716 4200 -3684
rect 4160 -3720 4200 -3716
rect 4240 1036 4280 1040
rect 4240 1004 4244 1036
rect 4276 1004 4280 1036
rect 4240 956 4280 1004
rect 4240 924 4244 956
rect 4276 924 4280 956
rect 4240 876 4280 924
rect 4240 844 4244 876
rect 4276 844 4280 876
rect 4240 796 4280 844
rect 4240 764 4244 796
rect 4276 764 4280 796
rect 4240 716 4280 764
rect 4240 684 4244 716
rect 4276 684 4280 716
rect 4240 636 4280 684
rect 4240 604 4244 636
rect 4276 604 4280 636
rect 4240 556 4280 604
rect 4240 524 4244 556
rect 4276 524 4280 556
rect 4240 476 4280 524
rect 4240 444 4244 476
rect 4276 444 4280 476
rect 4240 396 4280 444
rect 4240 364 4244 396
rect 4276 364 4280 396
rect 4240 316 4280 364
rect 4240 284 4244 316
rect 4276 284 4280 316
rect 4240 236 4280 284
rect 4240 204 4244 236
rect 4276 204 4280 236
rect 4240 156 4280 204
rect 4240 124 4244 156
rect 4276 124 4280 156
rect 4240 76 4280 124
rect 4240 44 4244 76
rect 4276 44 4280 76
rect 4240 -4 4280 44
rect 4240 -36 4244 -4
rect 4276 -36 4280 -4
rect 4240 -84 4280 -36
rect 4240 -116 4244 -84
rect 4276 -116 4280 -84
rect 4240 -164 4280 -116
rect 4240 -196 4244 -164
rect 4276 -196 4280 -164
rect 4240 -244 4280 -196
rect 4240 -276 4244 -244
rect 4276 -276 4280 -244
rect 4240 -324 4280 -276
rect 4240 -356 4244 -324
rect 4276 -356 4280 -324
rect 4240 -404 4280 -356
rect 4240 -436 4244 -404
rect 4276 -436 4280 -404
rect 4240 -484 4280 -436
rect 4240 -516 4244 -484
rect 4276 -516 4280 -484
rect 4240 -564 4280 -516
rect 4240 -596 4244 -564
rect 4276 -596 4280 -564
rect 4240 -644 4280 -596
rect 4240 -676 4244 -644
rect 4276 -676 4280 -644
rect 4240 -724 4280 -676
rect 4240 -756 4244 -724
rect 4276 -756 4280 -724
rect 4240 -804 4280 -756
rect 4240 -836 4244 -804
rect 4276 -836 4280 -804
rect 4240 -884 4280 -836
rect 4240 -916 4244 -884
rect 4276 -916 4280 -884
rect 4240 -964 4280 -916
rect 4240 -996 4244 -964
rect 4276 -996 4280 -964
rect 4240 -1044 4280 -996
rect 4240 -1076 4244 -1044
rect 4276 -1076 4280 -1044
rect 4240 -1124 4280 -1076
rect 4240 -1156 4244 -1124
rect 4276 -1156 4280 -1124
rect 4240 -1204 4280 -1156
rect 4240 -1236 4244 -1204
rect 4276 -1236 4280 -1204
rect 4240 -1284 4280 -1236
rect 4240 -1316 4244 -1284
rect 4276 -1316 4280 -1284
rect 4240 -1364 4280 -1316
rect 4240 -1396 4244 -1364
rect 4276 -1396 4280 -1364
rect 4240 -1444 4280 -1396
rect 4240 -1476 4244 -1444
rect 4276 -1476 4280 -1444
rect 4240 -1524 4280 -1476
rect 4240 -1556 4244 -1524
rect 4276 -1556 4280 -1524
rect 4240 -1604 4280 -1556
rect 4240 -1636 4244 -1604
rect 4276 -1636 4280 -1604
rect 4240 -1684 4280 -1636
rect 4240 -1716 4244 -1684
rect 4276 -1716 4280 -1684
rect 4240 -1764 4280 -1716
rect 4240 -1796 4244 -1764
rect 4276 -1796 4280 -1764
rect 4240 -1844 4280 -1796
rect 4240 -1876 4244 -1844
rect 4276 -1876 4280 -1844
rect 4240 -1924 4280 -1876
rect 4240 -1956 4244 -1924
rect 4276 -1956 4280 -1924
rect 4240 -2004 4280 -1956
rect 4240 -2036 4244 -2004
rect 4276 -2036 4280 -2004
rect 4240 -2084 4280 -2036
rect 4240 -2116 4244 -2084
rect 4276 -2116 4280 -2084
rect 4240 -2164 4280 -2116
rect 4240 -2196 4244 -2164
rect 4276 -2196 4280 -2164
rect 4240 -2244 4280 -2196
rect 4240 -2276 4244 -2244
rect 4276 -2276 4280 -2244
rect 4240 -2324 4280 -2276
rect 4240 -2356 4244 -2324
rect 4276 -2356 4280 -2324
rect 4240 -2404 4280 -2356
rect 4240 -2436 4244 -2404
rect 4276 -2436 4280 -2404
rect 4240 -2484 4280 -2436
rect 4240 -2516 4244 -2484
rect 4276 -2516 4280 -2484
rect 4240 -2564 4280 -2516
rect 4240 -2596 4244 -2564
rect 4276 -2596 4280 -2564
rect 4240 -2644 4280 -2596
rect 4240 -2676 4244 -2644
rect 4276 -2676 4280 -2644
rect 4240 -2724 4280 -2676
rect 4240 -2756 4244 -2724
rect 4276 -2756 4280 -2724
rect 4240 -2804 4280 -2756
rect 4240 -2836 4244 -2804
rect 4276 -2836 4280 -2804
rect 4240 -2884 4280 -2836
rect 4240 -2916 4244 -2884
rect 4276 -2916 4280 -2884
rect 4240 -2964 4280 -2916
rect 4240 -2996 4244 -2964
rect 4276 -2996 4280 -2964
rect 4240 -3044 4280 -2996
rect 4240 -3076 4244 -3044
rect 4276 -3076 4280 -3044
rect 4240 -3124 4280 -3076
rect 4240 -3156 4244 -3124
rect 4276 -3156 4280 -3124
rect 4240 -3204 4280 -3156
rect 4240 -3236 4244 -3204
rect 4276 -3236 4280 -3204
rect 4240 -3284 4280 -3236
rect 4240 -3316 4244 -3284
rect 4276 -3316 4280 -3284
rect 4240 -3364 4280 -3316
rect 4240 -3396 4244 -3364
rect 4276 -3396 4280 -3364
rect 4240 -3444 4280 -3396
rect 4240 -3476 4244 -3444
rect 4276 -3476 4280 -3444
rect 4240 -3524 4280 -3476
rect 4240 -3556 4244 -3524
rect 4276 -3556 4280 -3524
rect 4240 -3604 4280 -3556
rect 4240 -3636 4244 -3604
rect 4276 -3636 4280 -3604
rect 4240 -3684 4280 -3636
rect 4240 -3716 4244 -3684
rect 4276 -3716 4280 -3684
rect 4240 -3720 4280 -3716
rect 4320 1036 4360 1040
rect 4320 1004 4324 1036
rect 4356 1004 4360 1036
rect 4320 956 4360 1004
rect 4320 924 4324 956
rect 4356 924 4360 956
rect 4320 876 4360 924
rect 4320 844 4324 876
rect 4356 844 4360 876
rect 4320 796 4360 844
rect 4320 764 4324 796
rect 4356 764 4360 796
rect 4320 716 4360 764
rect 4320 684 4324 716
rect 4356 684 4360 716
rect 4320 636 4360 684
rect 4320 604 4324 636
rect 4356 604 4360 636
rect 4320 556 4360 604
rect 4320 524 4324 556
rect 4356 524 4360 556
rect 4320 476 4360 524
rect 4320 444 4324 476
rect 4356 444 4360 476
rect 4320 396 4360 444
rect 4320 364 4324 396
rect 4356 364 4360 396
rect 4320 316 4360 364
rect 4320 284 4324 316
rect 4356 284 4360 316
rect 4320 236 4360 284
rect 4320 204 4324 236
rect 4356 204 4360 236
rect 4320 156 4360 204
rect 4320 124 4324 156
rect 4356 124 4360 156
rect 4320 76 4360 124
rect 4320 44 4324 76
rect 4356 44 4360 76
rect 4320 -4 4360 44
rect 4320 -36 4324 -4
rect 4356 -36 4360 -4
rect 4320 -84 4360 -36
rect 4320 -116 4324 -84
rect 4356 -116 4360 -84
rect 4320 -164 4360 -116
rect 4320 -196 4324 -164
rect 4356 -196 4360 -164
rect 4320 -244 4360 -196
rect 4320 -276 4324 -244
rect 4356 -276 4360 -244
rect 4320 -324 4360 -276
rect 4320 -356 4324 -324
rect 4356 -356 4360 -324
rect 4320 -404 4360 -356
rect 4320 -436 4324 -404
rect 4356 -436 4360 -404
rect 4320 -484 4360 -436
rect 4320 -516 4324 -484
rect 4356 -516 4360 -484
rect 4320 -564 4360 -516
rect 4320 -596 4324 -564
rect 4356 -596 4360 -564
rect 4320 -644 4360 -596
rect 4320 -676 4324 -644
rect 4356 -676 4360 -644
rect 4320 -724 4360 -676
rect 4320 -756 4324 -724
rect 4356 -756 4360 -724
rect 4320 -804 4360 -756
rect 4320 -836 4324 -804
rect 4356 -836 4360 -804
rect 4320 -884 4360 -836
rect 4320 -916 4324 -884
rect 4356 -916 4360 -884
rect 4320 -964 4360 -916
rect 4320 -996 4324 -964
rect 4356 -996 4360 -964
rect 4320 -1044 4360 -996
rect 4320 -1076 4324 -1044
rect 4356 -1076 4360 -1044
rect 4320 -1124 4360 -1076
rect 4320 -1156 4324 -1124
rect 4356 -1156 4360 -1124
rect 4320 -1204 4360 -1156
rect 4320 -1236 4324 -1204
rect 4356 -1236 4360 -1204
rect 4320 -1284 4360 -1236
rect 4320 -1316 4324 -1284
rect 4356 -1316 4360 -1284
rect 4320 -1364 4360 -1316
rect 4320 -1396 4324 -1364
rect 4356 -1396 4360 -1364
rect 4320 -1444 4360 -1396
rect 4320 -1476 4324 -1444
rect 4356 -1476 4360 -1444
rect 4320 -1524 4360 -1476
rect 4320 -1556 4324 -1524
rect 4356 -1556 4360 -1524
rect 4320 -1604 4360 -1556
rect 4320 -1636 4324 -1604
rect 4356 -1636 4360 -1604
rect 4320 -1684 4360 -1636
rect 4320 -1716 4324 -1684
rect 4356 -1716 4360 -1684
rect 4320 -1764 4360 -1716
rect 4320 -1796 4324 -1764
rect 4356 -1796 4360 -1764
rect 4320 -1844 4360 -1796
rect 4320 -1876 4324 -1844
rect 4356 -1876 4360 -1844
rect 4320 -1924 4360 -1876
rect 4320 -1956 4324 -1924
rect 4356 -1956 4360 -1924
rect 4320 -2004 4360 -1956
rect 4320 -2036 4324 -2004
rect 4356 -2036 4360 -2004
rect 4320 -2084 4360 -2036
rect 4320 -2116 4324 -2084
rect 4356 -2116 4360 -2084
rect 4320 -2164 4360 -2116
rect 4320 -2196 4324 -2164
rect 4356 -2196 4360 -2164
rect 4320 -2244 4360 -2196
rect 4320 -2276 4324 -2244
rect 4356 -2276 4360 -2244
rect 4320 -2324 4360 -2276
rect 4320 -2356 4324 -2324
rect 4356 -2356 4360 -2324
rect 4320 -2404 4360 -2356
rect 4320 -2436 4324 -2404
rect 4356 -2436 4360 -2404
rect 4320 -2484 4360 -2436
rect 4320 -2516 4324 -2484
rect 4356 -2516 4360 -2484
rect 4320 -2564 4360 -2516
rect 4320 -2596 4324 -2564
rect 4356 -2596 4360 -2564
rect 4320 -2644 4360 -2596
rect 4320 -2676 4324 -2644
rect 4356 -2676 4360 -2644
rect 4320 -2724 4360 -2676
rect 4320 -2756 4324 -2724
rect 4356 -2756 4360 -2724
rect 4320 -2804 4360 -2756
rect 4320 -2836 4324 -2804
rect 4356 -2836 4360 -2804
rect 4320 -2884 4360 -2836
rect 4320 -2916 4324 -2884
rect 4356 -2916 4360 -2884
rect 4320 -2964 4360 -2916
rect 4320 -2996 4324 -2964
rect 4356 -2996 4360 -2964
rect 4320 -3044 4360 -2996
rect 4320 -3076 4324 -3044
rect 4356 -3076 4360 -3044
rect 4320 -3124 4360 -3076
rect 4320 -3156 4324 -3124
rect 4356 -3156 4360 -3124
rect 4320 -3204 4360 -3156
rect 4320 -3236 4324 -3204
rect 4356 -3236 4360 -3204
rect 4320 -3284 4360 -3236
rect 4320 -3316 4324 -3284
rect 4356 -3316 4360 -3284
rect 4320 -3364 4360 -3316
rect 4320 -3396 4324 -3364
rect 4356 -3396 4360 -3364
rect 4320 -3444 4360 -3396
rect 4320 -3476 4324 -3444
rect 4356 -3476 4360 -3444
rect 4320 -3524 4360 -3476
rect 4320 -3556 4324 -3524
rect 4356 -3556 4360 -3524
rect 4320 -3604 4360 -3556
rect 4320 -3636 4324 -3604
rect 4356 -3636 4360 -3604
rect 4320 -3684 4360 -3636
rect 4320 -3716 4324 -3684
rect 4356 -3716 4360 -3684
rect 4320 -3720 4360 -3716
rect 4400 1036 4440 1040
rect 4400 1004 4404 1036
rect 4436 1004 4440 1036
rect 4400 956 4440 1004
rect 4400 924 4404 956
rect 4436 924 4440 956
rect 4400 876 4440 924
rect 4400 844 4404 876
rect 4436 844 4440 876
rect 4400 796 4440 844
rect 4400 764 4404 796
rect 4436 764 4440 796
rect 4400 716 4440 764
rect 4400 684 4404 716
rect 4436 684 4440 716
rect 4400 636 4440 684
rect 4400 604 4404 636
rect 4436 604 4440 636
rect 4400 556 4440 604
rect 4400 524 4404 556
rect 4436 524 4440 556
rect 4400 476 4440 524
rect 4400 444 4404 476
rect 4436 444 4440 476
rect 4400 396 4440 444
rect 4400 364 4404 396
rect 4436 364 4440 396
rect 4400 316 4440 364
rect 4400 284 4404 316
rect 4436 284 4440 316
rect 4400 236 4440 284
rect 4400 204 4404 236
rect 4436 204 4440 236
rect 4400 156 4440 204
rect 4400 124 4404 156
rect 4436 124 4440 156
rect 4400 76 4440 124
rect 4400 44 4404 76
rect 4436 44 4440 76
rect 4400 -4 4440 44
rect 4400 -36 4404 -4
rect 4436 -36 4440 -4
rect 4400 -84 4440 -36
rect 4400 -116 4404 -84
rect 4436 -116 4440 -84
rect 4400 -164 4440 -116
rect 4400 -196 4404 -164
rect 4436 -196 4440 -164
rect 4400 -244 4440 -196
rect 4400 -276 4404 -244
rect 4436 -276 4440 -244
rect 4400 -324 4440 -276
rect 4400 -356 4404 -324
rect 4436 -356 4440 -324
rect 4400 -404 4440 -356
rect 4400 -436 4404 -404
rect 4436 -436 4440 -404
rect 4400 -484 4440 -436
rect 4400 -516 4404 -484
rect 4436 -516 4440 -484
rect 4400 -564 4440 -516
rect 4400 -596 4404 -564
rect 4436 -596 4440 -564
rect 4400 -644 4440 -596
rect 4400 -676 4404 -644
rect 4436 -676 4440 -644
rect 4400 -724 4440 -676
rect 4400 -756 4404 -724
rect 4436 -756 4440 -724
rect 4400 -804 4440 -756
rect 4400 -836 4404 -804
rect 4436 -836 4440 -804
rect 4400 -884 4440 -836
rect 4400 -916 4404 -884
rect 4436 -916 4440 -884
rect 4400 -964 4440 -916
rect 4400 -996 4404 -964
rect 4436 -996 4440 -964
rect 4400 -1044 4440 -996
rect 4400 -1076 4404 -1044
rect 4436 -1076 4440 -1044
rect 4400 -1124 4440 -1076
rect 4400 -1156 4404 -1124
rect 4436 -1156 4440 -1124
rect 4400 -1204 4440 -1156
rect 4400 -1236 4404 -1204
rect 4436 -1236 4440 -1204
rect 4400 -1284 4440 -1236
rect 4400 -1316 4404 -1284
rect 4436 -1316 4440 -1284
rect 4400 -1364 4440 -1316
rect 4400 -1396 4404 -1364
rect 4436 -1396 4440 -1364
rect 4400 -1444 4440 -1396
rect 4400 -1476 4404 -1444
rect 4436 -1476 4440 -1444
rect 4400 -1524 4440 -1476
rect 4400 -1556 4404 -1524
rect 4436 -1556 4440 -1524
rect 4400 -1604 4440 -1556
rect 4400 -1636 4404 -1604
rect 4436 -1636 4440 -1604
rect 4400 -1684 4440 -1636
rect 4400 -1716 4404 -1684
rect 4436 -1716 4440 -1684
rect 4400 -1764 4440 -1716
rect 4400 -1796 4404 -1764
rect 4436 -1796 4440 -1764
rect 4400 -1844 4440 -1796
rect 4400 -1876 4404 -1844
rect 4436 -1876 4440 -1844
rect 4400 -1924 4440 -1876
rect 4400 -1956 4404 -1924
rect 4436 -1956 4440 -1924
rect 4400 -2004 4440 -1956
rect 4400 -2036 4404 -2004
rect 4436 -2036 4440 -2004
rect 4400 -2084 4440 -2036
rect 4400 -2116 4404 -2084
rect 4436 -2116 4440 -2084
rect 4400 -2164 4440 -2116
rect 4400 -2196 4404 -2164
rect 4436 -2196 4440 -2164
rect 4400 -2244 4440 -2196
rect 4400 -2276 4404 -2244
rect 4436 -2276 4440 -2244
rect 4400 -2324 4440 -2276
rect 4400 -2356 4404 -2324
rect 4436 -2356 4440 -2324
rect 4400 -2404 4440 -2356
rect 4400 -2436 4404 -2404
rect 4436 -2436 4440 -2404
rect 4400 -2484 4440 -2436
rect 4400 -2516 4404 -2484
rect 4436 -2516 4440 -2484
rect 4400 -2564 4440 -2516
rect 4400 -2596 4404 -2564
rect 4436 -2596 4440 -2564
rect 4400 -2644 4440 -2596
rect 4400 -2676 4404 -2644
rect 4436 -2676 4440 -2644
rect 4400 -2724 4440 -2676
rect 4400 -2756 4404 -2724
rect 4436 -2756 4440 -2724
rect 4400 -2804 4440 -2756
rect 4400 -2836 4404 -2804
rect 4436 -2836 4440 -2804
rect 4400 -2884 4440 -2836
rect 4400 -2916 4404 -2884
rect 4436 -2916 4440 -2884
rect 4400 -2964 4440 -2916
rect 4400 -2996 4404 -2964
rect 4436 -2996 4440 -2964
rect 4400 -3044 4440 -2996
rect 4400 -3076 4404 -3044
rect 4436 -3076 4440 -3044
rect 4400 -3124 4440 -3076
rect 4400 -3156 4404 -3124
rect 4436 -3156 4440 -3124
rect 4400 -3204 4440 -3156
rect 4400 -3236 4404 -3204
rect 4436 -3236 4440 -3204
rect 4400 -3284 4440 -3236
rect 4400 -3316 4404 -3284
rect 4436 -3316 4440 -3284
rect 4400 -3364 4440 -3316
rect 4400 -3396 4404 -3364
rect 4436 -3396 4440 -3364
rect 4400 -3444 4440 -3396
rect 4400 -3476 4404 -3444
rect 4436 -3476 4440 -3444
rect 4400 -3524 4440 -3476
rect 4400 -3556 4404 -3524
rect 4436 -3556 4440 -3524
rect 4400 -3604 4440 -3556
rect 4400 -3636 4404 -3604
rect 4436 -3636 4440 -3604
rect 4400 -3684 4440 -3636
rect 4400 -3716 4404 -3684
rect 4436 -3716 4440 -3684
rect 4400 -3720 4440 -3716
rect 4480 1036 4520 1040
rect 4480 1004 4484 1036
rect 4516 1004 4520 1036
rect 4480 956 4520 1004
rect 4480 924 4484 956
rect 4516 924 4520 956
rect 4480 876 4520 924
rect 4480 844 4484 876
rect 4516 844 4520 876
rect 4480 796 4520 844
rect 4480 764 4484 796
rect 4516 764 4520 796
rect 4480 716 4520 764
rect 4480 684 4484 716
rect 4516 684 4520 716
rect 4480 636 4520 684
rect 4480 604 4484 636
rect 4516 604 4520 636
rect 4480 556 4520 604
rect 4480 524 4484 556
rect 4516 524 4520 556
rect 4480 476 4520 524
rect 4480 444 4484 476
rect 4516 444 4520 476
rect 4480 396 4520 444
rect 4480 364 4484 396
rect 4516 364 4520 396
rect 4480 316 4520 364
rect 4480 284 4484 316
rect 4516 284 4520 316
rect 4480 236 4520 284
rect 4480 204 4484 236
rect 4516 204 4520 236
rect 4480 156 4520 204
rect 4480 124 4484 156
rect 4516 124 4520 156
rect 4480 76 4520 124
rect 4480 44 4484 76
rect 4516 44 4520 76
rect 4480 -4 4520 44
rect 4480 -36 4484 -4
rect 4516 -36 4520 -4
rect 4480 -84 4520 -36
rect 4480 -116 4484 -84
rect 4516 -116 4520 -84
rect 4480 -164 4520 -116
rect 4480 -196 4484 -164
rect 4516 -196 4520 -164
rect 4480 -244 4520 -196
rect 4480 -276 4484 -244
rect 4516 -276 4520 -244
rect 4480 -324 4520 -276
rect 4480 -356 4484 -324
rect 4516 -356 4520 -324
rect 4480 -404 4520 -356
rect 4480 -436 4484 -404
rect 4516 -436 4520 -404
rect 4480 -484 4520 -436
rect 4480 -516 4484 -484
rect 4516 -516 4520 -484
rect 4480 -564 4520 -516
rect 4480 -596 4484 -564
rect 4516 -596 4520 -564
rect 4480 -644 4520 -596
rect 4480 -676 4484 -644
rect 4516 -676 4520 -644
rect 4480 -724 4520 -676
rect 4480 -756 4484 -724
rect 4516 -756 4520 -724
rect 4480 -804 4520 -756
rect 4480 -836 4484 -804
rect 4516 -836 4520 -804
rect 4480 -884 4520 -836
rect 4480 -916 4484 -884
rect 4516 -916 4520 -884
rect 4480 -964 4520 -916
rect 4480 -996 4484 -964
rect 4516 -996 4520 -964
rect 4480 -1044 4520 -996
rect 4480 -1076 4484 -1044
rect 4516 -1076 4520 -1044
rect 4480 -1124 4520 -1076
rect 4480 -1156 4484 -1124
rect 4516 -1156 4520 -1124
rect 4480 -1204 4520 -1156
rect 4480 -1236 4484 -1204
rect 4516 -1236 4520 -1204
rect 4480 -1284 4520 -1236
rect 4480 -1316 4484 -1284
rect 4516 -1316 4520 -1284
rect 4480 -1364 4520 -1316
rect 4480 -1396 4484 -1364
rect 4516 -1396 4520 -1364
rect 4480 -1444 4520 -1396
rect 4480 -1476 4484 -1444
rect 4516 -1476 4520 -1444
rect 4480 -1524 4520 -1476
rect 4480 -1556 4484 -1524
rect 4516 -1556 4520 -1524
rect 4480 -1604 4520 -1556
rect 4480 -1636 4484 -1604
rect 4516 -1636 4520 -1604
rect 4480 -1684 4520 -1636
rect 4480 -1716 4484 -1684
rect 4516 -1716 4520 -1684
rect 4480 -1764 4520 -1716
rect 4480 -1796 4484 -1764
rect 4516 -1796 4520 -1764
rect 4480 -1844 4520 -1796
rect 4480 -1876 4484 -1844
rect 4516 -1876 4520 -1844
rect 4480 -1924 4520 -1876
rect 4480 -1956 4484 -1924
rect 4516 -1956 4520 -1924
rect 4480 -2004 4520 -1956
rect 4480 -2036 4484 -2004
rect 4516 -2036 4520 -2004
rect 4480 -2084 4520 -2036
rect 4480 -2116 4484 -2084
rect 4516 -2116 4520 -2084
rect 4480 -2164 4520 -2116
rect 4480 -2196 4484 -2164
rect 4516 -2196 4520 -2164
rect 4480 -2244 4520 -2196
rect 4480 -2276 4484 -2244
rect 4516 -2276 4520 -2244
rect 4480 -2324 4520 -2276
rect 4480 -2356 4484 -2324
rect 4516 -2356 4520 -2324
rect 4480 -2404 4520 -2356
rect 4480 -2436 4484 -2404
rect 4516 -2436 4520 -2404
rect 4480 -2484 4520 -2436
rect 4480 -2516 4484 -2484
rect 4516 -2516 4520 -2484
rect 4480 -2564 4520 -2516
rect 4480 -2596 4484 -2564
rect 4516 -2596 4520 -2564
rect 4480 -2644 4520 -2596
rect 4480 -2676 4484 -2644
rect 4516 -2676 4520 -2644
rect 4480 -2724 4520 -2676
rect 4480 -2756 4484 -2724
rect 4516 -2756 4520 -2724
rect 4480 -2804 4520 -2756
rect 4480 -2836 4484 -2804
rect 4516 -2836 4520 -2804
rect 4480 -2884 4520 -2836
rect 4480 -2916 4484 -2884
rect 4516 -2916 4520 -2884
rect 4480 -2964 4520 -2916
rect 4480 -2996 4484 -2964
rect 4516 -2996 4520 -2964
rect 4480 -3044 4520 -2996
rect 4480 -3076 4484 -3044
rect 4516 -3076 4520 -3044
rect 4480 -3124 4520 -3076
rect 4480 -3156 4484 -3124
rect 4516 -3156 4520 -3124
rect 4480 -3204 4520 -3156
rect 4480 -3236 4484 -3204
rect 4516 -3236 4520 -3204
rect 4480 -3284 4520 -3236
rect 4480 -3316 4484 -3284
rect 4516 -3316 4520 -3284
rect 4480 -3364 4520 -3316
rect 4480 -3396 4484 -3364
rect 4516 -3396 4520 -3364
rect 4480 -3444 4520 -3396
rect 4480 -3476 4484 -3444
rect 4516 -3476 4520 -3444
rect 4480 -3524 4520 -3476
rect 4480 -3556 4484 -3524
rect 4516 -3556 4520 -3524
rect 4480 -3604 4520 -3556
rect 4480 -3636 4484 -3604
rect 4516 -3636 4520 -3604
rect 4480 -3684 4520 -3636
rect 4480 -3716 4484 -3684
rect 4516 -3716 4520 -3684
rect 4480 -3720 4520 -3716
rect 4560 1036 4600 1040
rect 4560 1004 4564 1036
rect 4596 1004 4600 1036
rect 4560 956 4600 1004
rect 4560 924 4564 956
rect 4596 924 4600 956
rect 4560 876 4600 924
rect 4560 844 4564 876
rect 4596 844 4600 876
rect 4560 796 4600 844
rect 4560 764 4564 796
rect 4596 764 4600 796
rect 4560 716 4600 764
rect 4560 684 4564 716
rect 4596 684 4600 716
rect 4560 636 4600 684
rect 4560 604 4564 636
rect 4596 604 4600 636
rect 4560 556 4600 604
rect 4560 524 4564 556
rect 4596 524 4600 556
rect 4560 476 4600 524
rect 4560 444 4564 476
rect 4596 444 4600 476
rect 4560 396 4600 444
rect 4560 364 4564 396
rect 4596 364 4600 396
rect 4560 316 4600 364
rect 4560 284 4564 316
rect 4596 284 4600 316
rect 4560 236 4600 284
rect 4560 204 4564 236
rect 4596 204 4600 236
rect 4560 156 4600 204
rect 4560 124 4564 156
rect 4596 124 4600 156
rect 4560 76 4600 124
rect 4560 44 4564 76
rect 4596 44 4600 76
rect 4560 -4 4600 44
rect 4560 -36 4564 -4
rect 4596 -36 4600 -4
rect 4560 -84 4600 -36
rect 4560 -116 4564 -84
rect 4596 -116 4600 -84
rect 4560 -164 4600 -116
rect 4560 -196 4564 -164
rect 4596 -196 4600 -164
rect 4560 -244 4600 -196
rect 4560 -276 4564 -244
rect 4596 -276 4600 -244
rect 4560 -324 4600 -276
rect 4560 -356 4564 -324
rect 4596 -356 4600 -324
rect 4560 -404 4600 -356
rect 4560 -436 4564 -404
rect 4596 -436 4600 -404
rect 4560 -484 4600 -436
rect 4560 -516 4564 -484
rect 4596 -516 4600 -484
rect 4560 -564 4600 -516
rect 4560 -596 4564 -564
rect 4596 -596 4600 -564
rect 4560 -644 4600 -596
rect 4560 -676 4564 -644
rect 4596 -676 4600 -644
rect 4560 -724 4600 -676
rect 4560 -756 4564 -724
rect 4596 -756 4600 -724
rect 4560 -804 4600 -756
rect 4560 -836 4564 -804
rect 4596 -836 4600 -804
rect 4560 -884 4600 -836
rect 4560 -916 4564 -884
rect 4596 -916 4600 -884
rect 4560 -964 4600 -916
rect 4560 -996 4564 -964
rect 4596 -996 4600 -964
rect 4560 -1044 4600 -996
rect 4560 -1076 4564 -1044
rect 4596 -1076 4600 -1044
rect 4560 -1124 4600 -1076
rect 4560 -1156 4564 -1124
rect 4596 -1156 4600 -1124
rect 4560 -1204 4600 -1156
rect 4560 -1236 4564 -1204
rect 4596 -1236 4600 -1204
rect 4560 -1284 4600 -1236
rect 4560 -1316 4564 -1284
rect 4596 -1316 4600 -1284
rect 4560 -1364 4600 -1316
rect 4560 -1396 4564 -1364
rect 4596 -1396 4600 -1364
rect 4560 -1444 4600 -1396
rect 4560 -1476 4564 -1444
rect 4596 -1476 4600 -1444
rect 4560 -1524 4600 -1476
rect 4560 -1556 4564 -1524
rect 4596 -1556 4600 -1524
rect 4560 -1604 4600 -1556
rect 4560 -1636 4564 -1604
rect 4596 -1636 4600 -1604
rect 4560 -1684 4600 -1636
rect 4560 -1716 4564 -1684
rect 4596 -1716 4600 -1684
rect 4560 -1764 4600 -1716
rect 4560 -1796 4564 -1764
rect 4596 -1796 4600 -1764
rect 4560 -1844 4600 -1796
rect 4560 -1876 4564 -1844
rect 4596 -1876 4600 -1844
rect 4560 -1924 4600 -1876
rect 4560 -1956 4564 -1924
rect 4596 -1956 4600 -1924
rect 4560 -2004 4600 -1956
rect 4560 -2036 4564 -2004
rect 4596 -2036 4600 -2004
rect 4560 -2084 4600 -2036
rect 4560 -2116 4564 -2084
rect 4596 -2116 4600 -2084
rect 4560 -2164 4600 -2116
rect 4560 -2196 4564 -2164
rect 4596 -2196 4600 -2164
rect 4560 -2244 4600 -2196
rect 4560 -2276 4564 -2244
rect 4596 -2276 4600 -2244
rect 4560 -2324 4600 -2276
rect 4560 -2356 4564 -2324
rect 4596 -2356 4600 -2324
rect 4560 -2404 4600 -2356
rect 4560 -2436 4564 -2404
rect 4596 -2436 4600 -2404
rect 4560 -2484 4600 -2436
rect 4560 -2516 4564 -2484
rect 4596 -2516 4600 -2484
rect 4560 -2564 4600 -2516
rect 4560 -2596 4564 -2564
rect 4596 -2596 4600 -2564
rect 4560 -2644 4600 -2596
rect 4560 -2676 4564 -2644
rect 4596 -2676 4600 -2644
rect 4560 -2724 4600 -2676
rect 4560 -2756 4564 -2724
rect 4596 -2756 4600 -2724
rect 4560 -2804 4600 -2756
rect 4560 -2836 4564 -2804
rect 4596 -2836 4600 -2804
rect 4560 -2884 4600 -2836
rect 4560 -2916 4564 -2884
rect 4596 -2916 4600 -2884
rect 4560 -2964 4600 -2916
rect 4560 -2996 4564 -2964
rect 4596 -2996 4600 -2964
rect 4560 -3044 4600 -2996
rect 4560 -3076 4564 -3044
rect 4596 -3076 4600 -3044
rect 4560 -3124 4600 -3076
rect 4560 -3156 4564 -3124
rect 4596 -3156 4600 -3124
rect 4560 -3204 4600 -3156
rect 4560 -3236 4564 -3204
rect 4596 -3236 4600 -3204
rect 4560 -3284 4600 -3236
rect 4560 -3316 4564 -3284
rect 4596 -3316 4600 -3284
rect 4560 -3364 4600 -3316
rect 4560 -3396 4564 -3364
rect 4596 -3396 4600 -3364
rect 4560 -3444 4600 -3396
rect 4560 -3476 4564 -3444
rect 4596 -3476 4600 -3444
rect 4560 -3524 4600 -3476
rect 4560 -3556 4564 -3524
rect 4596 -3556 4600 -3524
rect 4560 -3604 4600 -3556
rect 4560 -3636 4564 -3604
rect 4596 -3636 4600 -3604
rect 4560 -3684 4600 -3636
rect 4560 -3716 4564 -3684
rect 4596 -3716 4600 -3684
rect 4560 -3720 4600 -3716
rect 4640 1036 4680 1040
rect 4640 1004 4644 1036
rect 4676 1004 4680 1036
rect 4640 956 4680 1004
rect 4640 924 4644 956
rect 4676 924 4680 956
rect 4640 876 4680 924
rect 4640 844 4644 876
rect 4676 844 4680 876
rect 4640 796 4680 844
rect 4640 764 4644 796
rect 4676 764 4680 796
rect 4640 716 4680 764
rect 4640 684 4644 716
rect 4676 684 4680 716
rect 4640 636 4680 684
rect 4640 604 4644 636
rect 4676 604 4680 636
rect 4640 556 4680 604
rect 4640 524 4644 556
rect 4676 524 4680 556
rect 4640 476 4680 524
rect 4640 444 4644 476
rect 4676 444 4680 476
rect 4640 396 4680 444
rect 4640 364 4644 396
rect 4676 364 4680 396
rect 4640 316 4680 364
rect 4640 284 4644 316
rect 4676 284 4680 316
rect 4640 236 4680 284
rect 4640 204 4644 236
rect 4676 204 4680 236
rect 4640 156 4680 204
rect 4640 124 4644 156
rect 4676 124 4680 156
rect 4640 76 4680 124
rect 4640 44 4644 76
rect 4676 44 4680 76
rect 4640 -4 4680 44
rect 4640 -36 4644 -4
rect 4676 -36 4680 -4
rect 4640 -84 4680 -36
rect 4640 -116 4644 -84
rect 4676 -116 4680 -84
rect 4640 -164 4680 -116
rect 4640 -196 4644 -164
rect 4676 -196 4680 -164
rect 4640 -244 4680 -196
rect 4640 -276 4644 -244
rect 4676 -276 4680 -244
rect 4640 -324 4680 -276
rect 4640 -356 4644 -324
rect 4676 -356 4680 -324
rect 4640 -404 4680 -356
rect 4640 -436 4644 -404
rect 4676 -436 4680 -404
rect 4640 -484 4680 -436
rect 4640 -516 4644 -484
rect 4676 -516 4680 -484
rect 4640 -564 4680 -516
rect 4640 -596 4644 -564
rect 4676 -596 4680 -564
rect 4640 -644 4680 -596
rect 4640 -676 4644 -644
rect 4676 -676 4680 -644
rect 4640 -724 4680 -676
rect 4640 -756 4644 -724
rect 4676 -756 4680 -724
rect 4640 -804 4680 -756
rect 4640 -836 4644 -804
rect 4676 -836 4680 -804
rect 4640 -884 4680 -836
rect 4640 -916 4644 -884
rect 4676 -916 4680 -884
rect 4640 -964 4680 -916
rect 4640 -996 4644 -964
rect 4676 -996 4680 -964
rect 4640 -1044 4680 -996
rect 4640 -1076 4644 -1044
rect 4676 -1076 4680 -1044
rect 4640 -1124 4680 -1076
rect 4640 -1156 4644 -1124
rect 4676 -1156 4680 -1124
rect 4640 -1204 4680 -1156
rect 4640 -1236 4644 -1204
rect 4676 -1236 4680 -1204
rect 4640 -1284 4680 -1236
rect 4640 -1316 4644 -1284
rect 4676 -1316 4680 -1284
rect 4640 -1364 4680 -1316
rect 4640 -1396 4644 -1364
rect 4676 -1396 4680 -1364
rect 4640 -1444 4680 -1396
rect 4640 -1476 4644 -1444
rect 4676 -1476 4680 -1444
rect 4640 -1524 4680 -1476
rect 4640 -1556 4644 -1524
rect 4676 -1556 4680 -1524
rect 4640 -1604 4680 -1556
rect 4640 -1636 4644 -1604
rect 4676 -1636 4680 -1604
rect 4640 -1684 4680 -1636
rect 4640 -1716 4644 -1684
rect 4676 -1716 4680 -1684
rect 4640 -1764 4680 -1716
rect 4640 -1796 4644 -1764
rect 4676 -1796 4680 -1764
rect 4640 -1844 4680 -1796
rect 4640 -1876 4644 -1844
rect 4676 -1876 4680 -1844
rect 4640 -1924 4680 -1876
rect 4640 -1956 4644 -1924
rect 4676 -1956 4680 -1924
rect 4640 -2004 4680 -1956
rect 4640 -2036 4644 -2004
rect 4676 -2036 4680 -2004
rect 4640 -2084 4680 -2036
rect 4640 -2116 4644 -2084
rect 4676 -2116 4680 -2084
rect 4640 -2164 4680 -2116
rect 4640 -2196 4644 -2164
rect 4676 -2196 4680 -2164
rect 4640 -2244 4680 -2196
rect 4640 -2276 4644 -2244
rect 4676 -2276 4680 -2244
rect 4640 -2324 4680 -2276
rect 4640 -2356 4644 -2324
rect 4676 -2356 4680 -2324
rect 4640 -2404 4680 -2356
rect 4640 -2436 4644 -2404
rect 4676 -2436 4680 -2404
rect 4640 -2484 4680 -2436
rect 4640 -2516 4644 -2484
rect 4676 -2516 4680 -2484
rect 4640 -2564 4680 -2516
rect 4640 -2596 4644 -2564
rect 4676 -2596 4680 -2564
rect 4640 -2644 4680 -2596
rect 4640 -2676 4644 -2644
rect 4676 -2676 4680 -2644
rect 4640 -2724 4680 -2676
rect 4640 -2756 4644 -2724
rect 4676 -2756 4680 -2724
rect 4640 -2804 4680 -2756
rect 4640 -2836 4644 -2804
rect 4676 -2836 4680 -2804
rect 4640 -2884 4680 -2836
rect 4640 -2916 4644 -2884
rect 4676 -2916 4680 -2884
rect 4640 -2964 4680 -2916
rect 4640 -2996 4644 -2964
rect 4676 -2996 4680 -2964
rect 4640 -3044 4680 -2996
rect 4640 -3076 4644 -3044
rect 4676 -3076 4680 -3044
rect 4640 -3124 4680 -3076
rect 4640 -3156 4644 -3124
rect 4676 -3156 4680 -3124
rect 4640 -3204 4680 -3156
rect 4640 -3236 4644 -3204
rect 4676 -3236 4680 -3204
rect 4640 -3284 4680 -3236
rect 4640 -3316 4644 -3284
rect 4676 -3316 4680 -3284
rect 4640 -3364 4680 -3316
rect 4640 -3396 4644 -3364
rect 4676 -3396 4680 -3364
rect 4640 -3444 4680 -3396
rect 4640 -3476 4644 -3444
rect 4676 -3476 4680 -3444
rect 4640 -3524 4680 -3476
rect 4640 -3556 4644 -3524
rect 4676 -3556 4680 -3524
rect 4640 -3604 4680 -3556
rect 4640 -3636 4644 -3604
rect 4676 -3636 4680 -3604
rect 4640 -3684 4680 -3636
rect 4640 -3716 4644 -3684
rect 4676 -3716 4680 -3684
rect 4640 -3720 4680 -3716
rect 4720 1036 4760 1040
rect 4720 1004 4724 1036
rect 4756 1004 4760 1036
rect 4720 956 4760 1004
rect 4720 924 4724 956
rect 4756 924 4760 956
rect 4720 876 4760 924
rect 4720 844 4724 876
rect 4756 844 4760 876
rect 4720 796 4760 844
rect 4720 764 4724 796
rect 4756 764 4760 796
rect 4720 716 4760 764
rect 4720 684 4724 716
rect 4756 684 4760 716
rect 4720 636 4760 684
rect 4720 604 4724 636
rect 4756 604 4760 636
rect 4720 556 4760 604
rect 4720 524 4724 556
rect 4756 524 4760 556
rect 4720 476 4760 524
rect 4720 444 4724 476
rect 4756 444 4760 476
rect 4720 396 4760 444
rect 4720 364 4724 396
rect 4756 364 4760 396
rect 4720 316 4760 364
rect 4720 284 4724 316
rect 4756 284 4760 316
rect 4720 236 4760 284
rect 4720 204 4724 236
rect 4756 204 4760 236
rect 4720 156 4760 204
rect 4720 124 4724 156
rect 4756 124 4760 156
rect 4720 76 4760 124
rect 4720 44 4724 76
rect 4756 44 4760 76
rect 4720 -4 4760 44
rect 4720 -36 4724 -4
rect 4756 -36 4760 -4
rect 4720 -84 4760 -36
rect 4720 -116 4724 -84
rect 4756 -116 4760 -84
rect 4720 -164 4760 -116
rect 4720 -196 4724 -164
rect 4756 -196 4760 -164
rect 4720 -244 4760 -196
rect 4720 -276 4724 -244
rect 4756 -276 4760 -244
rect 4720 -324 4760 -276
rect 4720 -356 4724 -324
rect 4756 -356 4760 -324
rect 4720 -404 4760 -356
rect 4720 -436 4724 -404
rect 4756 -436 4760 -404
rect 4720 -484 4760 -436
rect 4720 -516 4724 -484
rect 4756 -516 4760 -484
rect 4720 -564 4760 -516
rect 4720 -596 4724 -564
rect 4756 -596 4760 -564
rect 4720 -644 4760 -596
rect 4720 -676 4724 -644
rect 4756 -676 4760 -644
rect 4720 -724 4760 -676
rect 4720 -756 4724 -724
rect 4756 -756 4760 -724
rect 4720 -804 4760 -756
rect 4720 -836 4724 -804
rect 4756 -836 4760 -804
rect 4720 -884 4760 -836
rect 4720 -916 4724 -884
rect 4756 -916 4760 -884
rect 4720 -964 4760 -916
rect 4720 -996 4724 -964
rect 4756 -996 4760 -964
rect 4720 -1044 4760 -996
rect 4720 -1076 4724 -1044
rect 4756 -1076 4760 -1044
rect 4720 -1124 4760 -1076
rect 4720 -1156 4724 -1124
rect 4756 -1156 4760 -1124
rect 4720 -1204 4760 -1156
rect 4720 -1236 4724 -1204
rect 4756 -1236 4760 -1204
rect 4720 -1284 4760 -1236
rect 4720 -1316 4724 -1284
rect 4756 -1316 4760 -1284
rect 4720 -1364 4760 -1316
rect 4720 -1396 4724 -1364
rect 4756 -1396 4760 -1364
rect 4720 -1444 4760 -1396
rect 4720 -1476 4724 -1444
rect 4756 -1476 4760 -1444
rect 4720 -1524 4760 -1476
rect 4720 -1556 4724 -1524
rect 4756 -1556 4760 -1524
rect 4720 -1604 4760 -1556
rect 4720 -1636 4724 -1604
rect 4756 -1636 4760 -1604
rect 4720 -1684 4760 -1636
rect 4720 -1716 4724 -1684
rect 4756 -1716 4760 -1684
rect 4720 -1764 4760 -1716
rect 4720 -1796 4724 -1764
rect 4756 -1796 4760 -1764
rect 4720 -1844 4760 -1796
rect 4720 -1876 4724 -1844
rect 4756 -1876 4760 -1844
rect 4720 -1924 4760 -1876
rect 4720 -1956 4724 -1924
rect 4756 -1956 4760 -1924
rect 4720 -2004 4760 -1956
rect 4720 -2036 4724 -2004
rect 4756 -2036 4760 -2004
rect 4720 -2084 4760 -2036
rect 4720 -2116 4724 -2084
rect 4756 -2116 4760 -2084
rect 4720 -2164 4760 -2116
rect 4720 -2196 4724 -2164
rect 4756 -2196 4760 -2164
rect 4720 -2244 4760 -2196
rect 4720 -2276 4724 -2244
rect 4756 -2276 4760 -2244
rect 4720 -2324 4760 -2276
rect 4720 -2356 4724 -2324
rect 4756 -2356 4760 -2324
rect 4720 -2404 4760 -2356
rect 4720 -2436 4724 -2404
rect 4756 -2436 4760 -2404
rect 4720 -2484 4760 -2436
rect 4720 -2516 4724 -2484
rect 4756 -2516 4760 -2484
rect 4720 -2564 4760 -2516
rect 4720 -2596 4724 -2564
rect 4756 -2596 4760 -2564
rect 4720 -2644 4760 -2596
rect 4720 -2676 4724 -2644
rect 4756 -2676 4760 -2644
rect 4720 -2724 4760 -2676
rect 4720 -2756 4724 -2724
rect 4756 -2756 4760 -2724
rect 4720 -2804 4760 -2756
rect 4720 -2836 4724 -2804
rect 4756 -2836 4760 -2804
rect 4720 -2884 4760 -2836
rect 4720 -2916 4724 -2884
rect 4756 -2916 4760 -2884
rect 4720 -2964 4760 -2916
rect 4720 -2996 4724 -2964
rect 4756 -2996 4760 -2964
rect 4720 -3044 4760 -2996
rect 4720 -3076 4724 -3044
rect 4756 -3076 4760 -3044
rect 4720 -3124 4760 -3076
rect 4720 -3156 4724 -3124
rect 4756 -3156 4760 -3124
rect 4720 -3204 4760 -3156
rect 4720 -3236 4724 -3204
rect 4756 -3236 4760 -3204
rect 4720 -3284 4760 -3236
rect 4720 -3316 4724 -3284
rect 4756 -3316 4760 -3284
rect 4720 -3364 4760 -3316
rect 4720 -3396 4724 -3364
rect 4756 -3396 4760 -3364
rect 4720 -3444 4760 -3396
rect 4720 -3476 4724 -3444
rect 4756 -3476 4760 -3444
rect 4720 -3524 4760 -3476
rect 4720 -3556 4724 -3524
rect 4756 -3556 4760 -3524
rect 4720 -3604 4760 -3556
rect 4720 -3636 4724 -3604
rect 4756 -3636 4760 -3604
rect 4720 -3684 4760 -3636
rect 4720 -3716 4724 -3684
rect 4756 -3716 4760 -3684
rect 4720 -3720 4760 -3716
rect 4800 1036 4840 1040
rect 4800 1004 4804 1036
rect 4836 1004 4840 1036
rect 4800 956 4840 1004
rect 4800 924 4804 956
rect 4836 924 4840 956
rect 4800 876 4840 924
rect 4800 844 4804 876
rect 4836 844 4840 876
rect 4800 796 4840 844
rect 4800 764 4804 796
rect 4836 764 4840 796
rect 4800 716 4840 764
rect 4800 684 4804 716
rect 4836 684 4840 716
rect 4800 636 4840 684
rect 4800 604 4804 636
rect 4836 604 4840 636
rect 4800 556 4840 604
rect 4800 524 4804 556
rect 4836 524 4840 556
rect 4800 476 4840 524
rect 4800 444 4804 476
rect 4836 444 4840 476
rect 4800 396 4840 444
rect 4800 364 4804 396
rect 4836 364 4840 396
rect 4800 316 4840 364
rect 4800 284 4804 316
rect 4836 284 4840 316
rect 4800 236 4840 284
rect 4800 204 4804 236
rect 4836 204 4840 236
rect 4800 156 4840 204
rect 4800 124 4804 156
rect 4836 124 4840 156
rect 4800 76 4840 124
rect 4800 44 4804 76
rect 4836 44 4840 76
rect 4800 -4 4840 44
rect 4800 -36 4804 -4
rect 4836 -36 4840 -4
rect 4800 -84 4840 -36
rect 4800 -116 4804 -84
rect 4836 -116 4840 -84
rect 4800 -164 4840 -116
rect 4800 -196 4804 -164
rect 4836 -196 4840 -164
rect 4800 -244 4840 -196
rect 4800 -276 4804 -244
rect 4836 -276 4840 -244
rect 4800 -324 4840 -276
rect 4800 -356 4804 -324
rect 4836 -356 4840 -324
rect 4800 -404 4840 -356
rect 4800 -436 4804 -404
rect 4836 -436 4840 -404
rect 4800 -484 4840 -436
rect 4800 -516 4804 -484
rect 4836 -516 4840 -484
rect 4800 -564 4840 -516
rect 4800 -596 4804 -564
rect 4836 -596 4840 -564
rect 4800 -644 4840 -596
rect 4800 -676 4804 -644
rect 4836 -676 4840 -644
rect 4800 -724 4840 -676
rect 4800 -756 4804 -724
rect 4836 -756 4840 -724
rect 4800 -804 4840 -756
rect 4800 -836 4804 -804
rect 4836 -836 4840 -804
rect 4800 -884 4840 -836
rect 4800 -916 4804 -884
rect 4836 -916 4840 -884
rect 4800 -964 4840 -916
rect 4800 -996 4804 -964
rect 4836 -996 4840 -964
rect 4800 -1044 4840 -996
rect 4800 -1076 4804 -1044
rect 4836 -1076 4840 -1044
rect 4800 -1124 4840 -1076
rect 4800 -1156 4804 -1124
rect 4836 -1156 4840 -1124
rect 4800 -1204 4840 -1156
rect 4800 -1236 4804 -1204
rect 4836 -1236 4840 -1204
rect 4800 -1284 4840 -1236
rect 4800 -1316 4804 -1284
rect 4836 -1316 4840 -1284
rect 4800 -1364 4840 -1316
rect 4800 -1396 4804 -1364
rect 4836 -1396 4840 -1364
rect 4800 -1444 4840 -1396
rect 4800 -1476 4804 -1444
rect 4836 -1476 4840 -1444
rect 4800 -1524 4840 -1476
rect 4800 -1556 4804 -1524
rect 4836 -1556 4840 -1524
rect 4800 -1604 4840 -1556
rect 4800 -1636 4804 -1604
rect 4836 -1636 4840 -1604
rect 4800 -1684 4840 -1636
rect 4800 -1716 4804 -1684
rect 4836 -1716 4840 -1684
rect 4800 -1764 4840 -1716
rect 4800 -1796 4804 -1764
rect 4836 -1796 4840 -1764
rect 4800 -1844 4840 -1796
rect 4800 -1876 4804 -1844
rect 4836 -1876 4840 -1844
rect 4800 -1924 4840 -1876
rect 4800 -1956 4804 -1924
rect 4836 -1956 4840 -1924
rect 4800 -2004 4840 -1956
rect 4800 -2036 4804 -2004
rect 4836 -2036 4840 -2004
rect 4800 -2084 4840 -2036
rect 4800 -2116 4804 -2084
rect 4836 -2116 4840 -2084
rect 4800 -2164 4840 -2116
rect 4800 -2196 4804 -2164
rect 4836 -2196 4840 -2164
rect 4800 -2244 4840 -2196
rect 4800 -2276 4804 -2244
rect 4836 -2276 4840 -2244
rect 4800 -2324 4840 -2276
rect 4800 -2356 4804 -2324
rect 4836 -2356 4840 -2324
rect 4800 -2404 4840 -2356
rect 4800 -2436 4804 -2404
rect 4836 -2436 4840 -2404
rect 4800 -2484 4840 -2436
rect 4800 -2516 4804 -2484
rect 4836 -2516 4840 -2484
rect 4800 -2564 4840 -2516
rect 4800 -2596 4804 -2564
rect 4836 -2596 4840 -2564
rect 4800 -2644 4840 -2596
rect 4800 -2676 4804 -2644
rect 4836 -2676 4840 -2644
rect 4800 -2724 4840 -2676
rect 4800 -2756 4804 -2724
rect 4836 -2756 4840 -2724
rect 4800 -2804 4840 -2756
rect 4800 -2836 4804 -2804
rect 4836 -2836 4840 -2804
rect 4800 -2884 4840 -2836
rect 4800 -2916 4804 -2884
rect 4836 -2916 4840 -2884
rect 4800 -2964 4840 -2916
rect 4800 -2996 4804 -2964
rect 4836 -2996 4840 -2964
rect 4800 -3044 4840 -2996
rect 4800 -3076 4804 -3044
rect 4836 -3076 4840 -3044
rect 4800 -3124 4840 -3076
rect 4800 -3156 4804 -3124
rect 4836 -3156 4840 -3124
rect 4800 -3204 4840 -3156
rect 4800 -3236 4804 -3204
rect 4836 -3236 4840 -3204
rect 4800 -3284 4840 -3236
rect 4800 -3316 4804 -3284
rect 4836 -3316 4840 -3284
rect 4800 -3364 4840 -3316
rect 4800 -3396 4804 -3364
rect 4836 -3396 4840 -3364
rect 4800 -3444 4840 -3396
rect 4800 -3476 4804 -3444
rect 4836 -3476 4840 -3444
rect 4800 -3524 4840 -3476
rect 4800 -3556 4804 -3524
rect 4836 -3556 4840 -3524
rect 4800 -3604 4840 -3556
rect 4800 -3636 4804 -3604
rect 4836 -3636 4840 -3604
rect 4800 -3684 4840 -3636
rect 4800 -3716 4804 -3684
rect 4836 -3716 4840 -3684
rect 4800 -3720 4840 -3716
rect 4880 1036 4920 1040
rect 4880 1004 4884 1036
rect 4916 1004 4920 1036
rect 4880 956 4920 1004
rect 4880 924 4884 956
rect 4916 924 4920 956
rect 4880 876 4920 924
rect 4880 844 4884 876
rect 4916 844 4920 876
rect 4880 796 4920 844
rect 4880 764 4884 796
rect 4916 764 4920 796
rect 4880 716 4920 764
rect 4880 684 4884 716
rect 4916 684 4920 716
rect 4880 636 4920 684
rect 4880 604 4884 636
rect 4916 604 4920 636
rect 4880 556 4920 604
rect 4880 524 4884 556
rect 4916 524 4920 556
rect 4880 476 4920 524
rect 4880 444 4884 476
rect 4916 444 4920 476
rect 4880 396 4920 444
rect 4880 364 4884 396
rect 4916 364 4920 396
rect 4880 316 4920 364
rect 4880 284 4884 316
rect 4916 284 4920 316
rect 4880 236 4920 284
rect 4880 204 4884 236
rect 4916 204 4920 236
rect 4880 156 4920 204
rect 4880 124 4884 156
rect 4916 124 4920 156
rect 4880 76 4920 124
rect 4880 44 4884 76
rect 4916 44 4920 76
rect 4880 -4 4920 44
rect 4880 -36 4884 -4
rect 4916 -36 4920 -4
rect 4880 -84 4920 -36
rect 4880 -116 4884 -84
rect 4916 -116 4920 -84
rect 4880 -164 4920 -116
rect 4880 -196 4884 -164
rect 4916 -196 4920 -164
rect 4880 -244 4920 -196
rect 4880 -276 4884 -244
rect 4916 -276 4920 -244
rect 4880 -324 4920 -276
rect 4880 -356 4884 -324
rect 4916 -356 4920 -324
rect 4880 -404 4920 -356
rect 4880 -436 4884 -404
rect 4916 -436 4920 -404
rect 4880 -484 4920 -436
rect 4880 -516 4884 -484
rect 4916 -516 4920 -484
rect 4880 -564 4920 -516
rect 4880 -596 4884 -564
rect 4916 -596 4920 -564
rect 4880 -644 4920 -596
rect 4880 -676 4884 -644
rect 4916 -676 4920 -644
rect 4880 -724 4920 -676
rect 4880 -756 4884 -724
rect 4916 -756 4920 -724
rect 4880 -804 4920 -756
rect 4880 -836 4884 -804
rect 4916 -836 4920 -804
rect 4880 -884 4920 -836
rect 4880 -916 4884 -884
rect 4916 -916 4920 -884
rect 4880 -964 4920 -916
rect 4880 -996 4884 -964
rect 4916 -996 4920 -964
rect 4880 -1044 4920 -996
rect 4880 -1076 4884 -1044
rect 4916 -1076 4920 -1044
rect 4880 -1124 4920 -1076
rect 4880 -1156 4884 -1124
rect 4916 -1156 4920 -1124
rect 4880 -1204 4920 -1156
rect 4880 -1236 4884 -1204
rect 4916 -1236 4920 -1204
rect 4880 -1284 4920 -1236
rect 4880 -1316 4884 -1284
rect 4916 -1316 4920 -1284
rect 4880 -1364 4920 -1316
rect 4880 -1396 4884 -1364
rect 4916 -1396 4920 -1364
rect 4880 -1444 4920 -1396
rect 4880 -1476 4884 -1444
rect 4916 -1476 4920 -1444
rect 4880 -1524 4920 -1476
rect 4880 -1556 4884 -1524
rect 4916 -1556 4920 -1524
rect 4880 -1604 4920 -1556
rect 4880 -1636 4884 -1604
rect 4916 -1636 4920 -1604
rect 4880 -1684 4920 -1636
rect 4880 -1716 4884 -1684
rect 4916 -1716 4920 -1684
rect 4880 -1764 4920 -1716
rect 4880 -1796 4884 -1764
rect 4916 -1796 4920 -1764
rect 4880 -1844 4920 -1796
rect 4880 -1876 4884 -1844
rect 4916 -1876 4920 -1844
rect 4880 -1924 4920 -1876
rect 4880 -1956 4884 -1924
rect 4916 -1956 4920 -1924
rect 4880 -2004 4920 -1956
rect 4880 -2036 4884 -2004
rect 4916 -2036 4920 -2004
rect 4880 -2084 4920 -2036
rect 4880 -2116 4884 -2084
rect 4916 -2116 4920 -2084
rect 4880 -2164 4920 -2116
rect 4880 -2196 4884 -2164
rect 4916 -2196 4920 -2164
rect 4880 -2244 4920 -2196
rect 4880 -2276 4884 -2244
rect 4916 -2276 4920 -2244
rect 4880 -2324 4920 -2276
rect 4880 -2356 4884 -2324
rect 4916 -2356 4920 -2324
rect 4880 -2404 4920 -2356
rect 4880 -2436 4884 -2404
rect 4916 -2436 4920 -2404
rect 4880 -2484 4920 -2436
rect 4880 -2516 4884 -2484
rect 4916 -2516 4920 -2484
rect 4880 -2564 4920 -2516
rect 4880 -2596 4884 -2564
rect 4916 -2596 4920 -2564
rect 4880 -2644 4920 -2596
rect 4880 -2676 4884 -2644
rect 4916 -2676 4920 -2644
rect 4880 -2724 4920 -2676
rect 4880 -2756 4884 -2724
rect 4916 -2756 4920 -2724
rect 4880 -2804 4920 -2756
rect 4880 -2836 4884 -2804
rect 4916 -2836 4920 -2804
rect 4880 -2884 4920 -2836
rect 4880 -2916 4884 -2884
rect 4916 -2916 4920 -2884
rect 4880 -2964 4920 -2916
rect 4880 -2996 4884 -2964
rect 4916 -2996 4920 -2964
rect 4880 -3044 4920 -2996
rect 4880 -3076 4884 -3044
rect 4916 -3076 4920 -3044
rect 4880 -3124 4920 -3076
rect 4880 -3156 4884 -3124
rect 4916 -3156 4920 -3124
rect 4880 -3204 4920 -3156
rect 4880 -3236 4884 -3204
rect 4916 -3236 4920 -3204
rect 4880 -3284 4920 -3236
rect 4880 -3316 4884 -3284
rect 4916 -3316 4920 -3284
rect 4880 -3364 4920 -3316
rect 4880 -3396 4884 -3364
rect 4916 -3396 4920 -3364
rect 4880 -3444 4920 -3396
rect 4880 -3476 4884 -3444
rect 4916 -3476 4920 -3444
rect 4880 -3524 4920 -3476
rect 4880 -3556 4884 -3524
rect 4916 -3556 4920 -3524
rect 4880 -3604 4920 -3556
rect 4880 -3636 4884 -3604
rect 4916 -3636 4920 -3604
rect 4880 -3684 4920 -3636
rect 4880 -3716 4884 -3684
rect 4916 -3716 4920 -3684
rect 4880 -3720 4920 -3716
rect 4960 1036 5000 1040
rect 4960 1004 4964 1036
rect 4996 1004 5000 1036
rect 4960 956 5000 1004
rect 4960 924 4964 956
rect 4996 924 5000 956
rect 4960 876 5000 924
rect 4960 844 4964 876
rect 4996 844 5000 876
rect 4960 796 5000 844
rect 4960 764 4964 796
rect 4996 764 5000 796
rect 4960 716 5000 764
rect 4960 684 4964 716
rect 4996 684 5000 716
rect 4960 636 5000 684
rect 4960 604 4964 636
rect 4996 604 5000 636
rect 4960 556 5000 604
rect 4960 524 4964 556
rect 4996 524 5000 556
rect 4960 476 5000 524
rect 4960 444 4964 476
rect 4996 444 5000 476
rect 4960 396 5000 444
rect 4960 364 4964 396
rect 4996 364 5000 396
rect 4960 316 5000 364
rect 4960 284 4964 316
rect 4996 284 5000 316
rect 4960 236 5000 284
rect 4960 204 4964 236
rect 4996 204 5000 236
rect 4960 156 5000 204
rect 4960 124 4964 156
rect 4996 124 5000 156
rect 4960 76 5000 124
rect 4960 44 4964 76
rect 4996 44 5000 76
rect 4960 -4 5000 44
rect 4960 -36 4964 -4
rect 4996 -36 5000 -4
rect 4960 -84 5000 -36
rect 4960 -116 4964 -84
rect 4996 -116 5000 -84
rect 4960 -164 5000 -116
rect 4960 -196 4964 -164
rect 4996 -196 5000 -164
rect 4960 -244 5000 -196
rect 4960 -276 4964 -244
rect 4996 -276 5000 -244
rect 4960 -324 5000 -276
rect 4960 -356 4964 -324
rect 4996 -356 5000 -324
rect 4960 -404 5000 -356
rect 4960 -436 4964 -404
rect 4996 -436 5000 -404
rect 4960 -484 5000 -436
rect 4960 -516 4964 -484
rect 4996 -516 5000 -484
rect 4960 -564 5000 -516
rect 4960 -596 4964 -564
rect 4996 -596 5000 -564
rect 4960 -644 5000 -596
rect 4960 -676 4964 -644
rect 4996 -676 5000 -644
rect 4960 -724 5000 -676
rect 4960 -756 4964 -724
rect 4996 -756 5000 -724
rect 4960 -804 5000 -756
rect 4960 -836 4964 -804
rect 4996 -836 5000 -804
rect 4960 -884 5000 -836
rect 4960 -916 4964 -884
rect 4996 -916 5000 -884
rect 4960 -964 5000 -916
rect 4960 -996 4964 -964
rect 4996 -996 5000 -964
rect 4960 -1044 5000 -996
rect 4960 -1076 4964 -1044
rect 4996 -1076 5000 -1044
rect 4960 -1124 5000 -1076
rect 4960 -1156 4964 -1124
rect 4996 -1156 5000 -1124
rect 4960 -1204 5000 -1156
rect 4960 -1236 4964 -1204
rect 4996 -1236 5000 -1204
rect 4960 -1284 5000 -1236
rect 4960 -1316 4964 -1284
rect 4996 -1316 5000 -1284
rect 4960 -1364 5000 -1316
rect 4960 -1396 4964 -1364
rect 4996 -1396 5000 -1364
rect 4960 -1444 5000 -1396
rect 4960 -1476 4964 -1444
rect 4996 -1476 5000 -1444
rect 4960 -1524 5000 -1476
rect 4960 -1556 4964 -1524
rect 4996 -1556 5000 -1524
rect 4960 -1604 5000 -1556
rect 4960 -1636 4964 -1604
rect 4996 -1636 5000 -1604
rect 4960 -1684 5000 -1636
rect 4960 -1716 4964 -1684
rect 4996 -1716 5000 -1684
rect 4960 -1764 5000 -1716
rect 4960 -1796 4964 -1764
rect 4996 -1796 5000 -1764
rect 4960 -1844 5000 -1796
rect 4960 -1876 4964 -1844
rect 4996 -1876 5000 -1844
rect 4960 -1924 5000 -1876
rect 4960 -1956 4964 -1924
rect 4996 -1956 5000 -1924
rect 4960 -2004 5000 -1956
rect 4960 -2036 4964 -2004
rect 4996 -2036 5000 -2004
rect 4960 -2084 5000 -2036
rect 4960 -2116 4964 -2084
rect 4996 -2116 5000 -2084
rect 4960 -2164 5000 -2116
rect 4960 -2196 4964 -2164
rect 4996 -2196 5000 -2164
rect 4960 -2244 5000 -2196
rect 4960 -2276 4964 -2244
rect 4996 -2276 5000 -2244
rect 4960 -2324 5000 -2276
rect 4960 -2356 4964 -2324
rect 4996 -2356 5000 -2324
rect 4960 -2404 5000 -2356
rect 4960 -2436 4964 -2404
rect 4996 -2436 5000 -2404
rect 4960 -2484 5000 -2436
rect 4960 -2516 4964 -2484
rect 4996 -2516 5000 -2484
rect 4960 -2564 5000 -2516
rect 4960 -2596 4964 -2564
rect 4996 -2596 5000 -2564
rect 4960 -2644 5000 -2596
rect 4960 -2676 4964 -2644
rect 4996 -2676 5000 -2644
rect 4960 -2724 5000 -2676
rect 4960 -2756 4964 -2724
rect 4996 -2756 5000 -2724
rect 4960 -2804 5000 -2756
rect 4960 -2836 4964 -2804
rect 4996 -2836 5000 -2804
rect 4960 -2884 5000 -2836
rect 4960 -2916 4964 -2884
rect 4996 -2916 5000 -2884
rect 4960 -2964 5000 -2916
rect 4960 -2996 4964 -2964
rect 4996 -2996 5000 -2964
rect 4960 -3044 5000 -2996
rect 4960 -3076 4964 -3044
rect 4996 -3076 5000 -3044
rect 4960 -3124 5000 -3076
rect 4960 -3156 4964 -3124
rect 4996 -3156 5000 -3124
rect 4960 -3204 5000 -3156
rect 4960 -3236 4964 -3204
rect 4996 -3236 5000 -3204
rect 4960 -3284 5000 -3236
rect 4960 -3316 4964 -3284
rect 4996 -3316 5000 -3284
rect 4960 -3364 5000 -3316
rect 4960 -3396 4964 -3364
rect 4996 -3396 5000 -3364
rect 4960 -3444 5000 -3396
rect 4960 -3476 4964 -3444
rect 4996 -3476 5000 -3444
rect 4960 -3524 5000 -3476
rect 4960 -3556 4964 -3524
rect 4996 -3556 5000 -3524
rect 4960 -3604 5000 -3556
rect 4960 -3636 4964 -3604
rect 4996 -3636 5000 -3604
rect 4960 -3684 5000 -3636
rect 4960 -3716 4964 -3684
rect 4996 -3716 5000 -3684
rect 4960 -3720 5000 -3716
rect 5040 1036 5080 1040
rect 5040 1004 5044 1036
rect 5076 1004 5080 1036
rect 5040 956 5080 1004
rect 5040 924 5044 956
rect 5076 924 5080 956
rect 5040 876 5080 924
rect 5040 844 5044 876
rect 5076 844 5080 876
rect 5040 796 5080 844
rect 5040 764 5044 796
rect 5076 764 5080 796
rect 5040 716 5080 764
rect 5040 684 5044 716
rect 5076 684 5080 716
rect 5040 636 5080 684
rect 5040 604 5044 636
rect 5076 604 5080 636
rect 5040 556 5080 604
rect 5040 524 5044 556
rect 5076 524 5080 556
rect 5040 476 5080 524
rect 5040 444 5044 476
rect 5076 444 5080 476
rect 5040 396 5080 444
rect 5040 364 5044 396
rect 5076 364 5080 396
rect 5040 316 5080 364
rect 5040 284 5044 316
rect 5076 284 5080 316
rect 5040 236 5080 284
rect 5040 204 5044 236
rect 5076 204 5080 236
rect 5040 156 5080 204
rect 5040 124 5044 156
rect 5076 124 5080 156
rect 5040 76 5080 124
rect 5040 44 5044 76
rect 5076 44 5080 76
rect 5040 -4 5080 44
rect 5040 -36 5044 -4
rect 5076 -36 5080 -4
rect 5040 -84 5080 -36
rect 5040 -116 5044 -84
rect 5076 -116 5080 -84
rect 5040 -164 5080 -116
rect 5040 -196 5044 -164
rect 5076 -196 5080 -164
rect 5040 -244 5080 -196
rect 5040 -276 5044 -244
rect 5076 -276 5080 -244
rect 5040 -324 5080 -276
rect 5040 -356 5044 -324
rect 5076 -356 5080 -324
rect 5040 -404 5080 -356
rect 5040 -436 5044 -404
rect 5076 -436 5080 -404
rect 5040 -484 5080 -436
rect 5040 -516 5044 -484
rect 5076 -516 5080 -484
rect 5040 -564 5080 -516
rect 5040 -596 5044 -564
rect 5076 -596 5080 -564
rect 5040 -644 5080 -596
rect 5040 -676 5044 -644
rect 5076 -676 5080 -644
rect 5040 -724 5080 -676
rect 5040 -756 5044 -724
rect 5076 -756 5080 -724
rect 5040 -804 5080 -756
rect 5040 -836 5044 -804
rect 5076 -836 5080 -804
rect 5040 -884 5080 -836
rect 5040 -916 5044 -884
rect 5076 -916 5080 -884
rect 5040 -964 5080 -916
rect 5040 -996 5044 -964
rect 5076 -996 5080 -964
rect 5040 -1044 5080 -996
rect 5040 -1076 5044 -1044
rect 5076 -1076 5080 -1044
rect 5040 -1124 5080 -1076
rect 5040 -1156 5044 -1124
rect 5076 -1156 5080 -1124
rect 5040 -1204 5080 -1156
rect 5040 -1236 5044 -1204
rect 5076 -1236 5080 -1204
rect 5040 -1284 5080 -1236
rect 5040 -1316 5044 -1284
rect 5076 -1316 5080 -1284
rect 5040 -1364 5080 -1316
rect 5040 -1396 5044 -1364
rect 5076 -1396 5080 -1364
rect 5040 -1444 5080 -1396
rect 5040 -1476 5044 -1444
rect 5076 -1476 5080 -1444
rect 5040 -1524 5080 -1476
rect 5040 -1556 5044 -1524
rect 5076 -1556 5080 -1524
rect 5040 -1604 5080 -1556
rect 5040 -1636 5044 -1604
rect 5076 -1636 5080 -1604
rect 5040 -1684 5080 -1636
rect 5040 -1716 5044 -1684
rect 5076 -1716 5080 -1684
rect 5040 -1764 5080 -1716
rect 5040 -1796 5044 -1764
rect 5076 -1796 5080 -1764
rect 5040 -1844 5080 -1796
rect 5040 -1876 5044 -1844
rect 5076 -1876 5080 -1844
rect 5040 -1924 5080 -1876
rect 5040 -1956 5044 -1924
rect 5076 -1956 5080 -1924
rect 5040 -2004 5080 -1956
rect 5040 -2036 5044 -2004
rect 5076 -2036 5080 -2004
rect 5040 -2084 5080 -2036
rect 5040 -2116 5044 -2084
rect 5076 -2116 5080 -2084
rect 5040 -2164 5080 -2116
rect 5040 -2196 5044 -2164
rect 5076 -2196 5080 -2164
rect 5040 -2244 5080 -2196
rect 5040 -2276 5044 -2244
rect 5076 -2276 5080 -2244
rect 5040 -2324 5080 -2276
rect 5040 -2356 5044 -2324
rect 5076 -2356 5080 -2324
rect 5040 -2404 5080 -2356
rect 5040 -2436 5044 -2404
rect 5076 -2436 5080 -2404
rect 5040 -2484 5080 -2436
rect 5040 -2516 5044 -2484
rect 5076 -2516 5080 -2484
rect 5040 -2564 5080 -2516
rect 5040 -2596 5044 -2564
rect 5076 -2596 5080 -2564
rect 5040 -2644 5080 -2596
rect 5040 -2676 5044 -2644
rect 5076 -2676 5080 -2644
rect 5040 -2724 5080 -2676
rect 5040 -2756 5044 -2724
rect 5076 -2756 5080 -2724
rect 5040 -2804 5080 -2756
rect 5040 -2836 5044 -2804
rect 5076 -2836 5080 -2804
rect 5040 -2884 5080 -2836
rect 5040 -2916 5044 -2884
rect 5076 -2916 5080 -2884
rect 5040 -2964 5080 -2916
rect 5040 -2996 5044 -2964
rect 5076 -2996 5080 -2964
rect 5040 -3044 5080 -2996
rect 5040 -3076 5044 -3044
rect 5076 -3076 5080 -3044
rect 5040 -3124 5080 -3076
rect 5040 -3156 5044 -3124
rect 5076 -3156 5080 -3124
rect 5040 -3204 5080 -3156
rect 5040 -3236 5044 -3204
rect 5076 -3236 5080 -3204
rect 5040 -3284 5080 -3236
rect 5040 -3316 5044 -3284
rect 5076 -3316 5080 -3284
rect 5040 -3364 5080 -3316
rect 5040 -3396 5044 -3364
rect 5076 -3396 5080 -3364
rect 5040 -3444 5080 -3396
rect 5040 -3476 5044 -3444
rect 5076 -3476 5080 -3444
rect 5040 -3524 5080 -3476
rect 5040 -3556 5044 -3524
rect 5076 -3556 5080 -3524
rect 5040 -3604 5080 -3556
rect 5040 -3636 5044 -3604
rect 5076 -3636 5080 -3604
rect 5040 -3684 5080 -3636
rect 5040 -3716 5044 -3684
rect 5076 -3716 5080 -3684
rect 5040 -3720 5080 -3716
rect 5120 1036 5160 1040
rect 5120 1004 5124 1036
rect 5156 1004 5160 1036
rect 5120 956 5160 1004
rect 5120 924 5124 956
rect 5156 924 5160 956
rect 5120 876 5160 924
rect 5120 844 5124 876
rect 5156 844 5160 876
rect 5120 796 5160 844
rect 5120 764 5124 796
rect 5156 764 5160 796
rect 5120 716 5160 764
rect 5120 684 5124 716
rect 5156 684 5160 716
rect 5120 636 5160 684
rect 5120 604 5124 636
rect 5156 604 5160 636
rect 5120 556 5160 604
rect 5120 524 5124 556
rect 5156 524 5160 556
rect 5120 476 5160 524
rect 5120 444 5124 476
rect 5156 444 5160 476
rect 5120 396 5160 444
rect 5120 364 5124 396
rect 5156 364 5160 396
rect 5120 316 5160 364
rect 5120 284 5124 316
rect 5156 284 5160 316
rect 5120 236 5160 284
rect 5120 204 5124 236
rect 5156 204 5160 236
rect 5120 156 5160 204
rect 5120 124 5124 156
rect 5156 124 5160 156
rect 5120 76 5160 124
rect 5120 44 5124 76
rect 5156 44 5160 76
rect 5120 -4 5160 44
rect 5120 -36 5124 -4
rect 5156 -36 5160 -4
rect 5120 -84 5160 -36
rect 5120 -116 5124 -84
rect 5156 -116 5160 -84
rect 5120 -164 5160 -116
rect 5120 -196 5124 -164
rect 5156 -196 5160 -164
rect 5120 -244 5160 -196
rect 5120 -276 5124 -244
rect 5156 -276 5160 -244
rect 5120 -324 5160 -276
rect 5120 -356 5124 -324
rect 5156 -356 5160 -324
rect 5120 -404 5160 -356
rect 5120 -436 5124 -404
rect 5156 -436 5160 -404
rect 5120 -484 5160 -436
rect 5120 -516 5124 -484
rect 5156 -516 5160 -484
rect 5120 -564 5160 -516
rect 5120 -596 5124 -564
rect 5156 -596 5160 -564
rect 5120 -644 5160 -596
rect 5120 -676 5124 -644
rect 5156 -676 5160 -644
rect 5120 -724 5160 -676
rect 5120 -756 5124 -724
rect 5156 -756 5160 -724
rect 5120 -804 5160 -756
rect 5120 -836 5124 -804
rect 5156 -836 5160 -804
rect 5120 -884 5160 -836
rect 5120 -916 5124 -884
rect 5156 -916 5160 -884
rect 5120 -964 5160 -916
rect 5120 -996 5124 -964
rect 5156 -996 5160 -964
rect 5120 -1044 5160 -996
rect 5120 -1076 5124 -1044
rect 5156 -1076 5160 -1044
rect 5120 -1124 5160 -1076
rect 5120 -1156 5124 -1124
rect 5156 -1156 5160 -1124
rect 5120 -1204 5160 -1156
rect 5120 -1236 5124 -1204
rect 5156 -1236 5160 -1204
rect 5120 -1284 5160 -1236
rect 5120 -1316 5124 -1284
rect 5156 -1316 5160 -1284
rect 5120 -1364 5160 -1316
rect 5120 -1396 5124 -1364
rect 5156 -1396 5160 -1364
rect 5120 -1444 5160 -1396
rect 5120 -1476 5124 -1444
rect 5156 -1476 5160 -1444
rect 5120 -1524 5160 -1476
rect 5120 -1556 5124 -1524
rect 5156 -1556 5160 -1524
rect 5120 -1604 5160 -1556
rect 5120 -1636 5124 -1604
rect 5156 -1636 5160 -1604
rect 5120 -1684 5160 -1636
rect 5120 -1716 5124 -1684
rect 5156 -1716 5160 -1684
rect 5120 -1764 5160 -1716
rect 5120 -1796 5124 -1764
rect 5156 -1796 5160 -1764
rect 5120 -1844 5160 -1796
rect 5120 -1876 5124 -1844
rect 5156 -1876 5160 -1844
rect 5120 -1924 5160 -1876
rect 5120 -1956 5124 -1924
rect 5156 -1956 5160 -1924
rect 5120 -2004 5160 -1956
rect 5120 -2036 5124 -2004
rect 5156 -2036 5160 -2004
rect 5120 -2084 5160 -2036
rect 5120 -2116 5124 -2084
rect 5156 -2116 5160 -2084
rect 5120 -2164 5160 -2116
rect 5120 -2196 5124 -2164
rect 5156 -2196 5160 -2164
rect 5120 -2244 5160 -2196
rect 5120 -2276 5124 -2244
rect 5156 -2276 5160 -2244
rect 5120 -2324 5160 -2276
rect 5120 -2356 5124 -2324
rect 5156 -2356 5160 -2324
rect 5120 -2404 5160 -2356
rect 5120 -2436 5124 -2404
rect 5156 -2436 5160 -2404
rect 5120 -2484 5160 -2436
rect 5120 -2516 5124 -2484
rect 5156 -2516 5160 -2484
rect 5120 -2564 5160 -2516
rect 5120 -2596 5124 -2564
rect 5156 -2596 5160 -2564
rect 5120 -2644 5160 -2596
rect 5120 -2676 5124 -2644
rect 5156 -2676 5160 -2644
rect 5120 -2724 5160 -2676
rect 5120 -2756 5124 -2724
rect 5156 -2756 5160 -2724
rect 5120 -2804 5160 -2756
rect 5120 -2836 5124 -2804
rect 5156 -2836 5160 -2804
rect 5120 -2884 5160 -2836
rect 5120 -2916 5124 -2884
rect 5156 -2916 5160 -2884
rect 5120 -2964 5160 -2916
rect 5120 -2996 5124 -2964
rect 5156 -2996 5160 -2964
rect 5120 -3044 5160 -2996
rect 5120 -3076 5124 -3044
rect 5156 -3076 5160 -3044
rect 5120 -3124 5160 -3076
rect 5120 -3156 5124 -3124
rect 5156 -3156 5160 -3124
rect 5120 -3204 5160 -3156
rect 5120 -3236 5124 -3204
rect 5156 -3236 5160 -3204
rect 5120 -3284 5160 -3236
rect 5120 -3316 5124 -3284
rect 5156 -3316 5160 -3284
rect 5120 -3364 5160 -3316
rect 5120 -3396 5124 -3364
rect 5156 -3396 5160 -3364
rect 5120 -3444 5160 -3396
rect 5120 -3476 5124 -3444
rect 5156 -3476 5160 -3444
rect 5120 -3524 5160 -3476
rect 5120 -3556 5124 -3524
rect 5156 -3556 5160 -3524
rect 5120 -3604 5160 -3556
rect 5120 -3636 5124 -3604
rect 5156 -3636 5160 -3604
rect 5120 -3684 5160 -3636
rect 5120 -3716 5124 -3684
rect 5156 -3716 5160 -3684
rect 5120 -3720 5160 -3716
rect 5200 1036 5240 1040
rect 5200 1004 5204 1036
rect 5236 1004 5240 1036
rect 5200 956 5240 1004
rect 5200 924 5204 956
rect 5236 924 5240 956
rect 5200 876 5240 924
rect 5200 844 5204 876
rect 5236 844 5240 876
rect 5200 796 5240 844
rect 5200 764 5204 796
rect 5236 764 5240 796
rect 5200 716 5240 764
rect 5200 684 5204 716
rect 5236 684 5240 716
rect 5200 636 5240 684
rect 5200 604 5204 636
rect 5236 604 5240 636
rect 5200 556 5240 604
rect 5200 524 5204 556
rect 5236 524 5240 556
rect 5200 476 5240 524
rect 5200 444 5204 476
rect 5236 444 5240 476
rect 5200 396 5240 444
rect 5200 364 5204 396
rect 5236 364 5240 396
rect 5200 316 5240 364
rect 5200 284 5204 316
rect 5236 284 5240 316
rect 5200 236 5240 284
rect 5200 204 5204 236
rect 5236 204 5240 236
rect 5200 156 5240 204
rect 5200 124 5204 156
rect 5236 124 5240 156
rect 5200 76 5240 124
rect 5200 44 5204 76
rect 5236 44 5240 76
rect 5200 -4 5240 44
rect 5200 -36 5204 -4
rect 5236 -36 5240 -4
rect 5200 -84 5240 -36
rect 5200 -116 5204 -84
rect 5236 -116 5240 -84
rect 5200 -164 5240 -116
rect 5200 -196 5204 -164
rect 5236 -196 5240 -164
rect 5200 -244 5240 -196
rect 5200 -276 5204 -244
rect 5236 -276 5240 -244
rect 5200 -324 5240 -276
rect 5200 -356 5204 -324
rect 5236 -356 5240 -324
rect 5200 -404 5240 -356
rect 5200 -436 5204 -404
rect 5236 -436 5240 -404
rect 5200 -484 5240 -436
rect 5200 -516 5204 -484
rect 5236 -516 5240 -484
rect 5200 -564 5240 -516
rect 5200 -596 5204 -564
rect 5236 -596 5240 -564
rect 5200 -644 5240 -596
rect 5200 -676 5204 -644
rect 5236 -676 5240 -644
rect 5200 -724 5240 -676
rect 5200 -756 5204 -724
rect 5236 -756 5240 -724
rect 5200 -804 5240 -756
rect 5200 -836 5204 -804
rect 5236 -836 5240 -804
rect 5200 -884 5240 -836
rect 5200 -916 5204 -884
rect 5236 -916 5240 -884
rect 5200 -964 5240 -916
rect 5200 -996 5204 -964
rect 5236 -996 5240 -964
rect 5200 -1044 5240 -996
rect 5200 -1076 5204 -1044
rect 5236 -1076 5240 -1044
rect 5200 -1124 5240 -1076
rect 5200 -1156 5204 -1124
rect 5236 -1156 5240 -1124
rect 5200 -1204 5240 -1156
rect 5200 -1236 5204 -1204
rect 5236 -1236 5240 -1204
rect 5200 -1284 5240 -1236
rect 5200 -1316 5204 -1284
rect 5236 -1316 5240 -1284
rect 5200 -1364 5240 -1316
rect 5200 -1396 5204 -1364
rect 5236 -1396 5240 -1364
rect 5200 -1444 5240 -1396
rect 5200 -1476 5204 -1444
rect 5236 -1476 5240 -1444
rect 5200 -1524 5240 -1476
rect 5200 -1556 5204 -1524
rect 5236 -1556 5240 -1524
rect 5200 -1604 5240 -1556
rect 5200 -1636 5204 -1604
rect 5236 -1636 5240 -1604
rect 5200 -1684 5240 -1636
rect 5200 -1716 5204 -1684
rect 5236 -1716 5240 -1684
rect 5200 -1764 5240 -1716
rect 5200 -1796 5204 -1764
rect 5236 -1796 5240 -1764
rect 5200 -1844 5240 -1796
rect 5200 -1876 5204 -1844
rect 5236 -1876 5240 -1844
rect 5200 -1924 5240 -1876
rect 5200 -1956 5204 -1924
rect 5236 -1956 5240 -1924
rect 5200 -2004 5240 -1956
rect 5200 -2036 5204 -2004
rect 5236 -2036 5240 -2004
rect 5200 -2084 5240 -2036
rect 5200 -2116 5204 -2084
rect 5236 -2116 5240 -2084
rect 5200 -2164 5240 -2116
rect 5200 -2196 5204 -2164
rect 5236 -2196 5240 -2164
rect 5200 -2244 5240 -2196
rect 5200 -2276 5204 -2244
rect 5236 -2276 5240 -2244
rect 5200 -2324 5240 -2276
rect 5200 -2356 5204 -2324
rect 5236 -2356 5240 -2324
rect 5200 -2404 5240 -2356
rect 5200 -2436 5204 -2404
rect 5236 -2436 5240 -2404
rect 5200 -2484 5240 -2436
rect 5200 -2516 5204 -2484
rect 5236 -2516 5240 -2484
rect 5200 -2564 5240 -2516
rect 5200 -2596 5204 -2564
rect 5236 -2596 5240 -2564
rect 5200 -2644 5240 -2596
rect 5200 -2676 5204 -2644
rect 5236 -2676 5240 -2644
rect 5200 -2724 5240 -2676
rect 5200 -2756 5204 -2724
rect 5236 -2756 5240 -2724
rect 5200 -2804 5240 -2756
rect 5200 -2836 5204 -2804
rect 5236 -2836 5240 -2804
rect 5200 -2884 5240 -2836
rect 5200 -2916 5204 -2884
rect 5236 -2916 5240 -2884
rect 5200 -2964 5240 -2916
rect 5200 -2996 5204 -2964
rect 5236 -2996 5240 -2964
rect 5200 -3044 5240 -2996
rect 5200 -3076 5204 -3044
rect 5236 -3076 5240 -3044
rect 5200 -3124 5240 -3076
rect 5200 -3156 5204 -3124
rect 5236 -3156 5240 -3124
rect 5200 -3204 5240 -3156
rect 5200 -3236 5204 -3204
rect 5236 -3236 5240 -3204
rect 5200 -3284 5240 -3236
rect 5200 -3316 5204 -3284
rect 5236 -3316 5240 -3284
rect 5200 -3364 5240 -3316
rect 5200 -3396 5204 -3364
rect 5236 -3396 5240 -3364
rect 5200 -3444 5240 -3396
rect 5200 -3476 5204 -3444
rect 5236 -3476 5240 -3444
rect 5200 -3524 5240 -3476
rect 5200 -3556 5204 -3524
rect 5236 -3556 5240 -3524
rect 5200 -3604 5240 -3556
rect 5200 -3636 5204 -3604
rect 5236 -3636 5240 -3604
rect 5200 -3684 5240 -3636
rect 5200 -3716 5204 -3684
rect 5236 -3716 5240 -3684
rect 5200 -3720 5240 -3716
rect 5280 1036 5320 1040
rect 5280 1004 5284 1036
rect 5316 1004 5320 1036
rect 5280 956 5320 1004
rect 5280 924 5284 956
rect 5316 924 5320 956
rect 5280 876 5320 924
rect 5280 844 5284 876
rect 5316 844 5320 876
rect 5280 796 5320 844
rect 5280 764 5284 796
rect 5316 764 5320 796
rect 5280 716 5320 764
rect 5280 684 5284 716
rect 5316 684 5320 716
rect 5280 636 5320 684
rect 5280 604 5284 636
rect 5316 604 5320 636
rect 5280 556 5320 604
rect 5280 524 5284 556
rect 5316 524 5320 556
rect 5280 476 5320 524
rect 5280 444 5284 476
rect 5316 444 5320 476
rect 5280 396 5320 444
rect 5280 364 5284 396
rect 5316 364 5320 396
rect 5280 316 5320 364
rect 5280 284 5284 316
rect 5316 284 5320 316
rect 5280 236 5320 284
rect 5280 204 5284 236
rect 5316 204 5320 236
rect 5280 156 5320 204
rect 5280 124 5284 156
rect 5316 124 5320 156
rect 5280 76 5320 124
rect 5280 44 5284 76
rect 5316 44 5320 76
rect 5280 -4 5320 44
rect 5280 -36 5284 -4
rect 5316 -36 5320 -4
rect 5280 -84 5320 -36
rect 5280 -116 5284 -84
rect 5316 -116 5320 -84
rect 5280 -164 5320 -116
rect 5280 -196 5284 -164
rect 5316 -196 5320 -164
rect 5280 -244 5320 -196
rect 5280 -276 5284 -244
rect 5316 -276 5320 -244
rect 5280 -324 5320 -276
rect 5280 -356 5284 -324
rect 5316 -356 5320 -324
rect 5280 -404 5320 -356
rect 5280 -436 5284 -404
rect 5316 -436 5320 -404
rect 5280 -484 5320 -436
rect 5280 -516 5284 -484
rect 5316 -516 5320 -484
rect 5280 -564 5320 -516
rect 5280 -596 5284 -564
rect 5316 -596 5320 -564
rect 5280 -644 5320 -596
rect 5280 -676 5284 -644
rect 5316 -676 5320 -644
rect 5280 -724 5320 -676
rect 5280 -756 5284 -724
rect 5316 -756 5320 -724
rect 5280 -804 5320 -756
rect 5280 -836 5284 -804
rect 5316 -836 5320 -804
rect 5280 -884 5320 -836
rect 5280 -916 5284 -884
rect 5316 -916 5320 -884
rect 5280 -964 5320 -916
rect 5280 -996 5284 -964
rect 5316 -996 5320 -964
rect 5280 -1044 5320 -996
rect 5280 -1076 5284 -1044
rect 5316 -1076 5320 -1044
rect 5280 -1124 5320 -1076
rect 5280 -1156 5284 -1124
rect 5316 -1156 5320 -1124
rect 5280 -1204 5320 -1156
rect 5280 -1236 5284 -1204
rect 5316 -1236 5320 -1204
rect 5280 -1284 5320 -1236
rect 5280 -1316 5284 -1284
rect 5316 -1316 5320 -1284
rect 5280 -1364 5320 -1316
rect 5280 -1396 5284 -1364
rect 5316 -1396 5320 -1364
rect 5280 -1444 5320 -1396
rect 5280 -1476 5284 -1444
rect 5316 -1476 5320 -1444
rect 5280 -1524 5320 -1476
rect 5280 -1556 5284 -1524
rect 5316 -1556 5320 -1524
rect 5280 -1604 5320 -1556
rect 5280 -1636 5284 -1604
rect 5316 -1636 5320 -1604
rect 5280 -1684 5320 -1636
rect 5280 -1716 5284 -1684
rect 5316 -1716 5320 -1684
rect 5280 -1764 5320 -1716
rect 5280 -1796 5284 -1764
rect 5316 -1796 5320 -1764
rect 5280 -1844 5320 -1796
rect 5280 -1876 5284 -1844
rect 5316 -1876 5320 -1844
rect 5280 -1924 5320 -1876
rect 5280 -1956 5284 -1924
rect 5316 -1956 5320 -1924
rect 5280 -2004 5320 -1956
rect 5280 -2036 5284 -2004
rect 5316 -2036 5320 -2004
rect 5280 -2084 5320 -2036
rect 5280 -2116 5284 -2084
rect 5316 -2116 5320 -2084
rect 5280 -2164 5320 -2116
rect 5280 -2196 5284 -2164
rect 5316 -2196 5320 -2164
rect 5280 -2244 5320 -2196
rect 5280 -2276 5284 -2244
rect 5316 -2276 5320 -2244
rect 5280 -2324 5320 -2276
rect 5280 -2356 5284 -2324
rect 5316 -2356 5320 -2324
rect 5280 -2404 5320 -2356
rect 5280 -2436 5284 -2404
rect 5316 -2436 5320 -2404
rect 5280 -2484 5320 -2436
rect 5280 -2516 5284 -2484
rect 5316 -2516 5320 -2484
rect 5280 -2564 5320 -2516
rect 5280 -2596 5284 -2564
rect 5316 -2596 5320 -2564
rect 5280 -2644 5320 -2596
rect 5280 -2676 5284 -2644
rect 5316 -2676 5320 -2644
rect 5280 -2724 5320 -2676
rect 5280 -2756 5284 -2724
rect 5316 -2756 5320 -2724
rect 5280 -2804 5320 -2756
rect 5280 -2836 5284 -2804
rect 5316 -2836 5320 -2804
rect 5280 -2884 5320 -2836
rect 5280 -2916 5284 -2884
rect 5316 -2916 5320 -2884
rect 5280 -2964 5320 -2916
rect 5280 -2996 5284 -2964
rect 5316 -2996 5320 -2964
rect 5280 -3044 5320 -2996
rect 5280 -3076 5284 -3044
rect 5316 -3076 5320 -3044
rect 5280 -3124 5320 -3076
rect 5280 -3156 5284 -3124
rect 5316 -3156 5320 -3124
rect 5280 -3204 5320 -3156
rect 5280 -3236 5284 -3204
rect 5316 -3236 5320 -3204
rect 5280 -3284 5320 -3236
rect 5280 -3316 5284 -3284
rect 5316 -3316 5320 -3284
rect 5280 -3364 5320 -3316
rect 5280 -3396 5284 -3364
rect 5316 -3396 5320 -3364
rect 5280 -3444 5320 -3396
rect 5280 -3476 5284 -3444
rect 5316 -3476 5320 -3444
rect 5280 -3524 5320 -3476
rect 5280 -3556 5284 -3524
rect 5316 -3556 5320 -3524
rect 5280 -3604 5320 -3556
rect 5280 -3636 5284 -3604
rect 5316 -3636 5320 -3604
rect 5280 -3684 5320 -3636
rect 5280 -3716 5284 -3684
rect 5316 -3716 5320 -3684
rect 5280 -3720 5320 -3716
rect 5360 1036 5400 1040
rect 5360 1004 5364 1036
rect 5396 1004 5400 1036
rect 5360 956 5400 1004
rect 5360 924 5364 956
rect 5396 924 5400 956
rect 5360 876 5400 924
rect 5360 844 5364 876
rect 5396 844 5400 876
rect 5360 796 5400 844
rect 5360 764 5364 796
rect 5396 764 5400 796
rect 5360 716 5400 764
rect 5360 684 5364 716
rect 5396 684 5400 716
rect 5360 636 5400 684
rect 5360 604 5364 636
rect 5396 604 5400 636
rect 5360 556 5400 604
rect 5360 524 5364 556
rect 5396 524 5400 556
rect 5360 476 5400 524
rect 5360 444 5364 476
rect 5396 444 5400 476
rect 5360 396 5400 444
rect 5360 364 5364 396
rect 5396 364 5400 396
rect 5360 316 5400 364
rect 5360 284 5364 316
rect 5396 284 5400 316
rect 5360 236 5400 284
rect 5360 204 5364 236
rect 5396 204 5400 236
rect 5360 156 5400 204
rect 5360 124 5364 156
rect 5396 124 5400 156
rect 5360 76 5400 124
rect 5360 44 5364 76
rect 5396 44 5400 76
rect 5360 -4 5400 44
rect 5360 -36 5364 -4
rect 5396 -36 5400 -4
rect 5360 -84 5400 -36
rect 5360 -116 5364 -84
rect 5396 -116 5400 -84
rect 5360 -164 5400 -116
rect 5360 -196 5364 -164
rect 5396 -196 5400 -164
rect 5360 -244 5400 -196
rect 5360 -276 5364 -244
rect 5396 -276 5400 -244
rect 5360 -324 5400 -276
rect 5360 -356 5364 -324
rect 5396 -356 5400 -324
rect 5360 -404 5400 -356
rect 5360 -436 5364 -404
rect 5396 -436 5400 -404
rect 5360 -484 5400 -436
rect 5360 -516 5364 -484
rect 5396 -516 5400 -484
rect 5360 -564 5400 -516
rect 5360 -596 5364 -564
rect 5396 -596 5400 -564
rect 5360 -644 5400 -596
rect 5360 -676 5364 -644
rect 5396 -676 5400 -644
rect 5360 -724 5400 -676
rect 5360 -756 5364 -724
rect 5396 -756 5400 -724
rect 5360 -804 5400 -756
rect 5360 -836 5364 -804
rect 5396 -836 5400 -804
rect 5360 -884 5400 -836
rect 5360 -916 5364 -884
rect 5396 -916 5400 -884
rect 5360 -964 5400 -916
rect 5360 -996 5364 -964
rect 5396 -996 5400 -964
rect 5360 -1044 5400 -996
rect 5360 -1076 5364 -1044
rect 5396 -1076 5400 -1044
rect 5360 -1124 5400 -1076
rect 5360 -1156 5364 -1124
rect 5396 -1156 5400 -1124
rect 5360 -1204 5400 -1156
rect 5360 -1236 5364 -1204
rect 5396 -1236 5400 -1204
rect 5360 -1284 5400 -1236
rect 5360 -1316 5364 -1284
rect 5396 -1316 5400 -1284
rect 5360 -1364 5400 -1316
rect 5360 -1396 5364 -1364
rect 5396 -1396 5400 -1364
rect 5360 -1444 5400 -1396
rect 5360 -1476 5364 -1444
rect 5396 -1476 5400 -1444
rect 5360 -1524 5400 -1476
rect 5360 -1556 5364 -1524
rect 5396 -1556 5400 -1524
rect 5360 -1604 5400 -1556
rect 5360 -1636 5364 -1604
rect 5396 -1636 5400 -1604
rect 5360 -1684 5400 -1636
rect 5360 -1716 5364 -1684
rect 5396 -1716 5400 -1684
rect 5360 -1764 5400 -1716
rect 5360 -1796 5364 -1764
rect 5396 -1796 5400 -1764
rect 5360 -1844 5400 -1796
rect 5360 -1876 5364 -1844
rect 5396 -1876 5400 -1844
rect 5360 -1924 5400 -1876
rect 5360 -1956 5364 -1924
rect 5396 -1956 5400 -1924
rect 5360 -2004 5400 -1956
rect 5360 -2036 5364 -2004
rect 5396 -2036 5400 -2004
rect 5360 -2084 5400 -2036
rect 5360 -2116 5364 -2084
rect 5396 -2116 5400 -2084
rect 5360 -2164 5400 -2116
rect 5360 -2196 5364 -2164
rect 5396 -2196 5400 -2164
rect 5360 -2244 5400 -2196
rect 5360 -2276 5364 -2244
rect 5396 -2276 5400 -2244
rect 5360 -2324 5400 -2276
rect 5360 -2356 5364 -2324
rect 5396 -2356 5400 -2324
rect 5360 -2404 5400 -2356
rect 5360 -2436 5364 -2404
rect 5396 -2436 5400 -2404
rect 5360 -2484 5400 -2436
rect 5360 -2516 5364 -2484
rect 5396 -2516 5400 -2484
rect 5360 -2564 5400 -2516
rect 5360 -2596 5364 -2564
rect 5396 -2596 5400 -2564
rect 5360 -2644 5400 -2596
rect 5360 -2676 5364 -2644
rect 5396 -2676 5400 -2644
rect 5360 -2724 5400 -2676
rect 5360 -2756 5364 -2724
rect 5396 -2756 5400 -2724
rect 5360 -2804 5400 -2756
rect 5360 -2836 5364 -2804
rect 5396 -2836 5400 -2804
rect 5360 -2884 5400 -2836
rect 5360 -2916 5364 -2884
rect 5396 -2916 5400 -2884
rect 5360 -2964 5400 -2916
rect 5360 -2996 5364 -2964
rect 5396 -2996 5400 -2964
rect 5360 -3044 5400 -2996
rect 5360 -3076 5364 -3044
rect 5396 -3076 5400 -3044
rect 5360 -3124 5400 -3076
rect 5360 -3156 5364 -3124
rect 5396 -3156 5400 -3124
rect 5360 -3204 5400 -3156
rect 5360 -3236 5364 -3204
rect 5396 -3236 5400 -3204
rect 5360 -3284 5400 -3236
rect 5360 -3316 5364 -3284
rect 5396 -3316 5400 -3284
rect 5360 -3364 5400 -3316
rect 5360 -3396 5364 -3364
rect 5396 -3396 5400 -3364
rect 5360 -3444 5400 -3396
rect 5360 -3476 5364 -3444
rect 5396 -3476 5400 -3444
rect 5360 -3524 5400 -3476
rect 5360 -3556 5364 -3524
rect 5396 -3556 5400 -3524
rect 5360 -3604 5400 -3556
rect 5360 -3636 5364 -3604
rect 5396 -3636 5400 -3604
rect 5360 -3684 5400 -3636
rect 5360 -3716 5364 -3684
rect 5396 -3716 5400 -3684
rect 5360 -3720 5400 -3716
rect 5440 1036 5480 1040
rect 5440 1004 5444 1036
rect 5476 1004 5480 1036
rect 5440 956 5480 1004
rect 5440 924 5444 956
rect 5476 924 5480 956
rect 5440 876 5480 924
rect 5440 844 5444 876
rect 5476 844 5480 876
rect 5440 796 5480 844
rect 5440 764 5444 796
rect 5476 764 5480 796
rect 5440 716 5480 764
rect 5440 684 5444 716
rect 5476 684 5480 716
rect 5440 636 5480 684
rect 5440 604 5444 636
rect 5476 604 5480 636
rect 5440 556 5480 604
rect 5440 524 5444 556
rect 5476 524 5480 556
rect 5440 476 5480 524
rect 5440 444 5444 476
rect 5476 444 5480 476
rect 5440 396 5480 444
rect 5440 364 5444 396
rect 5476 364 5480 396
rect 5440 316 5480 364
rect 5440 284 5444 316
rect 5476 284 5480 316
rect 5440 236 5480 284
rect 5440 204 5444 236
rect 5476 204 5480 236
rect 5440 156 5480 204
rect 5440 124 5444 156
rect 5476 124 5480 156
rect 5440 76 5480 124
rect 5440 44 5444 76
rect 5476 44 5480 76
rect 5440 -4 5480 44
rect 5440 -36 5444 -4
rect 5476 -36 5480 -4
rect 5440 -84 5480 -36
rect 5440 -116 5444 -84
rect 5476 -116 5480 -84
rect 5440 -164 5480 -116
rect 5440 -196 5444 -164
rect 5476 -196 5480 -164
rect 5440 -244 5480 -196
rect 5440 -276 5444 -244
rect 5476 -276 5480 -244
rect 5440 -324 5480 -276
rect 5440 -356 5444 -324
rect 5476 -356 5480 -324
rect 5440 -404 5480 -356
rect 5440 -436 5444 -404
rect 5476 -436 5480 -404
rect 5440 -484 5480 -436
rect 5440 -516 5444 -484
rect 5476 -516 5480 -484
rect 5440 -564 5480 -516
rect 5440 -596 5444 -564
rect 5476 -596 5480 -564
rect 5440 -644 5480 -596
rect 5440 -676 5444 -644
rect 5476 -676 5480 -644
rect 5440 -724 5480 -676
rect 5440 -756 5444 -724
rect 5476 -756 5480 -724
rect 5440 -804 5480 -756
rect 5440 -836 5444 -804
rect 5476 -836 5480 -804
rect 5440 -884 5480 -836
rect 5440 -916 5444 -884
rect 5476 -916 5480 -884
rect 5440 -964 5480 -916
rect 5440 -996 5444 -964
rect 5476 -996 5480 -964
rect 5440 -1044 5480 -996
rect 5440 -1076 5444 -1044
rect 5476 -1076 5480 -1044
rect 5440 -1124 5480 -1076
rect 5440 -1156 5444 -1124
rect 5476 -1156 5480 -1124
rect 5440 -1204 5480 -1156
rect 5440 -1236 5444 -1204
rect 5476 -1236 5480 -1204
rect 5440 -1284 5480 -1236
rect 5440 -1316 5444 -1284
rect 5476 -1316 5480 -1284
rect 5440 -1364 5480 -1316
rect 5440 -1396 5444 -1364
rect 5476 -1396 5480 -1364
rect 5440 -1444 5480 -1396
rect 5440 -1476 5444 -1444
rect 5476 -1476 5480 -1444
rect 5440 -1524 5480 -1476
rect 5440 -1556 5444 -1524
rect 5476 -1556 5480 -1524
rect 5440 -1604 5480 -1556
rect 5440 -1636 5444 -1604
rect 5476 -1636 5480 -1604
rect 5440 -1684 5480 -1636
rect 5440 -1716 5444 -1684
rect 5476 -1716 5480 -1684
rect 5440 -1764 5480 -1716
rect 5440 -1796 5444 -1764
rect 5476 -1796 5480 -1764
rect 5440 -1844 5480 -1796
rect 5440 -1876 5444 -1844
rect 5476 -1876 5480 -1844
rect 5440 -1924 5480 -1876
rect 5440 -1956 5444 -1924
rect 5476 -1956 5480 -1924
rect 5440 -2004 5480 -1956
rect 5440 -2036 5444 -2004
rect 5476 -2036 5480 -2004
rect 5440 -2084 5480 -2036
rect 5440 -2116 5444 -2084
rect 5476 -2116 5480 -2084
rect 5440 -2164 5480 -2116
rect 5440 -2196 5444 -2164
rect 5476 -2196 5480 -2164
rect 5440 -2244 5480 -2196
rect 5440 -2276 5444 -2244
rect 5476 -2276 5480 -2244
rect 5440 -2324 5480 -2276
rect 5440 -2356 5444 -2324
rect 5476 -2356 5480 -2324
rect 5440 -2404 5480 -2356
rect 5440 -2436 5444 -2404
rect 5476 -2436 5480 -2404
rect 5440 -2484 5480 -2436
rect 5440 -2516 5444 -2484
rect 5476 -2516 5480 -2484
rect 5440 -2564 5480 -2516
rect 5440 -2596 5444 -2564
rect 5476 -2596 5480 -2564
rect 5440 -2644 5480 -2596
rect 5440 -2676 5444 -2644
rect 5476 -2676 5480 -2644
rect 5440 -2724 5480 -2676
rect 5440 -2756 5444 -2724
rect 5476 -2756 5480 -2724
rect 5440 -2804 5480 -2756
rect 5440 -2836 5444 -2804
rect 5476 -2836 5480 -2804
rect 5440 -2884 5480 -2836
rect 5440 -2916 5444 -2884
rect 5476 -2916 5480 -2884
rect 5440 -2964 5480 -2916
rect 5440 -2996 5444 -2964
rect 5476 -2996 5480 -2964
rect 5440 -3044 5480 -2996
rect 5440 -3076 5444 -3044
rect 5476 -3076 5480 -3044
rect 5440 -3124 5480 -3076
rect 5440 -3156 5444 -3124
rect 5476 -3156 5480 -3124
rect 5440 -3204 5480 -3156
rect 5440 -3236 5444 -3204
rect 5476 -3236 5480 -3204
rect 5440 -3284 5480 -3236
rect 5440 -3316 5444 -3284
rect 5476 -3316 5480 -3284
rect 5440 -3364 5480 -3316
rect 5440 -3396 5444 -3364
rect 5476 -3396 5480 -3364
rect 5440 -3444 5480 -3396
rect 5440 -3476 5444 -3444
rect 5476 -3476 5480 -3444
rect 5440 -3524 5480 -3476
rect 5440 -3556 5444 -3524
rect 5476 -3556 5480 -3524
rect 5440 -3604 5480 -3556
rect 5440 -3636 5444 -3604
rect 5476 -3636 5480 -3604
rect 5440 -3684 5480 -3636
rect 5440 -3716 5444 -3684
rect 5476 -3716 5480 -3684
rect 5440 -3720 5480 -3716
rect 5520 1036 5560 1040
rect 5520 1004 5524 1036
rect 5556 1004 5560 1036
rect 5520 956 5560 1004
rect 5520 924 5524 956
rect 5556 924 5560 956
rect 5520 876 5560 924
rect 5520 844 5524 876
rect 5556 844 5560 876
rect 5520 796 5560 844
rect 5520 764 5524 796
rect 5556 764 5560 796
rect 5520 716 5560 764
rect 5520 684 5524 716
rect 5556 684 5560 716
rect 5520 636 5560 684
rect 5520 604 5524 636
rect 5556 604 5560 636
rect 5520 556 5560 604
rect 5520 524 5524 556
rect 5556 524 5560 556
rect 5520 476 5560 524
rect 5520 444 5524 476
rect 5556 444 5560 476
rect 5520 396 5560 444
rect 5520 364 5524 396
rect 5556 364 5560 396
rect 5520 316 5560 364
rect 5520 284 5524 316
rect 5556 284 5560 316
rect 5520 236 5560 284
rect 5520 204 5524 236
rect 5556 204 5560 236
rect 5520 156 5560 204
rect 5520 124 5524 156
rect 5556 124 5560 156
rect 5520 76 5560 124
rect 5520 44 5524 76
rect 5556 44 5560 76
rect 5520 -4 5560 44
rect 5520 -36 5524 -4
rect 5556 -36 5560 -4
rect 5520 -84 5560 -36
rect 5520 -116 5524 -84
rect 5556 -116 5560 -84
rect 5520 -164 5560 -116
rect 5520 -196 5524 -164
rect 5556 -196 5560 -164
rect 5520 -244 5560 -196
rect 5520 -276 5524 -244
rect 5556 -276 5560 -244
rect 5520 -324 5560 -276
rect 5520 -356 5524 -324
rect 5556 -356 5560 -324
rect 5520 -404 5560 -356
rect 5520 -436 5524 -404
rect 5556 -436 5560 -404
rect 5520 -484 5560 -436
rect 5520 -516 5524 -484
rect 5556 -516 5560 -484
rect 5520 -564 5560 -516
rect 5520 -596 5524 -564
rect 5556 -596 5560 -564
rect 5520 -644 5560 -596
rect 5520 -676 5524 -644
rect 5556 -676 5560 -644
rect 5520 -724 5560 -676
rect 5520 -756 5524 -724
rect 5556 -756 5560 -724
rect 5520 -804 5560 -756
rect 5520 -836 5524 -804
rect 5556 -836 5560 -804
rect 5520 -884 5560 -836
rect 5520 -916 5524 -884
rect 5556 -916 5560 -884
rect 5520 -964 5560 -916
rect 5520 -996 5524 -964
rect 5556 -996 5560 -964
rect 5520 -1044 5560 -996
rect 5520 -1076 5524 -1044
rect 5556 -1076 5560 -1044
rect 5520 -1124 5560 -1076
rect 5520 -1156 5524 -1124
rect 5556 -1156 5560 -1124
rect 5520 -1204 5560 -1156
rect 5520 -1236 5524 -1204
rect 5556 -1236 5560 -1204
rect 5520 -1284 5560 -1236
rect 5520 -1316 5524 -1284
rect 5556 -1316 5560 -1284
rect 5520 -1364 5560 -1316
rect 5520 -1396 5524 -1364
rect 5556 -1396 5560 -1364
rect 5520 -1444 5560 -1396
rect 5520 -1476 5524 -1444
rect 5556 -1476 5560 -1444
rect 5520 -1524 5560 -1476
rect 5520 -1556 5524 -1524
rect 5556 -1556 5560 -1524
rect 5520 -1604 5560 -1556
rect 5520 -1636 5524 -1604
rect 5556 -1636 5560 -1604
rect 5520 -1684 5560 -1636
rect 5520 -1716 5524 -1684
rect 5556 -1716 5560 -1684
rect 5520 -1764 5560 -1716
rect 5520 -1796 5524 -1764
rect 5556 -1796 5560 -1764
rect 5520 -1844 5560 -1796
rect 5520 -1876 5524 -1844
rect 5556 -1876 5560 -1844
rect 5520 -1924 5560 -1876
rect 5520 -1956 5524 -1924
rect 5556 -1956 5560 -1924
rect 5520 -2004 5560 -1956
rect 5520 -2036 5524 -2004
rect 5556 -2036 5560 -2004
rect 5520 -2084 5560 -2036
rect 5520 -2116 5524 -2084
rect 5556 -2116 5560 -2084
rect 5520 -2164 5560 -2116
rect 5520 -2196 5524 -2164
rect 5556 -2196 5560 -2164
rect 5520 -2244 5560 -2196
rect 5520 -2276 5524 -2244
rect 5556 -2276 5560 -2244
rect 5520 -2324 5560 -2276
rect 5520 -2356 5524 -2324
rect 5556 -2356 5560 -2324
rect 5520 -2404 5560 -2356
rect 5520 -2436 5524 -2404
rect 5556 -2436 5560 -2404
rect 5520 -2484 5560 -2436
rect 5520 -2516 5524 -2484
rect 5556 -2516 5560 -2484
rect 5520 -2564 5560 -2516
rect 5520 -2596 5524 -2564
rect 5556 -2596 5560 -2564
rect 5520 -2644 5560 -2596
rect 5520 -2676 5524 -2644
rect 5556 -2676 5560 -2644
rect 5520 -2724 5560 -2676
rect 5520 -2756 5524 -2724
rect 5556 -2756 5560 -2724
rect 5520 -2804 5560 -2756
rect 5520 -2836 5524 -2804
rect 5556 -2836 5560 -2804
rect 5520 -2884 5560 -2836
rect 5520 -2916 5524 -2884
rect 5556 -2916 5560 -2884
rect 5520 -2964 5560 -2916
rect 5520 -2996 5524 -2964
rect 5556 -2996 5560 -2964
rect 5520 -3044 5560 -2996
rect 5520 -3076 5524 -3044
rect 5556 -3076 5560 -3044
rect 5520 -3124 5560 -3076
rect 5520 -3156 5524 -3124
rect 5556 -3156 5560 -3124
rect 5520 -3204 5560 -3156
rect 5520 -3236 5524 -3204
rect 5556 -3236 5560 -3204
rect 5520 -3284 5560 -3236
rect 5520 -3316 5524 -3284
rect 5556 -3316 5560 -3284
rect 5520 -3364 5560 -3316
rect 5520 -3396 5524 -3364
rect 5556 -3396 5560 -3364
rect 5520 -3444 5560 -3396
rect 5520 -3476 5524 -3444
rect 5556 -3476 5560 -3444
rect 5520 -3524 5560 -3476
rect 5520 -3556 5524 -3524
rect 5556 -3556 5560 -3524
rect 5520 -3604 5560 -3556
rect 5520 -3636 5524 -3604
rect 5556 -3636 5560 -3604
rect 5520 -3684 5560 -3636
rect 5520 -3716 5524 -3684
rect 5556 -3716 5560 -3684
rect 5520 -3720 5560 -3716
rect 5600 1036 5640 1040
rect 5600 1004 5604 1036
rect 5636 1004 5640 1036
rect 5600 956 5640 1004
rect 5600 924 5604 956
rect 5636 924 5640 956
rect 5600 876 5640 924
rect 5600 844 5604 876
rect 5636 844 5640 876
rect 5600 796 5640 844
rect 5600 764 5604 796
rect 5636 764 5640 796
rect 5600 716 5640 764
rect 5600 684 5604 716
rect 5636 684 5640 716
rect 5600 636 5640 684
rect 5600 604 5604 636
rect 5636 604 5640 636
rect 5600 556 5640 604
rect 5600 524 5604 556
rect 5636 524 5640 556
rect 5600 476 5640 524
rect 5600 444 5604 476
rect 5636 444 5640 476
rect 5600 396 5640 444
rect 5600 364 5604 396
rect 5636 364 5640 396
rect 5600 316 5640 364
rect 5600 284 5604 316
rect 5636 284 5640 316
rect 5600 236 5640 284
rect 5600 204 5604 236
rect 5636 204 5640 236
rect 5600 156 5640 204
rect 5600 124 5604 156
rect 5636 124 5640 156
rect 5600 76 5640 124
rect 5600 44 5604 76
rect 5636 44 5640 76
rect 5600 -4 5640 44
rect 5600 -36 5604 -4
rect 5636 -36 5640 -4
rect 5600 -84 5640 -36
rect 5600 -116 5604 -84
rect 5636 -116 5640 -84
rect 5600 -164 5640 -116
rect 5600 -196 5604 -164
rect 5636 -196 5640 -164
rect 5600 -244 5640 -196
rect 5600 -276 5604 -244
rect 5636 -276 5640 -244
rect 5600 -324 5640 -276
rect 5600 -356 5604 -324
rect 5636 -356 5640 -324
rect 5600 -404 5640 -356
rect 5600 -436 5604 -404
rect 5636 -436 5640 -404
rect 5600 -484 5640 -436
rect 5600 -516 5604 -484
rect 5636 -516 5640 -484
rect 5600 -564 5640 -516
rect 5600 -596 5604 -564
rect 5636 -596 5640 -564
rect 5600 -644 5640 -596
rect 5600 -676 5604 -644
rect 5636 -676 5640 -644
rect 5600 -724 5640 -676
rect 5600 -756 5604 -724
rect 5636 -756 5640 -724
rect 5600 -804 5640 -756
rect 5600 -836 5604 -804
rect 5636 -836 5640 -804
rect 5600 -884 5640 -836
rect 5600 -916 5604 -884
rect 5636 -916 5640 -884
rect 5600 -964 5640 -916
rect 5600 -996 5604 -964
rect 5636 -996 5640 -964
rect 5600 -1044 5640 -996
rect 5600 -1076 5604 -1044
rect 5636 -1076 5640 -1044
rect 5600 -1124 5640 -1076
rect 5600 -1156 5604 -1124
rect 5636 -1156 5640 -1124
rect 5600 -1204 5640 -1156
rect 5600 -1236 5604 -1204
rect 5636 -1236 5640 -1204
rect 5600 -1284 5640 -1236
rect 5600 -1316 5604 -1284
rect 5636 -1316 5640 -1284
rect 5600 -1364 5640 -1316
rect 5600 -1396 5604 -1364
rect 5636 -1396 5640 -1364
rect 5600 -1444 5640 -1396
rect 5600 -1476 5604 -1444
rect 5636 -1476 5640 -1444
rect 5600 -1524 5640 -1476
rect 5600 -1556 5604 -1524
rect 5636 -1556 5640 -1524
rect 5600 -1604 5640 -1556
rect 5600 -1636 5604 -1604
rect 5636 -1636 5640 -1604
rect 5600 -1684 5640 -1636
rect 5600 -1716 5604 -1684
rect 5636 -1716 5640 -1684
rect 5600 -1764 5640 -1716
rect 5600 -1796 5604 -1764
rect 5636 -1796 5640 -1764
rect 5600 -1844 5640 -1796
rect 5600 -1876 5604 -1844
rect 5636 -1876 5640 -1844
rect 5600 -1924 5640 -1876
rect 5600 -1956 5604 -1924
rect 5636 -1956 5640 -1924
rect 5600 -2004 5640 -1956
rect 5600 -2036 5604 -2004
rect 5636 -2036 5640 -2004
rect 5600 -2084 5640 -2036
rect 5600 -2116 5604 -2084
rect 5636 -2116 5640 -2084
rect 5600 -2164 5640 -2116
rect 5600 -2196 5604 -2164
rect 5636 -2196 5640 -2164
rect 5600 -2244 5640 -2196
rect 5600 -2276 5604 -2244
rect 5636 -2276 5640 -2244
rect 5600 -2324 5640 -2276
rect 5600 -2356 5604 -2324
rect 5636 -2356 5640 -2324
rect 5600 -2404 5640 -2356
rect 5600 -2436 5604 -2404
rect 5636 -2436 5640 -2404
rect 5600 -2484 5640 -2436
rect 5600 -2516 5604 -2484
rect 5636 -2516 5640 -2484
rect 5600 -2564 5640 -2516
rect 5600 -2596 5604 -2564
rect 5636 -2596 5640 -2564
rect 5600 -2644 5640 -2596
rect 5600 -2676 5604 -2644
rect 5636 -2676 5640 -2644
rect 5600 -2724 5640 -2676
rect 5600 -2756 5604 -2724
rect 5636 -2756 5640 -2724
rect 5600 -2804 5640 -2756
rect 5600 -2836 5604 -2804
rect 5636 -2836 5640 -2804
rect 5600 -2884 5640 -2836
rect 5600 -2916 5604 -2884
rect 5636 -2916 5640 -2884
rect 5600 -2964 5640 -2916
rect 5600 -2996 5604 -2964
rect 5636 -2996 5640 -2964
rect 5600 -3044 5640 -2996
rect 5600 -3076 5604 -3044
rect 5636 -3076 5640 -3044
rect 5600 -3124 5640 -3076
rect 5600 -3156 5604 -3124
rect 5636 -3156 5640 -3124
rect 5600 -3204 5640 -3156
rect 5600 -3236 5604 -3204
rect 5636 -3236 5640 -3204
rect 5600 -3284 5640 -3236
rect 5600 -3316 5604 -3284
rect 5636 -3316 5640 -3284
rect 5600 -3364 5640 -3316
rect 5600 -3396 5604 -3364
rect 5636 -3396 5640 -3364
rect 5600 -3444 5640 -3396
rect 5600 -3476 5604 -3444
rect 5636 -3476 5640 -3444
rect 5600 -3524 5640 -3476
rect 5600 -3556 5604 -3524
rect 5636 -3556 5640 -3524
rect 5600 -3604 5640 -3556
rect 5600 -3636 5604 -3604
rect 5636 -3636 5640 -3604
rect 5600 -3684 5640 -3636
rect 5600 -3716 5604 -3684
rect 5636 -3716 5640 -3684
rect 5600 -3720 5640 -3716
rect 5680 1036 5720 1040
rect 5680 1004 5684 1036
rect 5716 1004 5720 1036
rect 5680 956 5720 1004
rect 5680 924 5684 956
rect 5716 924 5720 956
rect 5680 876 5720 924
rect 5680 844 5684 876
rect 5716 844 5720 876
rect 5680 796 5720 844
rect 5680 764 5684 796
rect 5716 764 5720 796
rect 5680 716 5720 764
rect 5680 684 5684 716
rect 5716 684 5720 716
rect 5680 636 5720 684
rect 5680 604 5684 636
rect 5716 604 5720 636
rect 5680 556 5720 604
rect 5680 524 5684 556
rect 5716 524 5720 556
rect 5680 476 5720 524
rect 5680 444 5684 476
rect 5716 444 5720 476
rect 5680 396 5720 444
rect 5680 364 5684 396
rect 5716 364 5720 396
rect 5680 316 5720 364
rect 5680 284 5684 316
rect 5716 284 5720 316
rect 5680 236 5720 284
rect 5680 204 5684 236
rect 5716 204 5720 236
rect 5680 156 5720 204
rect 5680 124 5684 156
rect 5716 124 5720 156
rect 5680 76 5720 124
rect 5680 44 5684 76
rect 5716 44 5720 76
rect 5680 -4 5720 44
rect 5680 -36 5684 -4
rect 5716 -36 5720 -4
rect 5680 -84 5720 -36
rect 5680 -116 5684 -84
rect 5716 -116 5720 -84
rect 5680 -164 5720 -116
rect 5680 -196 5684 -164
rect 5716 -196 5720 -164
rect 5680 -244 5720 -196
rect 5680 -276 5684 -244
rect 5716 -276 5720 -244
rect 5680 -324 5720 -276
rect 5680 -356 5684 -324
rect 5716 -356 5720 -324
rect 5680 -404 5720 -356
rect 5680 -436 5684 -404
rect 5716 -436 5720 -404
rect 5680 -484 5720 -436
rect 5680 -516 5684 -484
rect 5716 -516 5720 -484
rect 5680 -564 5720 -516
rect 5680 -596 5684 -564
rect 5716 -596 5720 -564
rect 5680 -644 5720 -596
rect 5680 -676 5684 -644
rect 5716 -676 5720 -644
rect 5680 -724 5720 -676
rect 5680 -756 5684 -724
rect 5716 -756 5720 -724
rect 5680 -804 5720 -756
rect 5680 -836 5684 -804
rect 5716 -836 5720 -804
rect 5680 -884 5720 -836
rect 5680 -916 5684 -884
rect 5716 -916 5720 -884
rect 5680 -964 5720 -916
rect 5680 -996 5684 -964
rect 5716 -996 5720 -964
rect 5680 -1044 5720 -996
rect 5680 -1076 5684 -1044
rect 5716 -1076 5720 -1044
rect 5680 -1124 5720 -1076
rect 5680 -1156 5684 -1124
rect 5716 -1156 5720 -1124
rect 5680 -1204 5720 -1156
rect 5680 -1236 5684 -1204
rect 5716 -1236 5720 -1204
rect 5680 -1284 5720 -1236
rect 5680 -1316 5684 -1284
rect 5716 -1316 5720 -1284
rect 5680 -1364 5720 -1316
rect 5680 -1396 5684 -1364
rect 5716 -1396 5720 -1364
rect 5680 -1444 5720 -1396
rect 5680 -1476 5684 -1444
rect 5716 -1476 5720 -1444
rect 5680 -1524 5720 -1476
rect 5680 -1556 5684 -1524
rect 5716 -1556 5720 -1524
rect 5680 -1604 5720 -1556
rect 5680 -1636 5684 -1604
rect 5716 -1636 5720 -1604
rect 5680 -1684 5720 -1636
rect 5680 -1716 5684 -1684
rect 5716 -1716 5720 -1684
rect 5680 -1764 5720 -1716
rect 5680 -1796 5684 -1764
rect 5716 -1796 5720 -1764
rect 5680 -1844 5720 -1796
rect 5680 -1876 5684 -1844
rect 5716 -1876 5720 -1844
rect 5680 -1924 5720 -1876
rect 5680 -1956 5684 -1924
rect 5716 -1956 5720 -1924
rect 5680 -2004 5720 -1956
rect 5680 -2036 5684 -2004
rect 5716 -2036 5720 -2004
rect 5680 -2084 5720 -2036
rect 5680 -2116 5684 -2084
rect 5716 -2116 5720 -2084
rect 5680 -2164 5720 -2116
rect 5680 -2196 5684 -2164
rect 5716 -2196 5720 -2164
rect 5680 -2244 5720 -2196
rect 5680 -2276 5684 -2244
rect 5716 -2276 5720 -2244
rect 5680 -2324 5720 -2276
rect 5680 -2356 5684 -2324
rect 5716 -2356 5720 -2324
rect 5680 -2404 5720 -2356
rect 5680 -2436 5684 -2404
rect 5716 -2436 5720 -2404
rect 5680 -2484 5720 -2436
rect 5680 -2516 5684 -2484
rect 5716 -2516 5720 -2484
rect 5680 -2564 5720 -2516
rect 5680 -2596 5684 -2564
rect 5716 -2596 5720 -2564
rect 5680 -2644 5720 -2596
rect 5680 -2676 5684 -2644
rect 5716 -2676 5720 -2644
rect 5680 -2724 5720 -2676
rect 5680 -2756 5684 -2724
rect 5716 -2756 5720 -2724
rect 5680 -2804 5720 -2756
rect 5680 -2836 5684 -2804
rect 5716 -2836 5720 -2804
rect 5680 -2884 5720 -2836
rect 5680 -2916 5684 -2884
rect 5716 -2916 5720 -2884
rect 5680 -2964 5720 -2916
rect 5680 -2996 5684 -2964
rect 5716 -2996 5720 -2964
rect 5680 -3044 5720 -2996
rect 5680 -3076 5684 -3044
rect 5716 -3076 5720 -3044
rect 5680 -3124 5720 -3076
rect 5680 -3156 5684 -3124
rect 5716 -3156 5720 -3124
rect 5680 -3204 5720 -3156
rect 5680 -3236 5684 -3204
rect 5716 -3236 5720 -3204
rect 5680 -3284 5720 -3236
rect 5680 -3316 5684 -3284
rect 5716 -3316 5720 -3284
rect 5680 -3364 5720 -3316
rect 5680 -3396 5684 -3364
rect 5716 -3396 5720 -3364
rect 5680 -3444 5720 -3396
rect 5680 -3476 5684 -3444
rect 5716 -3476 5720 -3444
rect 5680 -3524 5720 -3476
rect 5680 -3556 5684 -3524
rect 5716 -3556 5720 -3524
rect 5680 -3604 5720 -3556
rect 5680 -3636 5684 -3604
rect 5716 -3636 5720 -3604
rect 5680 -3684 5720 -3636
rect 5680 -3716 5684 -3684
rect 5716 -3716 5720 -3684
rect 5680 -3720 5720 -3716
rect 5760 1036 5800 1040
rect 5760 1004 5764 1036
rect 5796 1004 5800 1036
rect 5760 956 5800 1004
rect 5760 924 5764 956
rect 5796 924 5800 956
rect 5760 876 5800 924
rect 5760 844 5764 876
rect 5796 844 5800 876
rect 5760 796 5800 844
rect 5760 764 5764 796
rect 5796 764 5800 796
rect 5760 716 5800 764
rect 5760 684 5764 716
rect 5796 684 5800 716
rect 5760 636 5800 684
rect 5760 604 5764 636
rect 5796 604 5800 636
rect 5760 556 5800 604
rect 5760 524 5764 556
rect 5796 524 5800 556
rect 5760 476 5800 524
rect 5760 444 5764 476
rect 5796 444 5800 476
rect 5760 396 5800 444
rect 5760 364 5764 396
rect 5796 364 5800 396
rect 5760 316 5800 364
rect 5760 284 5764 316
rect 5796 284 5800 316
rect 5760 236 5800 284
rect 5760 204 5764 236
rect 5796 204 5800 236
rect 5760 156 5800 204
rect 5760 124 5764 156
rect 5796 124 5800 156
rect 5760 76 5800 124
rect 5760 44 5764 76
rect 5796 44 5800 76
rect 5760 -4 5800 44
rect 5760 -36 5764 -4
rect 5796 -36 5800 -4
rect 5760 -84 5800 -36
rect 5760 -116 5764 -84
rect 5796 -116 5800 -84
rect 5760 -164 5800 -116
rect 5760 -196 5764 -164
rect 5796 -196 5800 -164
rect 5760 -244 5800 -196
rect 5760 -276 5764 -244
rect 5796 -276 5800 -244
rect 5760 -324 5800 -276
rect 5760 -356 5764 -324
rect 5796 -356 5800 -324
rect 5760 -404 5800 -356
rect 5760 -436 5764 -404
rect 5796 -436 5800 -404
rect 5760 -484 5800 -436
rect 5760 -516 5764 -484
rect 5796 -516 5800 -484
rect 5760 -564 5800 -516
rect 5760 -596 5764 -564
rect 5796 -596 5800 -564
rect 5760 -644 5800 -596
rect 5760 -676 5764 -644
rect 5796 -676 5800 -644
rect 5760 -724 5800 -676
rect 5760 -756 5764 -724
rect 5796 -756 5800 -724
rect 5760 -804 5800 -756
rect 5760 -836 5764 -804
rect 5796 -836 5800 -804
rect 5760 -884 5800 -836
rect 5760 -916 5764 -884
rect 5796 -916 5800 -884
rect 5760 -964 5800 -916
rect 5760 -996 5764 -964
rect 5796 -996 5800 -964
rect 5760 -1044 5800 -996
rect 5760 -1076 5764 -1044
rect 5796 -1076 5800 -1044
rect 5760 -1124 5800 -1076
rect 5760 -1156 5764 -1124
rect 5796 -1156 5800 -1124
rect 5760 -1204 5800 -1156
rect 5760 -1236 5764 -1204
rect 5796 -1236 5800 -1204
rect 5760 -1284 5800 -1236
rect 5760 -1316 5764 -1284
rect 5796 -1316 5800 -1284
rect 5760 -1364 5800 -1316
rect 5760 -1396 5764 -1364
rect 5796 -1396 5800 -1364
rect 5760 -1444 5800 -1396
rect 5760 -1476 5764 -1444
rect 5796 -1476 5800 -1444
rect 5760 -1524 5800 -1476
rect 5760 -1556 5764 -1524
rect 5796 -1556 5800 -1524
rect 5760 -1604 5800 -1556
rect 5760 -1636 5764 -1604
rect 5796 -1636 5800 -1604
rect 5760 -1684 5800 -1636
rect 5760 -1716 5764 -1684
rect 5796 -1716 5800 -1684
rect 5760 -1764 5800 -1716
rect 5760 -1796 5764 -1764
rect 5796 -1796 5800 -1764
rect 5760 -1844 5800 -1796
rect 5760 -1876 5764 -1844
rect 5796 -1876 5800 -1844
rect 5760 -1924 5800 -1876
rect 5760 -1956 5764 -1924
rect 5796 -1956 5800 -1924
rect 5760 -2004 5800 -1956
rect 5760 -2036 5764 -2004
rect 5796 -2036 5800 -2004
rect 5760 -2084 5800 -2036
rect 5760 -2116 5764 -2084
rect 5796 -2116 5800 -2084
rect 5760 -2164 5800 -2116
rect 5760 -2196 5764 -2164
rect 5796 -2196 5800 -2164
rect 5760 -2244 5800 -2196
rect 5760 -2276 5764 -2244
rect 5796 -2276 5800 -2244
rect 5760 -2324 5800 -2276
rect 5760 -2356 5764 -2324
rect 5796 -2356 5800 -2324
rect 5760 -2404 5800 -2356
rect 5760 -2436 5764 -2404
rect 5796 -2436 5800 -2404
rect 5760 -2484 5800 -2436
rect 5760 -2516 5764 -2484
rect 5796 -2516 5800 -2484
rect 5760 -2564 5800 -2516
rect 5760 -2596 5764 -2564
rect 5796 -2596 5800 -2564
rect 5760 -2644 5800 -2596
rect 5760 -2676 5764 -2644
rect 5796 -2676 5800 -2644
rect 5760 -2724 5800 -2676
rect 5760 -2756 5764 -2724
rect 5796 -2756 5800 -2724
rect 5760 -2804 5800 -2756
rect 5760 -2836 5764 -2804
rect 5796 -2836 5800 -2804
rect 5760 -2884 5800 -2836
rect 5760 -2916 5764 -2884
rect 5796 -2916 5800 -2884
rect 5760 -2964 5800 -2916
rect 5760 -2996 5764 -2964
rect 5796 -2996 5800 -2964
rect 5760 -3044 5800 -2996
rect 5760 -3076 5764 -3044
rect 5796 -3076 5800 -3044
rect 5760 -3124 5800 -3076
rect 5760 -3156 5764 -3124
rect 5796 -3156 5800 -3124
rect 5760 -3204 5800 -3156
rect 5760 -3236 5764 -3204
rect 5796 -3236 5800 -3204
rect 5760 -3284 5800 -3236
rect 5760 -3316 5764 -3284
rect 5796 -3316 5800 -3284
rect 5760 -3364 5800 -3316
rect 5760 -3396 5764 -3364
rect 5796 -3396 5800 -3364
rect 5760 -3444 5800 -3396
rect 5760 -3476 5764 -3444
rect 5796 -3476 5800 -3444
rect 5760 -3524 5800 -3476
rect 5760 -3556 5764 -3524
rect 5796 -3556 5800 -3524
rect 5760 -3604 5800 -3556
rect 5760 -3636 5764 -3604
rect 5796 -3636 5800 -3604
rect 5760 -3684 5800 -3636
rect 5760 -3716 5764 -3684
rect 5796 -3716 5800 -3684
rect 5760 -3720 5800 -3716
rect 5840 1036 5880 1040
rect 5840 1004 5844 1036
rect 5876 1004 5880 1036
rect 5840 956 5880 1004
rect 5840 924 5844 956
rect 5876 924 5880 956
rect 5840 876 5880 924
rect 5840 844 5844 876
rect 5876 844 5880 876
rect 5840 796 5880 844
rect 5840 764 5844 796
rect 5876 764 5880 796
rect 5840 716 5880 764
rect 5840 684 5844 716
rect 5876 684 5880 716
rect 5840 636 5880 684
rect 5840 604 5844 636
rect 5876 604 5880 636
rect 5840 556 5880 604
rect 5840 524 5844 556
rect 5876 524 5880 556
rect 5840 476 5880 524
rect 5840 444 5844 476
rect 5876 444 5880 476
rect 5840 396 5880 444
rect 5840 364 5844 396
rect 5876 364 5880 396
rect 5840 316 5880 364
rect 5840 284 5844 316
rect 5876 284 5880 316
rect 5840 236 5880 284
rect 5840 204 5844 236
rect 5876 204 5880 236
rect 5840 156 5880 204
rect 5840 124 5844 156
rect 5876 124 5880 156
rect 5840 76 5880 124
rect 5840 44 5844 76
rect 5876 44 5880 76
rect 5840 -4 5880 44
rect 5840 -36 5844 -4
rect 5876 -36 5880 -4
rect 5840 -84 5880 -36
rect 5840 -116 5844 -84
rect 5876 -116 5880 -84
rect 5840 -164 5880 -116
rect 5840 -196 5844 -164
rect 5876 -196 5880 -164
rect 5840 -244 5880 -196
rect 5840 -276 5844 -244
rect 5876 -276 5880 -244
rect 5840 -324 5880 -276
rect 5840 -356 5844 -324
rect 5876 -356 5880 -324
rect 5840 -404 5880 -356
rect 5840 -436 5844 -404
rect 5876 -436 5880 -404
rect 5840 -484 5880 -436
rect 5840 -516 5844 -484
rect 5876 -516 5880 -484
rect 5840 -564 5880 -516
rect 5840 -596 5844 -564
rect 5876 -596 5880 -564
rect 5840 -644 5880 -596
rect 5840 -676 5844 -644
rect 5876 -676 5880 -644
rect 5840 -724 5880 -676
rect 5840 -756 5844 -724
rect 5876 -756 5880 -724
rect 5840 -804 5880 -756
rect 5840 -836 5844 -804
rect 5876 -836 5880 -804
rect 5840 -884 5880 -836
rect 5840 -916 5844 -884
rect 5876 -916 5880 -884
rect 5840 -964 5880 -916
rect 5840 -996 5844 -964
rect 5876 -996 5880 -964
rect 5840 -1044 5880 -996
rect 5840 -1076 5844 -1044
rect 5876 -1076 5880 -1044
rect 5840 -1124 5880 -1076
rect 5840 -1156 5844 -1124
rect 5876 -1156 5880 -1124
rect 5840 -1204 5880 -1156
rect 5840 -1236 5844 -1204
rect 5876 -1236 5880 -1204
rect 5840 -1284 5880 -1236
rect 5840 -1316 5844 -1284
rect 5876 -1316 5880 -1284
rect 5840 -1364 5880 -1316
rect 5840 -1396 5844 -1364
rect 5876 -1396 5880 -1364
rect 5840 -1444 5880 -1396
rect 5840 -1476 5844 -1444
rect 5876 -1476 5880 -1444
rect 5840 -1524 5880 -1476
rect 5840 -1556 5844 -1524
rect 5876 -1556 5880 -1524
rect 5840 -1604 5880 -1556
rect 5840 -1636 5844 -1604
rect 5876 -1636 5880 -1604
rect 5840 -1684 5880 -1636
rect 5840 -1716 5844 -1684
rect 5876 -1716 5880 -1684
rect 5840 -1764 5880 -1716
rect 5840 -1796 5844 -1764
rect 5876 -1796 5880 -1764
rect 5840 -1844 5880 -1796
rect 5840 -1876 5844 -1844
rect 5876 -1876 5880 -1844
rect 5840 -1924 5880 -1876
rect 5840 -1956 5844 -1924
rect 5876 -1956 5880 -1924
rect 5840 -2004 5880 -1956
rect 5840 -2036 5844 -2004
rect 5876 -2036 5880 -2004
rect 5840 -2084 5880 -2036
rect 5840 -2116 5844 -2084
rect 5876 -2116 5880 -2084
rect 5840 -2164 5880 -2116
rect 5840 -2196 5844 -2164
rect 5876 -2196 5880 -2164
rect 5840 -2244 5880 -2196
rect 5840 -2276 5844 -2244
rect 5876 -2276 5880 -2244
rect 5840 -2324 5880 -2276
rect 5840 -2356 5844 -2324
rect 5876 -2356 5880 -2324
rect 5840 -2404 5880 -2356
rect 5840 -2436 5844 -2404
rect 5876 -2436 5880 -2404
rect 5840 -2484 5880 -2436
rect 5840 -2516 5844 -2484
rect 5876 -2516 5880 -2484
rect 5840 -2564 5880 -2516
rect 5840 -2596 5844 -2564
rect 5876 -2596 5880 -2564
rect 5840 -2644 5880 -2596
rect 5840 -2676 5844 -2644
rect 5876 -2676 5880 -2644
rect 5840 -2724 5880 -2676
rect 5840 -2756 5844 -2724
rect 5876 -2756 5880 -2724
rect 5840 -2804 5880 -2756
rect 5840 -2836 5844 -2804
rect 5876 -2836 5880 -2804
rect 5840 -2884 5880 -2836
rect 5840 -2916 5844 -2884
rect 5876 -2916 5880 -2884
rect 5840 -2964 5880 -2916
rect 5840 -2996 5844 -2964
rect 5876 -2996 5880 -2964
rect 5840 -3044 5880 -2996
rect 5840 -3076 5844 -3044
rect 5876 -3076 5880 -3044
rect 5840 -3124 5880 -3076
rect 5840 -3156 5844 -3124
rect 5876 -3156 5880 -3124
rect 5840 -3204 5880 -3156
rect 5840 -3236 5844 -3204
rect 5876 -3236 5880 -3204
rect 5840 -3284 5880 -3236
rect 5840 -3316 5844 -3284
rect 5876 -3316 5880 -3284
rect 5840 -3364 5880 -3316
rect 5840 -3396 5844 -3364
rect 5876 -3396 5880 -3364
rect 5840 -3444 5880 -3396
rect 5840 -3476 5844 -3444
rect 5876 -3476 5880 -3444
rect 5840 -3524 5880 -3476
rect 5840 -3556 5844 -3524
rect 5876 -3556 5880 -3524
rect 5840 -3604 5880 -3556
rect 5840 -3636 5844 -3604
rect 5876 -3636 5880 -3604
rect 5840 -3684 5880 -3636
rect 5840 -3716 5844 -3684
rect 5876 -3716 5880 -3684
rect 5840 -3720 5880 -3716
rect 5920 1036 5960 1040
rect 5920 1004 5924 1036
rect 5956 1004 5960 1036
rect 5920 956 5960 1004
rect 5920 924 5924 956
rect 5956 924 5960 956
rect 5920 876 5960 924
rect 5920 844 5924 876
rect 5956 844 5960 876
rect 5920 796 5960 844
rect 5920 764 5924 796
rect 5956 764 5960 796
rect 5920 716 5960 764
rect 5920 684 5924 716
rect 5956 684 5960 716
rect 5920 636 5960 684
rect 5920 604 5924 636
rect 5956 604 5960 636
rect 5920 556 5960 604
rect 5920 524 5924 556
rect 5956 524 5960 556
rect 5920 476 5960 524
rect 5920 444 5924 476
rect 5956 444 5960 476
rect 5920 396 5960 444
rect 5920 364 5924 396
rect 5956 364 5960 396
rect 5920 316 5960 364
rect 5920 284 5924 316
rect 5956 284 5960 316
rect 5920 236 5960 284
rect 5920 204 5924 236
rect 5956 204 5960 236
rect 5920 156 5960 204
rect 5920 124 5924 156
rect 5956 124 5960 156
rect 5920 76 5960 124
rect 5920 44 5924 76
rect 5956 44 5960 76
rect 5920 -4 5960 44
rect 5920 -36 5924 -4
rect 5956 -36 5960 -4
rect 5920 -84 5960 -36
rect 5920 -116 5924 -84
rect 5956 -116 5960 -84
rect 5920 -164 5960 -116
rect 5920 -196 5924 -164
rect 5956 -196 5960 -164
rect 5920 -244 5960 -196
rect 5920 -276 5924 -244
rect 5956 -276 5960 -244
rect 5920 -324 5960 -276
rect 5920 -356 5924 -324
rect 5956 -356 5960 -324
rect 5920 -404 5960 -356
rect 5920 -436 5924 -404
rect 5956 -436 5960 -404
rect 5920 -484 5960 -436
rect 5920 -516 5924 -484
rect 5956 -516 5960 -484
rect 5920 -564 5960 -516
rect 5920 -596 5924 -564
rect 5956 -596 5960 -564
rect 5920 -644 5960 -596
rect 5920 -676 5924 -644
rect 5956 -676 5960 -644
rect 5920 -724 5960 -676
rect 5920 -756 5924 -724
rect 5956 -756 5960 -724
rect 5920 -804 5960 -756
rect 5920 -836 5924 -804
rect 5956 -836 5960 -804
rect 5920 -884 5960 -836
rect 5920 -916 5924 -884
rect 5956 -916 5960 -884
rect 5920 -964 5960 -916
rect 5920 -996 5924 -964
rect 5956 -996 5960 -964
rect 5920 -1044 5960 -996
rect 5920 -1076 5924 -1044
rect 5956 -1076 5960 -1044
rect 5920 -1124 5960 -1076
rect 5920 -1156 5924 -1124
rect 5956 -1156 5960 -1124
rect 5920 -1204 5960 -1156
rect 5920 -1236 5924 -1204
rect 5956 -1236 5960 -1204
rect 5920 -1284 5960 -1236
rect 5920 -1316 5924 -1284
rect 5956 -1316 5960 -1284
rect 5920 -1364 5960 -1316
rect 5920 -1396 5924 -1364
rect 5956 -1396 5960 -1364
rect 5920 -1444 5960 -1396
rect 5920 -1476 5924 -1444
rect 5956 -1476 5960 -1444
rect 5920 -1524 5960 -1476
rect 5920 -1556 5924 -1524
rect 5956 -1556 5960 -1524
rect 5920 -1604 5960 -1556
rect 5920 -1636 5924 -1604
rect 5956 -1636 5960 -1604
rect 5920 -1684 5960 -1636
rect 5920 -1716 5924 -1684
rect 5956 -1716 5960 -1684
rect 5920 -1764 5960 -1716
rect 5920 -1796 5924 -1764
rect 5956 -1796 5960 -1764
rect 5920 -1844 5960 -1796
rect 5920 -1876 5924 -1844
rect 5956 -1876 5960 -1844
rect 5920 -1924 5960 -1876
rect 5920 -1956 5924 -1924
rect 5956 -1956 5960 -1924
rect 5920 -2004 5960 -1956
rect 5920 -2036 5924 -2004
rect 5956 -2036 5960 -2004
rect 5920 -2084 5960 -2036
rect 5920 -2116 5924 -2084
rect 5956 -2116 5960 -2084
rect 5920 -2164 5960 -2116
rect 5920 -2196 5924 -2164
rect 5956 -2196 5960 -2164
rect 5920 -2244 5960 -2196
rect 5920 -2276 5924 -2244
rect 5956 -2276 5960 -2244
rect 5920 -2324 5960 -2276
rect 5920 -2356 5924 -2324
rect 5956 -2356 5960 -2324
rect 5920 -2404 5960 -2356
rect 5920 -2436 5924 -2404
rect 5956 -2436 5960 -2404
rect 5920 -2484 5960 -2436
rect 5920 -2516 5924 -2484
rect 5956 -2516 5960 -2484
rect 5920 -2564 5960 -2516
rect 5920 -2596 5924 -2564
rect 5956 -2596 5960 -2564
rect 5920 -2644 5960 -2596
rect 5920 -2676 5924 -2644
rect 5956 -2676 5960 -2644
rect 5920 -2724 5960 -2676
rect 5920 -2756 5924 -2724
rect 5956 -2756 5960 -2724
rect 5920 -2804 5960 -2756
rect 5920 -2836 5924 -2804
rect 5956 -2836 5960 -2804
rect 5920 -2884 5960 -2836
rect 5920 -2916 5924 -2884
rect 5956 -2916 5960 -2884
rect 5920 -2964 5960 -2916
rect 5920 -2996 5924 -2964
rect 5956 -2996 5960 -2964
rect 5920 -3044 5960 -2996
rect 5920 -3076 5924 -3044
rect 5956 -3076 5960 -3044
rect 5920 -3124 5960 -3076
rect 5920 -3156 5924 -3124
rect 5956 -3156 5960 -3124
rect 5920 -3204 5960 -3156
rect 5920 -3236 5924 -3204
rect 5956 -3236 5960 -3204
rect 5920 -3284 5960 -3236
rect 5920 -3316 5924 -3284
rect 5956 -3316 5960 -3284
rect 5920 -3364 5960 -3316
rect 5920 -3396 5924 -3364
rect 5956 -3396 5960 -3364
rect 5920 -3444 5960 -3396
rect 5920 -3476 5924 -3444
rect 5956 -3476 5960 -3444
rect 5920 -3524 5960 -3476
rect 5920 -3556 5924 -3524
rect 5956 -3556 5960 -3524
rect 5920 -3604 5960 -3556
rect 5920 -3636 5924 -3604
rect 5956 -3636 5960 -3604
rect 5920 -3684 5960 -3636
rect 5920 -3716 5924 -3684
rect 5956 -3716 5960 -3684
rect 5920 -3720 5960 -3716
rect 6000 1036 6040 1040
rect 6000 1004 6004 1036
rect 6036 1004 6040 1036
rect 6000 956 6040 1004
rect 6000 924 6004 956
rect 6036 924 6040 956
rect 6000 876 6040 924
rect 6000 844 6004 876
rect 6036 844 6040 876
rect 6000 796 6040 844
rect 6000 764 6004 796
rect 6036 764 6040 796
rect 6000 716 6040 764
rect 6000 684 6004 716
rect 6036 684 6040 716
rect 6000 636 6040 684
rect 6000 604 6004 636
rect 6036 604 6040 636
rect 6000 556 6040 604
rect 6000 524 6004 556
rect 6036 524 6040 556
rect 6000 476 6040 524
rect 6000 444 6004 476
rect 6036 444 6040 476
rect 6000 396 6040 444
rect 6000 364 6004 396
rect 6036 364 6040 396
rect 6000 316 6040 364
rect 6000 284 6004 316
rect 6036 284 6040 316
rect 6000 236 6040 284
rect 6000 204 6004 236
rect 6036 204 6040 236
rect 6000 156 6040 204
rect 6000 124 6004 156
rect 6036 124 6040 156
rect 6000 76 6040 124
rect 6000 44 6004 76
rect 6036 44 6040 76
rect 6000 -4 6040 44
rect 6000 -36 6004 -4
rect 6036 -36 6040 -4
rect 6000 -84 6040 -36
rect 6000 -116 6004 -84
rect 6036 -116 6040 -84
rect 6000 -164 6040 -116
rect 6000 -196 6004 -164
rect 6036 -196 6040 -164
rect 6000 -244 6040 -196
rect 6000 -276 6004 -244
rect 6036 -276 6040 -244
rect 6000 -324 6040 -276
rect 6000 -356 6004 -324
rect 6036 -356 6040 -324
rect 6000 -404 6040 -356
rect 6000 -436 6004 -404
rect 6036 -436 6040 -404
rect 6000 -484 6040 -436
rect 6000 -516 6004 -484
rect 6036 -516 6040 -484
rect 6000 -564 6040 -516
rect 6000 -596 6004 -564
rect 6036 -596 6040 -564
rect 6000 -644 6040 -596
rect 6000 -676 6004 -644
rect 6036 -676 6040 -644
rect 6000 -724 6040 -676
rect 6000 -756 6004 -724
rect 6036 -756 6040 -724
rect 6000 -804 6040 -756
rect 6000 -836 6004 -804
rect 6036 -836 6040 -804
rect 6000 -884 6040 -836
rect 6000 -916 6004 -884
rect 6036 -916 6040 -884
rect 6000 -964 6040 -916
rect 6000 -996 6004 -964
rect 6036 -996 6040 -964
rect 6000 -1044 6040 -996
rect 6000 -1076 6004 -1044
rect 6036 -1076 6040 -1044
rect 6000 -1124 6040 -1076
rect 6000 -1156 6004 -1124
rect 6036 -1156 6040 -1124
rect 6000 -1204 6040 -1156
rect 6000 -1236 6004 -1204
rect 6036 -1236 6040 -1204
rect 6000 -1284 6040 -1236
rect 6000 -1316 6004 -1284
rect 6036 -1316 6040 -1284
rect 6000 -1364 6040 -1316
rect 6000 -1396 6004 -1364
rect 6036 -1396 6040 -1364
rect 6000 -1444 6040 -1396
rect 6000 -1476 6004 -1444
rect 6036 -1476 6040 -1444
rect 6000 -1524 6040 -1476
rect 6000 -1556 6004 -1524
rect 6036 -1556 6040 -1524
rect 6000 -1604 6040 -1556
rect 6000 -1636 6004 -1604
rect 6036 -1636 6040 -1604
rect 6000 -1684 6040 -1636
rect 6000 -1716 6004 -1684
rect 6036 -1716 6040 -1684
rect 6000 -1764 6040 -1716
rect 6000 -1796 6004 -1764
rect 6036 -1796 6040 -1764
rect 6000 -1844 6040 -1796
rect 6000 -1876 6004 -1844
rect 6036 -1876 6040 -1844
rect 6000 -1924 6040 -1876
rect 6000 -1956 6004 -1924
rect 6036 -1956 6040 -1924
rect 6000 -2004 6040 -1956
rect 6000 -2036 6004 -2004
rect 6036 -2036 6040 -2004
rect 6000 -2084 6040 -2036
rect 6000 -2116 6004 -2084
rect 6036 -2116 6040 -2084
rect 6000 -2164 6040 -2116
rect 6000 -2196 6004 -2164
rect 6036 -2196 6040 -2164
rect 6000 -2244 6040 -2196
rect 6000 -2276 6004 -2244
rect 6036 -2276 6040 -2244
rect 6000 -2324 6040 -2276
rect 6000 -2356 6004 -2324
rect 6036 -2356 6040 -2324
rect 6000 -2404 6040 -2356
rect 6000 -2436 6004 -2404
rect 6036 -2436 6040 -2404
rect 6000 -2484 6040 -2436
rect 6000 -2516 6004 -2484
rect 6036 -2516 6040 -2484
rect 6000 -2564 6040 -2516
rect 6000 -2596 6004 -2564
rect 6036 -2596 6040 -2564
rect 6000 -2644 6040 -2596
rect 6000 -2676 6004 -2644
rect 6036 -2676 6040 -2644
rect 6000 -2724 6040 -2676
rect 6000 -2756 6004 -2724
rect 6036 -2756 6040 -2724
rect 6000 -2804 6040 -2756
rect 6000 -2836 6004 -2804
rect 6036 -2836 6040 -2804
rect 6000 -2884 6040 -2836
rect 6000 -2916 6004 -2884
rect 6036 -2916 6040 -2884
rect 6000 -2964 6040 -2916
rect 6000 -2996 6004 -2964
rect 6036 -2996 6040 -2964
rect 6000 -3044 6040 -2996
rect 6000 -3076 6004 -3044
rect 6036 -3076 6040 -3044
rect 6000 -3124 6040 -3076
rect 6000 -3156 6004 -3124
rect 6036 -3156 6040 -3124
rect 6000 -3204 6040 -3156
rect 6000 -3236 6004 -3204
rect 6036 -3236 6040 -3204
rect 6000 -3284 6040 -3236
rect 6000 -3316 6004 -3284
rect 6036 -3316 6040 -3284
rect 6000 -3364 6040 -3316
rect 6000 -3396 6004 -3364
rect 6036 -3396 6040 -3364
rect 6000 -3444 6040 -3396
rect 6000 -3476 6004 -3444
rect 6036 -3476 6040 -3444
rect 6000 -3524 6040 -3476
rect 6000 -3556 6004 -3524
rect 6036 -3556 6040 -3524
rect 6000 -3604 6040 -3556
rect 6000 -3636 6004 -3604
rect 6036 -3636 6040 -3604
rect 6000 -3684 6040 -3636
rect 6000 -3716 6004 -3684
rect 6036 -3716 6040 -3684
rect 6000 -3720 6040 -3716
rect 6080 1036 6120 1040
rect 6080 1004 6084 1036
rect 6116 1004 6120 1036
rect 6080 956 6120 1004
rect 6080 924 6084 956
rect 6116 924 6120 956
rect 6080 876 6120 924
rect 6080 844 6084 876
rect 6116 844 6120 876
rect 6080 796 6120 844
rect 6080 764 6084 796
rect 6116 764 6120 796
rect 6080 716 6120 764
rect 6080 684 6084 716
rect 6116 684 6120 716
rect 6080 636 6120 684
rect 6080 604 6084 636
rect 6116 604 6120 636
rect 6080 556 6120 604
rect 6080 524 6084 556
rect 6116 524 6120 556
rect 6080 476 6120 524
rect 6080 444 6084 476
rect 6116 444 6120 476
rect 6080 396 6120 444
rect 6080 364 6084 396
rect 6116 364 6120 396
rect 6080 316 6120 364
rect 6080 284 6084 316
rect 6116 284 6120 316
rect 6080 236 6120 284
rect 6080 204 6084 236
rect 6116 204 6120 236
rect 6080 156 6120 204
rect 6080 124 6084 156
rect 6116 124 6120 156
rect 6080 76 6120 124
rect 6080 44 6084 76
rect 6116 44 6120 76
rect 6080 -4 6120 44
rect 6080 -36 6084 -4
rect 6116 -36 6120 -4
rect 6080 -84 6120 -36
rect 6080 -116 6084 -84
rect 6116 -116 6120 -84
rect 6080 -164 6120 -116
rect 6080 -196 6084 -164
rect 6116 -196 6120 -164
rect 6080 -244 6120 -196
rect 6080 -276 6084 -244
rect 6116 -276 6120 -244
rect 6080 -324 6120 -276
rect 6080 -356 6084 -324
rect 6116 -356 6120 -324
rect 6080 -404 6120 -356
rect 6080 -436 6084 -404
rect 6116 -436 6120 -404
rect 6080 -484 6120 -436
rect 6080 -516 6084 -484
rect 6116 -516 6120 -484
rect 6080 -564 6120 -516
rect 6080 -596 6084 -564
rect 6116 -596 6120 -564
rect 6080 -644 6120 -596
rect 6080 -676 6084 -644
rect 6116 -676 6120 -644
rect 6080 -724 6120 -676
rect 6080 -756 6084 -724
rect 6116 -756 6120 -724
rect 6080 -804 6120 -756
rect 6080 -836 6084 -804
rect 6116 -836 6120 -804
rect 6080 -884 6120 -836
rect 6080 -916 6084 -884
rect 6116 -916 6120 -884
rect 6080 -964 6120 -916
rect 6080 -996 6084 -964
rect 6116 -996 6120 -964
rect 6080 -1044 6120 -996
rect 6080 -1076 6084 -1044
rect 6116 -1076 6120 -1044
rect 6080 -1124 6120 -1076
rect 6080 -1156 6084 -1124
rect 6116 -1156 6120 -1124
rect 6080 -1204 6120 -1156
rect 6080 -1236 6084 -1204
rect 6116 -1236 6120 -1204
rect 6080 -1284 6120 -1236
rect 6080 -1316 6084 -1284
rect 6116 -1316 6120 -1284
rect 6080 -1364 6120 -1316
rect 6080 -1396 6084 -1364
rect 6116 -1396 6120 -1364
rect 6080 -1444 6120 -1396
rect 6080 -1476 6084 -1444
rect 6116 -1476 6120 -1444
rect 6080 -1524 6120 -1476
rect 6080 -1556 6084 -1524
rect 6116 -1556 6120 -1524
rect 6080 -1604 6120 -1556
rect 6080 -1636 6084 -1604
rect 6116 -1636 6120 -1604
rect 6080 -1684 6120 -1636
rect 6080 -1716 6084 -1684
rect 6116 -1716 6120 -1684
rect 6080 -1764 6120 -1716
rect 6080 -1796 6084 -1764
rect 6116 -1796 6120 -1764
rect 6080 -1844 6120 -1796
rect 6080 -1876 6084 -1844
rect 6116 -1876 6120 -1844
rect 6080 -1924 6120 -1876
rect 6080 -1956 6084 -1924
rect 6116 -1956 6120 -1924
rect 6080 -2004 6120 -1956
rect 6080 -2036 6084 -2004
rect 6116 -2036 6120 -2004
rect 6080 -2084 6120 -2036
rect 6080 -2116 6084 -2084
rect 6116 -2116 6120 -2084
rect 6080 -2164 6120 -2116
rect 6080 -2196 6084 -2164
rect 6116 -2196 6120 -2164
rect 6080 -2244 6120 -2196
rect 6080 -2276 6084 -2244
rect 6116 -2276 6120 -2244
rect 6080 -2324 6120 -2276
rect 6080 -2356 6084 -2324
rect 6116 -2356 6120 -2324
rect 6080 -2404 6120 -2356
rect 6080 -2436 6084 -2404
rect 6116 -2436 6120 -2404
rect 6080 -2484 6120 -2436
rect 6080 -2516 6084 -2484
rect 6116 -2516 6120 -2484
rect 6080 -2564 6120 -2516
rect 6080 -2596 6084 -2564
rect 6116 -2596 6120 -2564
rect 6080 -2644 6120 -2596
rect 6080 -2676 6084 -2644
rect 6116 -2676 6120 -2644
rect 6080 -2724 6120 -2676
rect 6080 -2756 6084 -2724
rect 6116 -2756 6120 -2724
rect 6080 -2804 6120 -2756
rect 6080 -2836 6084 -2804
rect 6116 -2836 6120 -2804
rect 6080 -2884 6120 -2836
rect 6080 -2916 6084 -2884
rect 6116 -2916 6120 -2884
rect 6080 -2964 6120 -2916
rect 6080 -2996 6084 -2964
rect 6116 -2996 6120 -2964
rect 6080 -3044 6120 -2996
rect 6080 -3076 6084 -3044
rect 6116 -3076 6120 -3044
rect 6080 -3124 6120 -3076
rect 6080 -3156 6084 -3124
rect 6116 -3156 6120 -3124
rect 6080 -3204 6120 -3156
rect 6080 -3236 6084 -3204
rect 6116 -3236 6120 -3204
rect 6080 -3284 6120 -3236
rect 6080 -3316 6084 -3284
rect 6116 -3316 6120 -3284
rect 6080 -3364 6120 -3316
rect 6080 -3396 6084 -3364
rect 6116 -3396 6120 -3364
rect 6080 -3444 6120 -3396
rect 6080 -3476 6084 -3444
rect 6116 -3476 6120 -3444
rect 6080 -3524 6120 -3476
rect 6080 -3556 6084 -3524
rect 6116 -3556 6120 -3524
rect 6080 -3604 6120 -3556
rect 6080 -3636 6084 -3604
rect 6116 -3636 6120 -3604
rect 6080 -3684 6120 -3636
rect 6080 -3716 6084 -3684
rect 6116 -3716 6120 -3684
rect 6080 -3720 6120 -3716
rect 6160 1036 6200 1040
rect 6160 1004 6164 1036
rect 6196 1004 6200 1036
rect 6160 956 6200 1004
rect 6160 924 6164 956
rect 6196 924 6200 956
rect 6160 876 6200 924
rect 6160 844 6164 876
rect 6196 844 6200 876
rect 6160 796 6200 844
rect 6160 764 6164 796
rect 6196 764 6200 796
rect 6160 716 6200 764
rect 6160 684 6164 716
rect 6196 684 6200 716
rect 6160 636 6200 684
rect 6160 604 6164 636
rect 6196 604 6200 636
rect 6160 556 6200 604
rect 6160 524 6164 556
rect 6196 524 6200 556
rect 6160 476 6200 524
rect 6160 444 6164 476
rect 6196 444 6200 476
rect 6160 396 6200 444
rect 6160 364 6164 396
rect 6196 364 6200 396
rect 6160 316 6200 364
rect 6160 284 6164 316
rect 6196 284 6200 316
rect 6160 236 6200 284
rect 6160 204 6164 236
rect 6196 204 6200 236
rect 6160 156 6200 204
rect 6160 124 6164 156
rect 6196 124 6200 156
rect 6160 76 6200 124
rect 6160 44 6164 76
rect 6196 44 6200 76
rect 6160 -4 6200 44
rect 6160 -36 6164 -4
rect 6196 -36 6200 -4
rect 6160 -84 6200 -36
rect 6160 -116 6164 -84
rect 6196 -116 6200 -84
rect 6160 -164 6200 -116
rect 6160 -196 6164 -164
rect 6196 -196 6200 -164
rect 6160 -244 6200 -196
rect 6160 -276 6164 -244
rect 6196 -276 6200 -244
rect 6160 -324 6200 -276
rect 6160 -356 6164 -324
rect 6196 -356 6200 -324
rect 6160 -404 6200 -356
rect 6160 -436 6164 -404
rect 6196 -436 6200 -404
rect 6160 -484 6200 -436
rect 6160 -516 6164 -484
rect 6196 -516 6200 -484
rect 6160 -564 6200 -516
rect 6160 -596 6164 -564
rect 6196 -596 6200 -564
rect 6160 -644 6200 -596
rect 6160 -676 6164 -644
rect 6196 -676 6200 -644
rect 6160 -724 6200 -676
rect 6160 -756 6164 -724
rect 6196 -756 6200 -724
rect 6160 -804 6200 -756
rect 6160 -836 6164 -804
rect 6196 -836 6200 -804
rect 6160 -884 6200 -836
rect 6160 -916 6164 -884
rect 6196 -916 6200 -884
rect 6160 -964 6200 -916
rect 6160 -996 6164 -964
rect 6196 -996 6200 -964
rect 6160 -1044 6200 -996
rect 6160 -1076 6164 -1044
rect 6196 -1076 6200 -1044
rect 6160 -1124 6200 -1076
rect 6160 -1156 6164 -1124
rect 6196 -1156 6200 -1124
rect 6160 -1204 6200 -1156
rect 6160 -1236 6164 -1204
rect 6196 -1236 6200 -1204
rect 6160 -1284 6200 -1236
rect 6160 -1316 6164 -1284
rect 6196 -1316 6200 -1284
rect 6160 -1364 6200 -1316
rect 6160 -1396 6164 -1364
rect 6196 -1396 6200 -1364
rect 6160 -1444 6200 -1396
rect 6160 -1476 6164 -1444
rect 6196 -1476 6200 -1444
rect 6160 -1524 6200 -1476
rect 6160 -1556 6164 -1524
rect 6196 -1556 6200 -1524
rect 6160 -1604 6200 -1556
rect 6160 -1636 6164 -1604
rect 6196 -1636 6200 -1604
rect 6160 -1684 6200 -1636
rect 6160 -1716 6164 -1684
rect 6196 -1716 6200 -1684
rect 6160 -1764 6200 -1716
rect 6160 -1796 6164 -1764
rect 6196 -1796 6200 -1764
rect 6160 -1844 6200 -1796
rect 6160 -1876 6164 -1844
rect 6196 -1876 6200 -1844
rect 6160 -1924 6200 -1876
rect 6160 -1956 6164 -1924
rect 6196 -1956 6200 -1924
rect 6160 -2004 6200 -1956
rect 6160 -2036 6164 -2004
rect 6196 -2036 6200 -2004
rect 6160 -2084 6200 -2036
rect 6160 -2116 6164 -2084
rect 6196 -2116 6200 -2084
rect 6160 -2164 6200 -2116
rect 6160 -2196 6164 -2164
rect 6196 -2196 6200 -2164
rect 6160 -2244 6200 -2196
rect 6160 -2276 6164 -2244
rect 6196 -2276 6200 -2244
rect 6160 -2324 6200 -2276
rect 6160 -2356 6164 -2324
rect 6196 -2356 6200 -2324
rect 6160 -2404 6200 -2356
rect 6160 -2436 6164 -2404
rect 6196 -2436 6200 -2404
rect 6160 -2484 6200 -2436
rect 6160 -2516 6164 -2484
rect 6196 -2516 6200 -2484
rect 6160 -2564 6200 -2516
rect 6160 -2596 6164 -2564
rect 6196 -2596 6200 -2564
rect 6160 -2644 6200 -2596
rect 6160 -2676 6164 -2644
rect 6196 -2676 6200 -2644
rect 6160 -2724 6200 -2676
rect 6160 -2756 6164 -2724
rect 6196 -2756 6200 -2724
rect 6160 -2804 6200 -2756
rect 6160 -2836 6164 -2804
rect 6196 -2836 6200 -2804
rect 6160 -2884 6200 -2836
rect 6160 -2916 6164 -2884
rect 6196 -2916 6200 -2884
rect 6160 -2964 6200 -2916
rect 6160 -2996 6164 -2964
rect 6196 -2996 6200 -2964
rect 6160 -3044 6200 -2996
rect 6160 -3076 6164 -3044
rect 6196 -3076 6200 -3044
rect 6160 -3124 6200 -3076
rect 6160 -3156 6164 -3124
rect 6196 -3156 6200 -3124
rect 6160 -3204 6200 -3156
rect 6160 -3236 6164 -3204
rect 6196 -3236 6200 -3204
rect 6160 -3284 6200 -3236
rect 6160 -3316 6164 -3284
rect 6196 -3316 6200 -3284
rect 6160 -3364 6200 -3316
rect 6160 -3396 6164 -3364
rect 6196 -3396 6200 -3364
rect 6160 -3444 6200 -3396
rect 6160 -3476 6164 -3444
rect 6196 -3476 6200 -3444
rect 6160 -3524 6200 -3476
rect 6160 -3556 6164 -3524
rect 6196 -3556 6200 -3524
rect 6160 -3604 6200 -3556
rect 6160 -3636 6164 -3604
rect 6196 -3636 6200 -3604
rect 6160 -3684 6200 -3636
rect 6160 -3716 6164 -3684
rect 6196 -3716 6200 -3684
rect 6160 -3720 6200 -3716
rect 6240 1036 6280 1040
rect 6240 1004 6244 1036
rect 6276 1004 6280 1036
rect 6240 956 6280 1004
rect 6240 924 6244 956
rect 6276 924 6280 956
rect 6240 876 6280 924
rect 6240 844 6244 876
rect 6276 844 6280 876
rect 6240 796 6280 844
rect 6240 764 6244 796
rect 6276 764 6280 796
rect 6240 716 6280 764
rect 6240 684 6244 716
rect 6276 684 6280 716
rect 6240 636 6280 684
rect 6240 604 6244 636
rect 6276 604 6280 636
rect 6240 556 6280 604
rect 6240 524 6244 556
rect 6276 524 6280 556
rect 6240 476 6280 524
rect 6240 444 6244 476
rect 6276 444 6280 476
rect 6240 396 6280 444
rect 6240 364 6244 396
rect 6276 364 6280 396
rect 6240 316 6280 364
rect 6240 284 6244 316
rect 6276 284 6280 316
rect 6240 236 6280 284
rect 6240 204 6244 236
rect 6276 204 6280 236
rect 6240 156 6280 204
rect 6240 124 6244 156
rect 6276 124 6280 156
rect 6240 76 6280 124
rect 6240 44 6244 76
rect 6276 44 6280 76
rect 6240 -4 6280 44
rect 6240 -36 6244 -4
rect 6276 -36 6280 -4
rect 6240 -84 6280 -36
rect 6240 -116 6244 -84
rect 6276 -116 6280 -84
rect 6240 -164 6280 -116
rect 6240 -196 6244 -164
rect 6276 -196 6280 -164
rect 6240 -244 6280 -196
rect 6240 -276 6244 -244
rect 6276 -276 6280 -244
rect 6240 -324 6280 -276
rect 6240 -356 6244 -324
rect 6276 -356 6280 -324
rect 6240 -404 6280 -356
rect 6240 -436 6244 -404
rect 6276 -436 6280 -404
rect 6240 -484 6280 -436
rect 6240 -516 6244 -484
rect 6276 -516 6280 -484
rect 6240 -564 6280 -516
rect 6240 -596 6244 -564
rect 6276 -596 6280 -564
rect 6240 -644 6280 -596
rect 6240 -676 6244 -644
rect 6276 -676 6280 -644
rect 6240 -724 6280 -676
rect 6240 -756 6244 -724
rect 6276 -756 6280 -724
rect 6240 -804 6280 -756
rect 6240 -836 6244 -804
rect 6276 -836 6280 -804
rect 6240 -884 6280 -836
rect 6240 -916 6244 -884
rect 6276 -916 6280 -884
rect 6240 -964 6280 -916
rect 6240 -996 6244 -964
rect 6276 -996 6280 -964
rect 6240 -1044 6280 -996
rect 6240 -1076 6244 -1044
rect 6276 -1076 6280 -1044
rect 6240 -1124 6280 -1076
rect 6240 -1156 6244 -1124
rect 6276 -1156 6280 -1124
rect 6240 -1204 6280 -1156
rect 6240 -1236 6244 -1204
rect 6276 -1236 6280 -1204
rect 6240 -1284 6280 -1236
rect 6240 -1316 6244 -1284
rect 6276 -1316 6280 -1284
rect 6240 -1364 6280 -1316
rect 6240 -1396 6244 -1364
rect 6276 -1396 6280 -1364
rect 6240 -1444 6280 -1396
rect 6240 -1476 6244 -1444
rect 6276 -1476 6280 -1444
rect 6240 -1524 6280 -1476
rect 6240 -1556 6244 -1524
rect 6276 -1556 6280 -1524
rect 6240 -1604 6280 -1556
rect 6240 -1636 6244 -1604
rect 6276 -1636 6280 -1604
rect 6240 -1684 6280 -1636
rect 6240 -1716 6244 -1684
rect 6276 -1716 6280 -1684
rect 6240 -1764 6280 -1716
rect 6240 -1796 6244 -1764
rect 6276 -1796 6280 -1764
rect 6240 -1844 6280 -1796
rect 6240 -1876 6244 -1844
rect 6276 -1876 6280 -1844
rect 6240 -1924 6280 -1876
rect 6240 -1956 6244 -1924
rect 6276 -1956 6280 -1924
rect 6240 -2004 6280 -1956
rect 6240 -2036 6244 -2004
rect 6276 -2036 6280 -2004
rect 6240 -2084 6280 -2036
rect 6240 -2116 6244 -2084
rect 6276 -2116 6280 -2084
rect 6240 -2164 6280 -2116
rect 6240 -2196 6244 -2164
rect 6276 -2196 6280 -2164
rect 6240 -2244 6280 -2196
rect 6240 -2276 6244 -2244
rect 6276 -2276 6280 -2244
rect 6240 -2324 6280 -2276
rect 6240 -2356 6244 -2324
rect 6276 -2356 6280 -2324
rect 6240 -2404 6280 -2356
rect 6240 -2436 6244 -2404
rect 6276 -2436 6280 -2404
rect 6240 -2484 6280 -2436
rect 6240 -2516 6244 -2484
rect 6276 -2516 6280 -2484
rect 6240 -2564 6280 -2516
rect 6240 -2596 6244 -2564
rect 6276 -2596 6280 -2564
rect 6240 -2644 6280 -2596
rect 6240 -2676 6244 -2644
rect 6276 -2676 6280 -2644
rect 6240 -2724 6280 -2676
rect 6240 -2756 6244 -2724
rect 6276 -2756 6280 -2724
rect 6240 -2804 6280 -2756
rect 6240 -2836 6244 -2804
rect 6276 -2836 6280 -2804
rect 6240 -2884 6280 -2836
rect 6240 -2916 6244 -2884
rect 6276 -2916 6280 -2884
rect 6240 -2964 6280 -2916
rect 6240 -2996 6244 -2964
rect 6276 -2996 6280 -2964
rect 6240 -3044 6280 -2996
rect 6240 -3076 6244 -3044
rect 6276 -3076 6280 -3044
rect 6240 -3124 6280 -3076
rect 6240 -3156 6244 -3124
rect 6276 -3156 6280 -3124
rect 6240 -3204 6280 -3156
rect 6240 -3236 6244 -3204
rect 6276 -3236 6280 -3204
rect 6240 -3284 6280 -3236
rect 6240 -3316 6244 -3284
rect 6276 -3316 6280 -3284
rect 6240 -3364 6280 -3316
rect 6240 -3396 6244 -3364
rect 6276 -3396 6280 -3364
rect 6240 -3444 6280 -3396
rect 6240 -3476 6244 -3444
rect 6276 -3476 6280 -3444
rect 6240 -3524 6280 -3476
rect 6240 -3556 6244 -3524
rect 6276 -3556 6280 -3524
rect 6240 -3604 6280 -3556
rect 6240 -3636 6244 -3604
rect 6276 -3636 6280 -3604
rect 6240 -3684 6280 -3636
rect 6240 -3716 6244 -3684
rect 6276 -3716 6280 -3684
rect 6240 -3720 6280 -3716
rect 6320 1036 6360 1040
rect 6320 1004 6324 1036
rect 6356 1004 6360 1036
rect 6320 956 6360 1004
rect 6320 924 6324 956
rect 6356 924 6360 956
rect 6320 876 6360 924
rect 6320 844 6324 876
rect 6356 844 6360 876
rect 6320 796 6360 844
rect 6320 764 6324 796
rect 6356 764 6360 796
rect 6320 716 6360 764
rect 6320 684 6324 716
rect 6356 684 6360 716
rect 6320 636 6360 684
rect 6320 604 6324 636
rect 6356 604 6360 636
rect 6320 556 6360 604
rect 6320 524 6324 556
rect 6356 524 6360 556
rect 6320 476 6360 524
rect 6320 444 6324 476
rect 6356 444 6360 476
rect 6320 396 6360 444
rect 6320 364 6324 396
rect 6356 364 6360 396
rect 6320 316 6360 364
rect 6320 284 6324 316
rect 6356 284 6360 316
rect 6320 236 6360 284
rect 6320 204 6324 236
rect 6356 204 6360 236
rect 6320 156 6360 204
rect 6320 124 6324 156
rect 6356 124 6360 156
rect 6320 76 6360 124
rect 6320 44 6324 76
rect 6356 44 6360 76
rect 6320 -4 6360 44
rect 6320 -36 6324 -4
rect 6356 -36 6360 -4
rect 6320 -84 6360 -36
rect 6320 -116 6324 -84
rect 6356 -116 6360 -84
rect 6320 -164 6360 -116
rect 6320 -196 6324 -164
rect 6356 -196 6360 -164
rect 6320 -244 6360 -196
rect 6320 -276 6324 -244
rect 6356 -276 6360 -244
rect 6320 -324 6360 -276
rect 6320 -356 6324 -324
rect 6356 -356 6360 -324
rect 6320 -404 6360 -356
rect 6320 -436 6324 -404
rect 6356 -436 6360 -404
rect 6320 -484 6360 -436
rect 6320 -516 6324 -484
rect 6356 -516 6360 -484
rect 6320 -564 6360 -516
rect 6320 -596 6324 -564
rect 6356 -596 6360 -564
rect 6320 -644 6360 -596
rect 6320 -676 6324 -644
rect 6356 -676 6360 -644
rect 6320 -724 6360 -676
rect 6320 -756 6324 -724
rect 6356 -756 6360 -724
rect 6320 -804 6360 -756
rect 6320 -836 6324 -804
rect 6356 -836 6360 -804
rect 6320 -884 6360 -836
rect 6320 -916 6324 -884
rect 6356 -916 6360 -884
rect 6320 -964 6360 -916
rect 6320 -996 6324 -964
rect 6356 -996 6360 -964
rect 6320 -1044 6360 -996
rect 6320 -1076 6324 -1044
rect 6356 -1076 6360 -1044
rect 6320 -1124 6360 -1076
rect 6320 -1156 6324 -1124
rect 6356 -1156 6360 -1124
rect 6320 -1204 6360 -1156
rect 6320 -1236 6324 -1204
rect 6356 -1236 6360 -1204
rect 6320 -1284 6360 -1236
rect 6320 -1316 6324 -1284
rect 6356 -1316 6360 -1284
rect 6320 -1364 6360 -1316
rect 6320 -1396 6324 -1364
rect 6356 -1396 6360 -1364
rect 6320 -1444 6360 -1396
rect 6320 -1476 6324 -1444
rect 6356 -1476 6360 -1444
rect 6320 -1524 6360 -1476
rect 6320 -1556 6324 -1524
rect 6356 -1556 6360 -1524
rect 6320 -1604 6360 -1556
rect 6320 -1636 6324 -1604
rect 6356 -1636 6360 -1604
rect 6320 -1684 6360 -1636
rect 6320 -1716 6324 -1684
rect 6356 -1716 6360 -1684
rect 6320 -1764 6360 -1716
rect 6320 -1796 6324 -1764
rect 6356 -1796 6360 -1764
rect 6320 -1844 6360 -1796
rect 6320 -1876 6324 -1844
rect 6356 -1876 6360 -1844
rect 6320 -1924 6360 -1876
rect 6320 -1956 6324 -1924
rect 6356 -1956 6360 -1924
rect 6320 -2004 6360 -1956
rect 6320 -2036 6324 -2004
rect 6356 -2036 6360 -2004
rect 6320 -2084 6360 -2036
rect 6320 -2116 6324 -2084
rect 6356 -2116 6360 -2084
rect 6320 -2164 6360 -2116
rect 6320 -2196 6324 -2164
rect 6356 -2196 6360 -2164
rect 6320 -2244 6360 -2196
rect 6320 -2276 6324 -2244
rect 6356 -2276 6360 -2244
rect 6320 -2324 6360 -2276
rect 6320 -2356 6324 -2324
rect 6356 -2356 6360 -2324
rect 6320 -2404 6360 -2356
rect 6320 -2436 6324 -2404
rect 6356 -2436 6360 -2404
rect 6320 -2484 6360 -2436
rect 6320 -2516 6324 -2484
rect 6356 -2516 6360 -2484
rect 6320 -2564 6360 -2516
rect 6320 -2596 6324 -2564
rect 6356 -2596 6360 -2564
rect 6320 -2644 6360 -2596
rect 6320 -2676 6324 -2644
rect 6356 -2676 6360 -2644
rect 6320 -2724 6360 -2676
rect 6320 -2756 6324 -2724
rect 6356 -2756 6360 -2724
rect 6320 -2804 6360 -2756
rect 6320 -2836 6324 -2804
rect 6356 -2836 6360 -2804
rect 6320 -2884 6360 -2836
rect 6320 -2916 6324 -2884
rect 6356 -2916 6360 -2884
rect 6320 -2964 6360 -2916
rect 6320 -2996 6324 -2964
rect 6356 -2996 6360 -2964
rect 6320 -3044 6360 -2996
rect 6320 -3076 6324 -3044
rect 6356 -3076 6360 -3044
rect 6320 -3124 6360 -3076
rect 6320 -3156 6324 -3124
rect 6356 -3156 6360 -3124
rect 6320 -3204 6360 -3156
rect 6320 -3236 6324 -3204
rect 6356 -3236 6360 -3204
rect 6320 -3284 6360 -3236
rect 6320 -3316 6324 -3284
rect 6356 -3316 6360 -3284
rect 6320 -3364 6360 -3316
rect 6320 -3396 6324 -3364
rect 6356 -3396 6360 -3364
rect 6320 -3444 6360 -3396
rect 6320 -3476 6324 -3444
rect 6356 -3476 6360 -3444
rect 6320 -3524 6360 -3476
rect 6320 -3556 6324 -3524
rect 6356 -3556 6360 -3524
rect 6320 -3604 6360 -3556
rect 6320 -3636 6324 -3604
rect 6356 -3636 6360 -3604
rect 6320 -3684 6360 -3636
rect 6320 -3716 6324 -3684
rect 6356 -3716 6360 -3684
rect 6320 -3720 6360 -3716
rect 6400 1036 6440 1040
rect 6400 1004 6404 1036
rect 6436 1004 6440 1036
rect 6400 956 6440 1004
rect 6400 924 6404 956
rect 6436 924 6440 956
rect 6400 876 6440 924
rect 6400 844 6404 876
rect 6436 844 6440 876
rect 6400 796 6440 844
rect 6400 764 6404 796
rect 6436 764 6440 796
rect 6400 716 6440 764
rect 6400 684 6404 716
rect 6436 684 6440 716
rect 6400 636 6440 684
rect 6400 604 6404 636
rect 6436 604 6440 636
rect 6400 556 6440 604
rect 6400 524 6404 556
rect 6436 524 6440 556
rect 6400 476 6440 524
rect 6400 444 6404 476
rect 6436 444 6440 476
rect 6400 396 6440 444
rect 6400 364 6404 396
rect 6436 364 6440 396
rect 6400 316 6440 364
rect 6400 284 6404 316
rect 6436 284 6440 316
rect 6400 236 6440 284
rect 6400 204 6404 236
rect 6436 204 6440 236
rect 6400 156 6440 204
rect 6400 124 6404 156
rect 6436 124 6440 156
rect 6400 76 6440 124
rect 6400 44 6404 76
rect 6436 44 6440 76
rect 6400 -4 6440 44
rect 6400 -36 6404 -4
rect 6436 -36 6440 -4
rect 6400 -84 6440 -36
rect 6400 -116 6404 -84
rect 6436 -116 6440 -84
rect 6400 -164 6440 -116
rect 6400 -196 6404 -164
rect 6436 -196 6440 -164
rect 6400 -244 6440 -196
rect 6400 -276 6404 -244
rect 6436 -276 6440 -244
rect 6400 -324 6440 -276
rect 6400 -356 6404 -324
rect 6436 -356 6440 -324
rect 6400 -404 6440 -356
rect 6400 -436 6404 -404
rect 6436 -436 6440 -404
rect 6400 -484 6440 -436
rect 6400 -516 6404 -484
rect 6436 -516 6440 -484
rect 6400 -564 6440 -516
rect 6400 -596 6404 -564
rect 6436 -596 6440 -564
rect 6400 -644 6440 -596
rect 6400 -676 6404 -644
rect 6436 -676 6440 -644
rect 6400 -724 6440 -676
rect 6400 -756 6404 -724
rect 6436 -756 6440 -724
rect 6400 -804 6440 -756
rect 6400 -836 6404 -804
rect 6436 -836 6440 -804
rect 6400 -884 6440 -836
rect 6400 -916 6404 -884
rect 6436 -916 6440 -884
rect 6400 -964 6440 -916
rect 6400 -996 6404 -964
rect 6436 -996 6440 -964
rect 6400 -1044 6440 -996
rect 6400 -1076 6404 -1044
rect 6436 -1076 6440 -1044
rect 6400 -1124 6440 -1076
rect 6400 -1156 6404 -1124
rect 6436 -1156 6440 -1124
rect 6400 -1204 6440 -1156
rect 6400 -1236 6404 -1204
rect 6436 -1236 6440 -1204
rect 6400 -1284 6440 -1236
rect 6400 -1316 6404 -1284
rect 6436 -1316 6440 -1284
rect 6400 -1364 6440 -1316
rect 6400 -1396 6404 -1364
rect 6436 -1396 6440 -1364
rect 6400 -1444 6440 -1396
rect 6400 -1476 6404 -1444
rect 6436 -1476 6440 -1444
rect 6400 -1524 6440 -1476
rect 6400 -1556 6404 -1524
rect 6436 -1556 6440 -1524
rect 6400 -1604 6440 -1556
rect 6400 -1636 6404 -1604
rect 6436 -1636 6440 -1604
rect 6400 -1684 6440 -1636
rect 6400 -1716 6404 -1684
rect 6436 -1716 6440 -1684
rect 6400 -1764 6440 -1716
rect 6400 -1796 6404 -1764
rect 6436 -1796 6440 -1764
rect 6400 -1844 6440 -1796
rect 6400 -1876 6404 -1844
rect 6436 -1876 6440 -1844
rect 6400 -1924 6440 -1876
rect 6400 -1956 6404 -1924
rect 6436 -1956 6440 -1924
rect 6400 -2004 6440 -1956
rect 6400 -2036 6404 -2004
rect 6436 -2036 6440 -2004
rect 6400 -2084 6440 -2036
rect 6400 -2116 6404 -2084
rect 6436 -2116 6440 -2084
rect 6400 -2164 6440 -2116
rect 6400 -2196 6404 -2164
rect 6436 -2196 6440 -2164
rect 6400 -2244 6440 -2196
rect 6400 -2276 6404 -2244
rect 6436 -2276 6440 -2244
rect 6400 -2324 6440 -2276
rect 6400 -2356 6404 -2324
rect 6436 -2356 6440 -2324
rect 6400 -2404 6440 -2356
rect 6400 -2436 6404 -2404
rect 6436 -2436 6440 -2404
rect 6400 -2484 6440 -2436
rect 6400 -2516 6404 -2484
rect 6436 -2516 6440 -2484
rect 6400 -2564 6440 -2516
rect 6400 -2596 6404 -2564
rect 6436 -2596 6440 -2564
rect 6400 -2644 6440 -2596
rect 6400 -2676 6404 -2644
rect 6436 -2676 6440 -2644
rect 6400 -2724 6440 -2676
rect 6400 -2756 6404 -2724
rect 6436 -2756 6440 -2724
rect 6400 -2804 6440 -2756
rect 6400 -2836 6404 -2804
rect 6436 -2836 6440 -2804
rect 6400 -2884 6440 -2836
rect 6400 -2916 6404 -2884
rect 6436 -2916 6440 -2884
rect 6400 -2964 6440 -2916
rect 6400 -2996 6404 -2964
rect 6436 -2996 6440 -2964
rect 6400 -3044 6440 -2996
rect 6400 -3076 6404 -3044
rect 6436 -3076 6440 -3044
rect 6400 -3124 6440 -3076
rect 6400 -3156 6404 -3124
rect 6436 -3156 6440 -3124
rect 6400 -3204 6440 -3156
rect 6400 -3236 6404 -3204
rect 6436 -3236 6440 -3204
rect 6400 -3284 6440 -3236
rect 6400 -3316 6404 -3284
rect 6436 -3316 6440 -3284
rect 6400 -3364 6440 -3316
rect 6400 -3396 6404 -3364
rect 6436 -3396 6440 -3364
rect 6400 -3444 6440 -3396
rect 6400 -3476 6404 -3444
rect 6436 -3476 6440 -3444
rect 6400 -3524 6440 -3476
rect 6400 -3556 6404 -3524
rect 6436 -3556 6440 -3524
rect 6400 -3604 6440 -3556
rect 6400 -3636 6404 -3604
rect 6436 -3636 6440 -3604
rect 6400 -3684 6440 -3636
rect 6400 -3716 6404 -3684
rect 6436 -3716 6440 -3684
rect 6400 -3720 6440 -3716
rect 6480 1036 6520 1040
rect 6480 1004 6484 1036
rect 6516 1004 6520 1036
rect 6480 956 6520 1004
rect 6480 924 6484 956
rect 6516 924 6520 956
rect 6480 876 6520 924
rect 6480 844 6484 876
rect 6516 844 6520 876
rect 6480 796 6520 844
rect 6480 764 6484 796
rect 6516 764 6520 796
rect 6480 716 6520 764
rect 6480 684 6484 716
rect 6516 684 6520 716
rect 6480 636 6520 684
rect 6480 604 6484 636
rect 6516 604 6520 636
rect 6480 556 6520 604
rect 6480 524 6484 556
rect 6516 524 6520 556
rect 6480 476 6520 524
rect 6480 444 6484 476
rect 6516 444 6520 476
rect 6480 396 6520 444
rect 6480 364 6484 396
rect 6516 364 6520 396
rect 6480 316 6520 364
rect 6480 284 6484 316
rect 6516 284 6520 316
rect 6480 236 6520 284
rect 6480 204 6484 236
rect 6516 204 6520 236
rect 6480 156 6520 204
rect 6480 124 6484 156
rect 6516 124 6520 156
rect 6480 76 6520 124
rect 6480 44 6484 76
rect 6516 44 6520 76
rect 6480 -4 6520 44
rect 6480 -36 6484 -4
rect 6516 -36 6520 -4
rect 6480 -84 6520 -36
rect 6480 -116 6484 -84
rect 6516 -116 6520 -84
rect 6480 -164 6520 -116
rect 6480 -196 6484 -164
rect 6516 -196 6520 -164
rect 6480 -244 6520 -196
rect 6480 -276 6484 -244
rect 6516 -276 6520 -244
rect 6480 -324 6520 -276
rect 6480 -356 6484 -324
rect 6516 -356 6520 -324
rect 6480 -404 6520 -356
rect 6480 -436 6484 -404
rect 6516 -436 6520 -404
rect 6480 -484 6520 -436
rect 6480 -516 6484 -484
rect 6516 -516 6520 -484
rect 6480 -564 6520 -516
rect 6480 -596 6484 -564
rect 6516 -596 6520 -564
rect 6480 -644 6520 -596
rect 6480 -676 6484 -644
rect 6516 -676 6520 -644
rect 6480 -724 6520 -676
rect 6480 -756 6484 -724
rect 6516 -756 6520 -724
rect 6480 -804 6520 -756
rect 6480 -836 6484 -804
rect 6516 -836 6520 -804
rect 6480 -884 6520 -836
rect 6480 -916 6484 -884
rect 6516 -916 6520 -884
rect 6480 -964 6520 -916
rect 6480 -996 6484 -964
rect 6516 -996 6520 -964
rect 6480 -1044 6520 -996
rect 6480 -1076 6484 -1044
rect 6516 -1076 6520 -1044
rect 6480 -1124 6520 -1076
rect 6480 -1156 6484 -1124
rect 6516 -1156 6520 -1124
rect 6480 -1204 6520 -1156
rect 6480 -1236 6484 -1204
rect 6516 -1236 6520 -1204
rect 6480 -1284 6520 -1236
rect 6480 -1316 6484 -1284
rect 6516 -1316 6520 -1284
rect 6480 -1364 6520 -1316
rect 6480 -1396 6484 -1364
rect 6516 -1396 6520 -1364
rect 6480 -1444 6520 -1396
rect 6480 -1476 6484 -1444
rect 6516 -1476 6520 -1444
rect 6480 -1524 6520 -1476
rect 6480 -1556 6484 -1524
rect 6516 -1556 6520 -1524
rect 6480 -1604 6520 -1556
rect 6480 -1636 6484 -1604
rect 6516 -1636 6520 -1604
rect 6480 -1684 6520 -1636
rect 6480 -1716 6484 -1684
rect 6516 -1716 6520 -1684
rect 6480 -1764 6520 -1716
rect 6480 -1796 6484 -1764
rect 6516 -1796 6520 -1764
rect 6480 -1844 6520 -1796
rect 6480 -1876 6484 -1844
rect 6516 -1876 6520 -1844
rect 6480 -1924 6520 -1876
rect 6480 -1956 6484 -1924
rect 6516 -1956 6520 -1924
rect 6480 -2004 6520 -1956
rect 6480 -2036 6484 -2004
rect 6516 -2036 6520 -2004
rect 6480 -2084 6520 -2036
rect 6480 -2116 6484 -2084
rect 6516 -2116 6520 -2084
rect 6480 -2164 6520 -2116
rect 6480 -2196 6484 -2164
rect 6516 -2196 6520 -2164
rect 6480 -2244 6520 -2196
rect 6480 -2276 6484 -2244
rect 6516 -2276 6520 -2244
rect 6480 -2324 6520 -2276
rect 6480 -2356 6484 -2324
rect 6516 -2356 6520 -2324
rect 6480 -2404 6520 -2356
rect 6480 -2436 6484 -2404
rect 6516 -2436 6520 -2404
rect 6480 -2484 6520 -2436
rect 6480 -2516 6484 -2484
rect 6516 -2516 6520 -2484
rect 6480 -2564 6520 -2516
rect 6480 -2596 6484 -2564
rect 6516 -2596 6520 -2564
rect 6480 -2644 6520 -2596
rect 6480 -2676 6484 -2644
rect 6516 -2676 6520 -2644
rect 6480 -2724 6520 -2676
rect 6480 -2756 6484 -2724
rect 6516 -2756 6520 -2724
rect 6480 -2804 6520 -2756
rect 6480 -2836 6484 -2804
rect 6516 -2836 6520 -2804
rect 6480 -2884 6520 -2836
rect 6480 -2916 6484 -2884
rect 6516 -2916 6520 -2884
rect 6480 -2964 6520 -2916
rect 6480 -2996 6484 -2964
rect 6516 -2996 6520 -2964
rect 6480 -3044 6520 -2996
rect 6480 -3076 6484 -3044
rect 6516 -3076 6520 -3044
rect 6480 -3124 6520 -3076
rect 6480 -3156 6484 -3124
rect 6516 -3156 6520 -3124
rect 6480 -3204 6520 -3156
rect 6480 -3236 6484 -3204
rect 6516 -3236 6520 -3204
rect 6480 -3284 6520 -3236
rect 6480 -3316 6484 -3284
rect 6516 -3316 6520 -3284
rect 6480 -3364 6520 -3316
rect 6480 -3396 6484 -3364
rect 6516 -3396 6520 -3364
rect 6480 -3444 6520 -3396
rect 6480 -3476 6484 -3444
rect 6516 -3476 6520 -3444
rect 6480 -3524 6520 -3476
rect 6480 -3556 6484 -3524
rect 6516 -3556 6520 -3524
rect 6480 -3604 6520 -3556
rect 6480 -3636 6484 -3604
rect 6516 -3636 6520 -3604
rect 6480 -3684 6520 -3636
rect 6480 -3716 6484 -3684
rect 6516 -3716 6520 -3684
rect 6480 -3720 6520 -3716
rect 6560 1036 6600 1040
rect 6560 1004 6564 1036
rect 6596 1004 6600 1036
rect 6560 956 6600 1004
rect 6560 924 6564 956
rect 6596 924 6600 956
rect 6560 876 6600 924
rect 6560 844 6564 876
rect 6596 844 6600 876
rect 6560 796 6600 844
rect 6560 764 6564 796
rect 6596 764 6600 796
rect 6560 716 6600 764
rect 6560 684 6564 716
rect 6596 684 6600 716
rect 6560 636 6600 684
rect 6560 604 6564 636
rect 6596 604 6600 636
rect 6560 556 6600 604
rect 6560 524 6564 556
rect 6596 524 6600 556
rect 6560 476 6600 524
rect 6560 444 6564 476
rect 6596 444 6600 476
rect 6560 396 6600 444
rect 6560 364 6564 396
rect 6596 364 6600 396
rect 6560 316 6600 364
rect 6560 284 6564 316
rect 6596 284 6600 316
rect 6560 236 6600 284
rect 6560 204 6564 236
rect 6596 204 6600 236
rect 6560 156 6600 204
rect 6560 124 6564 156
rect 6596 124 6600 156
rect 6560 76 6600 124
rect 6560 44 6564 76
rect 6596 44 6600 76
rect 6560 -4 6600 44
rect 6560 -36 6564 -4
rect 6596 -36 6600 -4
rect 6560 -84 6600 -36
rect 6560 -116 6564 -84
rect 6596 -116 6600 -84
rect 6560 -164 6600 -116
rect 6560 -196 6564 -164
rect 6596 -196 6600 -164
rect 6560 -244 6600 -196
rect 6560 -276 6564 -244
rect 6596 -276 6600 -244
rect 6560 -324 6600 -276
rect 6560 -356 6564 -324
rect 6596 -356 6600 -324
rect 6560 -404 6600 -356
rect 6560 -436 6564 -404
rect 6596 -436 6600 -404
rect 6560 -484 6600 -436
rect 6560 -516 6564 -484
rect 6596 -516 6600 -484
rect 6560 -564 6600 -516
rect 6560 -596 6564 -564
rect 6596 -596 6600 -564
rect 6560 -644 6600 -596
rect 6560 -676 6564 -644
rect 6596 -676 6600 -644
rect 6560 -724 6600 -676
rect 6560 -756 6564 -724
rect 6596 -756 6600 -724
rect 6560 -804 6600 -756
rect 6560 -836 6564 -804
rect 6596 -836 6600 -804
rect 6560 -884 6600 -836
rect 6560 -916 6564 -884
rect 6596 -916 6600 -884
rect 6560 -964 6600 -916
rect 6560 -996 6564 -964
rect 6596 -996 6600 -964
rect 6560 -1044 6600 -996
rect 6560 -1076 6564 -1044
rect 6596 -1076 6600 -1044
rect 6560 -1124 6600 -1076
rect 6560 -1156 6564 -1124
rect 6596 -1156 6600 -1124
rect 6560 -1204 6600 -1156
rect 6560 -1236 6564 -1204
rect 6596 -1236 6600 -1204
rect 6560 -1284 6600 -1236
rect 6560 -1316 6564 -1284
rect 6596 -1316 6600 -1284
rect 6560 -1364 6600 -1316
rect 6560 -1396 6564 -1364
rect 6596 -1396 6600 -1364
rect 6560 -1444 6600 -1396
rect 6560 -1476 6564 -1444
rect 6596 -1476 6600 -1444
rect 6560 -1524 6600 -1476
rect 6560 -1556 6564 -1524
rect 6596 -1556 6600 -1524
rect 6560 -1604 6600 -1556
rect 6560 -1636 6564 -1604
rect 6596 -1636 6600 -1604
rect 6560 -1684 6600 -1636
rect 6560 -1716 6564 -1684
rect 6596 -1716 6600 -1684
rect 6560 -1764 6600 -1716
rect 6560 -1796 6564 -1764
rect 6596 -1796 6600 -1764
rect 6560 -1844 6600 -1796
rect 6560 -1876 6564 -1844
rect 6596 -1876 6600 -1844
rect 6560 -1924 6600 -1876
rect 6560 -1956 6564 -1924
rect 6596 -1956 6600 -1924
rect 6560 -2004 6600 -1956
rect 6560 -2036 6564 -2004
rect 6596 -2036 6600 -2004
rect 6560 -2084 6600 -2036
rect 6560 -2116 6564 -2084
rect 6596 -2116 6600 -2084
rect 6560 -2164 6600 -2116
rect 6560 -2196 6564 -2164
rect 6596 -2196 6600 -2164
rect 6560 -2244 6600 -2196
rect 6560 -2276 6564 -2244
rect 6596 -2276 6600 -2244
rect 6560 -2324 6600 -2276
rect 6560 -2356 6564 -2324
rect 6596 -2356 6600 -2324
rect 6560 -2404 6600 -2356
rect 6560 -2436 6564 -2404
rect 6596 -2436 6600 -2404
rect 6560 -2484 6600 -2436
rect 6560 -2516 6564 -2484
rect 6596 -2516 6600 -2484
rect 6560 -2564 6600 -2516
rect 6560 -2596 6564 -2564
rect 6596 -2596 6600 -2564
rect 6560 -2644 6600 -2596
rect 6560 -2676 6564 -2644
rect 6596 -2676 6600 -2644
rect 6560 -2724 6600 -2676
rect 6560 -2756 6564 -2724
rect 6596 -2756 6600 -2724
rect 6560 -2804 6600 -2756
rect 6560 -2836 6564 -2804
rect 6596 -2836 6600 -2804
rect 6560 -2884 6600 -2836
rect 6560 -2916 6564 -2884
rect 6596 -2916 6600 -2884
rect 6560 -2964 6600 -2916
rect 6560 -2996 6564 -2964
rect 6596 -2996 6600 -2964
rect 6560 -3044 6600 -2996
rect 6560 -3076 6564 -3044
rect 6596 -3076 6600 -3044
rect 6560 -3124 6600 -3076
rect 6560 -3156 6564 -3124
rect 6596 -3156 6600 -3124
rect 6560 -3204 6600 -3156
rect 6560 -3236 6564 -3204
rect 6596 -3236 6600 -3204
rect 6560 -3284 6600 -3236
rect 6560 -3316 6564 -3284
rect 6596 -3316 6600 -3284
rect 6560 -3364 6600 -3316
rect 6560 -3396 6564 -3364
rect 6596 -3396 6600 -3364
rect 6560 -3444 6600 -3396
rect 6560 -3476 6564 -3444
rect 6596 -3476 6600 -3444
rect 6560 -3524 6600 -3476
rect 6560 -3556 6564 -3524
rect 6596 -3556 6600 -3524
rect 6560 -3604 6600 -3556
rect 6560 -3636 6564 -3604
rect 6596 -3636 6600 -3604
rect 6560 -3684 6600 -3636
rect 6560 -3716 6564 -3684
rect 6596 -3716 6600 -3684
rect 6560 -3720 6600 -3716
rect 6640 1036 6680 1040
rect 6640 1004 6644 1036
rect 6676 1004 6680 1036
rect 6640 956 6680 1004
rect 6640 924 6644 956
rect 6676 924 6680 956
rect 6640 876 6680 924
rect 6640 844 6644 876
rect 6676 844 6680 876
rect 6640 796 6680 844
rect 6640 764 6644 796
rect 6676 764 6680 796
rect 6640 716 6680 764
rect 6640 684 6644 716
rect 6676 684 6680 716
rect 6640 636 6680 684
rect 6640 604 6644 636
rect 6676 604 6680 636
rect 6640 556 6680 604
rect 6640 524 6644 556
rect 6676 524 6680 556
rect 6640 476 6680 524
rect 6640 444 6644 476
rect 6676 444 6680 476
rect 6640 396 6680 444
rect 6640 364 6644 396
rect 6676 364 6680 396
rect 6640 316 6680 364
rect 6640 284 6644 316
rect 6676 284 6680 316
rect 6640 236 6680 284
rect 6640 204 6644 236
rect 6676 204 6680 236
rect 6640 156 6680 204
rect 6640 124 6644 156
rect 6676 124 6680 156
rect 6640 76 6680 124
rect 6640 44 6644 76
rect 6676 44 6680 76
rect 6640 -4 6680 44
rect 6640 -36 6644 -4
rect 6676 -36 6680 -4
rect 6640 -84 6680 -36
rect 6640 -116 6644 -84
rect 6676 -116 6680 -84
rect 6640 -164 6680 -116
rect 6640 -196 6644 -164
rect 6676 -196 6680 -164
rect 6640 -244 6680 -196
rect 6640 -276 6644 -244
rect 6676 -276 6680 -244
rect 6640 -324 6680 -276
rect 6640 -356 6644 -324
rect 6676 -356 6680 -324
rect 6640 -404 6680 -356
rect 6640 -436 6644 -404
rect 6676 -436 6680 -404
rect 6640 -484 6680 -436
rect 6640 -516 6644 -484
rect 6676 -516 6680 -484
rect 6640 -564 6680 -516
rect 6640 -596 6644 -564
rect 6676 -596 6680 -564
rect 6640 -644 6680 -596
rect 6640 -676 6644 -644
rect 6676 -676 6680 -644
rect 6640 -724 6680 -676
rect 6640 -756 6644 -724
rect 6676 -756 6680 -724
rect 6640 -804 6680 -756
rect 6640 -836 6644 -804
rect 6676 -836 6680 -804
rect 6640 -884 6680 -836
rect 6640 -916 6644 -884
rect 6676 -916 6680 -884
rect 6640 -964 6680 -916
rect 6640 -996 6644 -964
rect 6676 -996 6680 -964
rect 6640 -1044 6680 -996
rect 6640 -1076 6644 -1044
rect 6676 -1076 6680 -1044
rect 6640 -1124 6680 -1076
rect 6640 -1156 6644 -1124
rect 6676 -1156 6680 -1124
rect 6640 -1204 6680 -1156
rect 6640 -1236 6644 -1204
rect 6676 -1236 6680 -1204
rect 6640 -1284 6680 -1236
rect 6640 -1316 6644 -1284
rect 6676 -1316 6680 -1284
rect 6640 -1364 6680 -1316
rect 6640 -1396 6644 -1364
rect 6676 -1396 6680 -1364
rect 6640 -1444 6680 -1396
rect 6640 -1476 6644 -1444
rect 6676 -1476 6680 -1444
rect 6640 -1524 6680 -1476
rect 6640 -1556 6644 -1524
rect 6676 -1556 6680 -1524
rect 6640 -1604 6680 -1556
rect 6640 -1636 6644 -1604
rect 6676 -1636 6680 -1604
rect 6640 -1684 6680 -1636
rect 6640 -1716 6644 -1684
rect 6676 -1716 6680 -1684
rect 6640 -1764 6680 -1716
rect 6640 -1796 6644 -1764
rect 6676 -1796 6680 -1764
rect 6640 -1844 6680 -1796
rect 6640 -1876 6644 -1844
rect 6676 -1876 6680 -1844
rect 6640 -1924 6680 -1876
rect 6640 -1956 6644 -1924
rect 6676 -1956 6680 -1924
rect 6640 -2004 6680 -1956
rect 6640 -2036 6644 -2004
rect 6676 -2036 6680 -2004
rect 6640 -2084 6680 -2036
rect 6640 -2116 6644 -2084
rect 6676 -2116 6680 -2084
rect 6640 -2164 6680 -2116
rect 6640 -2196 6644 -2164
rect 6676 -2196 6680 -2164
rect 6640 -2244 6680 -2196
rect 6640 -2276 6644 -2244
rect 6676 -2276 6680 -2244
rect 6640 -2324 6680 -2276
rect 6640 -2356 6644 -2324
rect 6676 -2356 6680 -2324
rect 6640 -2404 6680 -2356
rect 6640 -2436 6644 -2404
rect 6676 -2436 6680 -2404
rect 6640 -2484 6680 -2436
rect 6640 -2516 6644 -2484
rect 6676 -2516 6680 -2484
rect 6640 -2564 6680 -2516
rect 6640 -2596 6644 -2564
rect 6676 -2596 6680 -2564
rect 6640 -2644 6680 -2596
rect 6640 -2676 6644 -2644
rect 6676 -2676 6680 -2644
rect 6640 -2724 6680 -2676
rect 6640 -2756 6644 -2724
rect 6676 -2756 6680 -2724
rect 6640 -2804 6680 -2756
rect 6640 -2836 6644 -2804
rect 6676 -2836 6680 -2804
rect 6640 -2884 6680 -2836
rect 6640 -2916 6644 -2884
rect 6676 -2916 6680 -2884
rect 6640 -2964 6680 -2916
rect 6640 -2996 6644 -2964
rect 6676 -2996 6680 -2964
rect 6640 -3044 6680 -2996
rect 6640 -3076 6644 -3044
rect 6676 -3076 6680 -3044
rect 6640 -3124 6680 -3076
rect 6640 -3156 6644 -3124
rect 6676 -3156 6680 -3124
rect 6640 -3204 6680 -3156
rect 6640 -3236 6644 -3204
rect 6676 -3236 6680 -3204
rect 6640 -3284 6680 -3236
rect 6640 -3316 6644 -3284
rect 6676 -3316 6680 -3284
rect 6640 -3364 6680 -3316
rect 6640 -3396 6644 -3364
rect 6676 -3396 6680 -3364
rect 6640 -3444 6680 -3396
rect 6640 -3476 6644 -3444
rect 6676 -3476 6680 -3444
rect 6640 -3524 6680 -3476
rect 6640 -3556 6644 -3524
rect 6676 -3556 6680 -3524
rect 6640 -3604 6680 -3556
rect 6640 -3636 6644 -3604
rect 6676 -3636 6680 -3604
rect 6640 -3684 6680 -3636
rect 6640 -3716 6644 -3684
rect 6676 -3716 6680 -3684
rect 6640 -3720 6680 -3716
rect 6720 1036 6760 1040
rect 6720 1004 6724 1036
rect 6756 1004 6760 1036
rect 6720 956 6760 1004
rect 6720 924 6724 956
rect 6756 924 6760 956
rect 6720 876 6760 924
rect 6720 844 6724 876
rect 6756 844 6760 876
rect 6720 796 6760 844
rect 6720 764 6724 796
rect 6756 764 6760 796
rect 6720 716 6760 764
rect 6720 684 6724 716
rect 6756 684 6760 716
rect 6720 636 6760 684
rect 6720 604 6724 636
rect 6756 604 6760 636
rect 6720 556 6760 604
rect 6720 524 6724 556
rect 6756 524 6760 556
rect 6720 476 6760 524
rect 6720 444 6724 476
rect 6756 444 6760 476
rect 6720 396 6760 444
rect 6720 364 6724 396
rect 6756 364 6760 396
rect 6720 316 6760 364
rect 6720 284 6724 316
rect 6756 284 6760 316
rect 6720 236 6760 284
rect 6720 204 6724 236
rect 6756 204 6760 236
rect 6720 156 6760 204
rect 6720 124 6724 156
rect 6756 124 6760 156
rect 6720 76 6760 124
rect 6720 44 6724 76
rect 6756 44 6760 76
rect 6720 -4 6760 44
rect 6720 -36 6724 -4
rect 6756 -36 6760 -4
rect 6720 -84 6760 -36
rect 6720 -116 6724 -84
rect 6756 -116 6760 -84
rect 6720 -164 6760 -116
rect 6720 -196 6724 -164
rect 6756 -196 6760 -164
rect 6720 -244 6760 -196
rect 6720 -276 6724 -244
rect 6756 -276 6760 -244
rect 6720 -324 6760 -276
rect 6720 -356 6724 -324
rect 6756 -356 6760 -324
rect 6720 -404 6760 -356
rect 6720 -436 6724 -404
rect 6756 -436 6760 -404
rect 6720 -484 6760 -436
rect 6720 -516 6724 -484
rect 6756 -516 6760 -484
rect 6720 -564 6760 -516
rect 6720 -596 6724 -564
rect 6756 -596 6760 -564
rect 6720 -644 6760 -596
rect 6720 -676 6724 -644
rect 6756 -676 6760 -644
rect 6720 -724 6760 -676
rect 6720 -756 6724 -724
rect 6756 -756 6760 -724
rect 6720 -804 6760 -756
rect 6720 -836 6724 -804
rect 6756 -836 6760 -804
rect 6720 -884 6760 -836
rect 6720 -916 6724 -884
rect 6756 -916 6760 -884
rect 6720 -964 6760 -916
rect 6720 -996 6724 -964
rect 6756 -996 6760 -964
rect 6720 -1044 6760 -996
rect 6720 -1076 6724 -1044
rect 6756 -1076 6760 -1044
rect 6720 -1124 6760 -1076
rect 6720 -1156 6724 -1124
rect 6756 -1156 6760 -1124
rect 6720 -1204 6760 -1156
rect 6720 -1236 6724 -1204
rect 6756 -1236 6760 -1204
rect 6720 -1284 6760 -1236
rect 6720 -1316 6724 -1284
rect 6756 -1316 6760 -1284
rect 6720 -1364 6760 -1316
rect 6720 -1396 6724 -1364
rect 6756 -1396 6760 -1364
rect 6720 -1444 6760 -1396
rect 6720 -1476 6724 -1444
rect 6756 -1476 6760 -1444
rect 6720 -1524 6760 -1476
rect 6720 -1556 6724 -1524
rect 6756 -1556 6760 -1524
rect 6720 -1604 6760 -1556
rect 6720 -1636 6724 -1604
rect 6756 -1636 6760 -1604
rect 6720 -1684 6760 -1636
rect 6720 -1716 6724 -1684
rect 6756 -1716 6760 -1684
rect 6720 -1764 6760 -1716
rect 6720 -1796 6724 -1764
rect 6756 -1796 6760 -1764
rect 6720 -1844 6760 -1796
rect 6720 -1876 6724 -1844
rect 6756 -1876 6760 -1844
rect 6720 -1924 6760 -1876
rect 6720 -1956 6724 -1924
rect 6756 -1956 6760 -1924
rect 6720 -2004 6760 -1956
rect 6720 -2036 6724 -2004
rect 6756 -2036 6760 -2004
rect 6720 -2084 6760 -2036
rect 6720 -2116 6724 -2084
rect 6756 -2116 6760 -2084
rect 6720 -2164 6760 -2116
rect 6720 -2196 6724 -2164
rect 6756 -2196 6760 -2164
rect 6720 -2244 6760 -2196
rect 6720 -2276 6724 -2244
rect 6756 -2276 6760 -2244
rect 6720 -2324 6760 -2276
rect 6720 -2356 6724 -2324
rect 6756 -2356 6760 -2324
rect 6720 -2404 6760 -2356
rect 6720 -2436 6724 -2404
rect 6756 -2436 6760 -2404
rect 6720 -2484 6760 -2436
rect 6720 -2516 6724 -2484
rect 6756 -2516 6760 -2484
rect 6720 -2564 6760 -2516
rect 6720 -2596 6724 -2564
rect 6756 -2596 6760 -2564
rect 6720 -2644 6760 -2596
rect 6720 -2676 6724 -2644
rect 6756 -2676 6760 -2644
rect 6720 -2724 6760 -2676
rect 6720 -2756 6724 -2724
rect 6756 -2756 6760 -2724
rect 6720 -2804 6760 -2756
rect 6720 -2836 6724 -2804
rect 6756 -2836 6760 -2804
rect 6720 -2884 6760 -2836
rect 6720 -2916 6724 -2884
rect 6756 -2916 6760 -2884
rect 6720 -2964 6760 -2916
rect 6720 -2996 6724 -2964
rect 6756 -2996 6760 -2964
rect 6720 -3044 6760 -2996
rect 6720 -3076 6724 -3044
rect 6756 -3076 6760 -3044
rect 6720 -3124 6760 -3076
rect 6720 -3156 6724 -3124
rect 6756 -3156 6760 -3124
rect 6720 -3204 6760 -3156
rect 6720 -3236 6724 -3204
rect 6756 -3236 6760 -3204
rect 6720 -3284 6760 -3236
rect 6720 -3316 6724 -3284
rect 6756 -3316 6760 -3284
rect 6720 -3364 6760 -3316
rect 6720 -3396 6724 -3364
rect 6756 -3396 6760 -3364
rect 6720 -3444 6760 -3396
rect 6720 -3476 6724 -3444
rect 6756 -3476 6760 -3444
rect 6720 -3524 6760 -3476
rect 6720 -3556 6724 -3524
rect 6756 -3556 6760 -3524
rect 6720 -3604 6760 -3556
rect 6720 -3636 6724 -3604
rect 6756 -3636 6760 -3604
rect 6720 -3684 6760 -3636
rect 6720 -3716 6724 -3684
rect 6756 -3716 6760 -3684
rect 6720 -3720 6760 -3716
rect 6800 1036 6840 1040
rect 6800 1004 6804 1036
rect 6836 1004 6840 1036
rect 6800 956 6840 1004
rect 6800 924 6804 956
rect 6836 924 6840 956
rect 6800 876 6840 924
rect 6800 844 6804 876
rect 6836 844 6840 876
rect 6800 796 6840 844
rect 6800 764 6804 796
rect 6836 764 6840 796
rect 6800 716 6840 764
rect 6800 684 6804 716
rect 6836 684 6840 716
rect 6800 636 6840 684
rect 6800 604 6804 636
rect 6836 604 6840 636
rect 6800 556 6840 604
rect 6800 524 6804 556
rect 6836 524 6840 556
rect 6800 476 6840 524
rect 6800 444 6804 476
rect 6836 444 6840 476
rect 6800 396 6840 444
rect 6800 364 6804 396
rect 6836 364 6840 396
rect 6800 316 6840 364
rect 6800 284 6804 316
rect 6836 284 6840 316
rect 6800 236 6840 284
rect 6800 204 6804 236
rect 6836 204 6840 236
rect 6800 156 6840 204
rect 6800 124 6804 156
rect 6836 124 6840 156
rect 6800 76 6840 124
rect 6800 44 6804 76
rect 6836 44 6840 76
rect 6800 -4 6840 44
rect 6800 -36 6804 -4
rect 6836 -36 6840 -4
rect 6800 -84 6840 -36
rect 6800 -116 6804 -84
rect 6836 -116 6840 -84
rect 6800 -164 6840 -116
rect 6800 -196 6804 -164
rect 6836 -196 6840 -164
rect 6800 -244 6840 -196
rect 6800 -276 6804 -244
rect 6836 -276 6840 -244
rect 6800 -324 6840 -276
rect 6800 -356 6804 -324
rect 6836 -356 6840 -324
rect 6800 -404 6840 -356
rect 6800 -436 6804 -404
rect 6836 -436 6840 -404
rect 6800 -484 6840 -436
rect 6800 -516 6804 -484
rect 6836 -516 6840 -484
rect 6800 -564 6840 -516
rect 6800 -596 6804 -564
rect 6836 -596 6840 -564
rect 6800 -644 6840 -596
rect 6800 -676 6804 -644
rect 6836 -676 6840 -644
rect 6800 -724 6840 -676
rect 6800 -756 6804 -724
rect 6836 -756 6840 -724
rect 6800 -804 6840 -756
rect 6800 -836 6804 -804
rect 6836 -836 6840 -804
rect 6800 -884 6840 -836
rect 6800 -916 6804 -884
rect 6836 -916 6840 -884
rect 6800 -964 6840 -916
rect 6800 -996 6804 -964
rect 6836 -996 6840 -964
rect 6800 -1044 6840 -996
rect 6800 -1076 6804 -1044
rect 6836 -1076 6840 -1044
rect 6800 -1124 6840 -1076
rect 6800 -1156 6804 -1124
rect 6836 -1156 6840 -1124
rect 6800 -1204 6840 -1156
rect 6800 -1236 6804 -1204
rect 6836 -1236 6840 -1204
rect 6800 -1284 6840 -1236
rect 6800 -1316 6804 -1284
rect 6836 -1316 6840 -1284
rect 6800 -1364 6840 -1316
rect 6800 -1396 6804 -1364
rect 6836 -1396 6840 -1364
rect 6800 -1444 6840 -1396
rect 6800 -1476 6804 -1444
rect 6836 -1476 6840 -1444
rect 6800 -1524 6840 -1476
rect 6800 -1556 6804 -1524
rect 6836 -1556 6840 -1524
rect 6800 -1604 6840 -1556
rect 6800 -1636 6804 -1604
rect 6836 -1636 6840 -1604
rect 6800 -1684 6840 -1636
rect 6800 -1716 6804 -1684
rect 6836 -1716 6840 -1684
rect 6800 -1764 6840 -1716
rect 6800 -1796 6804 -1764
rect 6836 -1796 6840 -1764
rect 6800 -1844 6840 -1796
rect 6800 -1876 6804 -1844
rect 6836 -1876 6840 -1844
rect 6800 -1924 6840 -1876
rect 6800 -1956 6804 -1924
rect 6836 -1956 6840 -1924
rect 6800 -2004 6840 -1956
rect 6800 -2036 6804 -2004
rect 6836 -2036 6840 -2004
rect 6800 -2084 6840 -2036
rect 6800 -2116 6804 -2084
rect 6836 -2116 6840 -2084
rect 6800 -2164 6840 -2116
rect 6800 -2196 6804 -2164
rect 6836 -2196 6840 -2164
rect 6800 -2244 6840 -2196
rect 6800 -2276 6804 -2244
rect 6836 -2276 6840 -2244
rect 6800 -2324 6840 -2276
rect 6800 -2356 6804 -2324
rect 6836 -2356 6840 -2324
rect 6800 -2404 6840 -2356
rect 6800 -2436 6804 -2404
rect 6836 -2436 6840 -2404
rect 6800 -2484 6840 -2436
rect 6800 -2516 6804 -2484
rect 6836 -2516 6840 -2484
rect 6800 -2564 6840 -2516
rect 6800 -2596 6804 -2564
rect 6836 -2596 6840 -2564
rect 6800 -2644 6840 -2596
rect 6800 -2676 6804 -2644
rect 6836 -2676 6840 -2644
rect 6800 -2724 6840 -2676
rect 6800 -2756 6804 -2724
rect 6836 -2756 6840 -2724
rect 6800 -2804 6840 -2756
rect 6800 -2836 6804 -2804
rect 6836 -2836 6840 -2804
rect 6800 -2884 6840 -2836
rect 6800 -2916 6804 -2884
rect 6836 -2916 6840 -2884
rect 6800 -2964 6840 -2916
rect 6800 -2996 6804 -2964
rect 6836 -2996 6840 -2964
rect 6800 -3044 6840 -2996
rect 6800 -3076 6804 -3044
rect 6836 -3076 6840 -3044
rect 6800 -3124 6840 -3076
rect 6800 -3156 6804 -3124
rect 6836 -3156 6840 -3124
rect 6800 -3204 6840 -3156
rect 6800 -3236 6804 -3204
rect 6836 -3236 6840 -3204
rect 6800 -3284 6840 -3236
rect 6800 -3316 6804 -3284
rect 6836 -3316 6840 -3284
rect 6800 -3364 6840 -3316
rect 6800 -3396 6804 -3364
rect 6836 -3396 6840 -3364
rect 6800 -3444 6840 -3396
rect 6800 -3476 6804 -3444
rect 6836 -3476 6840 -3444
rect 6800 -3524 6840 -3476
rect 6800 -3556 6804 -3524
rect 6836 -3556 6840 -3524
rect 6800 -3604 6840 -3556
rect 6800 -3636 6804 -3604
rect 6836 -3636 6840 -3604
rect 6800 -3684 6840 -3636
rect 6800 -3716 6804 -3684
rect 6836 -3716 6840 -3684
rect 6800 -3720 6840 -3716
rect 6880 1036 6920 1040
rect 6880 1004 6884 1036
rect 6916 1004 6920 1036
rect 6880 956 6920 1004
rect 6880 924 6884 956
rect 6916 924 6920 956
rect 6880 876 6920 924
rect 6880 844 6884 876
rect 6916 844 6920 876
rect 6880 796 6920 844
rect 6880 764 6884 796
rect 6916 764 6920 796
rect 6880 716 6920 764
rect 6880 684 6884 716
rect 6916 684 6920 716
rect 6880 636 6920 684
rect 6880 604 6884 636
rect 6916 604 6920 636
rect 6880 556 6920 604
rect 6880 524 6884 556
rect 6916 524 6920 556
rect 6880 476 6920 524
rect 6880 444 6884 476
rect 6916 444 6920 476
rect 6880 396 6920 444
rect 6880 364 6884 396
rect 6916 364 6920 396
rect 6880 316 6920 364
rect 6880 284 6884 316
rect 6916 284 6920 316
rect 6880 236 6920 284
rect 6880 204 6884 236
rect 6916 204 6920 236
rect 6880 156 6920 204
rect 6880 124 6884 156
rect 6916 124 6920 156
rect 6880 76 6920 124
rect 6880 44 6884 76
rect 6916 44 6920 76
rect 6880 -4 6920 44
rect 6880 -36 6884 -4
rect 6916 -36 6920 -4
rect 6880 -84 6920 -36
rect 6880 -116 6884 -84
rect 6916 -116 6920 -84
rect 6880 -164 6920 -116
rect 6880 -196 6884 -164
rect 6916 -196 6920 -164
rect 6880 -244 6920 -196
rect 6880 -276 6884 -244
rect 6916 -276 6920 -244
rect 6880 -324 6920 -276
rect 6880 -356 6884 -324
rect 6916 -356 6920 -324
rect 6880 -404 6920 -356
rect 6880 -436 6884 -404
rect 6916 -436 6920 -404
rect 6880 -484 6920 -436
rect 6880 -516 6884 -484
rect 6916 -516 6920 -484
rect 6880 -564 6920 -516
rect 6880 -596 6884 -564
rect 6916 -596 6920 -564
rect 6880 -644 6920 -596
rect 6880 -676 6884 -644
rect 6916 -676 6920 -644
rect 6880 -724 6920 -676
rect 6880 -756 6884 -724
rect 6916 -756 6920 -724
rect 6880 -804 6920 -756
rect 6880 -836 6884 -804
rect 6916 -836 6920 -804
rect 6880 -884 6920 -836
rect 6880 -916 6884 -884
rect 6916 -916 6920 -884
rect 6880 -964 6920 -916
rect 6880 -996 6884 -964
rect 6916 -996 6920 -964
rect 6880 -1044 6920 -996
rect 6880 -1076 6884 -1044
rect 6916 -1076 6920 -1044
rect 6880 -1124 6920 -1076
rect 6880 -1156 6884 -1124
rect 6916 -1156 6920 -1124
rect 6880 -1204 6920 -1156
rect 6880 -1236 6884 -1204
rect 6916 -1236 6920 -1204
rect 6880 -1284 6920 -1236
rect 6880 -1316 6884 -1284
rect 6916 -1316 6920 -1284
rect 6880 -1364 6920 -1316
rect 6880 -1396 6884 -1364
rect 6916 -1396 6920 -1364
rect 6880 -1444 6920 -1396
rect 6880 -1476 6884 -1444
rect 6916 -1476 6920 -1444
rect 6880 -1524 6920 -1476
rect 6880 -1556 6884 -1524
rect 6916 -1556 6920 -1524
rect 6880 -1604 6920 -1556
rect 6880 -1636 6884 -1604
rect 6916 -1636 6920 -1604
rect 6880 -1684 6920 -1636
rect 6880 -1716 6884 -1684
rect 6916 -1716 6920 -1684
rect 6880 -1764 6920 -1716
rect 6880 -1796 6884 -1764
rect 6916 -1796 6920 -1764
rect 6880 -1844 6920 -1796
rect 6880 -1876 6884 -1844
rect 6916 -1876 6920 -1844
rect 6880 -1924 6920 -1876
rect 6880 -1956 6884 -1924
rect 6916 -1956 6920 -1924
rect 6880 -2004 6920 -1956
rect 6880 -2036 6884 -2004
rect 6916 -2036 6920 -2004
rect 6880 -2084 6920 -2036
rect 6880 -2116 6884 -2084
rect 6916 -2116 6920 -2084
rect 6880 -2164 6920 -2116
rect 6880 -2196 6884 -2164
rect 6916 -2196 6920 -2164
rect 6880 -2244 6920 -2196
rect 6880 -2276 6884 -2244
rect 6916 -2276 6920 -2244
rect 6880 -2324 6920 -2276
rect 6880 -2356 6884 -2324
rect 6916 -2356 6920 -2324
rect 6880 -2404 6920 -2356
rect 6880 -2436 6884 -2404
rect 6916 -2436 6920 -2404
rect 6880 -2484 6920 -2436
rect 6880 -2516 6884 -2484
rect 6916 -2516 6920 -2484
rect 6880 -2564 6920 -2516
rect 6880 -2596 6884 -2564
rect 6916 -2596 6920 -2564
rect 6880 -2644 6920 -2596
rect 6880 -2676 6884 -2644
rect 6916 -2676 6920 -2644
rect 6880 -2724 6920 -2676
rect 6880 -2756 6884 -2724
rect 6916 -2756 6920 -2724
rect 6880 -2804 6920 -2756
rect 6880 -2836 6884 -2804
rect 6916 -2836 6920 -2804
rect 6880 -2884 6920 -2836
rect 6880 -2916 6884 -2884
rect 6916 -2916 6920 -2884
rect 6880 -2964 6920 -2916
rect 6880 -2996 6884 -2964
rect 6916 -2996 6920 -2964
rect 6880 -3044 6920 -2996
rect 6880 -3076 6884 -3044
rect 6916 -3076 6920 -3044
rect 6880 -3124 6920 -3076
rect 6880 -3156 6884 -3124
rect 6916 -3156 6920 -3124
rect 6880 -3204 6920 -3156
rect 6880 -3236 6884 -3204
rect 6916 -3236 6920 -3204
rect 6880 -3284 6920 -3236
rect 6880 -3316 6884 -3284
rect 6916 -3316 6920 -3284
rect 6880 -3364 6920 -3316
rect 6880 -3396 6884 -3364
rect 6916 -3396 6920 -3364
rect 6880 -3444 6920 -3396
rect 6880 -3476 6884 -3444
rect 6916 -3476 6920 -3444
rect 6880 -3524 6920 -3476
rect 6880 -3556 6884 -3524
rect 6916 -3556 6920 -3524
rect 6880 -3604 6920 -3556
rect 6880 -3636 6884 -3604
rect 6916 -3636 6920 -3604
rect 6880 -3684 6920 -3636
rect 6880 -3716 6884 -3684
rect 6916 -3716 6920 -3684
rect 6880 -3720 6920 -3716
rect 6960 1036 7000 1040
rect 6960 1004 6964 1036
rect 6996 1004 7000 1036
rect 6960 956 7000 1004
rect 6960 924 6964 956
rect 6996 924 7000 956
rect 6960 876 7000 924
rect 6960 844 6964 876
rect 6996 844 7000 876
rect 6960 796 7000 844
rect 6960 764 6964 796
rect 6996 764 7000 796
rect 6960 716 7000 764
rect 6960 684 6964 716
rect 6996 684 7000 716
rect 6960 636 7000 684
rect 6960 604 6964 636
rect 6996 604 7000 636
rect 6960 556 7000 604
rect 6960 524 6964 556
rect 6996 524 7000 556
rect 6960 476 7000 524
rect 6960 444 6964 476
rect 6996 444 7000 476
rect 6960 396 7000 444
rect 6960 364 6964 396
rect 6996 364 7000 396
rect 6960 316 7000 364
rect 6960 284 6964 316
rect 6996 284 7000 316
rect 6960 236 7000 284
rect 6960 204 6964 236
rect 6996 204 7000 236
rect 6960 156 7000 204
rect 6960 124 6964 156
rect 6996 124 7000 156
rect 6960 76 7000 124
rect 6960 44 6964 76
rect 6996 44 7000 76
rect 6960 -4 7000 44
rect 6960 -36 6964 -4
rect 6996 -36 7000 -4
rect 6960 -84 7000 -36
rect 6960 -116 6964 -84
rect 6996 -116 7000 -84
rect 6960 -164 7000 -116
rect 6960 -196 6964 -164
rect 6996 -196 7000 -164
rect 6960 -244 7000 -196
rect 6960 -276 6964 -244
rect 6996 -276 7000 -244
rect 6960 -324 7000 -276
rect 6960 -356 6964 -324
rect 6996 -356 7000 -324
rect 6960 -404 7000 -356
rect 6960 -436 6964 -404
rect 6996 -436 7000 -404
rect 6960 -484 7000 -436
rect 6960 -516 6964 -484
rect 6996 -516 7000 -484
rect 6960 -564 7000 -516
rect 6960 -596 6964 -564
rect 6996 -596 7000 -564
rect 6960 -644 7000 -596
rect 6960 -676 6964 -644
rect 6996 -676 7000 -644
rect 6960 -724 7000 -676
rect 6960 -756 6964 -724
rect 6996 -756 7000 -724
rect 6960 -804 7000 -756
rect 6960 -836 6964 -804
rect 6996 -836 7000 -804
rect 6960 -884 7000 -836
rect 6960 -916 6964 -884
rect 6996 -916 7000 -884
rect 6960 -964 7000 -916
rect 6960 -996 6964 -964
rect 6996 -996 7000 -964
rect 6960 -1044 7000 -996
rect 6960 -1076 6964 -1044
rect 6996 -1076 7000 -1044
rect 6960 -1124 7000 -1076
rect 6960 -1156 6964 -1124
rect 6996 -1156 7000 -1124
rect 6960 -1204 7000 -1156
rect 6960 -1236 6964 -1204
rect 6996 -1236 7000 -1204
rect 6960 -1284 7000 -1236
rect 6960 -1316 6964 -1284
rect 6996 -1316 7000 -1284
rect 6960 -1364 7000 -1316
rect 6960 -1396 6964 -1364
rect 6996 -1396 7000 -1364
rect 6960 -1444 7000 -1396
rect 6960 -1476 6964 -1444
rect 6996 -1476 7000 -1444
rect 6960 -1524 7000 -1476
rect 6960 -1556 6964 -1524
rect 6996 -1556 7000 -1524
rect 6960 -1604 7000 -1556
rect 6960 -1636 6964 -1604
rect 6996 -1636 7000 -1604
rect 6960 -1684 7000 -1636
rect 6960 -1716 6964 -1684
rect 6996 -1716 7000 -1684
rect 6960 -1764 7000 -1716
rect 6960 -1796 6964 -1764
rect 6996 -1796 7000 -1764
rect 6960 -1844 7000 -1796
rect 6960 -1876 6964 -1844
rect 6996 -1876 7000 -1844
rect 6960 -1924 7000 -1876
rect 6960 -1956 6964 -1924
rect 6996 -1956 7000 -1924
rect 6960 -2004 7000 -1956
rect 6960 -2036 6964 -2004
rect 6996 -2036 7000 -2004
rect 6960 -2084 7000 -2036
rect 6960 -2116 6964 -2084
rect 6996 -2116 7000 -2084
rect 6960 -2164 7000 -2116
rect 6960 -2196 6964 -2164
rect 6996 -2196 7000 -2164
rect 6960 -2244 7000 -2196
rect 6960 -2276 6964 -2244
rect 6996 -2276 7000 -2244
rect 6960 -2324 7000 -2276
rect 6960 -2356 6964 -2324
rect 6996 -2356 7000 -2324
rect 6960 -2404 7000 -2356
rect 6960 -2436 6964 -2404
rect 6996 -2436 7000 -2404
rect 6960 -2484 7000 -2436
rect 6960 -2516 6964 -2484
rect 6996 -2516 7000 -2484
rect 6960 -2564 7000 -2516
rect 6960 -2596 6964 -2564
rect 6996 -2596 7000 -2564
rect 6960 -2644 7000 -2596
rect 6960 -2676 6964 -2644
rect 6996 -2676 7000 -2644
rect 6960 -2724 7000 -2676
rect 6960 -2756 6964 -2724
rect 6996 -2756 7000 -2724
rect 6960 -2804 7000 -2756
rect 6960 -2836 6964 -2804
rect 6996 -2836 7000 -2804
rect 6960 -2884 7000 -2836
rect 6960 -2916 6964 -2884
rect 6996 -2916 7000 -2884
rect 6960 -2964 7000 -2916
rect 6960 -2996 6964 -2964
rect 6996 -2996 7000 -2964
rect 6960 -3044 7000 -2996
rect 6960 -3076 6964 -3044
rect 6996 -3076 7000 -3044
rect 6960 -3124 7000 -3076
rect 6960 -3156 6964 -3124
rect 6996 -3156 7000 -3124
rect 6960 -3204 7000 -3156
rect 6960 -3236 6964 -3204
rect 6996 -3236 7000 -3204
rect 6960 -3284 7000 -3236
rect 6960 -3316 6964 -3284
rect 6996 -3316 7000 -3284
rect 6960 -3364 7000 -3316
rect 6960 -3396 6964 -3364
rect 6996 -3396 7000 -3364
rect 6960 -3444 7000 -3396
rect 6960 -3476 6964 -3444
rect 6996 -3476 7000 -3444
rect 6960 -3524 7000 -3476
rect 6960 -3556 6964 -3524
rect 6996 -3556 7000 -3524
rect 6960 -3604 7000 -3556
rect 6960 -3636 6964 -3604
rect 6996 -3636 7000 -3604
rect 6960 -3684 7000 -3636
rect 6960 -3716 6964 -3684
rect 6996 -3716 7000 -3684
rect 6960 -3720 7000 -3716
rect 7040 1036 7080 1040
rect 7040 1004 7044 1036
rect 7076 1004 7080 1036
rect 7040 956 7080 1004
rect 7040 924 7044 956
rect 7076 924 7080 956
rect 7040 876 7080 924
rect 7040 844 7044 876
rect 7076 844 7080 876
rect 7040 796 7080 844
rect 7040 764 7044 796
rect 7076 764 7080 796
rect 7040 716 7080 764
rect 7040 684 7044 716
rect 7076 684 7080 716
rect 7040 636 7080 684
rect 7040 604 7044 636
rect 7076 604 7080 636
rect 7040 556 7080 604
rect 7040 524 7044 556
rect 7076 524 7080 556
rect 7040 476 7080 524
rect 7040 444 7044 476
rect 7076 444 7080 476
rect 7040 396 7080 444
rect 7040 364 7044 396
rect 7076 364 7080 396
rect 7040 316 7080 364
rect 7040 284 7044 316
rect 7076 284 7080 316
rect 7040 236 7080 284
rect 7040 204 7044 236
rect 7076 204 7080 236
rect 7040 156 7080 204
rect 7040 124 7044 156
rect 7076 124 7080 156
rect 7040 76 7080 124
rect 7040 44 7044 76
rect 7076 44 7080 76
rect 7040 -4 7080 44
rect 7040 -36 7044 -4
rect 7076 -36 7080 -4
rect 7040 -84 7080 -36
rect 7040 -116 7044 -84
rect 7076 -116 7080 -84
rect 7040 -164 7080 -116
rect 7040 -196 7044 -164
rect 7076 -196 7080 -164
rect 7040 -244 7080 -196
rect 7040 -276 7044 -244
rect 7076 -276 7080 -244
rect 7040 -324 7080 -276
rect 7040 -356 7044 -324
rect 7076 -356 7080 -324
rect 7040 -404 7080 -356
rect 7040 -436 7044 -404
rect 7076 -436 7080 -404
rect 7040 -484 7080 -436
rect 7040 -516 7044 -484
rect 7076 -516 7080 -484
rect 7040 -564 7080 -516
rect 7040 -596 7044 -564
rect 7076 -596 7080 -564
rect 7040 -644 7080 -596
rect 7040 -676 7044 -644
rect 7076 -676 7080 -644
rect 7040 -724 7080 -676
rect 7040 -756 7044 -724
rect 7076 -756 7080 -724
rect 7040 -804 7080 -756
rect 7040 -836 7044 -804
rect 7076 -836 7080 -804
rect 7040 -884 7080 -836
rect 7040 -916 7044 -884
rect 7076 -916 7080 -884
rect 7040 -964 7080 -916
rect 7040 -996 7044 -964
rect 7076 -996 7080 -964
rect 7040 -1044 7080 -996
rect 7040 -1076 7044 -1044
rect 7076 -1076 7080 -1044
rect 7040 -1124 7080 -1076
rect 7040 -1156 7044 -1124
rect 7076 -1156 7080 -1124
rect 7040 -1204 7080 -1156
rect 7040 -1236 7044 -1204
rect 7076 -1236 7080 -1204
rect 7040 -1284 7080 -1236
rect 7040 -1316 7044 -1284
rect 7076 -1316 7080 -1284
rect 7040 -1364 7080 -1316
rect 7040 -1396 7044 -1364
rect 7076 -1396 7080 -1364
rect 7040 -1444 7080 -1396
rect 7040 -1476 7044 -1444
rect 7076 -1476 7080 -1444
rect 7040 -1524 7080 -1476
rect 7040 -1556 7044 -1524
rect 7076 -1556 7080 -1524
rect 7040 -1604 7080 -1556
rect 7040 -1636 7044 -1604
rect 7076 -1636 7080 -1604
rect 7040 -1684 7080 -1636
rect 7040 -1716 7044 -1684
rect 7076 -1716 7080 -1684
rect 7040 -1764 7080 -1716
rect 7040 -1796 7044 -1764
rect 7076 -1796 7080 -1764
rect 7040 -1844 7080 -1796
rect 7040 -1876 7044 -1844
rect 7076 -1876 7080 -1844
rect 7040 -1924 7080 -1876
rect 7040 -1956 7044 -1924
rect 7076 -1956 7080 -1924
rect 7040 -2004 7080 -1956
rect 7040 -2036 7044 -2004
rect 7076 -2036 7080 -2004
rect 7040 -2084 7080 -2036
rect 7040 -2116 7044 -2084
rect 7076 -2116 7080 -2084
rect 7040 -2164 7080 -2116
rect 7040 -2196 7044 -2164
rect 7076 -2196 7080 -2164
rect 7040 -2244 7080 -2196
rect 7040 -2276 7044 -2244
rect 7076 -2276 7080 -2244
rect 7040 -2324 7080 -2276
rect 7040 -2356 7044 -2324
rect 7076 -2356 7080 -2324
rect 7040 -2404 7080 -2356
rect 7040 -2436 7044 -2404
rect 7076 -2436 7080 -2404
rect 7040 -2484 7080 -2436
rect 7040 -2516 7044 -2484
rect 7076 -2516 7080 -2484
rect 7040 -2564 7080 -2516
rect 7040 -2596 7044 -2564
rect 7076 -2596 7080 -2564
rect 7040 -2644 7080 -2596
rect 7040 -2676 7044 -2644
rect 7076 -2676 7080 -2644
rect 7040 -2724 7080 -2676
rect 7040 -2756 7044 -2724
rect 7076 -2756 7080 -2724
rect 7040 -2804 7080 -2756
rect 7040 -2836 7044 -2804
rect 7076 -2836 7080 -2804
rect 7040 -2884 7080 -2836
rect 7040 -2916 7044 -2884
rect 7076 -2916 7080 -2884
rect 7040 -2964 7080 -2916
rect 7040 -2996 7044 -2964
rect 7076 -2996 7080 -2964
rect 7040 -3044 7080 -2996
rect 7040 -3076 7044 -3044
rect 7076 -3076 7080 -3044
rect 7040 -3124 7080 -3076
rect 7040 -3156 7044 -3124
rect 7076 -3156 7080 -3124
rect 7040 -3204 7080 -3156
rect 7040 -3236 7044 -3204
rect 7076 -3236 7080 -3204
rect 7040 -3284 7080 -3236
rect 7040 -3316 7044 -3284
rect 7076 -3316 7080 -3284
rect 7040 -3364 7080 -3316
rect 7040 -3396 7044 -3364
rect 7076 -3396 7080 -3364
rect 7040 -3444 7080 -3396
rect 7040 -3476 7044 -3444
rect 7076 -3476 7080 -3444
rect 7040 -3524 7080 -3476
rect 7040 -3556 7044 -3524
rect 7076 -3556 7080 -3524
rect 7040 -3604 7080 -3556
rect 7040 -3636 7044 -3604
rect 7076 -3636 7080 -3604
rect 7040 -3684 7080 -3636
rect 7040 -3716 7044 -3684
rect 7076 -3716 7080 -3684
rect 7040 -3720 7080 -3716
rect 7120 1036 7160 1040
rect 7120 1004 7124 1036
rect 7156 1004 7160 1036
rect 7120 956 7160 1004
rect 7120 924 7124 956
rect 7156 924 7160 956
rect 7120 876 7160 924
rect 7120 844 7124 876
rect 7156 844 7160 876
rect 7120 796 7160 844
rect 7120 764 7124 796
rect 7156 764 7160 796
rect 7120 716 7160 764
rect 7120 684 7124 716
rect 7156 684 7160 716
rect 7120 636 7160 684
rect 7120 604 7124 636
rect 7156 604 7160 636
rect 7120 556 7160 604
rect 7120 524 7124 556
rect 7156 524 7160 556
rect 7120 476 7160 524
rect 7120 444 7124 476
rect 7156 444 7160 476
rect 7120 396 7160 444
rect 7120 364 7124 396
rect 7156 364 7160 396
rect 7120 316 7160 364
rect 7120 284 7124 316
rect 7156 284 7160 316
rect 7120 236 7160 284
rect 7120 204 7124 236
rect 7156 204 7160 236
rect 7120 156 7160 204
rect 7120 124 7124 156
rect 7156 124 7160 156
rect 7120 76 7160 124
rect 7120 44 7124 76
rect 7156 44 7160 76
rect 7120 -4 7160 44
rect 7120 -36 7124 -4
rect 7156 -36 7160 -4
rect 7120 -84 7160 -36
rect 7120 -116 7124 -84
rect 7156 -116 7160 -84
rect 7120 -164 7160 -116
rect 7120 -196 7124 -164
rect 7156 -196 7160 -164
rect 7120 -244 7160 -196
rect 7120 -276 7124 -244
rect 7156 -276 7160 -244
rect 7120 -324 7160 -276
rect 7120 -356 7124 -324
rect 7156 -356 7160 -324
rect 7120 -404 7160 -356
rect 7120 -436 7124 -404
rect 7156 -436 7160 -404
rect 7120 -484 7160 -436
rect 7120 -516 7124 -484
rect 7156 -516 7160 -484
rect 7120 -564 7160 -516
rect 7120 -596 7124 -564
rect 7156 -596 7160 -564
rect 7120 -644 7160 -596
rect 7120 -676 7124 -644
rect 7156 -676 7160 -644
rect 7120 -724 7160 -676
rect 7120 -756 7124 -724
rect 7156 -756 7160 -724
rect 7120 -804 7160 -756
rect 7120 -836 7124 -804
rect 7156 -836 7160 -804
rect 7120 -884 7160 -836
rect 7120 -916 7124 -884
rect 7156 -916 7160 -884
rect 7120 -964 7160 -916
rect 7120 -996 7124 -964
rect 7156 -996 7160 -964
rect 7120 -1044 7160 -996
rect 7120 -1076 7124 -1044
rect 7156 -1076 7160 -1044
rect 7120 -1124 7160 -1076
rect 7120 -1156 7124 -1124
rect 7156 -1156 7160 -1124
rect 7120 -1204 7160 -1156
rect 7120 -1236 7124 -1204
rect 7156 -1236 7160 -1204
rect 7120 -1284 7160 -1236
rect 7120 -1316 7124 -1284
rect 7156 -1316 7160 -1284
rect 7120 -1364 7160 -1316
rect 7120 -1396 7124 -1364
rect 7156 -1396 7160 -1364
rect 7120 -1444 7160 -1396
rect 7120 -1476 7124 -1444
rect 7156 -1476 7160 -1444
rect 7120 -1524 7160 -1476
rect 7120 -1556 7124 -1524
rect 7156 -1556 7160 -1524
rect 7120 -1604 7160 -1556
rect 7120 -1636 7124 -1604
rect 7156 -1636 7160 -1604
rect 7120 -1684 7160 -1636
rect 7120 -1716 7124 -1684
rect 7156 -1716 7160 -1684
rect 7120 -1764 7160 -1716
rect 7120 -1796 7124 -1764
rect 7156 -1796 7160 -1764
rect 7120 -1844 7160 -1796
rect 7120 -1876 7124 -1844
rect 7156 -1876 7160 -1844
rect 7120 -1924 7160 -1876
rect 7120 -1956 7124 -1924
rect 7156 -1956 7160 -1924
rect 7120 -2004 7160 -1956
rect 7120 -2036 7124 -2004
rect 7156 -2036 7160 -2004
rect 7120 -2084 7160 -2036
rect 7120 -2116 7124 -2084
rect 7156 -2116 7160 -2084
rect 7120 -2164 7160 -2116
rect 7120 -2196 7124 -2164
rect 7156 -2196 7160 -2164
rect 7120 -2244 7160 -2196
rect 7120 -2276 7124 -2244
rect 7156 -2276 7160 -2244
rect 7120 -2324 7160 -2276
rect 7120 -2356 7124 -2324
rect 7156 -2356 7160 -2324
rect 7120 -2404 7160 -2356
rect 7120 -2436 7124 -2404
rect 7156 -2436 7160 -2404
rect 7120 -2484 7160 -2436
rect 7120 -2516 7124 -2484
rect 7156 -2516 7160 -2484
rect 7120 -2564 7160 -2516
rect 7120 -2596 7124 -2564
rect 7156 -2596 7160 -2564
rect 7120 -2644 7160 -2596
rect 7120 -2676 7124 -2644
rect 7156 -2676 7160 -2644
rect 7120 -2724 7160 -2676
rect 7120 -2756 7124 -2724
rect 7156 -2756 7160 -2724
rect 7120 -2804 7160 -2756
rect 7120 -2836 7124 -2804
rect 7156 -2836 7160 -2804
rect 7120 -2884 7160 -2836
rect 7120 -2916 7124 -2884
rect 7156 -2916 7160 -2884
rect 7120 -2964 7160 -2916
rect 7120 -2996 7124 -2964
rect 7156 -2996 7160 -2964
rect 7120 -3044 7160 -2996
rect 7120 -3076 7124 -3044
rect 7156 -3076 7160 -3044
rect 7120 -3124 7160 -3076
rect 7120 -3156 7124 -3124
rect 7156 -3156 7160 -3124
rect 7120 -3204 7160 -3156
rect 7120 -3236 7124 -3204
rect 7156 -3236 7160 -3204
rect 7120 -3284 7160 -3236
rect 7120 -3316 7124 -3284
rect 7156 -3316 7160 -3284
rect 7120 -3364 7160 -3316
rect 7120 -3396 7124 -3364
rect 7156 -3396 7160 -3364
rect 7120 -3444 7160 -3396
rect 7120 -3476 7124 -3444
rect 7156 -3476 7160 -3444
rect 7120 -3524 7160 -3476
rect 7120 -3556 7124 -3524
rect 7156 -3556 7160 -3524
rect 7120 -3604 7160 -3556
rect 7120 -3636 7124 -3604
rect 7156 -3636 7160 -3604
rect 7120 -3684 7160 -3636
rect 7120 -3716 7124 -3684
rect 7156 -3716 7160 -3684
rect 7120 -3720 7160 -3716
rect 7200 1036 7240 1040
rect 7200 1004 7204 1036
rect 7236 1004 7240 1036
rect 7200 956 7240 1004
rect 7200 924 7204 956
rect 7236 924 7240 956
rect 7200 876 7240 924
rect 7200 844 7204 876
rect 7236 844 7240 876
rect 7200 796 7240 844
rect 7200 764 7204 796
rect 7236 764 7240 796
rect 7200 716 7240 764
rect 7200 684 7204 716
rect 7236 684 7240 716
rect 7200 636 7240 684
rect 7200 604 7204 636
rect 7236 604 7240 636
rect 7200 556 7240 604
rect 7200 524 7204 556
rect 7236 524 7240 556
rect 7200 476 7240 524
rect 7200 444 7204 476
rect 7236 444 7240 476
rect 7200 396 7240 444
rect 7200 364 7204 396
rect 7236 364 7240 396
rect 7200 316 7240 364
rect 7200 284 7204 316
rect 7236 284 7240 316
rect 7200 236 7240 284
rect 7200 204 7204 236
rect 7236 204 7240 236
rect 7200 156 7240 204
rect 7200 124 7204 156
rect 7236 124 7240 156
rect 7200 76 7240 124
rect 7200 44 7204 76
rect 7236 44 7240 76
rect 7200 -4 7240 44
rect 7200 -36 7204 -4
rect 7236 -36 7240 -4
rect 7200 -84 7240 -36
rect 7200 -116 7204 -84
rect 7236 -116 7240 -84
rect 7200 -164 7240 -116
rect 7200 -196 7204 -164
rect 7236 -196 7240 -164
rect 7200 -244 7240 -196
rect 7200 -276 7204 -244
rect 7236 -276 7240 -244
rect 7200 -324 7240 -276
rect 7200 -356 7204 -324
rect 7236 -356 7240 -324
rect 7200 -404 7240 -356
rect 7200 -436 7204 -404
rect 7236 -436 7240 -404
rect 7200 -484 7240 -436
rect 7200 -516 7204 -484
rect 7236 -516 7240 -484
rect 7200 -564 7240 -516
rect 7200 -596 7204 -564
rect 7236 -596 7240 -564
rect 7200 -644 7240 -596
rect 7200 -676 7204 -644
rect 7236 -676 7240 -644
rect 7200 -724 7240 -676
rect 7200 -756 7204 -724
rect 7236 -756 7240 -724
rect 7200 -804 7240 -756
rect 7200 -836 7204 -804
rect 7236 -836 7240 -804
rect 7200 -884 7240 -836
rect 7200 -916 7204 -884
rect 7236 -916 7240 -884
rect 7200 -964 7240 -916
rect 7200 -996 7204 -964
rect 7236 -996 7240 -964
rect 7200 -1044 7240 -996
rect 7200 -1076 7204 -1044
rect 7236 -1076 7240 -1044
rect 7200 -1124 7240 -1076
rect 7200 -1156 7204 -1124
rect 7236 -1156 7240 -1124
rect 7200 -1204 7240 -1156
rect 7200 -1236 7204 -1204
rect 7236 -1236 7240 -1204
rect 7200 -1284 7240 -1236
rect 7200 -1316 7204 -1284
rect 7236 -1316 7240 -1284
rect 7200 -1364 7240 -1316
rect 7200 -1396 7204 -1364
rect 7236 -1396 7240 -1364
rect 7200 -1444 7240 -1396
rect 7200 -1476 7204 -1444
rect 7236 -1476 7240 -1444
rect 7200 -1524 7240 -1476
rect 7200 -1556 7204 -1524
rect 7236 -1556 7240 -1524
rect 7200 -1604 7240 -1556
rect 7200 -1636 7204 -1604
rect 7236 -1636 7240 -1604
rect 7200 -1684 7240 -1636
rect 7200 -1716 7204 -1684
rect 7236 -1716 7240 -1684
rect 7200 -1764 7240 -1716
rect 7200 -1796 7204 -1764
rect 7236 -1796 7240 -1764
rect 7200 -1844 7240 -1796
rect 7200 -1876 7204 -1844
rect 7236 -1876 7240 -1844
rect 7200 -1924 7240 -1876
rect 7200 -1956 7204 -1924
rect 7236 -1956 7240 -1924
rect 7200 -2004 7240 -1956
rect 7200 -2036 7204 -2004
rect 7236 -2036 7240 -2004
rect 7200 -2084 7240 -2036
rect 7200 -2116 7204 -2084
rect 7236 -2116 7240 -2084
rect 7200 -2164 7240 -2116
rect 7200 -2196 7204 -2164
rect 7236 -2196 7240 -2164
rect 7200 -2244 7240 -2196
rect 7200 -2276 7204 -2244
rect 7236 -2276 7240 -2244
rect 7200 -2324 7240 -2276
rect 7200 -2356 7204 -2324
rect 7236 -2356 7240 -2324
rect 7200 -2404 7240 -2356
rect 7200 -2436 7204 -2404
rect 7236 -2436 7240 -2404
rect 7200 -2484 7240 -2436
rect 7200 -2516 7204 -2484
rect 7236 -2516 7240 -2484
rect 7200 -2564 7240 -2516
rect 7200 -2596 7204 -2564
rect 7236 -2596 7240 -2564
rect 7200 -2644 7240 -2596
rect 7200 -2676 7204 -2644
rect 7236 -2676 7240 -2644
rect 7200 -2724 7240 -2676
rect 7200 -2756 7204 -2724
rect 7236 -2756 7240 -2724
rect 7200 -2804 7240 -2756
rect 7200 -2836 7204 -2804
rect 7236 -2836 7240 -2804
rect 7200 -2884 7240 -2836
rect 7200 -2916 7204 -2884
rect 7236 -2916 7240 -2884
rect 7200 -2964 7240 -2916
rect 7200 -2996 7204 -2964
rect 7236 -2996 7240 -2964
rect 7200 -3044 7240 -2996
rect 7200 -3076 7204 -3044
rect 7236 -3076 7240 -3044
rect 7200 -3124 7240 -3076
rect 7200 -3156 7204 -3124
rect 7236 -3156 7240 -3124
rect 7200 -3204 7240 -3156
rect 7200 -3236 7204 -3204
rect 7236 -3236 7240 -3204
rect 7200 -3284 7240 -3236
rect 7200 -3316 7204 -3284
rect 7236 -3316 7240 -3284
rect 7200 -3364 7240 -3316
rect 7200 -3396 7204 -3364
rect 7236 -3396 7240 -3364
rect 7200 -3444 7240 -3396
rect 7200 -3476 7204 -3444
rect 7236 -3476 7240 -3444
rect 7200 -3524 7240 -3476
rect 7200 -3556 7204 -3524
rect 7236 -3556 7240 -3524
rect 7200 -3604 7240 -3556
rect 7200 -3636 7204 -3604
rect 7236 -3636 7240 -3604
rect 7200 -3684 7240 -3636
rect 7200 -3716 7204 -3684
rect 7236 -3716 7240 -3684
rect 7200 -3720 7240 -3716
rect 7280 1036 7320 1040
rect 7280 1004 7284 1036
rect 7316 1004 7320 1036
rect 7280 956 7320 1004
rect 7280 924 7284 956
rect 7316 924 7320 956
rect 7280 876 7320 924
rect 7280 844 7284 876
rect 7316 844 7320 876
rect 7280 796 7320 844
rect 7280 764 7284 796
rect 7316 764 7320 796
rect 7280 716 7320 764
rect 7280 684 7284 716
rect 7316 684 7320 716
rect 7280 636 7320 684
rect 7280 604 7284 636
rect 7316 604 7320 636
rect 7280 556 7320 604
rect 7280 524 7284 556
rect 7316 524 7320 556
rect 7280 476 7320 524
rect 7280 444 7284 476
rect 7316 444 7320 476
rect 7280 396 7320 444
rect 7280 364 7284 396
rect 7316 364 7320 396
rect 7280 316 7320 364
rect 7280 284 7284 316
rect 7316 284 7320 316
rect 7280 236 7320 284
rect 7280 204 7284 236
rect 7316 204 7320 236
rect 7280 156 7320 204
rect 7280 124 7284 156
rect 7316 124 7320 156
rect 7280 76 7320 124
rect 7280 44 7284 76
rect 7316 44 7320 76
rect 7280 -4 7320 44
rect 7280 -36 7284 -4
rect 7316 -36 7320 -4
rect 7280 -84 7320 -36
rect 7280 -116 7284 -84
rect 7316 -116 7320 -84
rect 7280 -164 7320 -116
rect 7280 -196 7284 -164
rect 7316 -196 7320 -164
rect 7280 -244 7320 -196
rect 7280 -276 7284 -244
rect 7316 -276 7320 -244
rect 7280 -324 7320 -276
rect 7280 -356 7284 -324
rect 7316 -356 7320 -324
rect 7280 -404 7320 -356
rect 7280 -436 7284 -404
rect 7316 -436 7320 -404
rect 7280 -484 7320 -436
rect 7280 -516 7284 -484
rect 7316 -516 7320 -484
rect 7280 -564 7320 -516
rect 7280 -596 7284 -564
rect 7316 -596 7320 -564
rect 7280 -644 7320 -596
rect 7280 -676 7284 -644
rect 7316 -676 7320 -644
rect 7280 -724 7320 -676
rect 7280 -756 7284 -724
rect 7316 -756 7320 -724
rect 7280 -804 7320 -756
rect 7280 -836 7284 -804
rect 7316 -836 7320 -804
rect 7280 -884 7320 -836
rect 7280 -916 7284 -884
rect 7316 -916 7320 -884
rect 7280 -964 7320 -916
rect 7280 -996 7284 -964
rect 7316 -996 7320 -964
rect 7280 -1044 7320 -996
rect 7280 -1076 7284 -1044
rect 7316 -1076 7320 -1044
rect 7280 -1124 7320 -1076
rect 7280 -1156 7284 -1124
rect 7316 -1156 7320 -1124
rect 7280 -1204 7320 -1156
rect 7280 -1236 7284 -1204
rect 7316 -1236 7320 -1204
rect 7280 -1284 7320 -1236
rect 7280 -1316 7284 -1284
rect 7316 -1316 7320 -1284
rect 7280 -1364 7320 -1316
rect 7280 -1396 7284 -1364
rect 7316 -1396 7320 -1364
rect 7280 -1444 7320 -1396
rect 7280 -1476 7284 -1444
rect 7316 -1476 7320 -1444
rect 7280 -1524 7320 -1476
rect 7280 -1556 7284 -1524
rect 7316 -1556 7320 -1524
rect 7280 -1604 7320 -1556
rect 7280 -1636 7284 -1604
rect 7316 -1636 7320 -1604
rect 7280 -1684 7320 -1636
rect 7280 -1716 7284 -1684
rect 7316 -1716 7320 -1684
rect 7280 -1764 7320 -1716
rect 7280 -1796 7284 -1764
rect 7316 -1796 7320 -1764
rect 7280 -1844 7320 -1796
rect 7280 -1876 7284 -1844
rect 7316 -1876 7320 -1844
rect 7280 -1924 7320 -1876
rect 7280 -1956 7284 -1924
rect 7316 -1956 7320 -1924
rect 7280 -2004 7320 -1956
rect 7280 -2036 7284 -2004
rect 7316 -2036 7320 -2004
rect 7280 -2084 7320 -2036
rect 7280 -2116 7284 -2084
rect 7316 -2116 7320 -2084
rect 7280 -2164 7320 -2116
rect 7280 -2196 7284 -2164
rect 7316 -2196 7320 -2164
rect 7280 -2244 7320 -2196
rect 7280 -2276 7284 -2244
rect 7316 -2276 7320 -2244
rect 7280 -2324 7320 -2276
rect 7280 -2356 7284 -2324
rect 7316 -2356 7320 -2324
rect 7280 -2404 7320 -2356
rect 7280 -2436 7284 -2404
rect 7316 -2436 7320 -2404
rect 7280 -2484 7320 -2436
rect 7280 -2516 7284 -2484
rect 7316 -2516 7320 -2484
rect 7280 -2564 7320 -2516
rect 7280 -2596 7284 -2564
rect 7316 -2596 7320 -2564
rect 7280 -2644 7320 -2596
rect 7280 -2676 7284 -2644
rect 7316 -2676 7320 -2644
rect 7280 -2724 7320 -2676
rect 7280 -2756 7284 -2724
rect 7316 -2756 7320 -2724
rect 7280 -2804 7320 -2756
rect 7280 -2836 7284 -2804
rect 7316 -2836 7320 -2804
rect 7280 -2884 7320 -2836
rect 7280 -2916 7284 -2884
rect 7316 -2916 7320 -2884
rect 7280 -2964 7320 -2916
rect 7280 -2996 7284 -2964
rect 7316 -2996 7320 -2964
rect 7280 -3044 7320 -2996
rect 7280 -3076 7284 -3044
rect 7316 -3076 7320 -3044
rect 7280 -3124 7320 -3076
rect 7280 -3156 7284 -3124
rect 7316 -3156 7320 -3124
rect 7280 -3204 7320 -3156
rect 7280 -3236 7284 -3204
rect 7316 -3236 7320 -3204
rect 7280 -3284 7320 -3236
rect 7280 -3316 7284 -3284
rect 7316 -3316 7320 -3284
rect 7280 -3364 7320 -3316
rect 7280 -3396 7284 -3364
rect 7316 -3396 7320 -3364
rect 7280 -3444 7320 -3396
rect 7280 -3476 7284 -3444
rect 7316 -3476 7320 -3444
rect 7280 -3524 7320 -3476
rect 7280 -3556 7284 -3524
rect 7316 -3556 7320 -3524
rect 7280 -3604 7320 -3556
rect 7280 -3636 7284 -3604
rect 7316 -3636 7320 -3604
rect 7280 -3684 7320 -3636
rect 7280 -3716 7284 -3684
rect 7316 -3716 7320 -3684
rect 7280 -3720 7320 -3716
rect 7360 1036 7400 1040
rect 7360 1004 7364 1036
rect 7396 1004 7400 1036
rect 7360 956 7400 1004
rect 7360 924 7364 956
rect 7396 924 7400 956
rect 7360 876 7400 924
rect 7360 844 7364 876
rect 7396 844 7400 876
rect 7360 796 7400 844
rect 7360 764 7364 796
rect 7396 764 7400 796
rect 7360 716 7400 764
rect 7360 684 7364 716
rect 7396 684 7400 716
rect 7360 636 7400 684
rect 7360 604 7364 636
rect 7396 604 7400 636
rect 7360 556 7400 604
rect 7360 524 7364 556
rect 7396 524 7400 556
rect 7360 476 7400 524
rect 7360 444 7364 476
rect 7396 444 7400 476
rect 7360 396 7400 444
rect 7360 364 7364 396
rect 7396 364 7400 396
rect 7360 316 7400 364
rect 7360 284 7364 316
rect 7396 284 7400 316
rect 7360 236 7400 284
rect 7360 204 7364 236
rect 7396 204 7400 236
rect 7360 156 7400 204
rect 7360 124 7364 156
rect 7396 124 7400 156
rect 7360 76 7400 124
rect 7360 44 7364 76
rect 7396 44 7400 76
rect 7360 -4 7400 44
rect 7360 -36 7364 -4
rect 7396 -36 7400 -4
rect 7360 -84 7400 -36
rect 7360 -116 7364 -84
rect 7396 -116 7400 -84
rect 7360 -164 7400 -116
rect 7360 -196 7364 -164
rect 7396 -196 7400 -164
rect 7360 -244 7400 -196
rect 7360 -276 7364 -244
rect 7396 -276 7400 -244
rect 7360 -324 7400 -276
rect 7360 -356 7364 -324
rect 7396 -356 7400 -324
rect 7360 -404 7400 -356
rect 7360 -436 7364 -404
rect 7396 -436 7400 -404
rect 7360 -484 7400 -436
rect 7360 -516 7364 -484
rect 7396 -516 7400 -484
rect 7360 -564 7400 -516
rect 7360 -596 7364 -564
rect 7396 -596 7400 -564
rect 7360 -644 7400 -596
rect 7360 -676 7364 -644
rect 7396 -676 7400 -644
rect 7360 -724 7400 -676
rect 7360 -756 7364 -724
rect 7396 -756 7400 -724
rect 7360 -804 7400 -756
rect 7360 -836 7364 -804
rect 7396 -836 7400 -804
rect 7360 -884 7400 -836
rect 7360 -916 7364 -884
rect 7396 -916 7400 -884
rect 7360 -964 7400 -916
rect 7360 -996 7364 -964
rect 7396 -996 7400 -964
rect 7360 -1044 7400 -996
rect 7360 -1076 7364 -1044
rect 7396 -1076 7400 -1044
rect 7360 -1124 7400 -1076
rect 7360 -1156 7364 -1124
rect 7396 -1156 7400 -1124
rect 7360 -1204 7400 -1156
rect 7360 -1236 7364 -1204
rect 7396 -1236 7400 -1204
rect 7360 -1284 7400 -1236
rect 7360 -1316 7364 -1284
rect 7396 -1316 7400 -1284
rect 7360 -1364 7400 -1316
rect 7360 -1396 7364 -1364
rect 7396 -1396 7400 -1364
rect 7360 -1444 7400 -1396
rect 7360 -1476 7364 -1444
rect 7396 -1476 7400 -1444
rect 7360 -1524 7400 -1476
rect 7360 -1556 7364 -1524
rect 7396 -1556 7400 -1524
rect 7360 -1604 7400 -1556
rect 7360 -1636 7364 -1604
rect 7396 -1636 7400 -1604
rect 7360 -1684 7400 -1636
rect 7360 -1716 7364 -1684
rect 7396 -1716 7400 -1684
rect 7360 -1764 7400 -1716
rect 7360 -1796 7364 -1764
rect 7396 -1796 7400 -1764
rect 7360 -1844 7400 -1796
rect 7360 -1876 7364 -1844
rect 7396 -1876 7400 -1844
rect 7360 -1924 7400 -1876
rect 7360 -1956 7364 -1924
rect 7396 -1956 7400 -1924
rect 7360 -2004 7400 -1956
rect 7360 -2036 7364 -2004
rect 7396 -2036 7400 -2004
rect 7360 -2084 7400 -2036
rect 7360 -2116 7364 -2084
rect 7396 -2116 7400 -2084
rect 7360 -2164 7400 -2116
rect 7360 -2196 7364 -2164
rect 7396 -2196 7400 -2164
rect 7360 -2244 7400 -2196
rect 7360 -2276 7364 -2244
rect 7396 -2276 7400 -2244
rect 7360 -2324 7400 -2276
rect 7360 -2356 7364 -2324
rect 7396 -2356 7400 -2324
rect 7360 -2404 7400 -2356
rect 7360 -2436 7364 -2404
rect 7396 -2436 7400 -2404
rect 7360 -2484 7400 -2436
rect 7360 -2516 7364 -2484
rect 7396 -2516 7400 -2484
rect 7360 -2564 7400 -2516
rect 7360 -2596 7364 -2564
rect 7396 -2596 7400 -2564
rect 7360 -2644 7400 -2596
rect 7360 -2676 7364 -2644
rect 7396 -2676 7400 -2644
rect 7360 -2724 7400 -2676
rect 7360 -2756 7364 -2724
rect 7396 -2756 7400 -2724
rect 7360 -2804 7400 -2756
rect 7360 -2836 7364 -2804
rect 7396 -2836 7400 -2804
rect 7360 -2884 7400 -2836
rect 7360 -2916 7364 -2884
rect 7396 -2916 7400 -2884
rect 7360 -2964 7400 -2916
rect 7360 -2996 7364 -2964
rect 7396 -2996 7400 -2964
rect 7360 -3044 7400 -2996
rect 7360 -3076 7364 -3044
rect 7396 -3076 7400 -3044
rect 7360 -3124 7400 -3076
rect 7360 -3156 7364 -3124
rect 7396 -3156 7400 -3124
rect 7360 -3204 7400 -3156
rect 7360 -3236 7364 -3204
rect 7396 -3236 7400 -3204
rect 7360 -3284 7400 -3236
rect 7360 -3316 7364 -3284
rect 7396 -3316 7400 -3284
rect 7360 -3364 7400 -3316
rect 7360 -3396 7364 -3364
rect 7396 -3396 7400 -3364
rect 7360 -3444 7400 -3396
rect 7360 -3476 7364 -3444
rect 7396 -3476 7400 -3444
rect 7360 -3524 7400 -3476
rect 7360 -3556 7364 -3524
rect 7396 -3556 7400 -3524
rect 7360 -3604 7400 -3556
rect 7360 -3636 7364 -3604
rect 7396 -3636 7400 -3604
rect 7360 -3684 7400 -3636
rect 7360 -3716 7364 -3684
rect 7396 -3716 7400 -3684
rect 7360 -3720 7400 -3716
rect 7440 1036 7480 1040
rect 7440 1004 7444 1036
rect 7476 1004 7480 1036
rect 7440 956 7480 1004
rect 7440 924 7444 956
rect 7476 924 7480 956
rect 7440 876 7480 924
rect 7440 844 7444 876
rect 7476 844 7480 876
rect 7440 796 7480 844
rect 7440 764 7444 796
rect 7476 764 7480 796
rect 7440 716 7480 764
rect 7440 684 7444 716
rect 7476 684 7480 716
rect 7440 636 7480 684
rect 7440 604 7444 636
rect 7476 604 7480 636
rect 7440 556 7480 604
rect 7440 524 7444 556
rect 7476 524 7480 556
rect 7440 476 7480 524
rect 7440 444 7444 476
rect 7476 444 7480 476
rect 7440 396 7480 444
rect 7440 364 7444 396
rect 7476 364 7480 396
rect 7440 316 7480 364
rect 7440 284 7444 316
rect 7476 284 7480 316
rect 7440 236 7480 284
rect 7440 204 7444 236
rect 7476 204 7480 236
rect 7440 156 7480 204
rect 7440 124 7444 156
rect 7476 124 7480 156
rect 7440 76 7480 124
rect 7440 44 7444 76
rect 7476 44 7480 76
rect 7440 -4 7480 44
rect 7440 -36 7444 -4
rect 7476 -36 7480 -4
rect 7440 -84 7480 -36
rect 7440 -116 7444 -84
rect 7476 -116 7480 -84
rect 7440 -164 7480 -116
rect 7440 -196 7444 -164
rect 7476 -196 7480 -164
rect 7440 -244 7480 -196
rect 7440 -276 7444 -244
rect 7476 -276 7480 -244
rect 7440 -324 7480 -276
rect 7440 -356 7444 -324
rect 7476 -356 7480 -324
rect 7440 -404 7480 -356
rect 7440 -436 7444 -404
rect 7476 -436 7480 -404
rect 7440 -484 7480 -436
rect 7440 -516 7444 -484
rect 7476 -516 7480 -484
rect 7440 -564 7480 -516
rect 7440 -596 7444 -564
rect 7476 -596 7480 -564
rect 7440 -644 7480 -596
rect 7440 -676 7444 -644
rect 7476 -676 7480 -644
rect 7440 -724 7480 -676
rect 7440 -756 7444 -724
rect 7476 -756 7480 -724
rect 7440 -804 7480 -756
rect 7440 -836 7444 -804
rect 7476 -836 7480 -804
rect 7440 -884 7480 -836
rect 7440 -916 7444 -884
rect 7476 -916 7480 -884
rect 7440 -964 7480 -916
rect 7440 -996 7444 -964
rect 7476 -996 7480 -964
rect 7440 -1044 7480 -996
rect 7440 -1076 7444 -1044
rect 7476 -1076 7480 -1044
rect 7440 -1124 7480 -1076
rect 7440 -1156 7444 -1124
rect 7476 -1156 7480 -1124
rect 7440 -1204 7480 -1156
rect 7440 -1236 7444 -1204
rect 7476 -1236 7480 -1204
rect 7440 -1284 7480 -1236
rect 7440 -1316 7444 -1284
rect 7476 -1316 7480 -1284
rect 7440 -1364 7480 -1316
rect 7440 -1396 7444 -1364
rect 7476 -1396 7480 -1364
rect 7440 -1444 7480 -1396
rect 7440 -1476 7444 -1444
rect 7476 -1476 7480 -1444
rect 7440 -1524 7480 -1476
rect 7440 -1556 7444 -1524
rect 7476 -1556 7480 -1524
rect 7440 -1604 7480 -1556
rect 7440 -1636 7444 -1604
rect 7476 -1636 7480 -1604
rect 7440 -1684 7480 -1636
rect 7440 -1716 7444 -1684
rect 7476 -1716 7480 -1684
rect 7440 -1764 7480 -1716
rect 7440 -1796 7444 -1764
rect 7476 -1796 7480 -1764
rect 7440 -1844 7480 -1796
rect 7440 -1876 7444 -1844
rect 7476 -1876 7480 -1844
rect 7440 -1924 7480 -1876
rect 7440 -1956 7444 -1924
rect 7476 -1956 7480 -1924
rect 7440 -2004 7480 -1956
rect 7440 -2036 7444 -2004
rect 7476 -2036 7480 -2004
rect 7440 -2084 7480 -2036
rect 7440 -2116 7444 -2084
rect 7476 -2116 7480 -2084
rect 7440 -2164 7480 -2116
rect 7440 -2196 7444 -2164
rect 7476 -2196 7480 -2164
rect 7440 -2244 7480 -2196
rect 7440 -2276 7444 -2244
rect 7476 -2276 7480 -2244
rect 7440 -2324 7480 -2276
rect 7440 -2356 7444 -2324
rect 7476 -2356 7480 -2324
rect 7440 -2404 7480 -2356
rect 7440 -2436 7444 -2404
rect 7476 -2436 7480 -2404
rect 7440 -2484 7480 -2436
rect 7440 -2516 7444 -2484
rect 7476 -2516 7480 -2484
rect 7440 -2564 7480 -2516
rect 7440 -2596 7444 -2564
rect 7476 -2596 7480 -2564
rect 7440 -2644 7480 -2596
rect 7440 -2676 7444 -2644
rect 7476 -2676 7480 -2644
rect 7440 -2724 7480 -2676
rect 7440 -2756 7444 -2724
rect 7476 -2756 7480 -2724
rect 7440 -2804 7480 -2756
rect 7440 -2836 7444 -2804
rect 7476 -2836 7480 -2804
rect 7440 -2884 7480 -2836
rect 7440 -2916 7444 -2884
rect 7476 -2916 7480 -2884
rect 7440 -2964 7480 -2916
rect 7440 -2996 7444 -2964
rect 7476 -2996 7480 -2964
rect 7440 -3044 7480 -2996
rect 7440 -3076 7444 -3044
rect 7476 -3076 7480 -3044
rect 7440 -3124 7480 -3076
rect 7440 -3156 7444 -3124
rect 7476 -3156 7480 -3124
rect 7440 -3204 7480 -3156
rect 7440 -3236 7444 -3204
rect 7476 -3236 7480 -3204
rect 7440 -3284 7480 -3236
rect 7440 -3316 7444 -3284
rect 7476 -3316 7480 -3284
rect 7440 -3364 7480 -3316
rect 7440 -3396 7444 -3364
rect 7476 -3396 7480 -3364
rect 7440 -3444 7480 -3396
rect 7440 -3476 7444 -3444
rect 7476 -3476 7480 -3444
rect 7440 -3524 7480 -3476
rect 7440 -3556 7444 -3524
rect 7476 -3556 7480 -3524
rect 7440 -3604 7480 -3556
rect 7440 -3636 7444 -3604
rect 7476 -3636 7480 -3604
rect 7440 -3684 7480 -3636
rect 7440 -3716 7444 -3684
rect 7476 -3716 7480 -3684
rect 7440 -3720 7480 -3716
rect 7520 1036 7560 1040
rect 7520 1004 7524 1036
rect 7556 1004 7560 1036
rect 7520 956 7560 1004
rect 7520 924 7524 956
rect 7556 924 7560 956
rect 7520 876 7560 924
rect 7520 844 7524 876
rect 7556 844 7560 876
rect 7520 796 7560 844
rect 7520 764 7524 796
rect 7556 764 7560 796
rect 7520 716 7560 764
rect 7520 684 7524 716
rect 7556 684 7560 716
rect 7520 636 7560 684
rect 7520 604 7524 636
rect 7556 604 7560 636
rect 7520 556 7560 604
rect 7520 524 7524 556
rect 7556 524 7560 556
rect 7520 476 7560 524
rect 7520 444 7524 476
rect 7556 444 7560 476
rect 7520 396 7560 444
rect 7520 364 7524 396
rect 7556 364 7560 396
rect 7520 316 7560 364
rect 7520 284 7524 316
rect 7556 284 7560 316
rect 7520 236 7560 284
rect 7520 204 7524 236
rect 7556 204 7560 236
rect 7520 156 7560 204
rect 7520 124 7524 156
rect 7556 124 7560 156
rect 7520 76 7560 124
rect 7520 44 7524 76
rect 7556 44 7560 76
rect 7520 -4 7560 44
rect 7520 -36 7524 -4
rect 7556 -36 7560 -4
rect 7520 -84 7560 -36
rect 7520 -116 7524 -84
rect 7556 -116 7560 -84
rect 7520 -164 7560 -116
rect 7520 -196 7524 -164
rect 7556 -196 7560 -164
rect 7520 -244 7560 -196
rect 7520 -276 7524 -244
rect 7556 -276 7560 -244
rect 7520 -324 7560 -276
rect 7520 -356 7524 -324
rect 7556 -356 7560 -324
rect 7520 -404 7560 -356
rect 7520 -436 7524 -404
rect 7556 -436 7560 -404
rect 7520 -484 7560 -436
rect 7520 -516 7524 -484
rect 7556 -516 7560 -484
rect 7520 -564 7560 -516
rect 7520 -596 7524 -564
rect 7556 -596 7560 -564
rect 7520 -644 7560 -596
rect 7520 -676 7524 -644
rect 7556 -676 7560 -644
rect 7520 -724 7560 -676
rect 7520 -756 7524 -724
rect 7556 -756 7560 -724
rect 7520 -804 7560 -756
rect 7520 -836 7524 -804
rect 7556 -836 7560 -804
rect 7520 -884 7560 -836
rect 7520 -916 7524 -884
rect 7556 -916 7560 -884
rect 7520 -964 7560 -916
rect 7520 -996 7524 -964
rect 7556 -996 7560 -964
rect 7520 -1044 7560 -996
rect 7520 -1076 7524 -1044
rect 7556 -1076 7560 -1044
rect 7520 -1124 7560 -1076
rect 7520 -1156 7524 -1124
rect 7556 -1156 7560 -1124
rect 7520 -1204 7560 -1156
rect 7520 -1236 7524 -1204
rect 7556 -1236 7560 -1204
rect 7520 -1284 7560 -1236
rect 7520 -1316 7524 -1284
rect 7556 -1316 7560 -1284
rect 7520 -1364 7560 -1316
rect 7520 -1396 7524 -1364
rect 7556 -1396 7560 -1364
rect 7520 -1444 7560 -1396
rect 7520 -1476 7524 -1444
rect 7556 -1476 7560 -1444
rect 7520 -1524 7560 -1476
rect 7520 -1556 7524 -1524
rect 7556 -1556 7560 -1524
rect 7520 -1604 7560 -1556
rect 7520 -1636 7524 -1604
rect 7556 -1636 7560 -1604
rect 7520 -1684 7560 -1636
rect 7520 -1716 7524 -1684
rect 7556 -1716 7560 -1684
rect 7520 -1764 7560 -1716
rect 7520 -1796 7524 -1764
rect 7556 -1796 7560 -1764
rect 7520 -1844 7560 -1796
rect 7520 -1876 7524 -1844
rect 7556 -1876 7560 -1844
rect 7520 -1924 7560 -1876
rect 7520 -1956 7524 -1924
rect 7556 -1956 7560 -1924
rect 7520 -2004 7560 -1956
rect 7520 -2036 7524 -2004
rect 7556 -2036 7560 -2004
rect 7520 -2084 7560 -2036
rect 7520 -2116 7524 -2084
rect 7556 -2116 7560 -2084
rect 7520 -2164 7560 -2116
rect 7520 -2196 7524 -2164
rect 7556 -2196 7560 -2164
rect 7520 -2244 7560 -2196
rect 7520 -2276 7524 -2244
rect 7556 -2276 7560 -2244
rect 7520 -2324 7560 -2276
rect 7520 -2356 7524 -2324
rect 7556 -2356 7560 -2324
rect 7520 -2404 7560 -2356
rect 7520 -2436 7524 -2404
rect 7556 -2436 7560 -2404
rect 7520 -2484 7560 -2436
rect 7520 -2516 7524 -2484
rect 7556 -2516 7560 -2484
rect 7520 -2564 7560 -2516
rect 7520 -2596 7524 -2564
rect 7556 -2596 7560 -2564
rect 7520 -2644 7560 -2596
rect 7520 -2676 7524 -2644
rect 7556 -2676 7560 -2644
rect 7520 -2724 7560 -2676
rect 7520 -2756 7524 -2724
rect 7556 -2756 7560 -2724
rect 7520 -2804 7560 -2756
rect 7520 -2836 7524 -2804
rect 7556 -2836 7560 -2804
rect 7520 -2884 7560 -2836
rect 7520 -2916 7524 -2884
rect 7556 -2916 7560 -2884
rect 7520 -2964 7560 -2916
rect 7520 -2996 7524 -2964
rect 7556 -2996 7560 -2964
rect 7520 -3044 7560 -2996
rect 7520 -3076 7524 -3044
rect 7556 -3076 7560 -3044
rect 7520 -3124 7560 -3076
rect 7520 -3156 7524 -3124
rect 7556 -3156 7560 -3124
rect 7520 -3204 7560 -3156
rect 7520 -3236 7524 -3204
rect 7556 -3236 7560 -3204
rect 7520 -3284 7560 -3236
rect 7520 -3316 7524 -3284
rect 7556 -3316 7560 -3284
rect 7520 -3364 7560 -3316
rect 7520 -3396 7524 -3364
rect 7556 -3396 7560 -3364
rect 7520 -3444 7560 -3396
rect 7520 -3476 7524 -3444
rect 7556 -3476 7560 -3444
rect 7520 -3524 7560 -3476
rect 7520 -3556 7524 -3524
rect 7556 -3556 7560 -3524
rect 7520 -3604 7560 -3556
rect 7520 -3636 7524 -3604
rect 7556 -3636 7560 -3604
rect 7520 -3684 7560 -3636
rect 7520 -3716 7524 -3684
rect 7556 -3716 7560 -3684
rect 7520 -3720 7560 -3716
rect 7600 1036 7640 1040
rect 7600 1004 7604 1036
rect 7636 1004 7640 1036
rect 7600 956 7640 1004
rect 7600 924 7604 956
rect 7636 924 7640 956
rect 7600 876 7640 924
rect 7600 844 7604 876
rect 7636 844 7640 876
rect 7600 796 7640 844
rect 7600 764 7604 796
rect 7636 764 7640 796
rect 7600 716 7640 764
rect 7600 684 7604 716
rect 7636 684 7640 716
rect 7600 636 7640 684
rect 7600 604 7604 636
rect 7636 604 7640 636
rect 7600 556 7640 604
rect 7600 524 7604 556
rect 7636 524 7640 556
rect 7600 476 7640 524
rect 7600 444 7604 476
rect 7636 444 7640 476
rect 7600 396 7640 444
rect 7600 364 7604 396
rect 7636 364 7640 396
rect 7600 316 7640 364
rect 7600 284 7604 316
rect 7636 284 7640 316
rect 7600 236 7640 284
rect 7600 204 7604 236
rect 7636 204 7640 236
rect 7600 156 7640 204
rect 7600 124 7604 156
rect 7636 124 7640 156
rect 7600 76 7640 124
rect 7600 44 7604 76
rect 7636 44 7640 76
rect 7600 -4 7640 44
rect 7600 -36 7604 -4
rect 7636 -36 7640 -4
rect 7600 -84 7640 -36
rect 7600 -116 7604 -84
rect 7636 -116 7640 -84
rect 7600 -164 7640 -116
rect 7600 -196 7604 -164
rect 7636 -196 7640 -164
rect 7600 -244 7640 -196
rect 7600 -276 7604 -244
rect 7636 -276 7640 -244
rect 7600 -324 7640 -276
rect 7600 -356 7604 -324
rect 7636 -356 7640 -324
rect 7600 -404 7640 -356
rect 7600 -436 7604 -404
rect 7636 -436 7640 -404
rect 7600 -484 7640 -436
rect 7600 -516 7604 -484
rect 7636 -516 7640 -484
rect 7600 -564 7640 -516
rect 7600 -596 7604 -564
rect 7636 -596 7640 -564
rect 7600 -644 7640 -596
rect 7600 -676 7604 -644
rect 7636 -676 7640 -644
rect 7600 -724 7640 -676
rect 7600 -756 7604 -724
rect 7636 -756 7640 -724
rect 7600 -804 7640 -756
rect 7600 -836 7604 -804
rect 7636 -836 7640 -804
rect 7600 -884 7640 -836
rect 7600 -916 7604 -884
rect 7636 -916 7640 -884
rect 7600 -964 7640 -916
rect 7600 -996 7604 -964
rect 7636 -996 7640 -964
rect 7600 -1044 7640 -996
rect 7600 -1076 7604 -1044
rect 7636 -1076 7640 -1044
rect 7600 -1124 7640 -1076
rect 7600 -1156 7604 -1124
rect 7636 -1156 7640 -1124
rect 7600 -1204 7640 -1156
rect 7600 -1236 7604 -1204
rect 7636 -1236 7640 -1204
rect 7600 -1284 7640 -1236
rect 7600 -1316 7604 -1284
rect 7636 -1316 7640 -1284
rect 7600 -1364 7640 -1316
rect 7600 -1396 7604 -1364
rect 7636 -1396 7640 -1364
rect 7600 -1444 7640 -1396
rect 7600 -1476 7604 -1444
rect 7636 -1476 7640 -1444
rect 7600 -1524 7640 -1476
rect 7600 -1556 7604 -1524
rect 7636 -1556 7640 -1524
rect 7600 -1604 7640 -1556
rect 7600 -1636 7604 -1604
rect 7636 -1636 7640 -1604
rect 7600 -1684 7640 -1636
rect 7600 -1716 7604 -1684
rect 7636 -1716 7640 -1684
rect 7600 -1764 7640 -1716
rect 7600 -1796 7604 -1764
rect 7636 -1796 7640 -1764
rect 7600 -1844 7640 -1796
rect 7600 -1876 7604 -1844
rect 7636 -1876 7640 -1844
rect 7600 -1924 7640 -1876
rect 7600 -1956 7604 -1924
rect 7636 -1956 7640 -1924
rect 7600 -2004 7640 -1956
rect 7600 -2036 7604 -2004
rect 7636 -2036 7640 -2004
rect 7600 -2084 7640 -2036
rect 7600 -2116 7604 -2084
rect 7636 -2116 7640 -2084
rect 7600 -2164 7640 -2116
rect 7600 -2196 7604 -2164
rect 7636 -2196 7640 -2164
rect 7600 -2244 7640 -2196
rect 7600 -2276 7604 -2244
rect 7636 -2276 7640 -2244
rect 7600 -2324 7640 -2276
rect 7600 -2356 7604 -2324
rect 7636 -2356 7640 -2324
rect 7600 -2404 7640 -2356
rect 7600 -2436 7604 -2404
rect 7636 -2436 7640 -2404
rect 7600 -2484 7640 -2436
rect 7600 -2516 7604 -2484
rect 7636 -2516 7640 -2484
rect 7600 -2564 7640 -2516
rect 7600 -2596 7604 -2564
rect 7636 -2596 7640 -2564
rect 7600 -2644 7640 -2596
rect 7600 -2676 7604 -2644
rect 7636 -2676 7640 -2644
rect 7600 -2724 7640 -2676
rect 7600 -2756 7604 -2724
rect 7636 -2756 7640 -2724
rect 7600 -2804 7640 -2756
rect 7600 -2836 7604 -2804
rect 7636 -2836 7640 -2804
rect 7600 -2884 7640 -2836
rect 7600 -2916 7604 -2884
rect 7636 -2916 7640 -2884
rect 7600 -2964 7640 -2916
rect 7600 -2996 7604 -2964
rect 7636 -2996 7640 -2964
rect 7600 -3044 7640 -2996
rect 7600 -3076 7604 -3044
rect 7636 -3076 7640 -3044
rect 7600 -3124 7640 -3076
rect 7600 -3156 7604 -3124
rect 7636 -3156 7640 -3124
rect 7600 -3204 7640 -3156
rect 7600 -3236 7604 -3204
rect 7636 -3236 7640 -3204
rect 7600 -3284 7640 -3236
rect 7600 -3316 7604 -3284
rect 7636 -3316 7640 -3284
rect 7600 -3364 7640 -3316
rect 7600 -3396 7604 -3364
rect 7636 -3396 7640 -3364
rect 7600 -3444 7640 -3396
rect 7600 -3476 7604 -3444
rect 7636 -3476 7640 -3444
rect 7600 -3524 7640 -3476
rect 7600 -3556 7604 -3524
rect 7636 -3556 7640 -3524
rect 7600 -3604 7640 -3556
rect 7600 -3636 7604 -3604
rect 7636 -3636 7640 -3604
rect 7600 -3684 7640 -3636
rect 7600 -3716 7604 -3684
rect 7636 -3716 7640 -3684
rect 7600 -3720 7640 -3716
rect 7680 1036 7720 1040
rect 7680 1004 7684 1036
rect 7716 1004 7720 1036
rect 7680 956 7720 1004
rect 7680 924 7684 956
rect 7716 924 7720 956
rect 7680 876 7720 924
rect 7680 844 7684 876
rect 7716 844 7720 876
rect 7680 796 7720 844
rect 7680 764 7684 796
rect 7716 764 7720 796
rect 7680 716 7720 764
rect 7680 684 7684 716
rect 7716 684 7720 716
rect 7680 636 7720 684
rect 7680 604 7684 636
rect 7716 604 7720 636
rect 7680 556 7720 604
rect 7680 524 7684 556
rect 7716 524 7720 556
rect 7680 476 7720 524
rect 7680 444 7684 476
rect 7716 444 7720 476
rect 7680 396 7720 444
rect 7680 364 7684 396
rect 7716 364 7720 396
rect 7680 316 7720 364
rect 7680 284 7684 316
rect 7716 284 7720 316
rect 7680 236 7720 284
rect 7680 204 7684 236
rect 7716 204 7720 236
rect 7680 156 7720 204
rect 7680 124 7684 156
rect 7716 124 7720 156
rect 7680 76 7720 124
rect 7680 44 7684 76
rect 7716 44 7720 76
rect 7680 -4 7720 44
rect 7680 -36 7684 -4
rect 7716 -36 7720 -4
rect 7680 -84 7720 -36
rect 7680 -116 7684 -84
rect 7716 -116 7720 -84
rect 7680 -164 7720 -116
rect 7680 -196 7684 -164
rect 7716 -196 7720 -164
rect 7680 -244 7720 -196
rect 7680 -276 7684 -244
rect 7716 -276 7720 -244
rect 7680 -324 7720 -276
rect 7680 -356 7684 -324
rect 7716 -356 7720 -324
rect 7680 -404 7720 -356
rect 7680 -436 7684 -404
rect 7716 -436 7720 -404
rect 7680 -484 7720 -436
rect 7680 -516 7684 -484
rect 7716 -516 7720 -484
rect 7680 -564 7720 -516
rect 7680 -596 7684 -564
rect 7716 -596 7720 -564
rect 7680 -644 7720 -596
rect 7680 -676 7684 -644
rect 7716 -676 7720 -644
rect 7680 -724 7720 -676
rect 7680 -756 7684 -724
rect 7716 -756 7720 -724
rect 7680 -804 7720 -756
rect 7680 -836 7684 -804
rect 7716 -836 7720 -804
rect 7680 -884 7720 -836
rect 7680 -916 7684 -884
rect 7716 -916 7720 -884
rect 7680 -964 7720 -916
rect 7680 -996 7684 -964
rect 7716 -996 7720 -964
rect 7680 -1044 7720 -996
rect 7680 -1076 7684 -1044
rect 7716 -1076 7720 -1044
rect 7680 -1124 7720 -1076
rect 7680 -1156 7684 -1124
rect 7716 -1156 7720 -1124
rect 7680 -1204 7720 -1156
rect 7680 -1236 7684 -1204
rect 7716 -1236 7720 -1204
rect 7680 -1284 7720 -1236
rect 7680 -1316 7684 -1284
rect 7716 -1316 7720 -1284
rect 7680 -1364 7720 -1316
rect 7680 -1396 7684 -1364
rect 7716 -1396 7720 -1364
rect 7680 -1444 7720 -1396
rect 7680 -1476 7684 -1444
rect 7716 -1476 7720 -1444
rect 7680 -1524 7720 -1476
rect 7680 -1556 7684 -1524
rect 7716 -1556 7720 -1524
rect 7680 -1604 7720 -1556
rect 7680 -1636 7684 -1604
rect 7716 -1636 7720 -1604
rect 7680 -1684 7720 -1636
rect 7680 -1716 7684 -1684
rect 7716 -1716 7720 -1684
rect 7680 -1764 7720 -1716
rect 7680 -1796 7684 -1764
rect 7716 -1796 7720 -1764
rect 7680 -1844 7720 -1796
rect 7680 -1876 7684 -1844
rect 7716 -1876 7720 -1844
rect 7680 -1924 7720 -1876
rect 7680 -1956 7684 -1924
rect 7716 -1956 7720 -1924
rect 7680 -2004 7720 -1956
rect 7680 -2036 7684 -2004
rect 7716 -2036 7720 -2004
rect 7680 -2084 7720 -2036
rect 7680 -2116 7684 -2084
rect 7716 -2116 7720 -2084
rect 7680 -2164 7720 -2116
rect 7680 -2196 7684 -2164
rect 7716 -2196 7720 -2164
rect 7680 -2244 7720 -2196
rect 7680 -2276 7684 -2244
rect 7716 -2276 7720 -2244
rect 7680 -2324 7720 -2276
rect 7680 -2356 7684 -2324
rect 7716 -2356 7720 -2324
rect 7680 -2404 7720 -2356
rect 7680 -2436 7684 -2404
rect 7716 -2436 7720 -2404
rect 7680 -2484 7720 -2436
rect 7680 -2516 7684 -2484
rect 7716 -2516 7720 -2484
rect 7680 -2564 7720 -2516
rect 7680 -2596 7684 -2564
rect 7716 -2596 7720 -2564
rect 7680 -2644 7720 -2596
rect 7680 -2676 7684 -2644
rect 7716 -2676 7720 -2644
rect 7680 -2724 7720 -2676
rect 7680 -2756 7684 -2724
rect 7716 -2756 7720 -2724
rect 7680 -2804 7720 -2756
rect 7680 -2836 7684 -2804
rect 7716 -2836 7720 -2804
rect 7680 -2884 7720 -2836
rect 7680 -2916 7684 -2884
rect 7716 -2916 7720 -2884
rect 7680 -2964 7720 -2916
rect 7680 -2996 7684 -2964
rect 7716 -2996 7720 -2964
rect 7680 -3044 7720 -2996
rect 7680 -3076 7684 -3044
rect 7716 -3076 7720 -3044
rect 7680 -3124 7720 -3076
rect 7680 -3156 7684 -3124
rect 7716 -3156 7720 -3124
rect 7680 -3204 7720 -3156
rect 7680 -3236 7684 -3204
rect 7716 -3236 7720 -3204
rect 7680 -3284 7720 -3236
rect 7680 -3316 7684 -3284
rect 7716 -3316 7720 -3284
rect 7680 -3364 7720 -3316
rect 7680 -3396 7684 -3364
rect 7716 -3396 7720 -3364
rect 7680 -3444 7720 -3396
rect 7680 -3476 7684 -3444
rect 7716 -3476 7720 -3444
rect 7680 -3524 7720 -3476
rect 7680 -3556 7684 -3524
rect 7716 -3556 7720 -3524
rect 7680 -3604 7720 -3556
rect 7680 -3636 7684 -3604
rect 7716 -3636 7720 -3604
rect 7680 -3684 7720 -3636
rect 7680 -3716 7684 -3684
rect 7716 -3716 7720 -3684
rect 7680 -3720 7720 -3716
rect 7760 1036 7800 1040
rect 7760 1004 7764 1036
rect 7796 1004 7800 1036
rect 7760 956 7800 1004
rect 7760 924 7764 956
rect 7796 924 7800 956
rect 7760 876 7800 924
rect 7760 844 7764 876
rect 7796 844 7800 876
rect 7760 796 7800 844
rect 7760 764 7764 796
rect 7796 764 7800 796
rect 7760 716 7800 764
rect 7760 684 7764 716
rect 7796 684 7800 716
rect 7760 636 7800 684
rect 7760 604 7764 636
rect 7796 604 7800 636
rect 7760 556 7800 604
rect 7760 524 7764 556
rect 7796 524 7800 556
rect 7760 476 7800 524
rect 7760 444 7764 476
rect 7796 444 7800 476
rect 7760 396 7800 444
rect 7760 364 7764 396
rect 7796 364 7800 396
rect 7760 316 7800 364
rect 7760 284 7764 316
rect 7796 284 7800 316
rect 7760 236 7800 284
rect 7760 204 7764 236
rect 7796 204 7800 236
rect 7760 156 7800 204
rect 7760 124 7764 156
rect 7796 124 7800 156
rect 7760 76 7800 124
rect 7760 44 7764 76
rect 7796 44 7800 76
rect 7760 -4 7800 44
rect 7760 -36 7764 -4
rect 7796 -36 7800 -4
rect 7760 -84 7800 -36
rect 7760 -116 7764 -84
rect 7796 -116 7800 -84
rect 7760 -164 7800 -116
rect 7760 -196 7764 -164
rect 7796 -196 7800 -164
rect 7760 -244 7800 -196
rect 7760 -276 7764 -244
rect 7796 -276 7800 -244
rect 7760 -324 7800 -276
rect 7760 -356 7764 -324
rect 7796 -356 7800 -324
rect 7760 -404 7800 -356
rect 7760 -436 7764 -404
rect 7796 -436 7800 -404
rect 7760 -484 7800 -436
rect 7760 -516 7764 -484
rect 7796 -516 7800 -484
rect 7760 -564 7800 -516
rect 7760 -596 7764 -564
rect 7796 -596 7800 -564
rect 7760 -644 7800 -596
rect 7760 -676 7764 -644
rect 7796 -676 7800 -644
rect 7760 -724 7800 -676
rect 7760 -756 7764 -724
rect 7796 -756 7800 -724
rect 7760 -804 7800 -756
rect 7760 -836 7764 -804
rect 7796 -836 7800 -804
rect 7760 -884 7800 -836
rect 7760 -916 7764 -884
rect 7796 -916 7800 -884
rect 7760 -964 7800 -916
rect 7760 -996 7764 -964
rect 7796 -996 7800 -964
rect 7760 -1044 7800 -996
rect 7760 -1076 7764 -1044
rect 7796 -1076 7800 -1044
rect 7760 -1124 7800 -1076
rect 7760 -1156 7764 -1124
rect 7796 -1156 7800 -1124
rect 7760 -1204 7800 -1156
rect 7760 -1236 7764 -1204
rect 7796 -1236 7800 -1204
rect 7760 -1284 7800 -1236
rect 7760 -1316 7764 -1284
rect 7796 -1316 7800 -1284
rect 7760 -1364 7800 -1316
rect 7760 -1396 7764 -1364
rect 7796 -1396 7800 -1364
rect 7760 -1444 7800 -1396
rect 7760 -1476 7764 -1444
rect 7796 -1476 7800 -1444
rect 7760 -1524 7800 -1476
rect 7760 -1556 7764 -1524
rect 7796 -1556 7800 -1524
rect 7760 -1604 7800 -1556
rect 7760 -1636 7764 -1604
rect 7796 -1636 7800 -1604
rect 7760 -1684 7800 -1636
rect 7760 -1716 7764 -1684
rect 7796 -1716 7800 -1684
rect 7760 -1764 7800 -1716
rect 7760 -1796 7764 -1764
rect 7796 -1796 7800 -1764
rect 7760 -1844 7800 -1796
rect 7760 -1876 7764 -1844
rect 7796 -1876 7800 -1844
rect 7760 -1924 7800 -1876
rect 7760 -1956 7764 -1924
rect 7796 -1956 7800 -1924
rect 7760 -2004 7800 -1956
rect 7760 -2036 7764 -2004
rect 7796 -2036 7800 -2004
rect 7760 -2084 7800 -2036
rect 7760 -2116 7764 -2084
rect 7796 -2116 7800 -2084
rect 7760 -2164 7800 -2116
rect 7760 -2196 7764 -2164
rect 7796 -2196 7800 -2164
rect 7760 -2244 7800 -2196
rect 7760 -2276 7764 -2244
rect 7796 -2276 7800 -2244
rect 7760 -2324 7800 -2276
rect 7760 -2356 7764 -2324
rect 7796 -2356 7800 -2324
rect 7760 -2404 7800 -2356
rect 7760 -2436 7764 -2404
rect 7796 -2436 7800 -2404
rect 7760 -2484 7800 -2436
rect 7760 -2516 7764 -2484
rect 7796 -2516 7800 -2484
rect 7760 -2564 7800 -2516
rect 7760 -2596 7764 -2564
rect 7796 -2596 7800 -2564
rect 7760 -2644 7800 -2596
rect 7760 -2676 7764 -2644
rect 7796 -2676 7800 -2644
rect 7760 -2724 7800 -2676
rect 7760 -2756 7764 -2724
rect 7796 -2756 7800 -2724
rect 7760 -2804 7800 -2756
rect 7760 -2836 7764 -2804
rect 7796 -2836 7800 -2804
rect 7760 -2884 7800 -2836
rect 7760 -2916 7764 -2884
rect 7796 -2916 7800 -2884
rect 7760 -2964 7800 -2916
rect 7760 -2996 7764 -2964
rect 7796 -2996 7800 -2964
rect 7760 -3044 7800 -2996
rect 7760 -3076 7764 -3044
rect 7796 -3076 7800 -3044
rect 7760 -3124 7800 -3076
rect 7760 -3156 7764 -3124
rect 7796 -3156 7800 -3124
rect 7760 -3204 7800 -3156
rect 7760 -3236 7764 -3204
rect 7796 -3236 7800 -3204
rect 7760 -3284 7800 -3236
rect 7760 -3316 7764 -3284
rect 7796 -3316 7800 -3284
rect 7760 -3364 7800 -3316
rect 7760 -3396 7764 -3364
rect 7796 -3396 7800 -3364
rect 7760 -3444 7800 -3396
rect 7760 -3476 7764 -3444
rect 7796 -3476 7800 -3444
rect 7760 -3524 7800 -3476
rect 7760 -3556 7764 -3524
rect 7796 -3556 7800 -3524
rect 7760 -3604 7800 -3556
rect 7760 -3636 7764 -3604
rect 7796 -3636 7800 -3604
rect 7760 -3684 7800 -3636
rect 7760 -3716 7764 -3684
rect 7796 -3716 7800 -3684
rect 7760 -3720 7800 -3716
rect 7840 1036 7880 1040
rect 7840 1004 7844 1036
rect 7876 1004 7880 1036
rect 7840 956 7880 1004
rect 7840 924 7844 956
rect 7876 924 7880 956
rect 7840 876 7880 924
rect 7840 844 7844 876
rect 7876 844 7880 876
rect 7840 796 7880 844
rect 7840 764 7844 796
rect 7876 764 7880 796
rect 7840 716 7880 764
rect 7840 684 7844 716
rect 7876 684 7880 716
rect 7840 636 7880 684
rect 7840 604 7844 636
rect 7876 604 7880 636
rect 7840 556 7880 604
rect 7840 524 7844 556
rect 7876 524 7880 556
rect 7840 476 7880 524
rect 7840 444 7844 476
rect 7876 444 7880 476
rect 7840 396 7880 444
rect 7840 364 7844 396
rect 7876 364 7880 396
rect 7840 316 7880 364
rect 7840 284 7844 316
rect 7876 284 7880 316
rect 7840 236 7880 284
rect 7840 204 7844 236
rect 7876 204 7880 236
rect 7840 156 7880 204
rect 7840 124 7844 156
rect 7876 124 7880 156
rect 7840 76 7880 124
rect 7840 44 7844 76
rect 7876 44 7880 76
rect 7840 -4 7880 44
rect 7840 -36 7844 -4
rect 7876 -36 7880 -4
rect 7840 -84 7880 -36
rect 7840 -116 7844 -84
rect 7876 -116 7880 -84
rect 7840 -164 7880 -116
rect 7840 -196 7844 -164
rect 7876 -196 7880 -164
rect 7840 -244 7880 -196
rect 7840 -276 7844 -244
rect 7876 -276 7880 -244
rect 7840 -324 7880 -276
rect 7840 -356 7844 -324
rect 7876 -356 7880 -324
rect 7840 -404 7880 -356
rect 7840 -436 7844 -404
rect 7876 -436 7880 -404
rect 7840 -484 7880 -436
rect 7840 -516 7844 -484
rect 7876 -516 7880 -484
rect 7840 -564 7880 -516
rect 7840 -596 7844 -564
rect 7876 -596 7880 -564
rect 7840 -644 7880 -596
rect 7840 -676 7844 -644
rect 7876 -676 7880 -644
rect 7840 -724 7880 -676
rect 7840 -756 7844 -724
rect 7876 -756 7880 -724
rect 7840 -804 7880 -756
rect 7840 -836 7844 -804
rect 7876 -836 7880 -804
rect 7840 -884 7880 -836
rect 7840 -916 7844 -884
rect 7876 -916 7880 -884
rect 7840 -964 7880 -916
rect 7840 -996 7844 -964
rect 7876 -996 7880 -964
rect 7840 -1044 7880 -996
rect 7840 -1076 7844 -1044
rect 7876 -1076 7880 -1044
rect 7840 -1124 7880 -1076
rect 7840 -1156 7844 -1124
rect 7876 -1156 7880 -1124
rect 7840 -1204 7880 -1156
rect 7840 -1236 7844 -1204
rect 7876 -1236 7880 -1204
rect 7840 -1284 7880 -1236
rect 7840 -1316 7844 -1284
rect 7876 -1316 7880 -1284
rect 7840 -1364 7880 -1316
rect 7840 -1396 7844 -1364
rect 7876 -1396 7880 -1364
rect 7840 -1444 7880 -1396
rect 7840 -1476 7844 -1444
rect 7876 -1476 7880 -1444
rect 7840 -1524 7880 -1476
rect 7840 -1556 7844 -1524
rect 7876 -1556 7880 -1524
rect 7840 -1604 7880 -1556
rect 7840 -1636 7844 -1604
rect 7876 -1636 7880 -1604
rect 7840 -1684 7880 -1636
rect 7840 -1716 7844 -1684
rect 7876 -1716 7880 -1684
rect 7840 -1764 7880 -1716
rect 7840 -1796 7844 -1764
rect 7876 -1796 7880 -1764
rect 7840 -1844 7880 -1796
rect 7840 -1876 7844 -1844
rect 7876 -1876 7880 -1844
rect 7840 -1924 7880 -1876
rect 7840 -1956 7844 -1924
rect 7876 -1956 7880 -1924
rect 7840 -2004 7880 -1956
rect 7840 -2036 7844 -2004
rect 7876 -2036 7880 -2004
rect 7840 -2084 7880 -2036
rect 7840 -2116 7844 -2084
rect 7876 -2116 7880 -2084
rect 7840 -2164 7880 -2116
rect 7840 -2196 7844 -2164
rect 7876 -2196 7880 -2164
rect 7840 -2244 7880 -2196
rect 7840 -2276 7844 -2244
rect 7876 -2276 7880 -2244
rect 7840 -2324 7880 -2276
rect 7840 -2356 7844 -2324
rect 7876 -2356 7880 -2324
rect 7840 -2404 7880 -2356
rect 7840 -2436 7844 -2404
rect 7876 -2436 7880 -2404
rect 7840 -2484 7880 -2436
rect 7840 -2516 7844 -2484
rect 7876 -2516 7880 -2484
rect 7840 -2564 7880 -2516
rect 7840 -2596 7844 -2564
rect 7876 -2596 7880 -2564
rect 7840 -2644 7880 -2596
rect 7840 -2676 7844 -2644
rect 7876 -2676 7880 -2644
rect 7840 -2724 7880 -2676
rect 7840 -2756 7844 -2724
rect 7876 -2756 7880 -2724
rect 7840 -2804 7880 -2756
rect 7840 -2836 7844 -2804
rect 7876 -2836 7880 -2804
rect 7840 -2884 7880 -2836
rect 7840 -2916 7844 -2884
rect 7876 -2916 7880 -2884
rect 7840 -2964 7880 -2916
rect 7840 -2996 7844 -2964
rect 7876 -2996 7880 -2964
rect 7840 -3044 7880 -2996
rect 7840 -3076 7844 -3044
rect 7876 -3076 7880 -3044
rect 7840 -3124 7880 -3076
rect 7840 -3156 7844 -3124
rect 7876 -3156 7880 -3124
rect 7840 -3204 7880 -3156
rect 7840 -3236 7844 -3204
rect 7876 -3236 7880 -3204
rect 7840 -3284 7880 -3236
rect 7840 -3316 7844 -3284
rect 7876 -3316 7880 -3284
rect 7840 -3364 7880 -3316
rect 7840 -3396 7844 -3364
rect 7876 -3396 7880 -3364
rect 7840 -3444 7880 -3396
rect 7840 -3476 7844 -3444
rect 7876 -3476 7880 -3444
rect 7840 -3524 7880 -3476
rect 7840 -3556 7844 -3524
rect 7876 -3556 7880 -3524
rect 7840 -3604 7880 -3556
rect 7840 -3636 7844 -3604
rect 7876 -3636 7880 -3604
rect 7840 -3684 7880 -3636
rect 7840 -3716 7844 -3684
rect 7876 -3716 7880 -3684
rect 7840 -3720 7880 -3716
rect 7920 1036 7960 1040
rect 7920 1004 7924 1036
rect 7956 1004 7960 1036
rect 7920 956 7960 1004
rect 7920 924 7924 956
rect 7956 924 7960 956
rect 7920 876 7960 924
rect 7920 844 7924 876
rect 7956 844 7960 876
rect 7920 796 7960 844
rect 7920 764 7924 796
rect 7956 764 7960 796
rect 7920 716 7960 764
rect 7920 684 7924 716
rect 7956 684 7960 716
rect 7920 636 7960 684
rect 7920 604 7924 636
rect 7956 604 7960 636
rect 7920 556 7960 604
rect 7920 524 7924 556
rect 7956 524 7960 556
rect 7920 476 7960 524
rect 7920 444 7924 476
rect 7956 444 7960 476
rect 7920 396 7960 444
rect 7920 364 7924 396
rect 7956 364 7960 396
rect 7920 316 7960 364
rect 7920 284 7924 316
rect 7956 284 7960 316
rect 7920 236 7960 284
rect 7920 204 7924 236
rect 7956 204 7960 236
rect 7920 156 7960 204
rect 7920 124 7924 156
rect 7956 124 7960 156
rect 7920 76 7960 124
rect 7920 44 7924 76
rect 7956 44 7960 76
rect 7920 -4 7960 44
rect 7920 -36 7924 -4
rect 7956 -36 7960 -4
rect 7920 -84 7960 -36
rect 7920 -116 7924 -84
rect 7956 -116 7960 -84
rect 7920 -164 7960 -116
rect 7920 -196 7924 -164
rect 7956 -196 7960 -164
rect 7920 -244 7960 -196
rect 7920 -276 7924 -244
rect 7956 -276 7960 -244
rect 7920 -324 7960 -276
rect 7920 -356 7924 -324
rect 7956 -356 7960 -324
rect 7920 -404 7960 -356
rect 7920 -436 7924 -404
rect 7956 -436 7960 -404
rect 7920 -484 7960 -436
rect 7920 -516 7924 -484
rect 7956 -516 7960 -484
rect 7920 -564 7960 -516
rect 7920 -596 7924 -564
rect 7956 -596 7960 -564
rect 7920 -644 7960 -596
rect 7920 -676 7924 -644
rect 7956 -676 7960 -644
rect 7920 -724 7960 -676
rect 7920 -756 7924 -724
rect 7956 -756 7960 -724
rect 7920 -804 7960 -756
rect 7920 -836 7924 -804
rect 7956 -836 7960 -804
rect 7920 -884 7960 -836
rect 7920 -916 7924 -884
rect 7956 -916 7960 -884
rect 7920 -964 7960 -916
rect 7920 -996 7924 -964
rect 7956 -996 7960 -964
rect 7920 -1044 7960 -996
rect 7920 -1076 7924 -1044
rect 7956 -1076 7960 -1044
rect 7920 -1124 7960 -1076
rect 7920 -1156 7924 -1124
rect 7956 -1156 7960 -1124
rect 7920 -1204 7960 -1156
rect 7920 -1236 7924 -1204
rect 7956 -1236 7960 -1204
rect 7920 -1284 7960 -1236
rect 7920 -1316 7924 -1284
rect 7956 -1316 7960 -1284
rect 7920 -1364 7960 -1316
rect 7920 -1396 7924 -1364
rect 7956 -1396 7960 -1364
rect 7920 -1444 7960 -1396
rect 7920 -1476 7924 -1444
rect 7956 -1476 7960 -1444
rect 7920 -1524 7960 -1476
rect 7920 -1556 7924 -1524
rect 7956 -1556 7960 -1524
rect 7920 -1604 7960 -1556
rect 7920 -1636 7924 -1604
rect 7956 -1636 7960 -1604
rect 7920 -1684 7960 -1636
rect 7920 -1716 7924 -1684
rect 7956 -1716 7960 -1684
rect 7920 -1764 7960 -1716
rect 7920 -1796 7924 -1764
rect 7956 -1796 7960 -1764
rect 7920 -1844 7960 -1796
rect 7920 -1876 7924 -1844
rect 7956 -1876 7960 -1844
rect 7920 -1924 7960 -1876
rect 7920 -1956 7924 -1924
rect 7956 -1956 7960 -1924
rect 7920 -2004 7960 -1956
rect 7920 -2036 7924 -2004
rect 7956 -2036 7960 -2004
rect 7920 -2084 7960 -2036
rect 7920 -2116 7924 -2084
rect 7956 -2116 7960 -2084
rect 7920 -2164 7960 -2116
rect 7920 -2196 7924 -2164
rect 7956 -2196 7960 -2164
rect 7920 -2244 7960 -2196
rect 7920 -2276 7924 -2244
rect 7956 -2276 7960 -2244
rect 7920 -2324 7960 -2276
rect 7920 -2356 7924 -2324
rect 7956 -2356 7960 -2324
rect 7920 -2404 7960 -2356
rect 7920 -2436 7924 -2404
rect 7956 -2436 7960 -2404
rect 7920 -2484 7960 -2436
rect 7920 -2516 7924 -2484
rect 7956 -2516 7960 -2484
rect 7920 -2564 7960 -2516
rect 7920 -2596 7924 -2564
rect 7956 -2596 7960 -2564
rect 7920 -2644 7960 -2596
rect 7920 -2676 7924 -2644
rect 7956 -2676 7960 -2644
rect 7920 -2724 7960 -2676
rect 7920 -2756 7924 -2724
rect 7956 -2756 7960 -2724
rect 7920 -2804 7960 -2756
rect 7920 -2836 7924 -2804
rect 7956 -2836 7960 -2804
rect 7920 -2884 7960 -2836
rect 7920 -2916 7924 -2884
rect 7956 -2916 7960 -2884
rect 7920 -2964 7960 -2916
rect 7920 -2996 7924 -2964
rect 7956 -2996 7960 -2964
rect 7920 -3044 7960 -2996
rect 7920 -3076 7924 -3044
rect 7956 -3076 7960 -3044
rect 7920 -3124 7960 -3076
rect 7920 -3156 7924 -3124
rect 7956 -3156 7960 -3124
rect 7920 -3204 7960 -3156
rect 7920 -3236 7924 -3204
rect 7956 -3236 7960 -3204
rect 7920 -3284 7960 -3236
rect 7920 -3316 7924 -3284
rect 7956 -3316 7960 -3284
rect 7920 -3364 7960 -3316
rect 7920 -3396 7924 -3364
rect 7956 -3396 7960 -3364
rect 7920 -3444 7960 -3396
rect 7920 -3476 7924 -3444
rect 7956 -3476 7960 -3444
rect 7920 -3524 7960 -3476
rect 7920 -3556 7924 -3524
rect 7956 -3556 7960 -3524
rect 7920 -3604 7960 -3556
rect 7920 -3636 7924 -3604
rect 7956 -3636 7960 -3604
rect 7920 -3684 7960 -3636
rect 7920 -3716 7924 -3684
rect 7956 -3716 7960 -3684
rect 7920 -3720 7960 -3716
rect 8000 1036 8040 1040
rect 8000 1004 8004 1036
rect 8036 1004 8040 1036
rect 8000 956 8040 1004
rect 8000 924 8004 956
rect 8036 924 8040 956
rect 8000 876 8040 924
rect 8000 844 8004 876
rect 8036 844 8040 876
rect 8000 796 8040 844
rect 8000 764 8004 796
rect 8036 764 8040 796
rect 8000 716 8040 764
rect 8000 684 8004 716
rect 8036 684 8040 716
rect 8000 636 8040 684
rect 8000 604 8004 636
rect 8036 604 8040 636
rect 8000 556 8040 604
rect 8000 524 8004 556
rect 8036 524 8040 556
rect 8000 476 8040 524
rect 8000 444 8004 476
rect 8036 444 8040 476
rect 8000 396 8040 444
rect 8000 364 8004 396
rect 8036 364 8040 396
rect 8000 316 8040 364
rect 8000 284 8004 316
rect 8036 284 8040 316
rect 8000 236 8040 284
rect 8000 204 8004 236
rect 8036 204 8040 236
rect 8000 156 8040 204
rect 8000 124 8004 156
rect 8036 124 8040 156
rect 8000 76 8040 124
rect 8000 44 8004 76
rect 8036 44 8040 76
rect 8000 -4 8040 44
rect 8000 -36 8004 -4
rect 8036 -36 8040 -4
rect 8000 -84 8040 -36
rect 8000 -116 8004 -84
rect 8036 -116 8040 -84
rect 8000 -164 8040 -116
rect 8000 -196 8004 -164
rect 8036 -196 8040 -164
rect 8000 -244 8040 -196
rect 8000 -276 8004 -244
rect 8036 -276 8040 -244
rect 8000 -324 8040 -276
rect 8000 -356 8004 -324
rect 8036 -356 8040 -324
rect 8000 -404 8040 -356
rect 8000 -436 8004 -404
rect 8036 -436 8040 -404
rect 8000 -484 8040 -436
rect 8000 -516 8004 -484
rect 8036 -516 8040 -484
rect 8000 -564 8040 -516
rect 8000 -596 8004 -564
rect 8036 -596 8040 -564
rect 8000 -644 8040 -596
rect 8000 -676 8004 -644
rect 8036 -676 8040 -644
rect 8000 -724 8040 -676
rect 8000 -756 8004 -724
rect 8036 -756 8040 -724
rect 8000 -804 8040 -756
rect 8000 -836 8004 -804
rect 8036 -836 8040 -804
rect 8000 -884 8040 -836
rect 8000 -916 8004 -884
rect 8036 -916 8040 -884
rect 8000 -964 8040 -916
rect 8000 -996 8004 -964
rect 8036 -996 8040 -964
rect 8000 -1044 8040 -996
rect 8000 -1076 8004 -1044
rect 8036 -1076 8040 -1044
rect 8000 -1124 8040 -1076
rect 8000 -1156 8004 -1124
rect 8036 -1156 8040 -1124
rect 8000 -1204 8040 -1156
rect 8000 -1236 8004 -1204
rect 8036 -1236 8040 -1204
rect 8000 -1284 8040 -1236
rect 8000 -1316 8004 -1284
rect 8036 -1316 8040 -1284
rect 8000 -1364 8040 -1316
rect 8000 -1396 8004 -1364
rect 8036 -1396 8040 -1364
rect 8000 -1444 8040 -1396
rect 8000 -1476 8004 -1444
rect 8036 -1476 8040 -1444
rect 8000 -1524 8040 -1476
rect 8000 -1556 8004 -1524
rect 8036 -1556 8040 -1524
rect 8000 -1604 8040 -1556
rect 8000 -1636 8004 -1604
rect 8036 -1636 8040 -1604
rect 8000 -1684 8040 -1636
rect 8000 -1716 8004 -1684
rect 8036 -1716 8040 -1684
rect 8000 -1764 8040 -1716
rect 8000 -1796 8004 -1764
rect 8036 -1796 8040 -1764
rect 8000 -1844 8040 -1796
rect 8000 -1876 8004 -1844
rect 8036 -1876 8040 -1844
rect 8000 -1924 8040 -1876
rect 8000 -1956 8004 -1924
rect 8036 -1956 8040 -1924
rect 8000 -2004 8040 -1956
rect 8000 -2036 8004 -2004
rect 8036 -2036 8040 -2004
rect 8000 -2084 8040 -2036
rect 8000 -2116 8004 -2084
rect 8036 -2116 8040 -2084
rect 8000 -2164 8040 -2116
rect 8000 -2196 8004 -2164
rect 8036 -2196 8040 -2164
rect 8000 -2244 8040 -2196
rect 8000 -2276 8004 -2244
rect 8036 -2276 8040 -2244
rect 8000 -2324 8040 -2276
rect 8000 -2356 8004 -2324
rect 8036 -2356 8040 -2324
rect 8000 -2404 8040 -2356
rect 8000 -2436 8004 -2404
rect 8036 -2436 8040 -2404
rect 8000 -2484 8040 -2436
rect 8000 -2516 8004 -2484
rect 8036 -2516 8040 -2484
rect 8000 -2564 8040 -2516
rect 8000 -2596 8004 -2564
rect 8036 -2596 8040 -2564
rect 8000 -2644 8040 -2596
rect 8000 -2676 8004 -2644
rect 8036 -2676 8040 -2644
rect 8000 -2724 8040 -2676
rect 8000 -2756 8004 -2724
rect 8036 -2756 8040 -2724
rect 8000 -2804 8040 -2756
rect 8000 -2836 8004 -2804
rect 8036 -2836 8040 -2804
rect 8000 -2884 8040 -2836
rect 8000 -2916 8004 -2884
rect 8036 -2916 8040 -2884
rect 8000 -2964 8040 -2916
rect 8000 -2996 8004 -2964
rect 8036 -2996 8040 -2964
rect 8000 -3044 8040 -2996
rect 8000 -3076 8004 -3044
rect 8036 -3076 8040 -3044
rect 8000 -3124 8040 -3076
rect 8000 -3156 8004 -3124
rect 8036 -3156 8040 -3124
rect 8000 -3204 8040 -3156
rect 8000 -3236 8004 -3204
rect 8036 -3236 8040 -3204
rect 8000 -3284 8040 -3236
rect 8000 -3316 8004 -3284
rect 8036 -3316 8040 -3284
rect 8000 -3364 8040 -3316
rect 8000 -3396 8004 -3364
rect 8036 -3396 8040 -3364
rect 8000 -3444 8040 -3396
rect 8000 -3476 8004 -3444
rect 8036 -3476 8040 -3444
rect 8000 -3524 8040 -3476
rect 8000 -3556 8004 -3524
rect 8036 -3556 8040 -3524
rect 8000 -3604 8040 -3556
rect 8000 -3636 8004 -3604
rect 8036 -3636 8040 -3604
rect 8000 -3684 8040 -3636
rect 8000 -3716 8004 -3684
rect 8036 -3716 8040 -3684
rect 8000 -3720 8040 -3716
rect 8080 1036 8120 1040
rect 8080 1004 8084 1036
rect 8116 1004 8120 1036
rect 8080 956 8120 1004
rect 8080 924 8084 956
rect 8116 924 8120 956
rect 8080 876 8120 924
rect 8080 844 8084 876
rect 8116 844 8120 876
rect 8080 796 8120 844
rect 8080 764 8084 796
rect 8116 764 8120 796
rect 8080 716 8120 764
rect 8080 684 8084 716
rect 8116 684 8120 716
rect 8080 636 8120 684
rect 8080 604 8084 636
rect 8116 604 8120 636
rect 8080 556 8120 604
rect 8080 524 8084 556
rect 8116 524 8120 556
rect 8080 476 8120 524
rect 8080 444 8084 476
rect 8116 444 8120 476
rect 8080 396 8120 444
rect 8080 364 8084 396
rect 8116 364 8120 396
rect 8080 316 8120 364
rect 8080 284 8084 316
rect 8116 284 8120 316
rect 8080 236 8120 284
rect 8080 204 8084 236
rect 8116 204 8120 236
rect 8080 156 8120 204
rect 8080 124 8084 156
rect 8116 124 8120 156
rect 8080 76 8120 124
rect 8080 44 8084 76
rect 8116 44 8120 76
rect 8080 -4 8120 44
rect 8080 -36 8084 -4
rect 8116 -36 8120 -4
rect 8080 -84 8120 -36
rect 8080 -116 8084 -84
rect 8116 -116 8120 -84
rect 8080 -164 8120 -116
rect 8080 -196 8084 -164
rect 8116 -196 8120 -164
rect 8080 -244 8120 -196
rect 8080 -276 8084 -244
rect 8116 -276 8120 -244
rect 8080 -324 8120 -276
rect 8080 -356 8084 -324
rect 8116 -356 8120 -324
rect 8080 -404 8120 -356
rect 8080 -436 8084 -404
rect 8116 -436 8120 -404
rect 8080 -484 8120 -436
rect 8080 -516 8084 -484
rect 8116 -516 8120 -484
rect 8080 -564 8120 -516
rect 8080 -596 8084 -564
rect 8116 -596 8120 -564
rect 8080 -644 8120 -596
rect 8080 -676 8084 -644
rect 8116 -676 8120 -644
rect 8080 -724 8120 -676
rect 8080 -756 8084 -724
rect 8116 -756 8120 -724
rect 8080 -804 8120 -756
rect 8080 -836 8084 -804
rect 8116 -836 8120 -804
rect 8080 -884 8120 -836
rect 8080 -916 8084 -884
rect 8116 -916 8120 -884
rect 8080 -964 8120 -916
rect 8080 -996 8084 -964
rect 8116 -996 8120 -964
rect 8080 -1044 8120 -996
rect 8080 -1076 8084 -1044
rect 8116 -1076 8120 -1044
rect 8080 -1124 8120 -1076
rect 8080 -1156 8084 -1124
rect 8116 -1156 8120 -1124
rect 8080 -1204 8120 -1156
rect 8080 -1236 8084 -1204
rect 8116 -1236 8120 -1204
rect 8080 -1284 8120 -1236
rect 8080 -1316 8084 -1284
rect 8116 -1316 8120 -1284
rect 8080 -1364 8120 -1316
rect 8080 -1396 8084 -1364
rect 8116 -1396 8120 -1364
rect 8080 -1444 8120 -1396
rect 8080 -1476 8084 -1444
rect 8116 -1476 8120 -1444
rect 8080 -1524 8120 -1476
rect 8080 -1556 8084 -1524
rect 8116 -1556 8120 -1524
rect 8080 -1604 8120 -1556
rect 8080 -1636 8084 -1604
rect 8116 -1636 8120 -1604
rect 8080 -1684 8120 -1636
rect 8080 -1716 8084 -1684
rect 8116 -1716 8120 -1684
rect 8080 -1764 8120 -1716
rect 8080 -1796 8084 -1764
rect 8116 -1796 8120 -1764
rect 8080 -1844 8120 -1796
rect 8080 -1876 8084 -1844
rect 8116 -1876 8120 -1844
rect 8080 -1924 8120 -1876
rect 8080 -1956 8084 -1924
rect 8116 -1956 8120 -1924
rect 8080 -2004 8120 -1956
rect 8080 -2036 8084 -2004
rect 8116 -2036 8120 -2004
rect 8080 -2084 8120 -2036
rect 8080 -2116 8084 -2084
rect 8116 -2116 8120 -2084
rect 8080 -2164 8120 -2116
rect 8080 -2196 8084 -2164
rect 8116 -2196 8120 -2164
rect 8080 -2244 8120 -2196
rect 8080 -2276 8084 -2244
rect 8116 -2276 8120 -2244
rect 8080 -2324 8120 -2276
rect 8080 -2356 8084 -2324
rect 8116 -2356 8120 -2324
rect 8080 -2404 8120 -2356
rect 8080 -2436 8084 -2404
rect 8116 -2436 8120 -2404
rect 8080 -2484 8120 -2436
rect 8080 -2516 8084 -2484
rect 8116 -2516 8120 -2484
rect 8080 -2564 8120 -2516
rect 8080 -2596 8084 -2564
rect 8116 -2596 8120 -2564
rect 8080 -2644 8120 -2596
rect 8080 -2676 8084 -2644
rect 8116 -2676 8120 -2644
rect 8080 -2724 8120 -2676
rect 8080 -2756 8084 -2724
rect 8116 -2756 8120 -2724
rect 8080 -2804 8120 -2756
rect 8080 -2836 8084 -2804
rect 8116 -2836 8120 -2804
rect 8080 -2884 8120 -2836
rect 8080 -2916 8084 -2884
rect 8116 -2916 8120 -2884
rect 8080 -2964 8120 -2916
rect 8080 -2996 8084 -2964
rect 8116 -2996 8120 -2964
rect 8080 -3044 8120 -2996
rect 8080 -3076 8084 -3044
rect 8116 -3076 8120 -3044
rect 8080 -3124 8120 -3076
rect 8080 -3156 8084 -3124
rect 8116 -3156 8120 -3124
rect 8080 -3204 8120 -3156
rect 8080 -3236 8084 -3204
rect 8116 -3236 8120 -3204
rect 8080 -3284 8120 -3236
rect 8080 -3316 8084 -3284
rect 8116 -3316 8120 -3284
rect 8080 -3364 8120 -3316
rect 8080 -3396 8084 -3364
rect 8116 -3396 8120 -3364
rect 8080 -3444 8120 -3396
rect 8080 -3476 8084 -3444
rect 8116 -3476 8120 -3444
rect 8080 -3524 8120 -3476
rect 8080 -3556 8084 -3524
rect 8116 -3556 8120 -3524
rect 8080 -3604 8120 -3556
rect 8080 -3636 8084 -3604
rect 8116 -3636 8120 -3604
rect 8080 -3684 8120 -3636
rect 8080 -3716 8084 -3684
rect 8116 -3716 8120 -3684
rect 8080 -3720 8120 -3716
rect 8160 1036 8200 1040
rect 8160 1004 8164 1036
rect 8196 1004 8200 1036
rect 8160 956 8200 1004
rect 8160 924 8164 956
rect 8196 924 8200 956
rect 8160 876 8200 924
rect 8160 844 8164 876
rect 8196 844 8200 876
rect 8160 796 8200 844
rect 8160 764 8164 796
rect 8196 764 8200 796
rect 8160 716 8200 764
rect 8160 684 8164 716
rect 8196 684 8200 716
rect 8160 636 8200 684
rect 8160 604 8164 636
rect 8196 604 8200 636
rect 8160 556 8200 604
rect 8160 524 8164 556
rect 8196 524 8200 556
rect 8160 476 8200 524
rect 8160 444 8164 476
rect 8196 444 8200 476
rect 8160 396 8200 444
rect 8160 364 8164 396
rect 8196 364 8200 396
rect 8160 316 8200 364
rect 8160 284 8164 316
rect 8196 284 8200 316
rect 8160 236 8200 284
rect 8160 204 8164 236
rect 8196 204 8200 236
rect 8160 156 8200 204
rect 8160 124 8164 156
rect 8196 124 8200 156
rect 8160 76 8200 124
rect 8160 44 8164 76
rect 8196 44 8200 76
rect 8160 -4 8200 44
rect 8160 -36 8164 -4
rect 8196 -36 8200 -4
rect 8160 -84 8200 -36
rect 8160 -116 8164 -84
rect 8196 -116 8200 -84
rect 8160 -164 8200 -116
rect 8160 -196 8164 -164
rect 8196 -196 8200 -164
rect 8160 -244 8200 -196
rect 8160 -276 8164 -244
rect 8196 -276 8200 -244
rect 8160 -324 8200 -276
rect 8160 -356 8164 -324
rect 8196 -356 8200 -324
rect 8160 -404 8200 -356
rect 8160 -436 8164 -404
rect 8196 -436 8200 -404
rect 8160 -484 8200 -436
rect 8160 -516 8164 -484
rect 8196 -516 8200 -484
rect 8160 -564 8200 -516
rect 8160 -596 8164 -564
rect 8196 -596 8200 -564
rect 8160 -644 8200 -596
rect 8160 -676 8164 -644
rect 8196 -676 8200 -644
rect 8160 -724 8200 -676
rect 8160 -756 8164 -724
rect 8196 -756 8200 -724
rect 8160 -804 8200 -756
rect 8160 -836 8164 -804
rect 8196 -836 8200 -804
rect 8160 -884 8200 -836
rect 8160 -916 8164 -884
rect 8196 -916 8200 -884
rect 8160 -964 8200 -916
rect 8160 -996 8164 -964
rect 8196 -996 8200 -964
rect 8160 -1044 8200 -996
rect 8160 -1076 8164 -1044
rect 8196 -1076 8200 -1044
rect 8160 -1124 8200 -1076
rect 8160 -1156 8164 -1124
rect 8196 -1156 8200 -1124
rect 8160 -1204 8200 -1156
rect 8160 -1236 8164 -1204
rect 8196 -1236 8200 -1204
rect 8160 -1284 8200 -1236
rect 8160 -1316 8164 -1284
rect 8196 -1316 8200 -1284
rect 8160 -1364 8200 -1316
rect 8160 -1396 8164 -1364
rect 8196 -1396 8200 -1364
rect 8160 -1444 8200 -1396
rect 8160 -1476 8164 -1444
rect 8196 -1476 8200 -1444
rect 8160 -1524 8200 -1476
rect 8160 -1556 8164 -1524
rect 8196 -1556 8200 -1524
rect 8160 -1604 8200 -1556
rect 8160 -1636 8164 -1604
rect 8196 -1636 8200 -1604
rect 8160 -1684 8200 -1636
rect 8160 -1716 8164 -1684
rect 8196 -1716 8200 -1684
rect 8160 -1764 8200 -1716
rect 8160 -1796 8164 -1764
rect 8196 -1796 8200 -1764
rect 8160 -1844 8200 -1796
rect 8160 -1876 8164 -1844
rect 8196 -1876 8200 -1844
rect 8160 -1924 8200 -1876
rect 8160 -1956 8164 -1924
rect 8196 -1956 8200 -1924
rect 8160 -2004 8200 -1956
rect 8160 -2036 8164 -2004
rect 8196 -2036 8200 -2004
rect 8160 -2084 8200 -2036
rect 8160 -2116 8164 -2084
rect 8196 -2116 8200 -2084
rect 8160 -2164 8200 -2116
rect 8160 -2196 8164 -2164
rect 8196 -2196 8200 -2164
rect 8160 -2244 8200 -2196
rect 8160 -2276 8164 -2244
rect 8196 -2276 8200 -2244
rect 8160 -2324 8200 -2276
rect 8160 -2356 8164 -2324
rect 8196 -2356 8200 -2324
rect 8160 -2404 8200 -2356
rect 8160 -2436 8164 -2404
rect 8196 -2436 8200 -2404
rect 8160 -2484 8200 -2436
rect 8160 -2516 8164 -2484
rect 8196 -2516 8200 -2484
rect 8160 -2564 8200 -2516
rect 8160 -2596 8164 -2564
rect 8196 -2596 8200 -2564
rect 8160 -2644 8200 -2596
rect 8160 -2676 8164 -2644
rect 8196 -2676 8200 -2644
rect 8160 -2724 8200 -2676
rect 8160 -2756 8164 -2724
rect 8196 -2756 8200 -2724
rect 8160 -2804 8200 -2756
rect 8160 -2836 8164 -2804
rect 8196 -2836 8200 -2804
rect 8160 -2884 8200 -2836
rect 8160 -2916 8164 -2884
rect 8196 -2916 8200 -2884
rect 8160 -2964 8200 -2916
rect 8160 -2996 8164 -2964
rect 8196 -2996 8200 -2964
rect 8160 -3044 8200 -2996
rect 8160 -3076 8164 -3044
rect 8196 -3076 8200 -3044
rect 8160 -3124 8200 -3076
rect 8160 -3156 8164 -3124
rect 8196 -3156 8200 -3124
rect 8160 -3204 8200 -3156
rect 8160 -3236 8164 -3204
rect 8196 -3236 8200 -3204
rect 8160 -3284 8200 -3236
rect 8160 -3316 8164 -3284
rect 8196 -3316 8200 -3284
rect 8160 -3364 8200 -3316
rect 8160 -3396 8164 -3364
rect 8196 -3396 8200 -3364
rect 8160 -3444 8200 -3396
rect 8160 -3476 8164 -3444
rect 8196 -3476 8200 -3444
rect 8160 -3524 8200 -3476
rect 8160 -3556 8164 -3524
rect 8196 -3556 8200 -3524
rect 8160 -3604 8200 -3556
rect 8160 -3636 8164 -3604
rect 8196 -3636 8200 -3604
rect 8160 -3684 8200 -3636
rect 8160 -3716 8164 -3684
rect 8196 -3716 8200 -3684
rect 8160 -3720 8200 -3716
rect 8240 1036 8280 1040
rect 8240 1004 8244 1036
rect 8276 1004 8280 1036
rect 8240 956 8280 1004
rect 8240 924 8244 956
rect 8276 924 8280 956
rect 8240 876 8280 924
rect 8240 844 8244 876
rect 8276 844 8280 876
rect 8240 796 8280 844
rect 8240 764 8244 796
rect 8276 764 8280 796
rect 8240 716 8280 764
rect 8240 684 8244 716
rect 8276 684 8280 716
rect 8240 636 8280 684
rect 8240 604 8244 636
rect 8276 604 8280 636
rect 8240 556 8280 604
rect 8240 524 8244 556
rect 8276 524 8280 556
rect 8240 476 8280 524
rect 8240 444 8244 476
rect 8276 444 8280 476
rect 8240 396 8280 444
rect 8240 364 8244 396
rect 8276 364 8280 396
rect 8240 316 8280 364
rect 8240 284 8244 316
rect 8276 284 8280 316
rect 8240 236 8280 284
rect 8240 204 8244 236
rect 8276 204 8280 236
rect 8240 156 8280 204
rect 8240 124 8244 156
rect 8276 124 8280 156
rect 8240 76 8280 124
rect 8240 44 8244 76
rect 8276 44 8280 76
rect 8240 -4 8280 44
rect 8240 -36 8244 -4
rect 8276 -36 8280 -4
rect 8240 -84 8280 -36
rect 8240 -116 8244 -84
rect 8276 -116 8280 -84
rect 8240 -164 8280 -116
rect 8240 -196 8244 -164
rect 8276 -196 8280 -164
rect 8240 -244 8280 -196
rect 8240 -276 8244 -244
rect 8276 -276 8280 -244
rect 8240 -324 8280 -276
rect 8240 -356 8244 -324
rect 8276 -356 8280 -324
rect 8240 -404 8280 -356
rect 8240 -436 8244 -404
rect 8276 -436 8280 -404
rect 8240 -484 8280 -436
rect 8240 -516 8244 -484
rect 8276 -516 8280 -484
rect 8240 -564 8280 -516
rect 8240 -596 8244 -564
rect 8276 -596 8280 -564
rect 8240 -644 8280 -596
rect 8240 -676 8244 -644
rect 8276 -676 8280 -644
rect 8240 -724 8280 -676
rect 8240 -756 8244 -724
rect 8276 -756 8280 -724
rect 8240 -804 8280 -756
rect 8240 -836 8244 -804
rect 8276 -836 8280 -804
rect 8240 -884 8280 -836
rect 8240 -916 8244 -884
rect 8276 -916 8280 -884
rect 8240 -964 8280 -916
rect 8240 -996 8244 -964
rect 8276 -996 8280 -964
rect 8240 -1044 8280 -996
rect 8240 -1076 8244 -1044
rect 8276 -1076 8280 -1044
rect 8240 -1124 8280 -1076
rect 8240 -1156 8244 -1124
rect 8276 -1156 8280 -1124
rect 8240 -1204 8280 -1156
rect 8240 -1236 8244 -1204
rect 8276 -1236 8280 -1204
rect 8240 -1284 8280 -1236
rect 8240 -1316 8244 -1284
rect 8276 -1316 8280 -1284
rect 8240 -1364 8280 -1316
rect 8240 -1396 8244 -1364
rect 8276 -1396 8280 -1364
rect 8240 -1444 8280 -1396
rect 8240 -1476 8244 -1444
rect 8276 -1476 8280 -1444
rect 8240 -1524 8280 -1476
rect 8240 -1556 8244 -1524
rect 8276 -1556 8280 -1524
rect 8240 -1604 8280 -1556
rect 8240 -1636 8244 -1604
rect 8276 -1636 8280 -1604
rect 8240 -1684 8280 -1636
rect 8240 -1716 8244 -1684
rect 8276 -1716 8280 -1684
rect 8240 -1764 8280 -1716
rect 8240 -1796 8244 -1764
rect 8276 -1796 8280 -1764
rect 8240 -1844 8280 -1796
rect 8240 -1876 8244 -1844
rect 8276 -1876 8280 -1844
rect 8240 -1924 8280 -1876
rect 8240 -1956 8244 -1924
rect 8276 -1956 8280 -1924
rect 8240 -2004 8280 -1956
rect 8240 -2036 8244 -2004
rect 8276 -2036 8280 -2004
rect 8240 -2084 8280 -2036
rect 8240 -2116 8244 -2084
rect 8276 -2116 8280 -2084
rect 8240 -2164 8280 -2116
rect 8240 -2196 8244 -2164
rect 8276 -2196 8280 -2164
rect 8240 -2244 8280 -2196
rect 8240 -2276 8244 -2244
rect 8276 -2276 8280 -2244
rect 8240 -2324 8280 -2276
rect 8240 -2356 8244 -2324
rect 8276 -2356 8280 -2324
rect 8240 -2404 8280 -2356
rect 8240 -2436 8244 -2404
rect 8276 -2436 8280 -2404
rect 8240 -2484 8280 -2436
rect 8240 -2516 8244 -2484
rect 8276 -2516 8280 -2484
rect 8240 -2564 8280 -2516
rect 8240 -2596 8244 -2564
rect 8276 -2596 8280 -2564
rect 8240 -2644 8280 -2596
rect 8240 -2676 8244 -2644
rect 8276 -2676 8280 -2644
rect 8240 -2724 8280 -2676
rect 8240 -2756 8244 -2724
rect 8276 -2756 8280 -2724
rect 8240 -2804 8280 -2756
rect 8240 -2836 8244 -2804
rect 8276 -2836 8280 -2804
rect 8240 -2884 8280 -2836
rect 8240 -2916 8244 -2884
rect 8276 -2916 8280 -2884
rect 8240 -2964 8280 -2916
rect 8240 -2996 8244 -2964
rect 8276 -2996 8280 -2964
rect 8240 -3044 8280 -2996
rect 8240 -3076 8244 -3044
rect 8276 -3076 8280 -3044
rect 8240 -3124 8280 -3076
rect 8240 -3156 8244 -3124
rect 8276 -3156 8280 -3124
rect 8240 -3204 8280 -3156
rect 8240 -3236 8244 -3204
rect 8276 -3236 8280 -3204
rect 8240 -3284 8280 -3236
rect 8240 -3316 8244 -3284
rect 8276 -3316 8280 -3284
rect 8240 -3364 8280 -3316
rect 8240 -3396 8244 -3364
rect 8276 -3396 8280 -3364
rect 8240 -3444 8280 -3396
rect 8240 -3476 8244 -3444
rect 8276 -3476 8280 -3444
rect 8240 -3524 8280 -3476
rect 8240 -3556 8244 -3524
rect 8276 -3556 8280 -3524
rect 8240 -3604 8280 -3556
rect 8240 -3636 8244 -3604
rect 8276 -3636 8280 -3604
rect 8240 -3684 8280 -3636
rect 8240 -3716 8244 -3684
rect 8276 -3716 8280 -3684
rect 8240 -3720 8280 -3716
rect 8320 1036 8360 1040
rect 8320 1004 8324 1036
rect 8356 1004 8360 1036
rect 8320 956 8360 1004
rect 8320 924 8324 956
rect 8356 924 8360 956
rect 8320 876 8360 924
rect 8320 844 8324 876
rect 8356 844 8360 876
rect 8320 796 8360 844
rect 8320 764 8324 796
rect 8356 764 8360 796
rect 8320 716 8360 764
rect 8320 684 8324 716
rect 8356 684 8360 716
rect 8320 636 8360 684
rect 8320 604 8324 636
rect 8356 604 8360 636
rect 8320 556 8360 604
rect 8320 524 8324 556
rect 8356 524 8360 556
rect 8320 476 8360 524
rect 8320 444 8324 476
rect 8356 444 8360 476
rect 8320 396 8360 444
rect 8320 364 8324 396
rect 8356 364 8360 396
rect 8320 316 8360 364
rect 8320 284 8324 316
rect 8356 284 8360 316
rect 8320 236 8360 284
rect 8320 204 8324 236
rect 8356 204 8360 236
rect 8320 156 8360 204
rect 8320 124 8324 156
rect 8356 124 8360 156
rect 8320 76 8360 124
rect 8320 44 8324 76
rect 8356 44 8360 76
rect 8320 -4 8360 44
rect 8320 -36 8324 -4
rect 8356 -36 8360 -4
rect 8320 -84 8360 -36
rect 8320 -116 8324 -84
rect 8356 -116 8360 -84
rect 8320 -164 8360 -116
rect 8320 -196 8324 -164
rect 8356 -196 8360 -164
rect 8320 -244 8360 -196
rect 8320 -276 8324 -244
rect 8356 -276 8360 -244
rect 8320 -324 8360 -276
rect 8320 -356 8324 -324
rect 8356 -356 8360 -324
rect 8320 -404 8360 -356
rect 8320 -436 8324 -404
rect 8356 -436 8360 -404
rect 8320 -484 8360 -436
rect 8320 -516 8324 -484
rect 8356 -516 8360 -484
rect 8320 -564 8360 -516
rect 8320 -596 8324 -564
rect 8356 -596 8360 -564
rect 8320 -644 8360 -596
rect 8320 -676 8324 -644
rect 8356 -676 8360 -644
rect 8320 -724 8360 -676
rect 8320 -756 8324 -724
rect 8356 -756 8360 -724
rect 8320 -804 8360 -756
rect 8320 -836 8324 -804
rect 8356 -836 8360 -804
rect 8320 -884 8360 -836
rect 8320 -916 8324 -884
rect 8356 -916 8360 -884
rect 8320 -964 8360 -916
rect 8320 -996 8324 -964
rect 8356 -996 8360 -964
rect 8320 -1044 8360 -996
rect 8320 -1076 8324 -1044
rect 8356 -1076 8360 -1044
rect 8320 -1124 8360 -1076
rect 8320 -1156 8324 -1124
rect 8356 -1156 8360 -1124
rect 8320 -1204 8360 -1156
rect 8320 -1236 8324 -1204
rect 8356 -1236 8360 -1204
rect 8320 -1284 8360 -1236
rect 8320 -1316 8324 -1284
rect 8356 -1316 8360 -1284
rect 8320 -1364 8360 -1316
rect 8320 -1396 8324 -1364
rect 8356 -1396 8360 -1364
rect 8320 -1444 8360 -1396
rect 8320 -1476 8324 -1444
rect 8356 -1476 8360 -1444
rect 8320 -1524 8360 -1476
rect 8320 -1556 8324 -1524
rect 8356 -1556 8360 -1524
rect 8320 -1604 8360 -1556
rect 8320 -1636 8324 -1604
rect 8356 -1636 8360 -1604
rect 8320 -1684 8360 -1636
rect 8320 -1716 8324 -1684
rect 8356 -1716 8360 -1684
rect 8320 -1764 8360 -1716
rect 8320 -1796 8324 -1764
rect 8356 -1796 8360 -1764
rect 8320 -1844 8360 -1796
rect 8320 -1876 8324 -1844
rect 8356 -1876 8360 -1844
rect 8320 -1924 8360 -1876
rect 8320 -1956 8324 -1924
rect 8356 -1956 8360 -1924
rect 8320 -2004 8360 -1956
rect 8320 -2036 8324 -2004
rect 8356 -2036 8360 -2004
rect 8320 -2084 8360 -2036
rect 8320 -2116 8324 -2084
rect 8356 -2116 8360 -2084
rect 8320 -2164 8360 -2116
rect 8320 -2196 8324 -2164
rect 8356 -2196 8360 -2164
rect 8320 -2244 8360 -2196
rect 8320 -2276 8324 -2244
rect 8356 -2276 8360 -2244
rect 8320 -2324 8360 -2276
rect 8320 -2356 8324 -2324
rect 8356 -2356 8360 -2324
rect 8320 -2404 8360 -2356
rect 8320 -2436 8324 -2404
rect 8356 -2436 8360 -2404
rect 8320 -2484 8360 -2436
rect 8320 -2516 8324 -2484
rect 8356 -2516 8360 -2484
rect 8320 -2564 8360 -2516
rect 8320 -2596 8324 -2564
rect 8356 -2596 8360 -2564
rect 8320 -2644 8360 -2596
rect 8320 -2676 8324 -2644
rect 8356 -2676 8360 -2644
rect 8320 -2724 8360 -2676
rect 8320 -2756 8324 -2724
rect 8356 -2756 8360 -2724
rect 8320 -2804 8360 -2756
rect 8320 -2836 8324 -2804
rect 8356 -2836 8360 -2804
rect 8320 -2884 8360 -2836
rect 8320 -2916 8324 -2884
rect 8356 -2916 8360 -2884
rect 8320 -2964 8360 -2916
rect 8320 -2996 8324 -2964
rect 8356 -2996 8360 -2964
rect 8320 -3044 8360 -2996
rect 8320 -3076 8324 -3044
rect 8356 -3076 8360 -3044
rect 8320 -3124 8360 -3076
rect 8320 -3156 8324 -3124
rect 8356 -3156 8360 -3124
rect 8320 -3204 8360 -3156
rect 8320 -3236 8324 -3204
rect 8356 -3236 8360 -3204
rect 8320 -3284 8360 -3236
rect 8320 -3316 8324 -3284
rect 8356 -3316 8360 -3284
rect 8320 -3364 8360 -3316
rect 8320 -3396 8324 -3364
rect 8356 -3396 8360 -3364
rect 8320 -3444 8360 -3396
rect 8320 -3476 8324 -3444
rect 8356 -3476 8360 -3444
rect 8320 -3524 8360 -3476
rect 8320 -3556 8324 -3524
rect 8356 -3556 8360 -3524
rect 8320 -3604 8360 -3556
rect 8320 -3636 8324 -3604
rect 8356 -3636 8360 -3604
rect 8320 -3684 8360 -3636
rect 8320 -3716 8324 -3684
rect 8356 -3716 8360 -3684
rect 8320 -3720 8360 -3716
rect 8400 1036 8440 1040
rect 8400 1004 8404 1036
rect 8436 1004 8440 1036
rect 8400 956 8440 1004
rect 8400 924 8404 956
rect 8436 924 8440 956
rect 8400 876 8440 924
rect 8400 844 8404 876
rect 8436 844 8440 876
rect 8400 796 8440 844
rect 8400 764 8404 796
rect 8436 764 8440 796
rect 8400 716 8440 764
rect 8400 684 8404 716
rect 8436 684 8440 716
rect 8400 636 8440 684
rect 8400 604 8404 636
rect 8436 604 8440 636
rect 8400 556 8440 604
rect 8400 524 8404 556
rect 8436 524 8440 556
rect 8400 476 8440 524
rect 8400 444 8404 476
rect 8436 444 8440 476
rect 8400 396 8440 444
rect 8400 364 8404 396
rect 8436 364 8440 396
rect 8400 316 8440 364
rect 8400 284 8404 316
rect 8436 284 8440 316
rect 8400 236 8440 284
rect 8400 204 8404 236
rect 8436 204 8440 236
rect 8400 156 8440 204
rect 8400 124 8404 156
rect 8436 124 8440 156
rect 8400 76 8440 124
rect 8400 44 8404 76
rect 8436 44 8440 76
rect 8400 -4 8440 44
rect 8400 -36 8404 -4
rect 8436 -36 8440 -4
rect 8400 -84 8440 -36
rect 8400 -116 8404 -84
rect 8436 -116 8440 -84
rect 8400 -164 8440 -116
rect 8400 -196 8404 -164
rect 8436 -196 8440 -164
rect 8400 -244 8440 -196
rect 8400 -276 8404 -244
rect 8436 -276 8440 -244
rect 8400 -324 8440 -276
rect 8400 -356 8404 -324
rect 8436 -356 8440 -324
rect 8400 -404 8440 -356
rect 8400 -436 8404 -404
rect 8436 -436 8440 -404
rect 8400 -484 8440 -436
rect 8400 -516 8404 -484
rect 8436 -516 8440 -484
rect 8400 -564 8440 -516
rect 8400 -596 8404 -564
rect 8436 -596 8440 -564
rect 8400 -644 8440 -596
rect 8400 -676 8404 -644
rect 8436 -676 8440 -644
rect 8400 -724 8440 -676
rect 8400 -756 8404 -724
rect 8436 -756 8440 -724
rect 8400 -804 8440 -756
rect 8400 -836 8404 -804
rect 8436 -836 8440 -804
rect 8400 -884 8440 -836
rect 8400 -916 8404 -884
rect 8436 -916 8440 -884
rect 8400 -964 8440 -916
rect 8400 -996 8404 -964
rect 8436 -996 8440 -964
rect 8400 -1044 8440 -996
rect 8400 -1076 8404 -1044
rect 8436 -1076 8440 -1044
rect 8400 -1124 8440 -1076
rect 8400 -1156 8404 -1124
rect 8436 -1156 8440 -1124
rect 8400 -1204 8440 -1156
rect 8400 -1236 8404 -1204
rect 8436 -1236 8440 -1204
rect 8400 -1284 8440 -1236
rect 8400 -1316 8404 -1284
rect 8436 -1316 8440 -1284
rect 8400 -1364 8440 -1316
rect 8400 -1396 8404 -1364
rect 8436 -1396 8440 -1364
rect 8400 -1444 8440 -1396
rect 8400 -1476 8404 -1444
rect 8436 -1476 8440 -1444
rect 8400 -1524 8440 -1476
rect 8400 -1556 8404 -1524
rect 8436 -1556 8440 -1524
rect 8400 -1604 8440 -1556
rect 8400 -1636 8404 -1604
rect 8436 -1636 8440 -1604
rect 8400 -1684 8440 -1636
rect 8400 -1716 8404 -1684
rect 8436 -1716 8440 -1684
rect 8400 -1764 8440 -1716
rect 8400 -1796 8404 -1764
rect 8436 -1796 8440 -1764
rect 8400 -1844 8440 -1796
rect 8400 -1876 8404 -1844
rect 8436 -1876 8440 -1844
rect 8400 -1924 8440 -1876
rect 8400 -1956 8404 -1924
rect 8436 -1956 8440 -1924
rect 8400 -2004 8440 -1956
rect 8400 -2036 8404 -2004
rect 8436 -2036 8440 -2004
rect 8400 -2084 8440 -2036
rect 8400 -2116 8404 -2084
rect 8436 -2116 8440 -2084
rect 8400 -2164 8440 -2116
rect 8400 -2196 8404 -2164
rect 8436 -2196 8440 -2164
rect 8400 -2244 8440 -2196
rect 8400 -2276 8404 -2244
rect 8436 -2276 8440 -2244
rect 8400 -2324 8440 -2276
rect 8400 -2356 8404 -2324
rect 8436 -2356 8440 -2324
rect 8400 -2404 8440 -2356
rect 8400 -2436 8404 -2404
rect 8436 -2436 8440 -2404
rect 8400 -2484 8440 -2436
rect 8400 -2516 8404 -2484
rect 8436 -2516 8440 -2484
rect 8400 -2564 8440 -2516
rect 8400 -2596 8404 -2564
rect 8436 -2596 8440 -2564
rect 8400 -2644 8440 -2596
rect 8400 -2676 8404 -2644
rect 8436 -2676 8440 -2644
rect 8400 -2724 8440 -2676
rect 8400 -2756 8404 -2724
rect 8436 -2756 8440 -2724
rect 8400 -2804 8440 -2756
rect 8400 -2836 8404 -2804
rect 8436 -2836 8440 -2804
rect 8400 -2884 8440 -2836
rect 8400 -2916 8404 -2884
rect 8436 -2916 8440 -2884
rect 8400 -2964 8440 -2916
rect 8400 -2996 8404 -2964
rect 8436 -2996 8440 -2964
rect 8400 -3044 8440 -2996
rect 8400 -3076 8404 -3044
rect 8436 -3076 8440 -3044
rect 8400 -3124 8440 -3076
rect 8400 -3156 8404 -3124
rect 8436 -3156 8440 -3124
rect 8400 -3204 8440 -3156
rect 8400 -3236 8404 -3204
rect 8436 -3236 8440 -3204
rect 8400 -3284 8440 -3236
rect 8400 -3316 8404 -3284
rect 8436 -3316 8440 -3284
rect 8400 -3364 8440 -3316
rect 8400 -3396 8404 -3364
rect 8436 -3396 8440 -3364
rect 8400 -3444 8440 -3396
rect 8400 -3476 8404 -3444
rect 8436 -3476 8440 -3444
rect 8400 -3524 8440 -3476
rect 8400 -3556 8404 -3524
rect 8436 -3556 8440 -3524
rect 8400 -3604 8440 -3556
rect 8400 -3636 8404 -3604
rect 8436 -3636 8440 -3604
rect 8400 -3684 8440 -3636
rect 8400 -3716 8404 -3684
rect 8436 -3716 8440 -3684
rect 8400 -3720 8440 -3716
rect 8480 1036 8520 1040
rect 8480 1004 8484 1036
rect 8516 1004 8520 1036
rect 8480 956 8520 1004
rect 8480 924 8484 956
rect 8516 924 8520 956
rect 8480 876 8520 924
rect 8480 844 8484 876
rect 8516 844 8520 876
rect 8480 796 8520 844
rect 8480 764 8484 796
rect 8516 764 8520 796
rect 8480 716 8520 764
rect 8480 684 8484 716
rect 8516 684 8520 716
rect 8480 636 8520 684
rect 8480 604 8484 636
rect 8516 604 8520 636
rect 8480 556 8520 604
rect 8480 524 8484 556
rect 8516 524 8520 556
rect 8480 476 8520 524
rect 8480 444 8484 476
rect 8516 444 8520 476
rect 8480 396 8520 444
rect 8480 364 8484 396
rect 8516 364 8520 396
rect 8480 316 8520 364
rect 8480 284 8484 316
rect 8516 284 8520 316
rect 8480 236 8520 284
rect 8480 204 8484 236
rect 8516 204 8520 236
rect 8480 156 8520 204
rect 8480 124 8484 156
rect 8516 124 8520 156
rect 8480 76 8520 124
rect 8480 44 8484 76
rect 8516 44 8520 76
rect 8480 -4 8520 44
rect 8480 -36 8484 -4
rect 8516 -36 8520 -4
rect 8480 -84 8520 -36
rect 8480 -116 8484 -84
rect 8516 -116 8520 -84
rect 8480 -164 8520 -116
rect 8480 -196 8484 -164
rect 8516 -196 8520 -164
rect 8480 -244 8520 -196
rect 8480 -276 8484 -244
rect 8516 -276 8520 -244
rect 8480 -324 8520 -276
rect 8480 -356 8484 -324
rect 8516 -356 8520 -324
rect 8480 -404 8520 -356
rect 8480 -436 8484 -404
rect 8516 -436 8520 -404
rect 8480 -484 8520 -436
rect 8480 -516 8484 -484
rect 8516 -516 8520 -484
rect 8480 -564 8520 -516
rect 8480 -596 8484 -564
rect 8516 -596 8520 -564
rect 8480 -644 8520 -596
rect 8480 -676 8484 -644
rect 8516 -676 8520 -644
rect 8480 -724 8520 -676
rect 8480 -756 8484 -724
rect 8516 -756 8520 -724
rect 8480 -804 8520 -756
rect 8480 -836 8484 -804
rect 8516 -836 8520 -804
rect 8480 -884 8520 -836
rect 8480 -916 8484 -884
rect 8516 -916 8520 -884
rect 8480 -964 8520 -916
rect 8480 -996 8484 -964
rect 8516 -996 8520 -964
rect 8480 -1044 8520 -996
rect 8480 -1076 8484 -1044
rect 8516 -1076 8520 -1044
rect 8480 -1124 8520 -1076
rect 8480 -1156 8484 -1124
rect 8516 -1156 8520 -1124
rect 8480 -1204 8520 -1156
rect 8480 -1236 8484 -1204
rect 8516 -1236 8520 -1204
rect 8480 -1284 8520 -1236
rect 8480 -1316 8484 -1284
rect 8516 -1316 8520 -1284
rect 8480 -1364 8520 -1316
rect 8480 -1396 8484 -1364
rect 8516 -1396 8520 -1364
rect 8480 -1444 8520 -1396
rect 8480 -1476 8484 -1444
rect 8516 -1476 8520 -1444
rect 8480 -1524 8520 -1476
rect 8480 -1556 8484 -1524
rect 8516 -1556 8520 -1524
rect 8480 -1604 8520 -1556
rect 8480 -1636 8484 -1604
rect 8516 -1636 8520 -1604
rect 8480 -1684 8520 -1636
rect 8480 -1716 8484 -1684
rect 8516 -1716 8520 -1684
rect 8480 -1764 8520 -1716
rect 8480 -1796 8484 -1764
rect 8516 -1796 8520 -1764
rect 8480 -1844 8520 -1796
rect 8480 -1876 8484 -1844
rect 8516 -1876 8520 -1844
rect 8480 -1924 8520 -1876
rect 8480 -1956 8484 -1924
rect 8516 -1956 8520 -1924
rect 8480 -2004 8520 -1956
rect 8480 -2036 8484 -2004
rect 8516 -2036 8520 -2004
rect 8480 -2084 8520 -2036
rect 8480 -2116 8484 -2084
rect 8516 -2116 8520 -2084
rect 8480 -2164 8520 -2116
rect 8480 -2196 8484 -2164
rect 8516 -2196 8520 -2164
rect 8480 -2244 8520 -2196
rect 8480 -2276 8484 -2244
rect 8516 -2276 8520 -2244
rect 8480 -2324 8520 -2276
rect 8480 -2356 8484 -2324
rect 8516 -2356 8520 -2324
rect 8480 -2404 8520 -2356
rect 8480 -2436 8484 -2404
rect 8516 -2436 8520 -2404
rect 8480 -2484 8520 -2436
rect 8480 -2516 8484 -2484
rect 8516 -2516 8520 -2484
rect 8480 -2564 8520 -2516
rect 8480 -2596 8484 -2564
rect 8516 -2596 8520 -2564
rect 8480 -2644 8520 -2596
rect 8480 -2676 8484 -2644
rect 8516 -2676 8520 -2644
rect 8480 -2724 8520 -2676
rect 8480 -2756 8484 -2724
rect 8516 -2756 8520 -2724
rect 8480 -2804 8520 -2756
rect 8480 -2836 8484 -2804
rect 8516 -2836 8520 -2804
rect 8480 -2884 8520 -2836
rect 8480 -2916 8484 -2884
rect 8516 -2916 8520 -2884
rect 8480 -2964 8520 -2916
rect 8480 -2996 8484 -2964
rect 8516 -2996 8520 -2964
rect 8480 -3044 8520 -2996
rect 8480 -3076 8484 -3044
rect 8516 -3076 8520 -3044
rect 8480 -3124 8520 -3076
rect 8480 -3156 8484 -3124
rect 8516 -3156 8520 -3124
rect 8480 -3204 8520 -3156
rect 8480 -3236 8484 -3204
rect 8516 -3236 8520 -3204
rect 8480 -3284 8520 -3236
rect 8480 -3316 8484 -3284
rect 8516 -3316 8520 -3284
rect 8480 -3364 8520 -3316
rect 8480 -3396 8484 -3364
rect 8516 -3396 8520 -3364
rect 8480 -3444 8520 -3396
rect 8480 -3476 8484 -3444
rect 8516 -3476 8520 -3444
rect 8480 -3524 8520 -3476
rect 8480 -3556 8484 -3524
rect 8516 -3556 8520 -3524
rect 8480 -3604 8520 -3556
rect 8480 -3636 8484 -3604
rect 8516 -3636 8520 -3604
rect 8480 -3684 8520 -3636
rect 8480 -3716 8484 -3684
rect 8516 -3716 8520 -3684
rect 8480 -3720 8520 -3716
rect 8560 1036 8600 1040
rect 8560 1004 8564 1036
rect 8596 1004 8600 1036
rect 8560 956 8600 1004
rect 8560 924 8564 956
rect 8596 924 8600 956
rect 8560 876 8600 924
rect 8560 844 8564 876
rect 8596 844 8600 876
rect 8560 796 8600 844
rect 8560 764 8564 796
rect 8596 764 8600 796
rect 8560 716 8600 764
rect 8560 684 8564 716
rect 8596 684 8600 716
rect 8560 636 8600 684
rect 8560 604 8564 636
rect 8596 604 8600 636
rect 8560 556 8600 604
rect 8560 524 8564 556
rect 8596 524 8600 556
rect 8560 476 8600 524
rect 8560 444 8564 476
rect 8596 444 8600 476
rect 8560 396 8600 444
rect 8560 364 8564 396
rect 8596 364 8600 396
rect 8560 316 8600 364
rect 8560 284 8564 316
rect 8596 284 8600 316
rect 8560 236 8600 284
rect 8560 204 8564 236
rect 8596 204 8600 236
rect 8560 156 8600 204
rect 8560 124 8564 156
rect 8596 124 8600 156
rect 8560 76 8600 124
rect 8560 44 8564 76
rect 8596 44 8600 76
rect 8560 -4 8600 44
rect 8560 -36 8564 -4
rect 8596 -36 8600 -4
rect 8560 -84 8600 -36
rect 8560 -116 8564 -84
rect 8596 -116 8600 -84
rect 8560 -164 8600 -116
rect 8560 -196 8564 -164
rect 8596 -196 8600 -164
rect 8560 -244 8600 -196
rect 8560 -276 8564 -244
rect 8596 -276 8600 -244
rect 8560 -324 8600 -276
rect 8560 -356 8564 -324
rect 8596 -356 8600 -324
rect 8560 -404 8600 -356
rect 8560 -436 8564 -404
rect 8596 -436 8600 -404
rect 8560 -484 8600 -436
rect 8560 -516 8564 -484
rect 8596 -516 8600 -484
rect 8560 -564 8600 -516
rect 8560 -596 8564 -564
rect 8596 -596 8600 -564
rect 8560 -644 8600 -596
rect 8560 -676 8564 -644
rect 8596 -676 8600 -644
rect 8560 -724 8600 -676
rect 8560 -756 8564 -724
rect 8596 -756 8600 -724
rect 8560 -804 8600 -756
rect 8560 -836 8564 -804
rect 8596 -836 8600 -804
rect 8560 -884 8600 -836
rect 8560 -916 8564 -884
rect 8596 -916 8600 -884
rect 8560 -964 8600 -916
rect 8560 -996 8564 -964
rect 8596 -996 8600 -964
rect 8560 -1044 8600 -996
rect 8560 -1076 8564 -1044
rect 8596 -1076 8600 -1044
rect 8560 -1124 8600 -1076
rect 8560 -1156 8564 -1124
rect 8596 -1156 8600 -1124
rect 8560 -1204 8600 -1156
rect 8560 -1236 8564 -1204
rect 8596 -1236 8600 -1204
rect 8560 -1284 8600 -1236
rect 8560 -1316 8564 -1284
rect 8596 -1316 8600 -1284
rect 8560 -1364 8600 -1316
rect 8560 -1396 8564 -1364
rect 8596 -1396 8600 -1364
rect 8560 -1444 8600 -1396
rect 8560 -1476 8564 -1444
rect 8596 -1476 8600 -1444
rect 8560 -1524 8600 -1476
rect 8560 -1556 8564 -1524
rect 8596 -1556 8600 -1524
rect 8560 -1604 8600 -1556
rect 8560 -1636 8564 -1604
rect 8596 -1636 8600 -1604
rect 8560 -1684 8600 -1636
rect 8560 -1716 8564 -1684
rect 8596 -1716 8600 -1684
rect 8560 -1764 8600 -1716
rect 8560 -1796 8564 -1764
rect 8596 -1796 8600 -1764
rect 8560 -1844 8600 -1796
rect 8560 -1876 8564 -1844
rect 8596 -1876 8600 -1844
rect 8560 -1924 8600 -1876
rect 8560 -1956 8564 -1924
rect 8596 -1956 8600 -1924
rect 8560 -2004 8600 -1956
rect 8560 -2036 8564 -2004
rect 8596 -2036 8600 -2004
rect 8560 -2084 8600 -2036
rect 8560 -2116 8564 -2084
rect 8596 -2116 8600 -2084
rect 8560 -2164 8600 -2116
rect 8560 -2196 8564 -2164
rect 8596 -2196 8600 -2164
rect 8560 -2244 8600 -2196
rect 8560 -2276 8564 -2244
rect 8596 -2276 8600 -2244
rect 8560 -2324 8600 -2276
rect 8560 -2356 8564 -2324
rect 8596 -2356 8600 -2324
rect 8560 -2404 8600 -2356
rect 8560 -2436 8564 -2404
rect 8596 -2436 8600 -2404
rect 8560 -2484 8600 -2436
rect 8560 -2516 8564 -2484
rect 8596 -2516 8600 -2484
rect 8560 -2564 8600 -2516
rect 8560 -2596 8564 -2564
rect 8596 -2596 8600 -2564
rect 8560 -2644 8600 -2596
rect 8560 -2676 8564 -2644
rect 8596 -2676 8600 -2644
rect 8560 -2724 8600 -2676
rect 8560 -2756 8564 -2724
rect 8596 -2756 8600 -2724
rect 8560 -2804 8600 -2756
rect 8560 -2836 8564 -2804
rect 8596 -2836 8600 -2804
rect 8560 -2884 8600 -2836
rect 8560 -2916 8564 -2884
rect 8596 -2916 8600 -2884
rect 8560 -2964 8600 -2916
rect 8560 -2996 8564 -2964
rect 8596 -2996 8600 -2964
rect 8560 -3044 8600 -2996
rect 8560 -3076 8564 -3044
rect 8596 -3076 8600 -3044
rect 8560 -3124 8600 -3076
rect 8560 -3156 8564 -3124
rect 8596 -3156 8600 -3124
rect 8560 -3204 8600 -3156
rect 8560 -3236 8564 -3204
rect 8596 -3236 8600 -3204
rect 8560 -3284 8600 -3236
rect 8560 -3316 8564 -3284
rect 8596 -3316 8600 -3284
rect 8560 -3364 8600 -3316
rect 8560 -3396 8564 -3364
rect 8596 -3396 8600 -3364
rect 8560 -3444 8600 -3396
rect 8560 -3476 8564 -3444
rect 8596 -3476 8600 -3444
rect 8560 -3524 8600 -3476
rect 8560 -3556 8564 -3524
rect 8596 -3556 8600 -3524
rect 8560 -3604 8600 -3556
rect 8560 -3636 8564 -3604
rect 8596 -3636 8600 -3604
rect 8560 -3684 8600 -3636
rect 8560 -3716 8564 -3684
rect 8596 -3716 8600 -3684
rect 8560 -3720 8600 -3716
rect 8640 1036 8680 1040
rect 8640 1004 8644 1036
rect 8676 1004 8680 1036
rect 8640 956 8680 1004
rect 8640 924 8644 956
rect 8676 924 8680 956
rect 8640 876 8680 924
rect 8640 844 8644 876
rect 8676 844 8680 876
rect 8640 796 8680 844
rect 8640 764 8644 796
rect 8676 764 8680 796
rect 8640 716 8680 764
rect 8640 684 8644 716
rect 8676 684 8680 716
rect 8640 636 8680 684
rect 8640 604 8644 636
rect 8676 604 8680 636
rect 8640 556 8680 604
rect 8640 524 8644 556
rect 8676 524 8680 556
rect 8640 476 8680 524
rect 8640 444 8644 476
rect 8676 444 8680 476
rect 8640 396 8680 444
rect 8640 364 8644 396
rect 8676 364 8680 396
rect 8640 316 8680 364
rect 8640 284 8644 316
rect 8676 284 8680 316
rect 8640 236 8680 284
rect 8640 204 8644 236
rect 8676 204 8680 236
rect 8640 156 8680 204
rect 8640 124 8644 156
rect 8676 124 8680 156
rect 8640 76 8680 124
rect 8640 44 8644 76
rect 8676 44 8680 76
rect 8640 -4 8680 44
rect 8640 -36 8644 -4
rect 8676 -36 8680 -4
rect 8640 -84 8680 -36
rect 8640 -116 8644 -84
rect 8676 -116 8680 -84
rect 8640 -164 8680 -116
rect 8640 -196 8644 -164
rect 8676 -196 8680 -164
rect 8640 -244 8680 -196
rect 8640 -276 8644 -244
rect 8676 -276 8680 -244
rect 8640 -324 8680 -276
rect 8640 -356 8644 -324
rect 8676 -356 8680 -324
rect 8640 -404 8680 -356
rect 8640 -436 8644 -404
rect 8676 -436 8680 -404
rect 8640 -484 8680 -436
rect 8640 -516 8644 -484
rect 8676 -516 8680 -484
rect 8640 -564 8680 -516
rect 8640 -596 8644 -564
rect 8676 -596 8680 -564
rect 8640 -644 8680 -596
rect 8640 -676 8644 -644
rect 8676 -676 8680 -644
rect 8640 -724 8680 -676
rect 8640 -756 8644 -724
rect 8676 -756 8680 -724
rect 8640 -804 8680 -756
rect 8640 -836 8644 -804
rect 8676 -836 8680 -804
rect 8640 -884 8680 -836
rect 8640 -916 8644 -884
rect 8676 -916 8680 -884
rect 8640 -964 8680 -916
rect 8640 -996 8644 -964
rect 8676 -996 8680 -964
rect 8640 -1044 8680 -996
rect 8640 -1076 8644 -1044
rect 8676 -1076 8680 -1044
rect 8640 -1124 8680 -1076
rect 8640 -1156 8644 -1124
rect 8676 -1156 8680 -1124
rect 8640 -1204 8680 -1156
rect 8640 -1236 8644 -1204
rect 8676 -1236 8680 -1204
rect 8640 -1284 8680 -1236
rect 8640 -1316 8644 -1284
rect 8676 -1316 8680 -1284
rect 8640 -1364 8680 -1316
rect 8640 -1396 8644 -1364
rect 8676 -1396 8680 -1364
rect 8640 -1444 8680 -1396
rect 8640 -1476 8644 -1444
rect 8676 -1476 8680 -1444
rect 8640 -1524 8680 -1476
rect 8640 -1556 8644 -1524
rect 8676 -1556 8680 -1524
rect 8640 -1604 8680 -1556
rect 8640 -1636 8644 -1604
rect 8676 -1636 8680 -1604
rect 8640 -1684 8680 -1636
rect 8640 -1716 8644 -1684
rect 8676 -1716 8680 -1684
rect 8640 -1764 8680 -1716
rect 8640 -1796 8644 -1764
rect 8676 -1796 8680 -1764
rect 8640 -1844 8680 -1796
rect 8640 -1876 8644 -1844
rect 8676 -1876 8680 -1844
rect 8640 -1924 8680 -1876
rect 8640 -1956 8644 -1924
rect 8676 -1956 8680 -1924
rect 8640 -2004 8680 -1956
rect 8640 -2036 8644 -2004
rect 8676 -2036 8680 -2004
rect 8640 -2084 8680 -2036
rect 8640 -2116 8644 -2084
rect 8676 -2116 8680 -2084
rect 8640 -2164 8680 -2116
rect 8640 -2196 8644 -2164
rect 8676 -2196 8680 -2164
rect 8640 -2244 8680 -2196
rect 8640 -2276 8644 -2244
rect 8676 -2276 8680 -2244
rect 8640 -2324 8680 -2276
rect 8640 -2356 8644 -2324
rect 8676 -2356 8680 -2324
rect 8640 -2404 8680 -2356
rect 8640 -2436 8644 -2404
rect 8676 -2436 8680 -2404
rect 8640 -2484 8680 -2436
rect 8640 -2516 8644 -2484
rect 8676 -2516 8680 -2484
rect 8640 -2564 8680 -2516
rect 8640 -2596 8644 -2564
rect 8676 -2596 8680 -2564
rect 8640 -2644 8680 -2596
rect 8640 -2676 8644 -2644
rect 8676 -2676 8680 -2644
rect 8640 -2724 8680 -2676
rect 8640 -2756 8644 -2724
rect 8676 -2756 8680 -2724
rect 8640 -2804 8680 -2756
rect 8640 -2836 8644 -2804
rect 8676 -2836 8680 -2804
rect 8640 -2884 8680 -2836
rect 8640 -2916 8644 -2884
rect 8676 -2916 8680 -2884
rect 8640 -2964 8680 -2916
rect 8640 -2996 8644 -2964
rect 8676 -2996 8680 -2964
rect 8640 -3044 8680 -2996
rect 8640 -3076 8644 -3044
rect 8676 -3076 8680 -3044
rect 8640 -3124 8680 -3076
rect 8640 -3156 8644 -3124
rect 8676 -3156 8680 -3124
rect 8640 -3204 8680 -3156
rect 8640 -3236 8644 -3204
rect 8676 -3236 8680 -3204
rect 8640 -3284 8680 -3236
rect 8640 -3316 8644 -3284
rect 8676 -3316 8680 -3284
rect 8640 -3364 8680 -3316
rect 8640 -3396 8644 -3364
rect 8676 -3396 8680 -3364
rect 8640 -3444 8680 -3396
rect 8640 -3476 8644 -3444
rect 8676 -3476 8680 -3444
rect 8640 -3524 8680 -3476
rect 8640 -3556 8644 -3524
rect 8676 -3556 8680 -3524
rect 8640 -3604 8680 -3556
rect 8640 -3636 8644 -3604
rect 8676 -3636 8680 -3604
rect 8640 -3684 8680 -3636
rect 8640 -3716 8644 -3684
rect 8676 -3716 8680 -3684
rect 8640 -3720 8680 -3716
rect 8720 1036 8760 1040
rect 8720 1004 8724 1036
rect 8756 1004 8760 1036
rect 8720 956 8760 1004
rect 8720 924 8724 956
rect 8756 924 8760 956
rect 8720 876 8760 924
rect 8720 844 8724 876
rect 8756 844 8760 876
rect 8720 796 8760 844
rect 8720 764 8724 796
rect 8756 764 8760 796
rect 8720 716 8760 764
rect 8720 684 8724 716
rect 8756 684 8760 716
rect 8720 636 8760 684
rect 8720 604 8724 636
rect 8756 604 8760 636
rect 8720 556 8760 604
rect 8720 524 8724 556
rect 8756 524 8760 556
rect 8720 476 8760 524
rect 8720 444 8724 476
rect 8756 444 8760 476
rect 8720 396 8760 444
rect 8720 364 8724 396
rect 8756 364 8760 396
rect 8720 316 8760 364
rect 8720 284 8724 316
rect 8756 284 8760 316
rect 8720 236 8760 284
rect 8720 204 8724 236
rect 8756 204 8760 236
rect 8720 156 8760 204
rect 8720 124 8724 156
rect 8756 124 8760 156
rect 8720 76 8760 124
rect 8720 44 8724 76
rect 8756 44 8760 76
rect 8720 -4 8760 44
rect 8720 -36 8724 -4
rect 8756 -36 8760 -4
rect 8720 -84 8760 -36
rect 8720 -116 8724 -84
rect 8756 -116 8760 -84
rect 8720 -164 8760 -116
rect 8720 -196 8724 -164
rect 8756 -196 8760 -164
rect 8720 -244 8760 -196
rect 8720 -276 8724 -244
rect 8756 -276 8760 -244
rect 8720 -324 8760 -276
rect 8720 -356 8724 -324
rect 8756 -356 8760 -324
rect 8720 -404 8760 -356
rect 8720 -436 8724 -404
rect 8756 -436 8760 -404
rect 8720 -484 8760 -436
rect 8720 -516 8724 -484
rect 8756 -516 8760 -484
rect 8720 -564 8760 -516
rect 8720 -596 8724 -564
rect 8756 -596 8760 -564
rect 8720 -644 8760 -596
rect 8720 -676 8724 -644
rect 8756 -676 8760 -644
rect 8720 -724 8760 -676
rect 8720 -756 8724 -724
rect 8756 -756 8760 -724
rect 8720 -804 8760 -756
rect 8720 -836 8724 -804
rect 8756 -836 8760 -804
rect 8720 -884 8760 -836
rect 8720 -916 8724 -884
rect 8756 -916 8760 -884
rect 8720 -964 8760 -916
rect 8720 -996 8724 -964
rect 8756 -996 8760 -964
rect 8720 -1044 8760 -996
rect 8720 -1076 8724 -1044
rect 8756 -1076 8760 -1044
rect 8720 -1124 8760 -1076
rect 8720 -1156 8724 -1124
rect 8756 -1156 8760 -1124
rect 8720 -1204 8760 -1156
rect 8720 -1236 8724 -1204
rect 8756 -1236 8760 -1204
rect 8720 -1284 8760 -1236
rect 8720 -1316 8724 -1284
rect 8756 -1316 8760 -1284
rect 8720 -1364 8760 -1316
rect 8720 -1396 8724 -1364
rect 8756 -1396 8760 -1364
rect 8720 -1444 8760 -1396
rect 8720 -1476 8724 -1444
rect 8756 -1476 8760 -1444
rect 8720 -1524 8760 -1476
rect 8720 -1556 8724 -1524
rect 8756 -1556 8760 -1524
rect 8720 -1604 8760 -1556
rect 8720 -1636 8724 -1604
rect 8756 -1636 8760 -1604
rect 8720 -1684 8760 -1636
rect 8720 -1716 8724 -1684
rect 8756 -1716 8760 -1684
rect 8720 -1764 8760 -1716
rect 8720 -1796 8724 -1764
rect 8756 -1796 8760 -1764
rect 8720 -1844 8760 -1796
rect 8720 -1876 8724 -1844
rect 8756 -1876 8760 -1844
rect 8720 -1924 8760 -1876
rect 8720 -1956 8724 -1924
rect 8756 -1956 8760 -1924
rect 8720 -2004 8760 -1956
rect 8720 -2036 8724 -2004
rect 8756 -2036 8760 -2004
rect 8720 -2084 8760 -2036
rect 8720 -2116 8724 -2084
rect 8756 -2116 8760 -2084
rect 8720 -2164 8760 -2116
rect 8720 -2196 8724 -2164
rect 8756 -2196 8760 -2164
rect 8720 -2244 8760 -2196
rect 8720 -2276 8724 -2244
rect 8756 -2276 8760 -2244
rect 8720 -2324 8760 -2276
rect 8720 -2356 8724 -2324
rect 8756 -2356 8760 -2324
rect 8720 -2404 8760 -2356
rect 8720 -2436 8724 -2404
rect 8756 -2436 8760 -2404
rect 8720 -2484 8760 -2436
rect 8720 -2516 8724 -2484
rect 8756 -2516 8760 -2484
rect 8720 -2564 8760 -2516
rect 8720 -2596 8724 -2564
rect 8756 -2596 8760 -2564
rect 8720 -2644 8760 -2596
rect 8720 -2676 8724 -2644
rect 8756 -2676 8760 -2644
rect 8720 -2724 8760 -2676
rect 8720 -2756 8724 -2724
rect 8756 -2756 8760 -2724
rect 8720 -2804 8760 -2756
rect 8720 -2836 8724 -2804
rect 8756 -2836 8760 -2804
rect 8720 -2884 8760 -2836
rect 8720 -2916 8724 -2884
rect 8756 -2916 8760 -2884
rect 8720 -2964 8760 -2916
rect 8720 -2996 8724 -2964
rect 8756 -2996 8760 -2964
rect 8720 -3044 8760 -2996
rect 8720 -3076 8724 -3044
rect 8756 -3076 8760 -3044
rect 8720 -3124 8760 -3076
rect 8720 -3156 8724 -3124
rect 8756 -3156 8760 -3124
rect 8720 -3204 8760 -3156
rect 8720 -3236 8724 -3204
rect 8756 -3236 8760 -3204
rect 8720 -3284 8760 -3236
rect 8720 -3316 8724 -3284
rect 8756 -3316 8760 -3284
rect 8720 -3364 8760 -3316
rect 8720 -3396 8724 -3364
rect 8756 -3396 8760 -3364
rect 8720 -3444 8760 -3396
rect 8720 -3476 8724 -3444
rect 8756 -3476 8760 -3444
rect 8720 -3524 8760 -3476
rect 8720 -3556 8724 -3524
rect 8756 -3556 8760 -3524
rect 8720 -3604 8760 -3556
rect 8720 -3636 8724 -3604
rect 8756 -3636 8760 -3604
rect 8720 -3684 8760 -3636
rect 8720 -3716 8724 -3684
rect 8756 -3716 8760 -3684
rect 8720 -3720 8760 -3716
rect 8800 1036 8840 1040
rect 8800 1004 8804 1036
rect 8836 1004 8840 1036
rect 8800 956 8840 1004
rect 8800 924 8804 956
rect 8836 924 8840 956
rect 8800 876 8840 924
rect 8800 844 8804 876
rect 8836 844 8840 876
rect 8800 796 8840 844
rect 8800 764 8804 796
rect 8836 764 8840 796
rect 8800 716 8840 764
rect 8800 684 8804 716
rect 8836 684 8840 716
rect 8800 636 8840 684
rect 8800 604 8804 636
rect 8836 604 8840 636
rect 8800 556 8840 604
rect 8800 524 8804 556
rect 8836 524 8840 556
rect 8800 476 8840 524
rect 8800 444 8804 476
rect 8836 444 8840 476
rect 8800 396 8840 444
rect 8800 364 8804 396
rect 8836 364 8840 396
rect 8800 316 8840 364
rect 8800 284 8804 316
rect 8836 284 8840 316
rect 8800 236 8840 284
rect 8800 204 8804 236
rect 8836 204 8840 236
rect 8800 156 8840 204
rect 8800 124 8804 156
rect 8836 124 8840 156
rect 8800 76 8840 124
rect 8800 44 8804 76
rect 8836 44 8840 76
rect 8800 -4 8840 44
rect 8800 -36 8804 -4
rect 8836 -36 8840 -4
rect 8800 -84 8840 -36
rect 8800 -116 8804 -84
rect 8836 -116 8840 -84
rect 8800 -164 8840 -116
rect 8800 -196 8804 -164
rect 8836 -196 8840 -164
rect 8800 -244 8840 -196
rect 8800 -276 8804 -244
rect 8836 -276 8840 -244
rect 8800 -324 8840 -276
rect 8800 -356 8804 -324
rect 8836 -356 8840 -324
rect 8800 -404 8840 -356
rect 8800 -436 8804 -404
rect 8836 -436 8840 -404
rect 8800 -484 8840 -436
rect 8800 -516 8804 -484
rect 8836 -516 8840 -484
rect 8800 -564 8840 -516
rect 8800 -596 8804 -564
rect 8836 -596 8840 -564
rect 8800 -644 8840 -596
rect 8800 -676 8804 -644
rect 8836 -676 8840 -644
rect 8800 -724 8840 -676
rect 8800 -756 8804 -724
rect 8836 -756 8840 -724
rect 8800 -804 8840 -756
rect 8800 -836 8804 -804
rect 8836 -836 8840 -804
rect 8800 -884 8840 -836
rect 8800 -916 8804 -884
rect 8836 -916 8840 -884
rect 8800 -964 8840 -916
rect 8800 -996 8804 -964
rect 8836 -996 8840 -964
rect 8800 -1044 8840 -996
rect 8800 -1076 8804 -1044
rect 8836 -1076 8840 -1044
rect 8800 -1124 8840 -1076
rect 8800 -1156 8804 -1124
rect 8836 -1156 8840 -1124
rect 8800 -1204 8840 -1156
rect 8800 -1236 8804 -1204
rect 8836 -1236 8840 -1204
rect 8800 -1284 8840 -1236
rect 8800 -1316 8804 -1284
rect 8836 -1316 8840 -1284
rect 8800 -1364 8840 -1316
rect 8800 -1396 8804 -1364
rect 8836 -1396 8840 -1364
rect 8800 -1444 8840 -1396
rect 8800 -1476 8804 -1444
rect 8836 -1476 8840 -1444
rect 8800 -1524 8840 -1476
rect 8800 -1556 8804 -1524
rect 8836 -1556 8840 -1524
rect 8800 -1604 8840 -1556
rect 8800 -1636 8804 -1604
rect 8836 -1636 8840 -1604
rect 8800 -1684 8840 -1636
rect 8800 -1716 8804 -1684
rect 8836 -1716 8840 -1684
rect 8800 -1764 8840 -1716
rect 8800 -1796 8804 -1764
rect 8836 -1796 8840 -1764
rect 8800 -1844 8840 -1796
rect 8800 -1876 8804 -1844
rect 8836 -1876 8840 -1844
rect 8800 -1924 8840 -1876
rect 8800 -1956 8804 -1924
rect 8836 -1956 8840 -1924
rect 8800 -2004 8840 -1956
rect 8800 -2036 8804 -2004
rect 8836 -2036 8840 -2004
rect 8800 -2084 8840 -2036
rect 8800 -2116 8804 -2084
rect 8836 -2116 8840 -2084
rect 8800 -2164 8840 -2116
rect 8800 -2196 8804 -2164
rect 8836 -2196 8840 -2164
rect 8800 -2244 8840 -2196
rect 8800 -2276 8804 -2244
rect 8836 -2276 8840 -2244
rect 8800 -2324 8840 -2276
rect 8800 -2356 8804 -2324
rect 8836 -2356 8840 -2324
rect 8800 -2404 8840 -2356
rect 8800 -2436 8804 -2404
rect 8836 -2436 8840 -2404
rect 8800 -2484 8840 -2436
rect 8800 -2516 8804 -2484
rect 8836 -2516 8840 -2484
rect 8800 -2564 8840 -2516
rect 8800 -2596 8804 -2564
rect 8836 -2596 8840 -2564
rect 8800 -2644 8840 -2596
rect 8800 -2676 8804 -2644
rect 8836 -2676 8840 -2644
rect 8800 -2724 8840 -2676
rect 8800 -2756 8804 -2724
rect 8836 -2756 8840 -2724
rect 8800 -2804 8840 -2756
rect 8800 -2836 8804 -2804
rect 8836 -2836 8840 -2804
rect 8800 -2884 8840 -2836
rect 8800 -2916 8804 -2884
rect 8836 -2916 8840 -2884
rect 8800 -2964 8840 -2916
rect 8800 -2996 8804 -2964
rect 8836 -2996 8840 -2964
rect 8800 -3044 8840 -2996
rect 8800 -3076 8804 -3044
rect 8836 -3076 8840 -3044
rect 8800 -3124 8840 -3076
rect 8800 -3156 8804 -3124
rect 8836 -3156 8840 -3124
rect 8800 -3204 8840 -3156
rect 8800 -3236 8804 -3204
rect 8836 -3236 8840 -3204
rect 8800 -3284 8840 -3236
rect 8800 -3316 8804 -3284
rect 8836 -3316 8840 -3284
rect 8800 -3364 8840 -3316
rect 8800 -3396 8804 -3364
rect 8836 -3396 8840 -3364
rect 8800 -3444 8840 -3396
rect 8800 -3476 8804 -3444
rect 8836 -3476 8840 -3444
rect 8800 -3524 8840 -3476
rect 8800 -3556 8804 -3524
rect 8836 -3556 8840 -3524
rect 8800 -3604 8840 -3556
rect 8800 -3636 8804 -3604
rect 8836 -3636 8840 -3604
rect 8800 -3684 8840 -3636
rect 8800 -3716 8804 -3684
rect 8836 -3716 8840 -3684
rect 8800 -3720 8840 -3716
rect 8880 1036 8920 1040
rect 8880 1004 8884 1036
rect 8916 1004 8920 1036
rect 8880 956 8920 1004
rect 8880 924 8884 956
rect 8916 924 8920 956
rect 8880 876 8920 924
rect 8880 844 8884 876
rect 8916 844 8920 876
rect 8880 796 8920 844
rect 8880 764 8884 796
rect 8916 764 8920 796
rect 8880 716 8920 764
rect 8880 684 8884 716
rect 8916 684 8920 716
rect 8880 636 8920 684
rect 8880 604 8884 636
rect 8916 604 8920 636
rect 8880 556 8920 604
rect 8880 524 8884 556
rect 8916 524 8920 556
rect 8880 476 8920 524
rect 8880 444 8884 476
rect 8916 444 8920 476
rect 8880 396 8920 444
rect 8880 364 8884 396
rect 8916 364 8920 396
rect 8880 316 8920 364
rect 8880 284 8884 316
rect 8916 284 8920 316
rect 8880 236 8920 284
rect 8880 204 8884 236
rect 8916 204 8920 236
rect 8880 156 8920 204
rect 8880 124 8884 156
rect 8916 124 8920 156
rect 8880 76 8920 124
rect 8880 44 8884 76
rect 8916 44 8920 76
rect 8880 -4 8920 44
rect 8880 -36 8884 -4
rect 8916 -36 8920 -4
rect 8880 -84 8920 -36
rect 8880 -116 8884 -84
rect 8916 -116 8920 -84
rect 8880 -164 8920 -116
rect 8880 -196 8884 -164
rect 8916 -196 8920 -164
rect 8880 -244 8920 -196
rect 8880 -276 8884 -244
rect 8916 -276 8920 -244
rect 8880 -324 8920 -276
rect 8880 -356 8884 -324
rect 8916 -356 8920 -324
rect 8880 -404 8920 -356
rect 8880 -436 8884 -404
rect 8916 -436 8920 -404
rect 8880 -484 8920 -436
rect 8880 -516 8884 -484
rect 8916 -516 8920 -484
rect 8880 -564 8920 -516
rect 8880 -596 8884 -564
rect 8916 -596 8920 -564
rect 8880 -644 8920 -596
rect 8880 -676 8884 -644
rect 8916 -676 8920 -644
rect 8880 -724 8920 -676
rect 8880 -756 8884 -724
rect 8916 -756 8920 -724
rect 8880 -804 8920 -756
rect 8880 -836 8884 -804
rect 8916 -836 8920 -804
rect 8880 -884 8920 -836
rect 8880 -916 8884 -884
rect 8916 -916 8920 -884
rect 8880 -964 8920 -916
rect 8880 -996 8884 -964
rect 8916 -996 8920 -964
rect 8880 -1044 8920 -996
rect 8880 -1076 8884 -1044
rect 8916 -1076 8920 -1044
rect 8880 -1124 8920 -1076
rect 8880 -1156 8884 -1124
rect 8916 -1156 8920 -1124
rect 8880 -1204 8920 -1156
rect 8880 -1236 8884 -1204
rect 8916 -1236 8920 -1204
rect 8880 -1284 8920 -1236
rect 8880 -1316 8884 -1284
rect 8916 -1316 8920 -1284
rect 8880 -1364 8920 -1316
rect 8880 -1396 8884 -1364
rect 8916 -1396 8920 -1364
rect 8880 -1444 8920 -1396
rect 8880 -1476 8884 -1444
rect 8916 -1476 8920 -1444
rect 8880 -1524 8920 -1476
rect 8880 -1556 8884 -1524
rect 8916 -1556 8920 -1524
rect 8880 -1604 8920 -1556
rect 8880 -1636 8884 -1604
rect 8916 -1636 8920 -1604
rect 8880 -1684 8920 -1636
rect 8880 -1716 8884 -1684
rect 8916 -1716 8920 -1684
rect 8880 -1764 8920 -1716
rect 8880 -1796 8884 -1764
rect 8916 -1796 8920 -1764
rect 8880 -1844 8920 -1796
rect 8880 -1876 8884 -1844
rect 8916 -1876 8920 -1844
rect 8880 -1924 8920 -1876
rect 8880 -1956 8884 -1924
rect 8916 -1956 8920 -1924
rect 8880 -2004 8920 -1956
rect 8880 -2036 8884 -2004
rect 8916 -2036 8920 -2004
rect 8880 -2084 8920 -2036
rect 8880 -2116 8884 -2084
rect 8916 -2116 8920 -2084
rect 8880 -2164 8920 -2116
rect 8880 -2196 8884 -2164
rect 8916 -2196 8920 -2164
rect 8880 -2244 8920 -2196
rect 8880 -2276 8884 -2244
rect 8916 -2276 8920 -2244
rect 8880 -2324 8920 -2276
rect 8880 -2356 8884 -2324
rect 8916 -2356 8920 -2324
rect 8880 -2404 8920 -2356
rect 8880 -2436 8884 -2404
rect 8916 -2436 8920 -2404
rect 8880 -2484 8920 -2436
rect 8880 -2516 8884 -2484
rect 8916 -2516 8920 -2484
rect 8880 -2564 8920 -2516
rect 8880 -2596 8884 -2564
rect 8916 -2596 8920 -2564
rect 8880 -2644 8920 -2596
rect 8880 -2676 8884 -2644
rect 8916 -2676 8920 -2644
rect 8880 -2724 8920 -2676
rect 8880 -2756 8884 -2724
rect 8916 -2756 8920 -2724
rect 8880 -2804 8920 -2756
rect 8880 -2836 8884 -2804
rect 8916 -2836 8920 -2804
rect 8880 -2884 8920 -2836
rect 8880 -2916 8884 -2884
rect 8916 -2916 8920 -2884
rect 8880 -2964 8920 -2916
rect 8880 -2996 8884 -2964
rect 8916 -2996 8920 -2964
rect 8880 -3044 8920 -2996
rect 8880 -3076 8884 -3044
rect 8916 -3076 8920 -3044
rect 8880 -3124 8920 -3076
rect 8880 -3156 8884 -3124
rect 8916 -3156 8920 -3124
rect 8880 -3204 8920 -3156
rect 8880 -3236 8884 -3204
rect 8916 -3236 8920 -3204
rect 8880 -3284 8920 -3236
rect 8880 -3316 8884 -3284
rect 8916 -3316 8920 -3284
rect 8880 -3364 8920 -3316
rect 8880 -3396 8884 -3364
rect 8916 -3396 8920 -3364
rect 8880 -3444 8920 -3396
rect 8880 -3476 8884 -3444
rect 8916 -3476 8920 -3444
rect 8880 -3524 8920 -3476
rect 8880 -3556 8884 -3524
rect 8916 -3556 8920 -3524
rect 8880 -3604 8920 -3556
rect 8880 -3636 8884 -3604
rect 8916 -3636 8920 -3604
rect 8880 -3684 8920 -3636
rect 8880 -3716 8884 -3684
rect 8916 -3716 8920 -3684
rect 8880 -3720 8920 -3716
rect 8960 1036 9000 1040
rect 8960 1004 8964 1036
rect 8996 1004 9000 1036
rect 8960 956 9000 1004
rect 8960 924 8964 956
rect 8996 924 9000 956
rect 8960 876 9000 924
rect 8960 844 8964 876
rect 8996 844 9000 876
rect 8960 796 9000 844
rect 8960 764 8964 796
rect 8996 764 9000 796
rect 8960 716 9000 764
rect 8960 684 8964 716
rect 8996 684 9000 716
rect 8960 636 9000 684
rect 8960 604 8964 636
rect 8996 604 9000 636
rect 8960 556 9000 604
rect 8960 524 8964 556
rect 8996 524 9000 556
rect 8960 476 9000 524
rect 8960 444 8964 476
rect 8996 444 9000 476
rect 8960 396 9000 444
rect 8960 364 8964 396
rect 8996 364 9000 396
rect 8960 316 9000 364
rect 8960 284 8964 316
rect 8996 284 9000 316
rect 8960 236 9000 284
rect 8960 204 8964 236
rect 8996 204 9000 236
rect 8960 156 9000 204
rect 8960 124 8964 156
rect 8996 124 9000 156
rect 8960 76 9000 124
rect 8960 44 8964 76
rect 8996 44 9000 76
rect 8960 -4 9000 44
rect 8960 -36 8964 -4
rect 8996 -36 9000 -4
rect 8960 -84 9000 -36
rect 8960 -116 8964 -84
rect 8996 -116 9000 -84
rect 8960 -164 9000 -116
rect 8960 -196 8964 -164
rect 8996 -196 9000 -164
rect 8960 -244 9000 -196
rect 8960 -276 8964 -244
rect 8996 -276 9000 -244
rect 8960 -324 9000 -276
rect 8960 -356 8964 -324
rect 8996 -356 9000 -324
rect 8960 -404 9000 -356
rect 8960 -436 8964 -404
rect 8996 -436 9000 -404
rect 8960 -484 9000 -436
rect 8960 -516 8964 -484
rect 8996 -516 9000 -484
rect 8960 -564 9000 -516
rect 8960 -596 8964 -564
rect 8996 -596 9000 -564
rect 8960 -644 9000 -596
rect 8960 -676 8964 -644
rect 8996 -676 9000 -644
rect 8960 -724 9000 -676
rect 8960 -756 8964 -724
rect 8996 -756 9000 -724
rect 8960 -804 9000 -756
rect 8960 -836 8964 -804
rect 8996 -836 9000 -804
rect 8960 -884 9000 -836
rect 8960 -916 8964 -884
rect 8996 -916 9000 -884
rect 8960 -964 9000 -916
rect 8960 -996 8964 -964
rect 8996 -996 9000 -964
rect 8960 -1044 9000 -996
rect 8960 -1076 8964 -1044
rect 8996 -1076 9000 -1044
rect 8960 -1124 9000 -1076
rect 8960 -1156 8964 -1124
rect 8996 -1156 9000 -1124
rect 8960 -1204 9000 -1156
rect 8960 -1236 8964 -1204
rect 8996 -1236 9000 -1204
rect 8960 -1284 9000 -1236
rect 8960 -1316 8964 -1284
rect 8996 -1316 9000 -1284
rect 8960 -1364 9000 -1316
rect 8960 -1396 8964 -1364
rect 8996 -1396 9000 -1364
rect 8960 -1444 9000 -1396
rect 8960 -1476 8964 -1444
rect 8996 -1476 9000 -1444
rect 8960 -1524 9000 -1476
rect 8960 -1556 8964 -1524
rect 8996 -1556 9000 -1524
rect 8960 -1604 9000 -1556
rect 8960 -1636 8964 -1604
rect 8996 -1636 9000 -1604
rect 8960 -1684 9000 -1636
rect 8960 -1716 8964 -1684
rect 8996 -1716 9000 -1684
rect 8960 -1764 9000 -1716
rect 8960 -1796 8964 -1764
rect 8996 -1796 9000 -1764
rect 8960 -1844 9000 -1796
rect 8960 -1876 8964 -1844
rect 8996 -1876 9000 -1844
rect 8960 -1924 9000 -1876
rect 8960 -1956 8964 -1924
rect 8996 -1956 9000 -1924
rect 8960 -2004 9000 -1956
rect 8960 -2036 8964 -2004
rect 8996 -2036 9000 -2004
rect 8960 -2084 9000 -2036
rect 8960 -2116 8964 -2084
rect 8996 -2116 9000 -2084
rect 8960 -2164 9000 -2116
rect 8960 -2196 8964 -2164
rect 8996 -2196 9000 -2164
rect 8960 -2244 9000 -2196
rect 8960 -2276 8964 -2244
rect 8996 -2276 9000 -2244
rect 8960 -2324 9000 -2276
rect 8960 -2356 8964 -2324
rect 8996 -2356 9000 -2324
rect 8960 -2404 9000 -2356
rect 8960 -2436 8964 -2404
rect 8996 -2436 9000 -2404
rect 8960 -2484 9000 -2436
rect 8960 -2516 8964 -2484
rect 8996 -2516 9000 -2484
rect 8960 -2564 9000 -2516
rect 8960 -2596 8964 -2564
rect 8996 -2596 9000 -2564
rect 8960 -2644 9000 -2596
rect 8960 -2676 8964 -2644
rect 8996 -2676 9000 -2644
rect 8960 -2724 9000 -2676
rect 8960 -2756 8964 -2724
rect 8996 -2756 9000 -2724
rect 8960 -2804 9000 -2756
rect 8960 -2836 8964 -2804
rect 8996 -2836 9000 -2804
rect 8960 -2884 9000 -2836
rect 8960 -2916 8964 -2884
rect 8996 -2916 9000 -2884
rect 8960 -2964 9000 -2916
rect 8960 -2996 8964 -2964
rect 8996 -2996 9000 -2964
rect 8960 -3044 9000 -2996
rect 8960 -3076 8964 -3044
rect 8996 -3076 9000 -3044
rect 8960 -3124 9000 -3076
rect 8960 -3156 8964 -3124
rect 8996 -3156 9000 -3124
rect 8960 -3204 9000 -3156
rect 8960 -3236 8964 -3204
rect 8996 -3236 9000 -3204
rect 8960 -3284 9000 -3236
rect 8960 -3316 8964 -3284
rect 8996 -3316 9000 -3284
rect 8960 -3364 9000 -3316
rect 8960 -3396 8964 -3364
rect 8996 -3396 9000 -3364
rect 8960 -3444 9000 -3396
rect 8960 -3476 8964 -3444
rect 8996 -3476 9000 -3444
rect 8960 -3524 9000 -3476
rect 8960 -3556 8964 -3524
rect 8996 -3556 9000 -3524
rect 8960 -3604 9000 -3556
rect 8960 -3636 8964 -3604
rect 8996 -3636 9000 -3604
rect 8960 -3684 9000 -3636
rect 8960 -3716 8964 -3684
rect 8996 -3716 9000 -3684
rect 8960 -3720 9000 -3716
rect 9040 1036 9080 1040
rect 9040 1004 9044 1036
rect 9076 1004 9080 1036
rect 9040 956 9080 1004
rect 9040 924 9044 956
rect 9076 924 9080 956
rect 9040 876 9080 924
rect 9040 844 9044 876
rect 9076 844 9080 876
rect 9040 796 9080 844
rect 9040 764 9044 796
rect 9076 764 9080 796
rect 9040 716 9080 764
rect 9040 684 9044 716
rect 9076 684 9080 716
rect 9040 636 9080 684
rect 9040 604 9044 636
rect 9076 604 9080 636
rect 9040 556 9080 604
rect 9040 524 9044 556
rect 9076 524 9080 556
rect 9040 476 9080 524
rect 9040 444 9044 476
rect 9076 444 9080 476
rect 9040 396 9080 444
rect 9040 364 9044 396
rect 9076 364 9080 396
rect 9040 316 9080 364
rect 9040 284 9044 316
rect 9076 284 9080 316
rect 9040 236 9080 284
rect 9040 204 9044 236
rect 9076 204 9080 236
rect 9040 156 9080 204
rect 9040 124 9044 156
rect 9076 124 9080 156
rect 9040 76 9080 124
rect 9040 44 9044 76
rect 9076 44 9080 76
rect 9040 -4 9080 44
rect 9040 -36 9044 -4
rect 9076 -36 9080 -4
rect 9040 -84 9080 -36
rect 9040 -116 9044 -84
rect 9076 -116 9080 -84
rect 9040 -164 9080 -116
rect 9040 -196 9044 -164
rect 9076 -196 9080 -164
rect 9040 -244 9080 -196
rect 9040 -276 9044 -244
rect 9076 -276 9080 -244
rect 9040 -324 9080 -276
rect 9040 -356 9044 -324
rect 9076 -356 9080 -324
rect 9040 -404 9080 -356
rect 9040 -436 9044 -404
rect 9076 -436 9080 -404
rect 9040 -484 9080 -436
rect 9040 -516 9044 -484
rect 9076 -516 9080 -484
rect 9040 -564 9080 -516
rect 9040 -596 9044 -564
rect 9076 -596 9080 -564
rect 9040 -644 9080 -596
rect 9040 -676 9044 -644
rect 9076 -676 9080 -644
rect 9040 -724 9080 -676
rect 9040 -756 9044 -724
rect 9076 -756 9080 -724
rect 9040 -804 9080 -756
rect 9040 -836 9044 -804
rect 9076 -836 9080 -804
rect 9040 -884 9080 -836
rect 9040 -916 9044 -884
rect 9076 -916 9080 -884
rect 9040 -964 9080 -916
rect 9040 -996 9044 -964
rect 9076 -996 9080 -964
rect 9040 -1044 9080 -996
rect 9040 -1076 9044 -1044
rect 9076 -1076 9080 -1044
rect 9040 -1124 9080 -1076
rect 9040 -1156 9044 -1124
rect 9076 -1156 9080 -1124
rect 9040 -1204 9080 -1156
rect 9040 -1236 9044 -1204
rect 9076 -1236 9080 -1204
rect 9040 -1284 9080 -1236
rect 9040 -1316 9044 -1284
rect 9076 -1316 9080 -1284
rect 9040 -1364 9080 -1316
rect 9040 -1396 9044 -1364
rect 9076 -1396 9080 -1364
rect 9040 -1444 9080 -1396
rect 9040 -1476 9044 -1444
rect 9076 -1476 9080 -1444
rect 9040 -1524 9080 -1476
rect 9040 -1556 9044 -1524
rect 9076 -1556 9080 -1524
rect 9040 -1604 9080 -1556
rect 9040 -1636 9044 -1604
rect 9076 -1636 9080 -1604
rect 9040 -1684 9080 -1636
rect 9040 -1716 9044 -1684
rect 9076 -1716 9080 -1684
rect 9040 -1764 9080 -1716
rect 9040 -1796 9044 -1764
rect 9076 -1796 9080 -1764
rect 9040 -1844 9080 -1796
rect 9040 -1876 9044 -1844
rect 9076 -1876 9080 -1844
rect 9040 -1924 9080 -1876
rect 9040 -1956 9044 -1924
rect 9076 -1956 9080 -1924
rect 9040 -2004 9080 -1956
rect 9040 -2036 9044 -2004
rect 9076 -2036 9080 -2004
rect 9040 -2084 9080 -2036
rect 9040 -2116 9044 -2084
rect 9076 -2116 9080 -2084
rect 9040 -2164 9080 -2116
rect 9040 -2196 9044 -2164
rect 9076 -2196 9080 -2164
rect 9040 -2244 9080 -2196
rect 9040 -2276 9044 -2244
rect 9076 -2276 9080 -2244
rect 9040 -2324 9080 -2276
rect 9040 -2356 9044 -2324
rect 9076 -2356 9080 -2324
rect 9040 -2404 9080 -2356
rect 9040 -2436 9044 -2404
rect 9076 -2436 9080 -2404
rect 9040 -2484 9080 -2436
rect 9040 -2516 9044 -2484
rect 9076 -2516 9080 -2484
rect 9040 -2564 9080 -2516
rect 9040 -2596 9044 -2564
rect 9076 -2596 9080 -2564
rect 9040 -2644 9080 -2596
rect 9040 -2676 9044 -2644
rect 9076 -2676 9080 -2644
rect 9040 -2724 9080 -2676
rect 9040 -2756 9044 -2724
rect 9076 -2756 9080 -2724
rect 9040 -2804 9080 -2756
rect 9040 -2836 9044 -2804
rect 9076 -2836 9080 -2804
rect 9040 -2884 9080 -2836
rect 9040 -2916 9044 -2884
rect 9076 -2916 9080 -2884
rect 9040 -2964 9080 -2916
rect 9040 -2996 9044 -2964
rect 9076 -2996 9080 -2964
rect 9040 -3044 9080 -2996
rect 9040 -3076 9044 -3044
rect 9076 -3076 9080 -3044
rect 9040 -3124 9080 -3076
rect 9040 -3156 9044 -3124
rect 9076 -3156 9080 -3124
rect 9040 -3204 9080 -3156
rect 9040 -3236 9044 -3204
rect 9076 -3236 9080 -3204
rect 9040 -3284 9080 -3236
rect 9040 -3316 9044 -3284
rect 9076 -3316 9080 -3284
rect 9040 -3364 9080 -3316
rect 9040 -3396 9044 -3364
rect 9076 -3396 9080 -3364
rect 9040 -3444 9080 -3396
rect 9040 -3476 9044 -3444
rect 9076 -3476 9080 -3444
rect 9040 -3524 9080 -3476
rect 9040 -3556 9044 -3524
rect 9076 -3556 9080 -3524
rect 9040 -3604 9080 -3556
rect 9040 -3636 9044 -3604
rect 9076 -3636 9080 -3604
rect 9040 -3684 9080 -3636
rect 9040 -3716 9044 -3684
rect 9076 -3716 9080 -3684
rect 9040 -3720 9080 -3716
rect 9120 1036 9160 1040
rect 9120 1004 9124 1036
rect 9156 1004 9160 1036
rect 9120 956 9160 1004
rect 9120 924 9124 956
rect 9156 924 9160 956
rect 9120 876 9160 924
rect 9120 844 9124 876
rect 9156 844 9160 876
rect 9120 796 9160 844
rect 9120 764 9124 796
rect 9156 764 9160 796
rect 9120 716 9160 764
rect 9120 684 9124 716
rect 9156 684 9160 716
rect 9120 636 9160 684
rect 9120 604 9124 636
rect 9156 604 9160 636
rect 9120 556 9160 604
rect 9120 524 9124 556
rect 9156 524 9160 556
rect 9120 476 9160 524
rect 9120 444 9124 476
rect 9156 444 9160 476
rect 9120 396 9160 444
rect 9120 364 9124 396
rect 9156 364 9160 396
rect 9120 316 9160 364
rect 9120 284 9124 316
rect 9156 284 9160 316
rect 9120 236 9160 284
rect 9120 204 9124 236
rect 9156 204 9160 236
rect 9120 156 9160 204
rect 9120 124 9124 156
rect 9156 124 9160 156
rect 9120 76 9160 124
rect 9120 44 9124 76
rect 9156 44 9160 76
rect 9120 -4 9160 44
rect 9120 -36 9124 -4
rect 9156 -36 9160 -4
rect 9120 -84 9160 -36
rect 9120 -116 9124 -84
rect 9156 -116 9160 -84
rect 9120 -164 9160 -116
rect 9120 -196 9124 -164
rect 9156 -196 9160 -164
rect 9120 -244 9160 -196
rect 9120 -276 9124 -244
rect 9156 -276 9160 -244
rect 9120 -324 9160 -276
rect 9120 -356 9124 -324
rect 9156 -356 9160 -324
rect 9120 -404 9160 -356
rect 9120 -436 9124 -404
rect 9156 -436 9160 -404
rect 9120 -484 9160 -436
rect 9120 -516 9124 -484
rect 9156 -516 9160 -484
rect 9120 -564 9160 -516
rect 9120 -596 9124 -564
rect 9156 -596 9160 -564
rect 9120 -644 9160 -596
rect 9120 -676 9124 -644
rect 9156 -676 9160 -644
rect 9120 -724 9160 -676
rect 9120 -756 9124 -724
rect 9156 -756 9160 -724
rect 9120 -804 9160 -756
rect 9120 -836 9124 -804
rect 9156 -836 9160 -804
rect 9120 -884 9160 -836
rect 9120 -916 9124 -884
rect 9156 -916 9160 -884
rect 9120 -964 9160 -916
rect 9120 -996 9124 -964
rect 9156 -996 9160 -964
rect 9120 -1044 9160 -996
rect 9120 -1076 9124 -1044
rect 9156 -1076 9160 -1044
rect 9120 -1124 9160 -1076
rect 9120 -1156 9124 -1124
rect 9156 -1156 9160 -1124
rect 9120 -1204 9160 -1156
rect 9120 -1236 9124 -1204
rect 9156 -1236 9160 -1204
rect 9120 -1284 9160 -1236
rect 9120 -1316 9124 -1284
rect 9156 -1316 9160 -1284
rect 9120 -1364 9160 -1316
rect 9120 -1396 9124 -1364
rect 9156 -1396 9160 -1364
rect 9120 -1444 9160 -1396
rect 9120 -1476 9124 -1444
rect 9156 -1476 9160 -1444
rect 9120 -1524 9160 -1476
rect 9120 -1556 9124 -1524
rect 9156 -1556 9160 -1524
rect 9120 -1604 9160 -1556
rect 9120 -1636 9124 -1604
rect 9156 -1636 9160 -1604
rect 9120 -1684 9160 -1636
rect 9120 -1716 9124 -1684
rect 9156 -1716 9160 -1684
rect 9120 -1764 9160 -1716
rect 9120 -1796 9124 -1764
rect 9156 -1796 9160 -1764
rect 9120 -1844 9160 -1796
rect 9120 -1876 9124 -1844
rect 9156 -1876 9160 -1844
rect 9120 -1924 9160 -1876
rect 9120 -1956 9124 -1924
rect 9156 -1956 9160 -1924
rect 9120 -2004 9160 -1956
rect 9120 -2036 9124 -2004
rect 9156 -2036 9160 -2004
rect 9120 -2084 9160 -2036
rect 9120 -2116 9124 -2084
rect 9156 -2116 9160 -2084
rect 9120 -2164 9160 -2116
rect 9120 -2196 9124 -2164
rect 9156 -2196 9160 -2164
rect 9120 -2244 9160 -2196
rect 9120 -2276 9124 -2244
rect 9156 -2276 9160 -2244
rect 9120 -2324 9160 -2276
rect 9120 -2356 9124 -2324
rect 9156 -2356 9160 -2324
rect 9120 -2404 9160 -2356
rect 9120 -2436 9124 -2404
rect 9156 -2436 9160 -2404
rect 9120 -2484 9160 -2436
rect 9120 -2516 9124 -2484
rect 9156 -2516 9160 -2484
rect 9120 -2564 9160 -2516
rect 9120 -2596 9124 -2564
rect 9156 -2596 9160 -2564
rect 9120 -2644 9160 -2596
rect 9120 -2676 9124 -2644
rect 9156 -2676 9160 -2644
rect 9120 -2724 9160 -2676
rect 9120 -2756 9124 -2724
rect 9156 -2756 9160 -2724
rect 9120 -2804 9160 -2756
rect 9120 -2836 9124 -2804
rect 9156 -2836 9160 -2804
rect 9120 -2884 9160 -2836
rect 9120 -2916 9124 -2884
rect 9156 -2916 9160 -2884
rect 9120 -2964 9160 -2916
rect 9120 -2996 9124 -2964
rect 9156 -2996 9160 -2964
rect 9120 -3044 9160 -2996
rect 9120 -3076 9124 -3044
rect 9156 -3076 9160 -3044
rect 9120 -3124 9160 -3076
rect 9120 -3156 9124 -3124
rect 9156 -3156 9160 -3124
rect 9120 -3204 9160 -3156
rect 9120 -3236 9124 -3204
rect 9156 -3236 9160 -3204
rect 9120 -3284 9160 -3236
rect 9120 -3316 9124 -3284
rect 9156 -3316 9160 -3284
rect 9120 -3364 9160 -3316
rect 9120 -3396 9124 -3364
rect 9156 -3396 9160 -3364
rect 9120 -3444 9160 -3396
rect 9120 -3476 9124 -3444
rect 9156 -3476 9160 -3444
rect 9120 -3524 9160 -3476
rect 9120 -3556 9124 -3524
rect 9156 -3556 9160 -3524
rect 9120 -3604 9160 -3556
rect 9120 -3636 9124 -3604
rect 9156 -3636 9160 -3604
rect 9120 -3684 9160 -3636
rect 9120 -3716 9124 -3684
rect 9156 -3716 9160 -3684
rect 9120 -3720 9160 -3716
rect 9200 1036 9240 1040
rect 9200 1004 9204 1036
rect 9236 1004 9240 1036
rect 9200 956 9240 1004
rect 9200 924 9204 956
rect 9236 924 9240 956
rect 9200 876 9240 924
rect 9200 844 9204 876
rect 9236 844 9240 876
rect 9200 796 9240 844
rect 9200 764 9204 796
rect 9236 764 9240 796
rect 9200 716 9240 764
rect 9200 684 9204 716
rect 9236 684 9240 716
rect 9200 636 9240 684
rect 9200 604 9204 636
rect 9236 604 9240 636
rect 9200 556 9240 604
rect 9200 524 9204 556
rect 9236 524 9240 556
rect 9200 476 9240 524
rect 9200 444 9204 476
rect 9236 444 9240 476
rect 9200 396 9240 444
rect 9200 364 9204 396
rect 9236 364 9240 396
rect 9200 316 9240 364
rect 9200 284 9204 316
rect 9236 284 9240 316
rect 9200 236 9240 284
rect 9200 204 9204 236
rect 9236 204 9240 236
rect 9200 156 9240 204
rect 9200 124 9204 156
rect 9236 124 9240 156
rect 9200 76 9240 124
rect 9200 44 9204 76
rect 9236 44 9240 76
rect 9200 -4 9240 44
rect 9200 -36 9204 -4
rect 9236 -36 9240 -4
rect 9200 -84 9240 -36
rect 9200 -116 9204 -84
rect 9236 -116 9240 -84
rect 9200 -164 9240 -116
rect 9200 -196 9204 -164
rect 9236 -196 9240 -164
rect 9200 -244 9240 -196
rect 9200 -276 9204 -244
rect 9236 -276 9240 -244
rect 9200 -324 9240 -276
rect 9200 -356 9204 -324
rect 9236 -356 9240 -324
rect 9200 -404 9240 -356
rect 9200 -436 9204 -404
rect 9236 -436 9240 -404
rect 9200 -484 9240 -436
rect 9200 -516 9204 -484
rect 9236 -516 9240 -484
rect 9200 -564 9240 -516
rect 9200 -596 9204 -564
rect 9236 -596 9240 -564
rect 9200 -644 9240 -596
rect 9200 -676 9204 -644
rect 9236 -676 9240 -644
rect 9200 -724 9240 -676
rect 9200 -756 9204 -724
rect 9236 -756 9240 -724
rect 9200 -804 9240 -756
rect 9200 -836 9204 -804
rect 9236 -836 9240 -804
rect 9200 -884 9240 -836
rect 9200 -916 9204 -884
rect 9236 -916 9240 -884
rect 9200 -964 9240 -916
rect 9200 -996 9204 -964
rect 9236 -996 9240 -964
rect 9200 -1044 9240 -996
rect 9200 -1076 9204 -1044
rect 9236 -1076 9240 -1044
rect 9200 -1124 9240 -1076
rect 9200 -1156 9204 -1124
rect 9236 -1156 9240 -1124
rect 9200 -1204 9240 -1156
rect 9200 -1236 9204 -1204
rect 9236 -1236 9240 -1204
rect 9200 -1284 9240 -1236
rect 9200 -1316 9204 -1284
rect 9236 -1316 9240 -1284
rect 9200 -1364 9240 -1316
rect 9200 -1396 9204 -1364
rect 9236 -1396 9240 -1364
rect 9200 -1444 9240 -1396
rect 9200 -1476 9204 -1444
rect 9236 -1476 9240 -1444
rect 9200 -1524 9240 -1476
rect 9200 -1556 9204 -1524
rect 9236 -1556 9240 -1524
rect 9200 -1604 9240 -1556
rect 9200 -1636 9204 -1604
rect 9236 -1636 9240 -1604
rect 9200 -1684 9240 -1636
rect 9200 -1716 9204 -1684
rect 9236 -1716 9240 -1684
rect 9200 -1764 9240 -1716
rect 9200 -1796 9204 -1764
rect 9236 -1796 9240 -1764
rect 9200 -1844 9240 -1796
rect 9200 -1876 9204 -1844
rect 9236 -1876 9240 -1844
rect 9200 -1924 9240 -1876
rect 9200 -1956 9204 -1924
rect 9236 -1956 9240 -1924
rect 9200 -2004 9240 -1956
rect 9200 -2036 9204 -2004
rect 9236 -2036 9240 -2004
rect 9200 -2084 9240 -2036
rect 9200 -2116 9204 -2084
rect 9236 -2116 9240 -2084
rect 9200 -2164 9240 -2116
rect 9200 -2196 9204 -2164
rect 9236 -2196 9240 -2164
rect 9200 -2244 9240 -2196
rect 9200 -2276 9204 -2244
rect 9236 -2276 9240 -2244
rect 9200 -2324 9240 -2276
rect 9200 -2356 9204 -2324
rect 9236 -2356 9240 -2324
rect 9200 -2404 9240 -2356
rect 9200 -2436 9204 -2404
rect 9236 -2436 9240 -2404
rect 9200 -2484 9240 -2436
rect 9200 -2516 9204 -2484
rect 9236 -2516 9240 -2484
rect 9200 -2564 9240 -2516
rect 9200 -2596 9204 -2564
rect 9236 -2596 9240 -2564
rect 9200 -2644 9240 -2596
rect 9200 -2676 9204 -2644
rect 9236 -2676 9240 -2644
rect 9200 -2724 9240 -2676
rect 9200 -2756 9204 -2724
rect 9236 -2756 9240 -2724
rect 9200 -2804 9240 -2756
rect 9200 -2836 9204 -2804
rect 9236 -2836 9240 -2804
rect 9200 -2884 9240 -2836
rect 9200 -2916 9204 -2884
rect 9236 -2916 9240 -2884
rect 9200 -2964 9240 -2916
rect 9200 -2996 9204 -2964
rect 9236 -2996 9240 -2964
rect 9200 -3044 9240 -2996
rect 9200 -3076 9204 -3044
rect 9236 -3076 9240 -3044
rect 9200 -3124 9240 -3076
rect 9200 -3156 9204 -3124
rect 9236 -3156 9240 -3124
rect 9200 -3204 9240 -3156
rect 9200 -3236 9204 -3204
rect 9236 -3236 9240 -3204
rect 9200 -3284 9240 -3236
rect 9200 -3316 9204 -3284
rect 9236 -3316 9240 -3284
rect 9200 -3364 9240 -3316
rect 9200 -3396 9204 -3364
rect 9236 -3396 9240 -3364
rect 9200 -3444 9240 -3396
rect 9200 -3476 9204 -3444
rect 9236 -3476 9240 -3444
rect 9200 -3524 9240 -3476
rect 9200 -3556 9204 -3524
rect 9236 -3556 9240 -3524
rect 9200 -3604 9240 -3556
rect 9200 -3636 9204 -3604
rect 9236 -3636 9240 -3604
rect 9200 -3684 9240 -3636
rect 9200 -3716 9204 -3684
rect 9236 -3716 9240 -3684
rect 9200 -3720 9240 -3716
rect 9280 1036 9320 1040
rect 9280 1004 9284 1036
rect 9316 1004 9320 1036
rect 9280 956 9320 1004
rect 9280 924 9284 956
rect 9316 924 9320 956
rect 9280 876 9320 924
rect 9280 844 9284 876
rect 9316 844 9320 876
rect 9280 796 9320 844
rect 9280 764 9284 796
rect 9316 764 9320 796
rect 9280 716 9320 764
rect 9280 684 9284 716
rect 9316 684 9320 716
rect 9280 636 9320 684
rect 9280 604 9284 636
rect 9316 604 9320 636
rect 9280 556 9320 604
rect 9280 524 9284 556
rect 9316 524 9320 556
rect 9280 476 9320 524
rect 9280 444 9284 476
rect 9316 444 9320 476
rect 9280 396 9320 444
rect 9280 364 9284 396
rect 9316 364 9320 396
rect 9280 316 9320 364
rect 9280 284 9284 316
rect 9316 284 9320 316
rect 9280 236 9320 284
rect 9280 204 9284 236
rect 9316 204 9320 236
rect 9280 156 9320 204
rect 9280 124 9284 156
rect 9316 124 9320 156
rect 9280 76 9320 124
rect 9280 44 9284 76
rect 9316 44 9320 76
rect 9280 -4 9320 44
rect 9280 -36 9284 -4
rect 9316 -36 9320 -4
rect 9280 -84 9320 -36
rect 9280 -116 9284 -84
rect 9316 -116 9320 -84
rect 9280 -164 9320 -116
rect 9280 -196 9284 -164
rect 9316 -196 9320 -164
rect 9280 -244 9320 -196
rect 9280 -276 9284 -244
rect 9316 -276 9320 -244
rect 9280 -324 9320 -276
rect 9280 -356 9284 -324
rect 9316 -356 9320 -324
rect 9280 -404 9320 -356
rect 9280 -436 9284 -404
rect 9316 -436 9320 -404
rect 9280 -484 9320 -436
rect 9280 -516 9284 -484
rect 9316 -516 9320 -484
rect 9280 -564 9320 -516
rect 9280 -596 9284 -564
rect 9316 -596 9320 -564
rect 9280 -644 9320 -596
rect 9280 -676 9284 -644
rect 9316 -676 9320 -644
rect 9280 -724 9320 -676
rect 9280 -756 9284 -724
rect 9316 -756 9320 -724
rect 9280 -804 9320 -756
rect 9280 -836 9284 -804
rect 9316 -836 9320 -804
rect 9280 -884 9320 -836
rect 9280 -916 9284 -884
rect 9316 -916 9320 -884
rect 9280 -964 9320 -916
rect 9280 -996 9284 -964
rect 9316 -996 9320 -964
rect 9280 -1044 9320 -996
rect 9280 -1076 9284 -1044
rect 9316 -1076 9320 -1044
rect 9280 -1124 9320 -1076
rect 9280 -1156 9284 -1124
rect 9316 -1156 9320 -1124
rect 9280 -1204 9320 -1156
rect 9280 -1236 9284 -1204
rect 9316 -1236 9320 -1204
rect 9280 -1284 9320 -1236
rect 9280 -1316 9284 -1284
rect 9316 -1316 9320 -1284
rect 9280 -1364 9320 -1316
rect 9280 -1396 9284 -1364
rect 9316 -1396 9320 -1364
rect 9280 -1444 9320 -1396
rect 9280 -1476 9284 -1444
rect 9316 -1476 9320 -1444
rect 9280 -1524 9320 -1476
rect 9280 -1556 9284 -1524
rect 9316 -1556 9320 -1524
rect 9280 -1604 9320 -1556
rect 9280 -1636 9284 -1604
rect 9316 -1636 9320 -1604
rect 9280 -1684 9320 -1636
rect 9280 -1716 9284 -1684
rect 9316 -1716 9320 -1684
rect 9280 -1764 9320 -1716
rect 9280 -1796 9284 -1764
rect 9316 -1796 9320 -1764
rect 9280 -1844 9320 -1796
rect 9280 -1876 9284 -1844
rect 9316 -1876 9320 -1844
rect 9280 -1924 9320 -1876
rect 9280 -1956 9284 -1924
rect 9316 -1956 9320 -1924
rect 9280 -2004 9320 -1956
rect 9280 -2036 9284 -2004
rect 9316 -2036 9320 -2004
rect 9280 -2084 9320 -2036
rect 9280 -2116 9284 -2084
rect 9316 -2116 9320 -2084
rect 9280 -2164 9320 -2116
rect 9280 -2196 9284 -2164
rect 9316 -2196 9320 -2164
rect 9280 -2244 9320 -2196
rect 9280 -2276 9284 -2244
rect 9316 -2276 9320 -2244
rect 9280 -2324 9320 -2276
rect 9280 -2356 9284 -2324
rect 9316 -2356 9320 -2324
rect 9280 -2404 9320 -2356
rect 9280 -2436 9284 -2404
rect 9316 -2436 9320 -2404
rect 9280 -2484 9320 -2436
rect 9280 -2516 9284 -2484
rect 9316 -2516 9320 -2484
rect 9280 -2564 9320 -2516
rect 9280 -2596 9284 -2564
rect 9316 -2596 9320 -2564
rect 9280 -2644 9320 -2596
rect 9280 -2676 9284 -2644
rect 9316 -2676 9320 -2644
rect 9280 -2724 9320 -2676
rect 9280 -2756 9284 -2724
rect 9316 -2756 9320 -2724
rect 9280 -2804 9320 -2756
rect 9280 -2836 9284 -2804
rect 9316 -2836 9320 -2804
rect 9280 -2884 9320 -2836
rect 9280 -2916 9284 -2884
rect 9316 -2916 9320 -2884
rect 9280 -2964 9320 -2916
rect 9280 -2996 9284 -2964
rect 9316 -2996 9320 -2964
rect 9280 -3044 9320 -2996
rect 9280 -3076 9284 -3044
rect 9316 -3076 9320 -3044
rect 9280 -3124 9320 -3076
rect 9280 -3156 9284 -3124
rect 9316 -3156 9320 -3124
rect 9280 -3204 9320 -3156
rect 9280 -3236 9284 -3204
rect 9316 -3236 9320 -3204
rect 9280 -3284 9320 -3236
rect 9280 -3316 9284 -3284
rect 9316 -3316 9320 -3284
rect 9280 -3364 9320 -3316
rect 9280 -3396 9284 -3364
rect 9316 -3396 9320 -3364
rect 9280 -3444 9320 -3396
rect 9280 -3476 9284 -3444
rect 9316 -3476 9320 -3444
rect 9280 -3524 9320 -3476
rect 9280 -3556 9284 -3524
rect 9316 -3556 9320 -3524
rect 9280 -3604 9320 -3556
rect 9280 -3636 9284 -3604
rect 9316 -3636 9320 -3604
rect 9280 -3684 9320 -3636
rect 9280 -3716 9284 -3684
rect 9316 -3716 9320 -3684
rect 9280 -3720 9320 -3716
rect 9360 1036 9400 1040
rect 9360 1004 9364 1036
rect 9396 1004 9400 1036
rect 9360 956 9400 1004
rect 9360 924 9364 956
rect 9396 924 9400 956
rect 9360 876 9400 924
rect 9360 844 9364 876
rect 9396 844 9400 876
rect 9360 796 9400 844
rect 9360 764 9364 796
rect 9396 764 9400 796
rect 9360 716 9400 764
rect 9360 684 9364 716
rect 9396 684 9400 716
rect 9360 636 9400 684
rect 9360 604 9364 636
rect 9396 604 9400 636
rect 9360 556 9400 604
rect 9360 524 9364 556
rect 9396 524 9400 556
rect 9360 476 9400 524
rect 9360 444 9364 476
rect 9396 444 9400 476
rect 9360 396 9400 444
rect 9360 364 9364 396
rect 9396 364 9400 396
rect 9360 316 9400 364
rect 9360 284 9364 316
rect 9396 284 9400 316
rect 9360 236 9400 284
rect 9360 204 9364 236
rect 9396 204 9400 236
rect 9360 156 9400 204
rect 9360 124 9364 156
rect 9396 124 9400 156
rect 9360 76 9400 124
rect 9360 44 9364 76
rect 9396 44 9400 76
rect 9360 -4 9400 44
rect 9360 -36 9364 -4
rect 9396 -36 9400 -4
rect 9360 -84 9400 -36
rect 9360 -116 9364 -84
rect 9396 -116 9400 -84
rect 9360 -164 9400 -116
rect 9360 -196 9364 -164
rect 9396 -196 9400 -164
rect 9360 -244 9400 -196
rect 9360 -276 9364 -244
rect 9396 -276 9400 -244
rect 9360 -324 9400 -276
rect 9360 -356 9364 -324
rect 9396 -356 9400 -324
rect 9360 -404 9400 -356
rect 9360 -436 9364 -404
rect 9396 -436 9400 -404
rect 9360 -484 9400 -436
rect 9360 -516 9364 -484
rect 9396 -516 9400 -484
rect 9360 -564 9400 -516
rect 9360 -596 9364 -564
rect 9396 -596 9400 -564
rect 9360 -644 9400 -596
rect 9360 -676 9364 -644
rect 9396 -676 9400 -644
rect 9360 -724 9400 -676
rect 9360 -756 9364 -724
rect 9396 -756 9400 -724
rect 9360 -804 9400 -756
rect 9360 -836 9364 -804
rect 9396 -836 9400 -804
rect 9360 -884 9400 -836
rect 9360 -916 9364 -884
rect 9396 -916 9400 -884
rect 9360 -964 9400 -916
rect 9360 -996 9364 -964
rect 9396 -996 9400 -964
rect 9360 -1044 9400 -996
rect 9360 -1076 9364 -1044
rect 9396 -1076 9400 -1044
rect 9360 -1124 9400 -1076
rect 9360 -1156 9364 -1124
rect 9396 -1156 9400 -1124
rect 9360 -1204 9400 -1156
rect 9360 -1236 9364 -1204
rect 9396 -1236 9400 -1204
rect 9360 -1284 9400 -1236
rect 9360 -1316 9364 -1284
rect 9396 -1316 9400 -1284
rect 9360 -1364 9400 -1316
rect 9360 -1396 9364 -1364
rect 9396 -1396 9400 -1364
rect 9360 -1444 9400 -1396
rect 9360 -1476 9364 -1444
rect 9396 -1476 9400 -1444
rect 9360 -1524 9400 -1476
rect 9360 -1556 9364 -1524
rect 9396 -1556 9400 -1524
rect 9360 -1604 9400 -1556
rect 9360 -1636 9364 -1604
rect 9396 -1636 9400 -1604
rect 9360 -1684 9400 -1636
rect 9360 -1716 9364 -1684
rect 9396 -1716 9400 -1684
rect 9360 -1764 9400 -1716
rect 9360 -1796 9364 -1764
rect 9396 -1796 9400 -1764
rect 9360 -1844 9400 -1796
rect 9360 -1876 9364 -1844
rect 9396 -1876 9400 -1844
rect 9360 -1924 9400 -1876
rect 9360 -1956 9364 -1924
rect 9396 -1956 9400 -1924
rect 9360 -2004 9400 -1956
rect 9360 -2036 9364 -2004
rect 9396 -2036 9400 -2004
rect 9360 -2084 9400 -2036
rect 9360 -2116 9364 -2084
rect 9396 -2116 9400 -2084
rect 9360 -2164 9400 -2116
rect 9360 -2196 9364 -2164
rect 9396 -2196 9400 -2164
rect 9360 -2244 9400 -2196
rect 9360 -2276 9364 -2244
rect 9396 -2276 9400 -2244
rect 9360 -2324 9400 -2276
rect 9360 -2356 9364 -2324
rect 9396 -2356 9400 -2324
rect 9360 -2404 9400 -2356
rect 9360 -2436 9364 -2404
rect 9396 -2436 9400 -2404
rect 9360 -2484 9400 -2436
rect 9360 -2516 9364 -2484
rect 9396 -2516 9400 -2484
rect 9360 -2564 9400 -2516
rect 9360 -2596 9364 -2564
rect 9396 -2596 9400 -2564
rect 9360 -2644 9400 -2596
rect 9360 -2676 9364 -2644
rect 9396 -2676 9400 -2644
rect 9360 -2724 9400 -2676
rect 9360 -2756 9364 -2724
rect 9396 -2756 9400 -2724
rect 9360 -2804 9400 -2756
rect 9360 -2836 9364 -2804
rect 9396 -2836 9400 -2804
rect 9360 -2884 9400 -2836
rect 9360 -2916 9364 -2884
rect 9396 -2916 9400 -2884
rect 9360 -2964 9400 -2916
rect 9360 -2996 9364 -2964
rect 9396 -2996 9400 -2964
rect 9360 -3044 9400 -2996
rect 9360 -3076 9364 -3044
rect 9396 -3076 9400 -3044
rect 9360 -3124 9400 -3076
rect 9360 -3156 9364 -3124
rect 9396 -3156 9400 -3124
rect 9360 -3204 9400 -3156
rect 9360 -3236 9364 -3204
rect 9396 -3236 9400 -3204
rect 9360 -3284 9400 -3236
rect 9360 -3316 9364 -3284
rect 9396 -3316 9400 -3284
rect 9360 -3364 9400 -3316
rect 9360 -3396 9364 -3364
rect 9396 -3396 9400 -3364
rect 9360 -3444 9400 -3396
rect 9360 -3476 9364 -3444
rect 9396 -3476 9400 -3444
rect 9360 -3524 9400 -3476
rect 9360 -3556 9364 -3524
rect 9396 -3556 9400 -3524
rect 9360 -3604 9400 -3556
rect 9360 -3636 9364 -3604
rect 9396 -3636 9400 -3604
rect 9360 -3684 9400 -3636
rect 9360 -3716 9364 -3684
rect 9396 -3716 9400 -3684
rect 9360 -3720 9400 -3716
rect 9440 1036 9480 1040
rect 9440 1004 9444 1036
rect 9476 1004 9480 1036
rect 9440 956 9480 1004
rect 9440 924 9444 956
rect 9476 924 9480 956
rect 9440 876 9480 924
rect 9440 844 9444 876
rect 9476 844 9480 876
rect 9440 796 9480 844
rect 9440 764 9444 796
rect 9476 764 9480 796
rect 9440 716 9480 764
rect 9440 684 9444 716
rect 9476 684 9480 716
rect 9440 636 9480 684
rect 9440 604 9444 636
rect 9476 604 9480 636
rect 9440 556 9480 604
rect 9440 524 9444 556
rect 9476 524 9480 556
rect 9440 476 9480 524
rect 9440 444 9444 476
rect 9476 444 9480 476
rect 9440 396 9480 444
rect 9440 364 9444 396
rect 9476 364 9480 396
rect 9440 316 9480 364
rect 9440 284 9444 316
rect 9476 284 9480 316
rect 9440 236 9480 284
rect 9440 204 9444 236
rect 9476 204 9480 236
rect 9440 156 9480 204
rect 9440 124 9444 156
rect 9476 124 9480 156
rect 9440 76 9480 124
rect 9440 44 9444 76
rect 9476 44 9480 76
rect 9440 -4 9480 44
rect 9440 -36 9444 -4
rect 9476 -36 9480 -4
rect 9440 -84 9480 -36
rect 9440 -116 9444 -84
rect 9476 -116 9480 -84
rect 9440 -164 9480 -116
rect 9440 -196 9444 -164
rect 9476 -196 9480 -164
rect 9440 -244 9480 -196
rect 9440 -276 9444 -244
rect 9476 -276 9480 -244
rect 9440 -324 9480 -276
rect 9440 -356 9444 -324
rect 9476 -356 9480 -324
rect 9440 -404 9480 -356
rect 9440 -436 9444 -404
rect 9476 -436 9480 -404
rect 9440 -484 9480 -436
rect 9440 -516 9444 -484
rect 9476 -516 9480 -484
rect 9440 -564 9480 -516
rect 9440 -596 9444 -564
rect 9476 -596 9480 -564
rect 9440 -644 9480 -596
rect 9440 -676 9444 -644
rect 9476 -676 9480 -644
rect 9440 -724 9480 -676
rect 9440 -756 9444 -724
rect 9476 -756 9480 -724
rect 9440 -804 9480 -756
rect 9440 -836 9444 -804
rect 9476 -836 9480 -804
rect 9440 -884 9480 -836
rect 9440 -916 9444 -884
rect 9476 -916 9480 -884
rect 9440 -964 9480 -916
rect 9440 -996 9444 -964
rect 9476 -996 9480 -964
rect 9440 -1044 9480 -996
rect 9440 -1076 9444 -1044
rect 9476 -1076 9480 -1044
rect 9440 -1124 9480 -1076
rect 9440 -1156 9444 -1124
rect 9476 -1156 9480 -1124
rect 9440 -1204 9480 -1156
rect 9440 -1236 9444 -1204
rect 9476 -1236 9480 -1204
rect 9440 -1284 9480 -1236
rect 9440 -1316 9444 -1284
rect 9476 -1316 9480 -1284
rect 9440 -1364 9480 -1316
rect 9440 -1396 9444 -1364
rect 9476 -1396 9480 -1364
rect 9440 -1444 9480 -1396
rect 9440 -1476 9444 -1444
rect 9476 -1476 9480 -1444
rect 9440 -1524 9480 -1476
rect 9440 -1556 9444 -1524
rect 9476 -1556 9480 -1524
rect 9440 -1604 9480 -1556
rect 9440 -1636 9444 -1604
rect 9476 -1636 9480 -1604
rect 9440 -1684 9480 -1636
rect 9440 -1716 9444 -1684
rect 9476 -1716 9480 -1684
rect 9440 -1764 9480 -1716
rect 9440 -1796 9444 -1764
rect 9476 -1796 9480 -1764
rect 9440 -1844 9480 -1796
rect 9440 -1876 9444 -1844
rect 9476 -1876 9480 -1844
rect 9440 -1924 9480 -1876
rect 9440 -1956 9444 -1924
rect 9476 -1956 9480 -1924
rect 9440 -2004 9480 -1956
rect 9440 -2036 9444 -2004
rect 9476 -2036 9480 -2004
rect 9440 -2084 9480 -2036
rect 9440 -2116 9444 -2084
rect 9476 -2116 9480 -2084
rect 9440 -2164 9480 -2116
rect 9440 -2196 9444 -2164
rect 9476 -2196 9480 -2164
rect 9440 -2244 9480 -2196
rect 9440 -2276 9444 -2244
rect 9476 -2276 9480 -2244
rect 9440 -2324 9480 -2276
rect 9440 -2356 9444 -2324
rect 9476 -2356 9480 -2324
rect 9440 -2404 9480 -2356
rect 9440 -2436 9444 -2404
rect 9476 -2436 9480 -2404
rect 9440 -2484 9480 -2436
rect 9440 -2516 9444 -2484
rect 9476 -2516 9480 -2484
rect 9440 -2564 9480 -2516
rect 9440 -2596 9444 -2564
rect 9476 -2596 9480 -2564
rect 9440 -2644 9480 -2596
rect 9440 -2676 9444 -2644
rect 9476 -2676 9480 -2644
rect 9440 -2724 9480 -2676
rect 9440 -2756 9444 -2724
rect 9476 -2756 9480 -2724
rect 9440 -2804 9480 -2756
rect 9440 -2836 9444 -2804
rect 9476 -2836 9480 -2804
rect 9440 -2884 9480 -2836
rect 9440 -2916 9444 -2884
rect 9476 -2916 9480 -2884
rect 9440 -2964 9480 -2916
rect 9440 -2996 9444 -2964
rect 9476 -2996 9480 -2964
rect 9440 -3044 9480 -2996
rect 9440 -3076 9444 -3044
rect 9476 -3076 9480 -3044
rect 9440 -3124 9480 -3076
rect 9440 -3156 9444 -3124
rect 9476 -3156 9480 -3124
rect 9440 -3204 9480 -3156
rect 9440 -3236 9444 -3204
rect 9476 -3236 9480 -3204
rect 9440 -3284 9480 -3236
rect 9440 -3316 9444 -3284
rect 9476 -3316 9480 -3284
rect 9440 -3364 9480 -3316
rect 9440 -3396 9444 -3364
rect 9476 -3396 9480 -3364
rect 9440 -3444 9480 -3396
rect 9440 -3476 9444 -3444
rect 9476 -3476 9480 -3444
rect 9440 -3524 9480 -3476
rect 9440 -3556 9444 -3524
rect 9476 -3556 9480 -3524
rect 9440 -3604 9480 -3556
rect 9440 -3636 9444 -3604
rect 9476 -3636 9480 -3604
rect 9440 -3684 9480 -3636
rect 9440 -3716 9444 -3684
rect 9476 -3716 9480 -3684
rect 9440 -3720 9480 -3716
rect 9520 1036 9560 1040
rect 9520 1004 9524 1036
rect 9556 1004 9560 1036
rect 9520 956 9560 1004
rect 9520 924 9524 956
rect 9556 924 9560 956
rect 9520 876 9560 924
rect 9520 844 9524 876
rect 9556 844 9560 876
rect 9520 796 9560 844
rect 9520 764 9524 796
rect 9556 764 9560 796
rect 9520 716 9560 764
rect 9520 684 9524 716
rect 9556 684 9560 716
rect 9520 636 9560 684
rect 9520 604 9524 636
rect 9556 604 9560 636
rect 9520 556 9560 604
rect 9520 524 9524 556
rect 9556 524 9560 556
rect 9520 476 9560 524
rect 9520 444 9524 476
rect 9556 444 9560 476
rect 9520 396 9560 444
rect 9520 364 9524 396
rect 9556 364 9560 396
rect 9520 316 9560 364
rect 9520 284 9524 316
rect 9556 284 9560 316
rect 9520 236 9560 284
rect 9520 204 9524 236
rect 9556 204 9560 236
rect 9520 156 9560 204
rect 9520 124 9524 156
rect 9556 124 9560 156
rect 9520 76 9560 124
rect 9520 44 9524 76
rect 9556 44 9560 76
rect 9520 -4 9560 44
rect 9520 -36 9524 -4
rect 9556 -36 9560 -4
rect 9520 -84 9560 -36
rect 9520 -116 9524 -84
rect 9556 -116 9560 -84
rect 9520 -164 9560 -116
rect 9520 -196 9524 -164
rect 9556 -196 9560 -164
rect 9520 -244 9560 -196
rect 9520 -276 9524 -244
rect 9556 -276 9560 -244
rect 9520 -324 9560 -276
rect 9520 -356 9524 -324
rect 9556 -356 9560 -324
rect 9520 -404 9560 -356
rect 9520 -436 9524 -404
rect 9556 -436 9560 -404
rect 9520 -484 9560 -436
rect 9520 -516 9524 -484
rect 9556 -516 9560 -484
rect 9520 -564 9560 -516
rect 9520 -596 9524 -564
rect 9556 -596 9560 -564
rect 9520 -644 9560 -596
rect 9520 -676 9524 -644
rect 9556 -676 9560 -644
rect 9520 -724 9560 -676
rect 9520 -756 9524 -724
rect 9556 -756 9560 -724
rect 9520 -804 9560 -756
rect 9520 -836 9524 -804
rect 9556 -836 9560 -804
rect 9520 -884 9560 -836
rect 9520 -916 9524 -884
rect 9556 -916 9560 -884
rect 9520 -964 9560 -916
rect 9520 -996 9524 -964
rect 9556 -996 9560 -964
rect 9520 -1044 9560 -996
rect 9520 -1076 9524 -1044
rect 9556 -1076 9560 -1044
rect 9520 -1124 9560 -1076
rect 9520 -1156 9524 -1124
rect 9556 -1156 9560 -1124
rect 9520 -1204 9560 -1156
rect 9520 -1236 9524 -1204
rect 9556 -1236 9560 -1204
rect 9520 -1284 9560 -1236
rect 9520 -1316 9524 -1284
rect 9556 -1316 9560 -1284
rect 9520 -1364 9560 -1316
rect 9520 -1396 9524 -1364
rect 9556 -1396 9560 -1364
rect 9520 -1444 9560 -1396
rect 9520 -1476 9524 -1444
rect 9556 -1476 9560 -1444
rect 9520 -1524 9560 -1476
rect 9520 -1556 9524 -1524
rect 9556 -1556 9560 -1524
rect 9520 -1604 9560 -1556
rect 9520 -1636 9524 -1604
rect 9556 -1636 9560 -1604
rect 9520 -1684 9560 -1636
rect 9520 -1716 9524 -1684
rect 9556 -1716 9560 -1684
rect 9520 -1764 9560 -1716
rect 9520 -1796 9524 -1764
rect 9556 -1796 9560 -1764
rect 9520 -1844 9560 -1796
rect 9520 -1876 9524 -1844
rect 9556 -1876 9560 -1844
rect 9520 -1924 9560 -1876
rect 9520 -1956 9524 -1924
rect 9556 -1956 9560 -1924
rect 9520 -2004 9560 -1956
rect 9520 -2036 9524 -2004
rect 9556 -2036 9560 -2004
rect 9520 -2084 9560 -2036
rect 9520 -2116 9524 -2084
rect 9556 -2116 9560 -2084
rect 9520 -2164 9560 -2116
rect 9520 -2196 9524 -2164
rect 9556 -2196 9560 -2164
rect 9520 -2244 9560 -2196
rect 9520 -2276 9524 -2244
rect 9556 -2276 9560 -2244
rect 9520 -2324 9560 -2276
rect 9520 -2356 9524 -2324
rect 9556 -2356 9560 -2324
rect 9520 -2404 9560 -2356
rect 9520 -2436 9524 -2404
rect 9556 -2436 9560 -2404
rect 9520 -2484 9560 -2436
rect 9520 -2516 9524 -2484
rect 9556 -2516 9560 -2484
rect 9520 -2564 9560 -2516
rect 9520 -2596 9524 -2564
rect 9556 -2596 9560 -2564
rect 9520 -2644 9560 -2596
rect 9520 -2676 9524 -2644
rect 9556 -2676 9560 -2644
rect 9520 -2724 9560 -2676
rect 9520 -2756 9524 -2724
rect 9556 -2756 9560 -2724
rect 9520 -2804 9560 -2756
rect 9520 -2836 9524 -2804
rect 9556 -2836 9560 -2804
rect 9520 -2884 9560 -2836
rect 9520 -2916 9524 -2884
rect 9556 -2916 9560 -2884
rect 9520 -2964 9560 -2916
rect 9520 -2996 9524 -2964
rect 9556 -2996 9560 -2964
rect 9520 -3044 9560 -2996
rect 9520 -3076 9524 -3044
rect 9556 -3076 9560 -3044
rect 9520 -3124 9560 -3076
rect 9520 -3156 9524 -3124
rect 9556 -3156 9560 -3124
rect 9520 -3204 9560 -3156
rect 9520 -3236 9524 -3204
rect 9556 -3236 9560 -3204
rect 9520 -3284 9560 -3236
rect 9520 -3316 9524 -3284
rect 9556 -3316 9560 -3284
rect 9520 -3364 9560 -3316
rect 9520 -3396 9524 -3364
rect 9556 -3396 9560 -3364
rect 9520 -3444 9560 -3396
rect 9520 -3476 9524 -3444
rect 9556 -3476 9560 -3444
rect 9520 -3524 9560 -3476
rect 9520 -3556 9524 -3524
rect 9556 -3556 9560 -3524
rect 9520 -3604 9560 -3556
rect 9520 -3636 9524 -3604
rect 9556 -3636 9560 -3604
rect 9520 -3684 9560 -3636
rect 9520 -3716 9524 -3684
rect 9556 -3716 9560 -3684
rect 9520 -3720 9560 -3716
rect 9600 1036 9640 1040
rect 9600 1004 9604 1036
rect 9636 1004 9640 1036
rect 9600 956 9640 1004
rect 9600 924 9604 956
rect 9636 924 9640 956
rect 9600 876 9640 924
rect 9600 844 9604 876
rect 9636 844 9640 876
rect 9600 796 9640 844
rect 9600 764 9604 796
rect 9636 764 9640 796
rect 9600 716 9640 764
rect 9600 684 9604 716
rect 9636 684 9640 716
rect 9600 636 9640 684
rect 9600 604 9604 636
rect 9636 604 9640 636
rect 9600 556 9640 604
rect 9600 524 9604 556
rect 9636 524 9640 556
rect 9600 476 9640 524
rect 9600 444 9604 476
rect 9636 444 9640 476
rect 9600 396 9640 444
rect 9600 364 9604 396
rect 9636 364 9640 396
rect 9600 316 9640 364
rect 9600 284 9604 316
rect 9636 284 9640 316
rect 9600 236 9640 284
rect 9600 204 9604 236
rect 9636 204 9640 236
rect 9600 156 9640 204
rect 9600 124 9604 156
rect 9636 124 9640 156
rect 9600 76 9640 124
rect 9600 44 9604 76
rect 9636 44 9640 76
rect 9600 -4 9640 44
rect 9600 -36 9604 -4
rect 9636 -36 9640 -4
rect 9600 -84 9640 -36
rect 9600 -116 9604 -84
rect 9636 -116 9640 -84
rect 9600 -164 9640 -116
rect 9600 -196 9604 -164
rect 9636 -196 9640 -164
rect 9600 -244 9640 -196
rect 9600 -276 9604 -244
rect 9636 -276 9640 -244
rect 9600 -324 9640 -276
rect 9600 -356 9604 -324
rect 9636 -356 9640 -324
rect 9600 -404 9640 -356
rect 9600 -436 9604 -404
rect 9636 -436 9640 -404
rect 9600 -484 9640 -436
rect 9600 -516 9604 -484
rect 9636 -516 9640 -484
rect 9600 -564 9640 -516
rect 9600 -596 9604 -564
rect 9636 -596 9640 -564
rect 9600 -644 9640 -596
rect 9600 -676 9604 -644
rect 9636 -676 9640 -644
rect 9600 -724 9640 -676
rect 9600 -756 9604 -724
rect 9636 -756 9640 -724
rect 9600 -804 9640 -756
rect 9600 -836 9604 -804
rect 9636 -836 9640 -804
rect 9600 -884 9640 -836
rect 9600 -916 9604 -884
rect 9636 -916 9640 -884
rect 9600 -964 9640 -916
rect 9600 -996 9604 -964
rect 9636 -996 9640 -964
rect 9600 -1044 9640 -996
rect 9600 -1076 9604 -1044
rect 9636 -1076 9640 -1044
rect 9600 -1124 9640 -1076
rect 9600 -1156 9604 -1124
rect 9636 -1156 9640 -1124
rect 9600 -1204 9640 -1156
rect 9600 -1236 9604 -1204
rect 9636 -1236 9640 -1204
rect 9600 -1284 9640 -1236
rect 9600 -1316 9604 -1284
rect 9636 -1316 9640 -1284
rect 9600 -1364 9640 -1316
rect 9600 -1396 9604 -1364
rect 9636 -1396 9640 -1364
rect 9600 -1444 9640 -1396
rect 9600 -1476 9604 -1444
rect 9636 -1476 9640 -1444
rect 9600 -1524 9640 -1476
rect 9600 -1556 9604 -1524
rect 9636 -1556 9640 -1524
rect 9600 -1604 9640 -1556
rect 9600 -1636 9604 -1604
rect 9636 -1636 9640 -1604
rect 9600 -1684 9640 -1636
rect 9600 -1716 9604 -1684
rect 9636 -1716 9640 -1684
rect 9600 -1764 9640 -1716
rect 9600 -1796 9604 -1764
rect 9636 -1796 9640 -1764
rect 9600 -1844 9640 -1796
rect 9600 -1876 9604 -1844
rect 9636 -1876 9640 -1844
rect 9600 -1924 9640 -1876
rect 9600 -1956 9604 -1924
rect 9636 -1956 9640 -1924
rect 9600 -2004 9640 -1956
rect 9600 -2036 9604 -2004
rect 9636 -2036 9640 -2004
rect 9600 -2084 9640 -2036
rect 9600 -2116 9604 -2084
rect 9636 -2116 9640 -2084
rect 9600 -2164 9640 -2116
rect 9600 -2196 9604 -2164
rect 9636 -2196 9640 -2164
rect 9600 -2244 9640 -2196
rect 9600 -2276 9604 -2244
rect 9636 -2276 9640 -2244
rect 9600 -2324 9640 -2276
rect 9600 -2356 9604 -2324
rect 9636 -2356 9640 -2324
rect 9600 -2404 9640 -2356
rect 9600 -2436 9604 -2404
rect 9636 -2436 9640 -2404
rect 9600 -2484 9640 -2436
rect 9600 -2516 9604 -2484
rect 9636 -2516 9640 -2484
rect 9600 -2564 9640 -2516
rect 9600 -2596 9604 -2564
rect 9636 -2596 9640 -2564
rect 9600 -2644 9640 -2596
rect 9600 -2676 9604 -2644
rect 9636 -2676 9640 -2644
rect 9600 -2724 9640 -2676
rect 9600 -2756 9604 -2724
rect 9636 -2756 9640 -2724
rect 9600 -2804 9640 -2756
rect 9600 -2836 9604 -2804
rect 9636 -2836 9640 -2804
rect 9600 -2884 9640 -2836
rect 9600 -2916 9604 -2884
rect 9636 -2916 9640 -2884
rect 9600 -2964 9640 -2916
rect 9600 -2996 9604 -2964
rect 9636 -2996 9640 -2964
rect 9600 -3044 9640 -2996
rect 9600 -3076 9604 -3044
rect 9636 -3076 9640 -3044
rect 9600 -3124 9640 -3076
rect 9600 -3156 9604 -3124
rect 9636 -3156 9640 -3124
rect 9600 -3204 9640 -3156
rect 9600 -3236 9604 -3204
rect 9636 -3236 9640 -3204
rect 9600 -3284 9640 -3236
rect 9600 -3316 9604 -3284
rect 9636 -3316 9640 -3284
rect 9600 -3364 9640 -3316
rect 9600 -3396 9604 -3364
rect 9636 -3396 9640 -3364
rect 9600 -3444 9640 -3396
rect 9600 -3476 9604 -3444
rect 9636 -3476 9640 -3444
rect 9600 -3524 9640 -3476
rect 9600 -3556 9604 -3524
rect 9636 -3556 9640 -3524
rect 9600 -3604 9640 -3556
rect 9600 -3636 9604 -3604
rect 9636 -3636 9640 -3604
rect 9600 -3684 9640 -3636
rect 9600 -3716 9604 -3684
rect 9636 -3716 9640 -3684
rect 9600 -3720 9640 -3716
rect 9680 1036 9720 1040
rect 9680 1004 9684 1036
rect 9716 1004 9720 1036
rect 9680 956 9720 1004
rect 9680 924 9684 956
rect 9716 924 9720 956
rect 9680 876 9720 924
rect 9680 844 9684 876
rect 9716 844 9720 876
rect 9680 796 9720 844
rect 9680 764 9684 796
rect 9716 764 9720 796
rect 9680 716 9720 764
rect 9680 684 9684 716
rect 9716 684 9720 716
rect 9680 636 9720 684
rect 9680 604 9684 636
rect 9716 604 9720 636
rect 9680 556 9720 604
rect 9680 524 9684 556
rect 9716 524 9720 556
rect 9680 476 9720 524
rect 9680 444 9684 476
rect 9716 444 9720 476
rect 9680 396 9720 444
rect 9680 364 9684 396
rect 9716 364 9720 396
rect 9680 316 9720 364
rect 9680 284 9684 316
rect 9716 284 9720 316
rect 9680 236 9720 284
rect 9680 204 9684 236
rect 9716 204 9720 236
rect 9680 156 9720 204
rect 9680 124 9684 156
rect 9716 124 9720 156
rect 9680 76 9720 124
rect 9680 44 9684 76
rect 9716 44 9720 76
rect 9680 -4 9720 44
rect 9680 -36 9684 -4
rect 9716 -36 9720 -4
rect 9680 -84 9720 -36
rect 9680 -116 9684 -84
rect 9716 -116 9720 -84
rect 9680 -164 9720 -116
rect 9680 -196 9684 -164
rect 9716 -196 9720 -164
rect 9680 -244 9720 -196
rect 9680 -276 9684 -244
rect 9716 -276 9720 -244
rect 9680 -324 9720 -276
rect 9680 -356 9684 -324
rect 9716 -356 9720 -324
rect 9680 -404 9720 -356
rect 9680 -436 9684 -404
rect 9716 -436 9720 -404
rect 9680 -484 9720 -436
rect 9680 -516 9684 -484
rect 9716 -516 9720 -484
rect 9680 -564 9720 -516
rect 9680 -596 9684 -564
rect 9716 -596 9720 -564
rect 9680 -644 9720 -596
rect 9680 -676 9684 -644
rect 9716 -676 9720 -644
rect 9680 -724 9720 -676
rect 9680 -756 9684 -724
rect 9716 -756 9720 -724
rect 9680 -804 9720 -756
rect 9680 -836 9684 -804
rect 9716 -836 9720 -804
rect 9680 -884 9720 -836
rect 9680 -916 9684 -884
rect 9716 -916 9720 -884
rect 9680 -964 9720 -916
rect 9680 -996 9684 -964
rect 9716 -996 9720 -964
rect 9680 -1044 9720 -996
rect 9680 -1076 9684 -1044
rect 9716 -1076 9720 -1044
rect 9680 -1124 9720 -1076
rect 9680 -1156 9684 -1124
rect 9716 -1156 9720 -1124
rect 9680 -1204 9720 -1156
rect 9680 -1236 9684 -1204
rect 9716 -1236 9720 -1204
rect 9680 -1284 9720 -1236
rect 9680 -1316 9684 -1284
rect 9716 -1316 9720 -1284
rect 9680 -1364 9720 -1316
rect 9680 -1396 9684 -1364
rect 9716 -1396 9720 -1364
rect 9680 -1444 9720 -1396
rect 9680 -1476 9684 -1444
rect 9716 -1476 9720 -1444
rect 9680 -1524 9720 -1476
rect 9680 -1556 9684 -1524
rect 9716 -1556 9720 -1524
rect 9680 -1604 9720 -1556
rect 9680 -1636 9684 -1604
rect 9716 -1636 9720 -1604
rect 9680 -1684 9720 -1636
rect 9680 -1716 9684 -1684
rect 9716 -1716 9720 -1684
rect 9680 -1764 9720 -1716
rect 9680 -1796 9684 -1764
rect 9716 -1796 9720 -1764
rect 9680 -1844 9720 -1796
rect 9680 -1876 9684 -1844
rect 9716 -1876 9720 -1844
rect 9680 -1924 9720 -1876
rect 9680 -1956 9684 -1924
rect 9716 -1956 9720 -1924
rect 9680 -2004 9720 -1956
rect 9680 -2036 9684 -2004
rect 9716 -2036 9720 -2004
rect 9680 -2084 9720 -2036
rect 9680 -2116 9684 -2084
rect 9716 -2116 9720 -2084
rect 9680 -2164 9720 -2116
rect 9680 -2196 9684 -2164
rect 9716 -2196 9720 -2164
rect 9680 -2244 9720 -2196
rect 9680 -2276 9684 -2244
rect 9716 -2276 9720 -2244
rect 9680 -2324 9720 -2276
rect 9680 -2356 9684 -2324
rect 9716 -2356 9720 -2324
rect 9680 -2404 9720 -2356
rect 9680 -2436 9684 -2404
rect 9716 -2436 9720 -2404
rect 9680 -2484 9720 -2436
rect 9680 -2516 9684 -2484
rect 9716 -2516 9720 -2484
rect 9680 -2564 9720 -2516
rect 9680 -2596 9684 -2564
rect 9716 -2596 9720 -2564
rect 9680 -2644 9720 -2596
rect 9680 -2676 9684 -2644
rect 9716 -2676 9720 -2644
rect 9680 -2724 9720 -2676
rect 9680 -2756 9684 -2724
rect 9716 -2756 9720 -2724
rect 9680 -2804 9720 -2756
rect 9680 -2836 9684 -2804
rect 9716 -2836 9720 -2804
rect 9680 -2884 9720 -2836
rect 9680 -2916 9684 -2884
rect 9716 -2916 9720 -2884
rect 9680 -2964 9720 -2916
rect 9680 -2996 9684 -2964
rect 9716 -2996 9720 -2964
rect 9680 -3044 9720 -2996
rect 9680 -3076 9684 -3044
rect 9716 -3076 9720 -3044
rect 9680 -3124 9720 -3076
rect 9680 -3156 9684 -3124
rect 9716 -3156 9720 -3124
rect 9680 -3204 9720 -3156
rect 9680 -3236 9684 -3204
rect 9716 -3236 9720 -3204
rect 9680 -3284 9720 -3236
rect 9680 -3316 9684 -3284
rect 9716 -3316 9720 -3284
rect 9680 -3364 9720 -3316
rect 9680 -3396 9684 -3364
rect 9716 -3396 9720 -3364
rect 9680 -3444 9720 -3396
rect 9680 -3476 9684 -3444
rect 9716 -3476 9720 -3444
rect 9680 -3524 9720 -3476
rect 9680 -3556 9684 -3524
rect 9716 -3556 9720 -3524
rect 9680 -3604 9720 -3556
rect 9680 -3636 9684 -3604
rect 9716 -3636 9720 -3604
rect 9680 -3684 9720 -3636
rect 9680 -3716 9684 -3684
rect 9716 -3716 9720 -3684
rect 9680 -3720 9720 -3716
rect 9760 1036 9800 1040
rect 9760 1004 9764 1036
rect 9796 1004 9800 1036
rect 9760 956 9800 1004
rect 9760 924 9764 956
rect 9796 924 9800 956
rect 9760 876 9800 924
rect 9760 844 9764 876
rect 9796 844 9800 876
rect 9760 796 9800 844
rect 9760 764 9764 796
rect 9796 764 9800 796
rect 9760 716 9800 764
rect 9760 684 9764 716
rect 9796 684 9800 716
rect 9760 636 9800 684
rect 9760 604 9764 636
rect 9796 604 9800 636
rect 9760 556 9800 604
rect 9760 524 9764 556
rect 9796 524 9800 556
rect 9760 476 9800 524
rect 9760 444 9764 476
rect 9796 444 9800 476
rect 9760 396 9800 444
rect 9760 364 9764 396
rect 9796 364 9800 396
rect 9760 316 9800 364
rect 9760 284 9764 316
rect 9796 284 9800 316
rect 9760 236 9800 284
rect 9760 204 9764 236
rect 9796 204 9800 236
rect 9760 156 9800 204
rect 9760 124 9764 156
rect 9796 124 9800 156
rect 9760 76 9800 124
rect 9760 44 9764 76
rect 9796 44 9800 76
rect 9760 -4 9800 44
rect 9760 -36 9764 -4
rect 9796 -36 9800 -4
rect 9760 -84 9800 -36
rect 9760 -116 9764 -84
rect 9796 -116 9800 -84
rect 9760 -164 9800 -116
rect 9760 -196 9764 -164
rect 9796 -196 9800 -164
rect 9760 -244 9800 -196
rect 9760 -276 9764 -244
rect 9796 -276 9800 -244
rect 9760 -324 9800 -276
rect 9760 -356 9764 -324
rect 9796 -356 9800 -324
rect 9760 -404 9800 -356
rect 9760 -436 9764 -404
rect 9796 -436 9800 -404
rect 9760 -484 9800 -436
rect 9760 -516 9764 -484
rect 9796 -516 9800 -484
rect 9760 -564 9800 -516
rect 9760 -596 9764 -564
rect 9796 -596 9800 -564
rect 9760 -644 9800 -596
rect 9760 -676 9764 -644
rect 9796 -676 9800 -644
rect 9760 -724 9800 -676
rect 9760 -756 9764 -724
rect 9796 -756 9800 -724
rect 9760 -804 9800 -756
rect 9760 -836 9764 -804
rect 9796 -836 9800 -804
rect 9760 -884 9800 -836
rect 9760 -916 9764 -884
rect 9796 -916 9800 -884
rect 9760 -964 9800 -916
rect 9760 -996 9764 -964
rect 9796 -996 9800 -964
rect 9760 -1044 9800 -996
rect 9760 -1076 9764 -1044
rect 9796 -1076 9800 -1044
rect 9760 -1124 9800 -1076
rect 9760 -1156 9764 -1124
rect 9796 -1156 9800 -1124
rect 9760 -1204 9800 -1156
rect 9760 -1236 9764 -1204
rect 9796 -1236 9800 -1204
rect 9760 -1284 9800 -1236
rect 9760 -1316 9764 -1284
rect 9796 -1316 9800 -1284
rect 9760 -1364 9800 -1316
rect 9760 -1396 9764 -1364
rect 9796 -1396 9800 -1364
rect 9760 -1444 9800 -1396
rect 9760 -1476 9764 -1444
rect 9796 -1476 9800 -1444
rect 9760 -1524 9800 -1476
rect 9760 -1556 9764 -1524
rect 9796 -1556 9800 -1524
rect 9760 -1604 9800 -1556
rect 9760 -1636 9764 -1604
rect 9796 -1636 9800 -1604
rect 9760 -1684 9800 -1636
rect 9760 -1716 9764 -1684
rect 9796 -1716 9800 -1684
rect 9760 -1764 9800 -1716
rect 9760 -1796 9764 -1764
rect 9796 -1796 9800 -1764
rect 9760 -1844 9800 -1796
rect 9760 -1876 9764 -1844
rect 9796 -1876 9800 -1844
rect 9760 -1924 9800 -1876
rect 9760 -1956 9764 -1924
rect 9796 -1956 9800 -1924
rect 9760 -2004 9800 -1956
rect 9760 -2036 9764 -2004
rect 9796 -2036 9800 -2004
rect 9760 -2084 9800 -2036
rect 9760 -2116 9764 -2084
rect 9796 -2116 9800 -2084
rect 9760 -2164 9800 -2116
rect 9760 -2196 9764 -2164
rect 9796 -2196 9800 -2164
rect 9760 -2244 9800 -2196
rect 9760 -2276 9764 -2244
rect 9796 -2276 9800 -2244
rect 9760 -2324 9800 -2276
rect 9760 -2356 9764 -2324
rect 9796 -2356 9800 -2324
rect 9760 -2404 9800 -2356
rect 9760 -2436 9764 -2404
rect 9796 -2436 9800 -2404
rect 9760 -2484 9800 -2436
rect 9760 -2516 9764 -2484
rect 9796 -2516 9800 -2484
rect 9760 -2564 9800 -2516
rect 9760 -2596 9764 -2564
rect 9796 -2596 9800 -2564
rect 9760 -2644 9800 -2596
rect 9760 -2676 9764 -2644
rect 9796 -2676 9800 -2644
rect 9760 -2724 9800 -2676
rect 9760 -2756 9764 -2724
rect 9796 -2756 9800 -2724
rect 9760 -2804 9800 -2756
rect 9760 -2836 9764 -2804
rect 9796 -2836 9800 -2804
rect 9760 -2884 9800 -2836
rect 9760 -2916 9764 -2884
rect 9796 -2916 9800 -2884
rect 9760 -2964 9800 -2916
rect 9760 -2996 9764 -2964
rect 9796 -2996 9800 -2964
rect 9760 -3044 9800 -2996
rect 9760 -3076 9764 -3044
rect 9796 -3076 9800 -3044
rect 9760 -3124 9800 -3076
rect 9760 -3156 9764 -3124
rect 9796 -3156 9800 -3124
rect 9760 -3204 9800 -3156
rect 9760 -3236 9764 -3204
rect 9796 -3236 9800 -3204
rect 9760 -3284 9800 -3236
rect 9760 -3316 9764 -3284
rect 9796 -3316 9800 -3284
rect 9760 -3364 9800 -3316
rect 9760 -3396 9764 -3364
rect 9796 -3396 9800 -3364
rect 9760 -3444 9800 -3396
rect 9760 -3476 9764 -3444
rect 9796 -3476 9800 -3444
rect 9760 -3524 9800 -3476
rect 9760 -3556 9764 -3524
rect 9796 -3556 9800 -3524
rect 9760 -3604 9800 -3556
rect 9760 -3636 9764 -3604
rect 9796 -3636 9800 -3604
rect 9760 -3684 9800 -3636
rect 9760 -3716 9764 -3684
rect 9796 -3716 9800 -3684
rect 9760 -3720 9800 -3716
rect 9840 1036 9880 1040
rect 9840 1004 9844 1036
rect 9876 1004 9880 1036
rect 9840 956 9880 1004
rect 9840 924 9844 956
rect 9876 924 9880 956
rect 9840 876 9880 924
rect 9840 844 9844 876
rect 9876 844 9880 876
rect 9840 796 9880 844
rect 9840 764 9844 796
rect 9876 764 9880 796
rect 9840 716 9880 764
rect 9840 684 9844 716
rect 9876 684 9880 716
rect 9840 636 9880 684
rect 9840 604 9844 636
rect 9876 604 9880 636
rect 9840 556 9880 604
rect 9840 524 9844 556
rect 9876 524 9880 556
rect 9840 476 9880 524
rect 9840 444 9844 476
rect 9876 444 9880 476
rect 9840 396 9880 444
rect 9840 364 9844 396
rect 9876 364 9880 396
rect 9840 316 9880 364
rect 9840 284 9844 316
rect 9876 284 9880 316
rect 9840 236 9880 284
rect 9840 204 9844 236
rect 9876 204 9880 236
rect 9840 156 9880 204
rect 9840 124 9844 156
rect 9876 124 9880 156
rect 9840 76 9880 124
rect 9840 44 9844 76
rect 9876 44 9880 76
rect 9840 -4 9880 44
rect 9840 -36 9844 -4
rect 9876 -36 9880 -4
rect 9840 -84 9880 -36
rect 9840 -116 9844 -84
rect 9876 -116 9880 -84
rect 9840 -164 9880 -116
rect 9840 -196 9844 -164
rect 9876 -196 9880 -164
rect 9840 -244 9880 -196
rect 9840 -276 9844 -244
rect 9876 -276 9880 -244
rect 9840 -324 9880 -276
rect 9840 -356 9844 -324
rect 9876 -356 9880 -324
rect 9840 -404 9880 -356
rect 9840 -436 9844 -404
rect 9876 -436 9880 -404
rect 9840 -484 9880 -436
rect 9840 -516 9844 -484
rect 9876 -516 9880 -484
rect 9840 -564 9880 -516
rect 9840 -596 9844 -564
rect 9876 -596 9880 -564
rect 9840 -644 9880 -596
rect 9840 -676 9844 -644
rect 9876 -676 9880 -644
rect 9840 -724 9880 -676
rect 9840 -756 9844 -724
rect 9876 -756 9880 -724
rect 9840 -804 9880 -756
rect 9840 -836 9844 -804
rect 9876 -836 9880 -804
rect 9840 -884 9880 -836
rect 9840 -916 9844 -884
rect 9876 -916 9880 -884
rect 9840 -964 9880 -916
rect 9840 -996 9844 -964
rect 9876 -996 9880 -964
rect 9840 -1044 9880 -996
rect 9840 -1076 9844 -1044
rect 9876 -1076 9880 -1044
rect 9840 -1124 9880 -1076
rect 9840 -1156 9844 -1124
rect 9876 -1156 9880 -1124
rect 9840 -1204 9880 -1156
rect 9840 -1236 9844 -1204
rect 9876 -1236 9880 -1204
rect 9840 -1284 9880 -1236
rect 9840 -1316 9844 -1284
rect 9876 -1316 9880 -1284
rect 9840 -1364 9880 -1316
rect 9840 -1396 9844 -1364
rect 9876 -1396 9880 -1364
rect 9840 -1444 9880 -1396
rect 9840 -1476 9844 -1444
rect 9876 -1476 9880 -1444
rect 9840 -1524 9880 -1476
rect 9840 -1556 9844 -1524
rect 9876 -1556 9880 -1524
rect 9840 -1604 9880 -1556
rect 9840 -1636 9844 -1604
rect 9876 -1636 9880 -1604
rect 9840 -1684 9880 -1636
rect 9840 -1716 9844 -1684
rect 9876 -1716 9880 -1684
rect 9840 -1764 9880 -1716
rect 9840 -1796 9844 -1764
rect 9876 -1796 9880 -1764
rect 9840 -1844 9880 -1796
rect 9840 -1876 9844 -1844
rect 9876 -1876 9880 -1844
rect 9840 -1924 9880 -1876
rect 9840 -1956 9844 -1924
rect 9876 -1956 9880 -1924
rect 9840 -2004 9880 -1956
rect 9840 -2036 9844 -2004
rect 9876 -2036 9880 -2004
rect 9840 -2084 9880 -2036
rect 9840 -2116 9844 -2084
rect 9876 -2116 9880 -2084
rect 9840 -2164 9880 -2116
rect 9840 -2196 9844 -2164
rect 9876 -2196 9880 -2164
rect 9840 -2244 9880 -2196
rect 9840 -2276 9844 -2244
rect 9876 -2276 9880 -2244
rect 9840 -2324 9880 -2276
rect 9840 -2356 9844 -2324
rect 9876 -2356 9880 -2324
rect 9840 -2404 9880 -2356
rect 9840 -2436 9844 -2404
rect 9876 -2436 9880 -2404
rect 9840 -2484 9880 -2436
rect 9840 -2516 9844 -2484
rect 9876 -2516 9880 -2484
rect 9840 -2564 9880 -2516
rect 9840 -2596 9844 -2564
rect 9876 -2596 9880 -2564
rect 9840 -2644 9880 -2596
rect 9840 -2676 9844 -2644
rect 9876 -2676 9880 -2644
rect 9840 -2724 9880 -2676
rect 9840 -2756 9844 -2724
rect 9876 -2756 9880 -2724
rect 9840 -2804 9880 -2756
rect 9840 -2836 9844 -2804
rect 9876 -2836 9880 -2804
rect 9840 -2884 9880 -2836
rect 9840 -2916 9844 -2884
rect 9876 -2916 9880 -2884
rect 9840 -2964 9880 -2916
rect 9840 -2996 9844 -2964
rect 9876 -2996 9880 -2964
rect 9840 -3044 9880 -2996
rect 9840 -3076 9844 -3044
rect 9876 -3076 9880 -3044
rect 9840 -3124 9880 -3076
rect 9840 -3156 9844 -3124
rect 9876 -3156 9880 -3124
rect 9840 -3204 9880 -3156
rect 9840 -3236 9844 -3204
rect 9876 -3236 9880 -3204
rect 9840 -3284 9880 -3236
rect 9840 -3316 9844 -3284
rect 9876 -3316 9880 -3284
rect 9840 -3364 9880 -3316
rect 9840 -3396 9844 -3364
rect 9876 -3396 9880 -3364
rect 9840 -3444 9880 -3396
rect 9840 -3476 9844 -3444
rect 9876 -3476 9880 -3444
rect 9840 -3524 9880 -3476
rect 9840 -3556 9844 -3524
rect 9876 -3556 9880 -3524
rect 9840 -3604 9880 -3556
rect 9840 -3636 9844 -3604
rect 9876 -3636 9880 -3604
rect 9840 -3684 9880 -3636
rect 9840 -3716 9844 -3684
rect 9876 -3716 9880 -3684
rect 9840 -3720 9880 -3716
rect 9920 1036 9960 1040
rect 9920 1004 9924 1036
rect 9956 1004 9960 1036
rect 9920 956 9960 1004
rect 9920 924 9924 956
rect 9956 924 9960 956
rect 9920 876 9960 924
rect 9920 844 9924 876
rect 9956 844 9960 876
rect 9920 796 9960 844
rect 9920 764 9924 796
rect 9956 764 9960 796
rect 9920 716 9960 764
rect 9920 684 9924 716
rect 9956 684 9960 716
rect 9920 636 9960 684
rect 9920 604 9924 636
rect 9956 604 9960 636
rect 9920 556 9960 604
rect 9920 524 9924 556
rect 9956 524 9960 556
rect 9920 476 9960 524
rect 9920 444 9924 476
rect 9956 444 9960 476
rect 9920 396 9960 444
rect 9920 364 9924 396
rect 9956 364 9960 396
rect 9920 316 9960 364
rect 9920 284 9924 316
rect 9956 284 9960 316
rect 9920 236 9960 284
rect 9920 204 9924 236
rect 9956 204 9960 236
rect 9920 156 9960 204
rect 9920 124 9924 156
rect 9956 124 9960 156
rect 9920 76 9960 124
rect 9920 44 9924 76
rect 9956 44 9960 76
rect 9920 -4 9960 44
rect 9920 -36 9924 -4
rect 9956 -36 9960 -4
rect 9920 -84 9960 -36
rect 9920 -116 9924 -84
rect 9956 -116 9960 -84
rect 9920 -164 9960 -116
rect 9920 -196 9924 -164
rect 9956 -196 9960 -164
rect 9920 -244 9960 -196
rect 9920 -276 9924 -244
rect 9956 -276 9960 -244
rect 9920 -324 9960 -276
rect 9920 -356 9924 -324
rect 9956 -356 9960 -324
rect 9920 -404 9960 -356
rect 9920 -436 9924 -404
rect 9956 -436 9960 -404
rect 9920 -484 9960 -436
rect 9920 -516 9924 -484
rect 9956 -516 9960 -484
rect 9920 -564 9960 -516
rect 9920 -596 9924 -564
rect 9956 -596 9960 -564
rect 9920 -644 9960 -596
rect 9920 -676 9924 -644
rect 9956 -676 9960 -644
rect 9920 -724 9960 -676
rect 9920 -756 9924 -724
rect 9956 -756 9960 -724
rect 9920 -804 9960 -756
rect 9920 -836 9924 -804
rect 9956 -836 9960 -804
rect 9920 -884 9960 -836
rect 9920 -916 9924 -884
rect 9956 -916 9960 -884
rect 9920 -964 9960 -916
rect 9920 -996 9924 -964
rect 9956 -996 9960 -964
rect 9920 -1044 9960 -996
rect 9920 -1076 9924 -1044
rect 9956 -1076 9960 -1044
rect 9920 -1124 9960 -1076
rect 9920 -1156 9924 -1124
rect 9956 -1156 9960 -1124
rect 9920 -1204 9960 -1156
rect 9920 -1236 9924 -1204
rect 9956 -1236 9960 -1204
rect 9920 -1284 9960 -1236
rect 9920 -1316 9924 -1284
rect 9956 -1316 9960 -1284
rect 9920 -1364 9960 -1316
rect 9920 -1396 9924 -1364
rect 9956 -1396 9960 -1364
rect 9920 -1444 9960 -1396
rect 9920 -1476 9924 -1444
rect 9956 -1476 9960 -1444
rect 9920 -1524 9960 -1476
rect 9920 -1556 9924 -1524
rect 9956 -1556 9960 -1524
rect 9920 -1604 9960 -1556
rect 9920 -1636 9924 -1604
rect 9956 -1636 9960 -1604
rect 9920 -1684 9960 -1636
rect 9920 -1716 9924 -1684
rect 9956 -1716 9960 -1684
rect 9920 -1764 9960 -1716
rect 9920 -1796 9924 -1764
rect 9956 -1796 9960 -1764
rect 9920 -1844 9960 -1796
rect 9920 -1876 9924 -1844
rect 9956 -1876 9960 -1844
rect 9920 -1924 9960 -1876
rect 9920 -1956 9924 -1924
rect 9956 -1956 9960 -1924
rect 9920 -2004 9960 -1956
rect 9920 -2036 9924 -2004
rect 9956 -2036 9960 -2004
rect 9920 -2084 9960 -2036
rect 9920 -2116 9924 -2084
rect 9956 -2116 9960 -2084
rect 9920 -2164 9960 -2116
rect 9920 -2196 9924 -2164
rect 9956 -2196 9960 -2164
rect 9920 -2244 9960 -2196
rect 9920 -2276 9924 -2244
rect 9956 -2276 9960 -2244
rect 9920 -2324 9960 -2276
rect 9920 -2356 9924 -2324
rect 9956 -2356 9960 -2324
rect 9920 -2404 9960 -2356
rect 9920 -2436 9924 -2404
rect 9956 -2436 9960 -2404
rect 9920 -2484 9960 -2436
rect 9920 -2516 9924 -2484
rect 9956 -2516 9960 -2484
rect 9920 -2564 9960 -2516
rect 9920 -2596 9924 -2564
rect 9956 -2596 9960 -2564
rect 9920 -2644 9960 -2596
rect 9920 -2676 9924 -2644
rect 9956 -2676 9960 -2644
rect 9920 -2724 9960 -2676
rect 9920 -2756 9924 -2724
rect 9956 -2756 9960 -2724
rect 9920 -2804 9960 -2756
rect 9920 -2836 9924 -2804
rect 9956 -2836 9960 -2804
rect 9920 -2884 9960 -2836
rect 9920 -2916 9924 -2884
rect 9956 -2916 9960 -2884
rect 9920 -2964 9960 -2916
rect 9920 -2996 9924 -2964
rect 9956 -2996 9960 -2964
rect 9920 -3044 9960 -2996
rect 9920 -3076 9924 -3044
rect 9956 -3076 9960 -3044
rect 9920 -3124 9960 -3076
rect 9920 -3156 9924 -3124
rect 9956 -3156 9960 -3124
rect 9920 -3204 9960 -3156
rect 9920 -3236 9924 -3204
rect 9956 -3236 9960 -3204
rect 9920 -3284 9960 -3236
rect 9920 -3316 9924 -3284
rect 9956 -3316 9960 -3284
rect 9920 -3364 9960 -3316
rect 9920 -3396 9924 -3364
rect 9956 -3396 9960 -3364
rect 9920 -3444 9960 -3396
rect 9920 -3476 9924 -3444
rect 9956 -3476 9960 -3444
rect 9920 -3524 9960 -3476
rect 9920 -3556 9924 -3524
rect 9956 -3556 9960 -3524
rect 9920 -3604 9960 -3556
rect 9920 -3636 9924 -3604
rect 9956 -3636 9960 -3604
rect 9920 -3684 9960 -3636
rect 9920 -3716 9924 -3684
rect 9956 -3716 9960 -3684
rect 9920 -3720 9960 -3716
rect 10000 1036 10040 1040
rect 10000 1004 10004 1036
rect 10036 1004 10040 1036
rect 10000 956 10040 1004
rect 10000 924 10004 956
rect 10036 924 10040 956
rect 10000 876 10040 924
rect 10000 844 10004 876
rect 10036 844 10040 876
rect 10000 796 10040 844
rect 10000 764 10004 796
rect 10036 764 10040 796
rect 10000 716 10040 764
rect 10000 684 10004 716
rect 10036 684 10040 716
rect 10000 636 10040 684
rect 10000 604 10004 636
rect 10036 604 10040 636
rect 10000 556 10040 604
rect 10000 524 10004 556
rect 10036 524 10040 556
rect 10000 476 10040 524
rect 10000 444 10004 476
rect 10036 444 10040 476
rect 10000 396 10040 444
rect 10000 364 10004 396
rect 10036 364 10040 396
rect 10000 316 10040 364
rect 10000 284 10004 316
rect 10036 284 10040 316
rect 10000 236 10040 284
rect 10000 204 10004 236
rect 10036 204 10040 236
rect 10000 156 10040 204
rect 10000 124 10004 156
rect 10036 124 10040 156
rect 10000 76 10040 124
rect 10000 44 10004 76
rect 10036 44 10040 76
rect 10000 -4 10040 44
rect 10000 -36 10004 -4
rect 10036 -36 10040 -4
rect 10000 -84 10040 -36
rect 10000 -116 10004 -84
rect 10036 -116 10040 -84
rect 10000 -164 10040 -116
rect 10000 -196 10004 -164
rect 10036 -196 10040 -164
rect 10000 -244 10040 -196
rect 10000 -276 10004 -244
rect 10036 -276 10040 -244
rect 10000 -324 10040 -276
rect 10000 -356 10004 -324
rect 10036 -356 10040 -324
rect 10000 -404 10040 -356
rect 10000 -436 10004 -404
rect 10036 -436 10040 -404
rect 10000 -484 10040 -436
rect 10000 -516 10004 -484
rect 10036 -516 10040 -484
rect 10000 -564 10040 -516
rect 10000 -596 10004 -564
rect 10036 -596 10040 -564
rect 10000 -644 10040 -596
rect 10000 -676 10004 -644
rect 10036 -676 10040 -644
rect 10000 -724 10040 -676
rect 10000 -756 10004 -724
rect 10036 -756 10040 -724
rect 10000 -804 10040 -756
rect 10000 -836 10004 -804
rect 10036 -836 10040 -804
rect 10000 -884 10040 -836
rect 10000 -916 10004 -884
rect 10036 -916 10040 -884
rect 10000 -964 10040 -916
rect 10000 -996 10004 -964
rect 10036 -996 10040 -964
rect 10000 -1044 10040 -996
rect 10000 -1076 10004 -1044
rect 10036 -1076 10040 -1044
rect 10000 -1124 10040 -1076
rect 10000 -1156 10004 -1124
rect 10036 -1156 10040 -1124
rect 10000 -1204 10040 -1156
rect 10000 -1236 10004 -1204
rect 10036 -1236 10040 -1204
rect 10000 -1284 10040 -1236
rect 10000 -1316 10004 -1284
rect 10036 -1316 10040 -1284
rect 10000 -1364 10040 -1316
rect 10000 -1396 10004 -1364
rect 10036 -1396 10040 -1364
rect 10000 -1444 10040 -1396
rect 10000 -1476 10004 -1444
rect 10036 -1476 10040 -1444
rect 10000 -1524 10040 -1476
rect 10000 -1556 10004 -1524
rect 10036 -1556 10040 -1524
rect 10000 -1604 10040 -1556
rect 10000 -1636 10004 -1604
rect 10036 -1636 10040 -1604
rect 10000 -1684 10040 -1636
rect 10000 -1716 10004 -1684
rect 10036 -1716 10040 -1684
rect 10000 -1764 10040 -1716
rect 10000 -1796 10004 -1764
rect 10036 -1796 10040 -1764
rect 10000 -1844 10040 -1796
rect 10000 -1876 10004 -1844
rect 10036 -1876 10040 -1844
rect 10000 -1924 10040 -1876
rect 10000 -1956 10004 -1924
rect 10036 -1956 10040 -1924
rect 10000 -2004 10040 -1956
rect 10000 -2036 10004 -2004
rect 10036 -2036 10040 -2004
rect 10000 -2084 10040 -2036
rect 10000 -2116 10004 -2084
rect 10036 -2116 10040 -2084
rect 10000 -2164 10040 -2116
rect 10000 -2196 10004 -2164
rect 10036 -2196 10040 -2164
rect 10000 -2244 10040 -2196
rect 10000 -2276 10004 -2244
rect 10036 -2276 10040 -2244
rect 10000 -2324 10040 -2276
rect 10000 -2356 10004 -2324
rect 10036 -2356 10040 -2324
rect 10000 -2404 10040 -2356
rect 10000 -2436 10004 -2404
rect 10036 -2436 10040 -2404
rect 10000 -2484 10040 -2436
rect 10000 -2516 10004 -2484
rect 10036 -2516 10040 -2484
rect 10000 -2564 10040 -2516
rect 10000 -2596 10004 -2564
rect 10036 -2596 10040 -2564
rect 10000 -2644 10040 -2596
rect 10000 -2676 10004 -2644
rect 10036 -2676 10040 -2644
rect 10000 -2724 10040 -2676
rect 10000 -2756 10004 -2724
rect 10036 -2756 10040 -2724
rect 10000 -2804 10040 -2756
rect 10000 -2836 10004 -2804
rect 10036 -2836 10040 -2804
rect 10000 -2884 10040 -2836
rect 10000 -2916 10004 -2884
rect 10036 -2916 10040 -2884
rect 10000 -2964 10040 -2916
rect 10000 -2996 10004 -2964
rect 10036 -2996 10040 -2964
rect 10000 -3044 10040 -2996
rect 10000 -3076 10004 -3044
rect 10036 -3076 10040 -3044
rect 10000 -3124 10040 -3076
rect 10000 -3156 10004 -3124
rect 10036 -3156 10040 -3124
rect 10000 -3204 10040 -3156
rect 10000 -3236 10004 -3204
rect 10036 -3236 10040 -3204
rect 10000 -3284 10040 -3236
rect 10000 -3316 10004 -3284
rect 10036 -3316 10040 -3284
rect 10000 -3364 10040 -3316
rect 10000 -3396 10004 -3364
rect 10036 -3396 10040 -3364
rect 10000 -3444 10040 -3396
rect 10000 -3476 10004 -3444
rect 10036 -3476 10040 -3444
rect 10000 -3524 10040 -3476
rect 10000 -3556 10004 -3524
rect 10036 -3556 10040 -3524
rect 10000 -3604 10040 -3556
rect 10000 -3636 10004 -3604
rect 10036 -3636 10040 -3604
rect 10000 -3684 10040 -3636
rect 10000 -3716 10004 -3684
rect 10036 -3716 10040 -3684
rect 10000 -3720 10040 -3716
rect 10080 1036 10120 1040
rect 10080 1004 10084 1036
rect 10116 1004 10120 1036
rect 10080 956 10120 1004
rect 10080 924 10084 956
rect 10116 924 10120 956
rect 10080 876 10120 924
rect 10080 844 10084 876
rect 10116 844 10120 876
rect 10080 796 10120 844
rect 10080 764 10084 796
rect 10116 764 10120 796
rect 10080 716 10120 764
rect 10080 684 10084 716
rect 10116 684 10120 716
rect 10080 636 10120 684
rect 10080 604 10084 636
rect 10116 604 10120 636
rect 10080 556 10120 604
rect 10080 524 10084 556
rect 10116 524 10120 556
rect 10080 476 10120 524
rect 10080 444 10084 476
rect 10116 444 10120 476
rect 10080 396 10120 444
rect 10080 364 10084 396
rect 10116 364 10120 396
rect 10080 316 10120 364
rect 10080 284 10084 316
rect 10116 284 10120 316
rect 10080 236 10120 284
rect 10080 204 10084 236
rect 10116 204 10120 236
rect 10080 156 10120 204
rect 10080 124 10084 156
rect 10116 124 10120 156
rect 10080 76 10120 124
rect 10080 44 10084 76
rect 10116 44 10120 76
rect 10080 -4 10120 44
rect 10080 -36 10084 -4
rect 10116 -36 10120 -4
rect 10080 -84 10120 -36
rect 10080 -116 10084 -84
rect 10116 -116 10120 -84
rect 10080 -164 10120 -116
rect 10080 -196 10084 -164
rect 10116 -196 10120 -164
rect 10080 -244 10120 -196
rect 10080 -276 10084 -244
rect 10116 -276 10120 -244
rect 10080 -324 10120 -276
rect 10080 -356 10084 -324
rect 10116 -356 10120 -324
rect 10080 -404 10120 -356
rect 10080 -436 10084 -404
rect 10116 -436 10120 -404
rect 10080 -484 10120 -436
rect 10080 -516 10084 -484
rect 10116 -516 10120 -484
rect 10080 -564 10120 -516
rect 10080 -596 10084 -564
rect 10116 -596 10120 -564
rect 10080 -644 10120 -596
rect 10080 -676 10084 -644
rect 10116 -676 10120 -644
rect 10080 -724 10120 -676
rect 10080 -756 10084 -724
rect 10116 -756 10120 -724
rect 10080 -804 10120 -756
rect 10080 -836 10084 -804
rect 10116 -836 10120 -804
rect 10080 -884 10120 -836
rect 10080 -916 10084 -884
rect 10116 -916 10120 -884
rect 10080 -964 10120 -916
rect 10080 -996 10084 -964
rect 10116 -996 10120 -964
rect 10080 -1044 10120 -996
rect 10080 -1076 10084 -1044
rect 10116 -1076 10120 -1044
rect 10080 -1124 10120 -1076
rect 10080 -1156 10084 -1124
rect 10116 -1156 10120 -1124
rect 10080 -1204 10120 -1156
rect 10080 -1236 10084 -1204
rect 10116 -1236 10120 -1204
rect 10080 -1284 10120 -1236
rect 10080 -1316 10084 -1284
rect 10116 -1316 10120 -1284
rect 10080 -1364 10120 -1316
rect 10080 -1396 10084 -1364
rect 10116 -1396 10120 -1364
rect 10080 -1444 10120 -1396
rect 10080 -1476 10084 -1444
rect 10116 -1476 10120 -1444
rect 10080 -1524 10120 -1476
rect 10080 -1556 10084 -1524
rect 10116 -1556 10120 -1524
rect 10080 -1604 10120 -1556
rect 10080 -1636 10084 -1604
rect 10116 -1636 10120 -1604
rect 10080 -1684 10120 -1636
rect 10080 -1716 10084 -1684
rect 10116 -1716 10120 -1684
rect 10080 -1764 10120 -1716
rect 10080 -1796 10084 -1764
rect 10116 -1796 10120 -1764
rect 10080 -1844 10120 -1796
rect 10080 -1876 10084 -1844
rect 10116 -1876 10120 -1844
rect 10080 -1924 10120 -1876
rect 10080 -1956 10084 -1924
rect 10116 -1956 10120 -1924
rect 10080 -2004 10120 -1956
rect 10080 -2036 10084 -2004
rect 10116 -2036 10120 -2004
rect 10080 -2084 10120 -2036
rect 10080 -2116 10084 -2084
rect 10116 -2116 10120 -2084
rect 10080 -2164 10120 -2116
rect 10080 -2196 10084 -2164
rect 10116 -2196 10120 -2164
rect 10080 -2244 10120 -2196
rect 10080 -2276 10084 -2244
rect 10116 -2276 10120 -2244
rect 10080 -2324 10120 -2276
rect 10080 -2356 10084 -2324
rect 10116 -2356 10120 -2324
rect 10080 -2404 10120 -2356
rect 10080 -2436 10084 -2404
rect 10116 -2436 10120 -2404
rect 10080 -2484 10120 -2436
rect 10080 -2516 10084 -2484
rect 10116 -2516 10120 -2484
rect 10080 -2564 10120 -2516
rect 10080 -2596 10084 -2564
rect 10116 -2596 10120 -2564
rect 10080 -2644 10120 -2596
rect 10080 -2676 10084 -2644
rect 10116 -2676 10120 -2644
rect 10080 -2724 10120 -2676
rect 10080 -2756 10084 -2724
rect 10116 -2756 10120 -2724
rect 10080 -2804 10120 -2756
rect 10080 -2836 10084 -2804
rect 10116 -2836 10120 -2804
rect 10080 -2884 10120 -2836
rect 10080 -2916 10084 -2884
rect 10116 -2916 10120 -2884
rect 10080 -2964 10120 -2916
rect 10080 -2996 10084 -2964
rect 10116 -2996 10120 -2964
rect 10080 -3044 10120 -2996
rect 10080 -3076 10084 -3044
rect 10116 -3076 10120 -3044
rect 10080 -3124 10120 -3076
rect 10080 -3156 10084 -3124
rect 10116 -3156 10120 -3124
rect 10080 -3204 10120 -3156
rect 10080 -3236 10084 -3204
rect 10116 -3236 10120 -3204
rect 10080 -3284 10120 -3236
rect 10080 -3316 10084 -3284
rect 10116 -3316 10120 -3284
rect 10080 -3364 10120 -3316
rect 10080 -3396 10084 -3364
rect 10116 -3396 10120 -3364
rect 10080 -3444 10120 -3396
rect 10080 -3476 10084 -3444
rect 10116 -3476 10120 -3444
rect 10080 -3524 10120 -3476
rect 10080 -3556 10084 -3524
rect 10116 -3556 10120 -3524
rect 10080 -3604 10120 -3556
rect 10080 -3636 10084 -3604
rect 10116 -3636 10120 -3604
rect 10080 -3684 10120 -3636
rect 10080 -3716 10084 -3684
rect 10116 -3716 10120 -3684
rect 10080 -3720 10120 -3716
rect 10160 1036 10200 1040
rect 10160 1004 10164 1036
rect 10196 1004 10200 1036
rect 10160 956 10200 1004
rect 10160 924 10164 956
rect 10196 924 10200 956
rect 10160 876 10200 924
rect 10160 844 10164 876
rect 10196 844 10200 876
rect 10160 796 10200 844
rect 10160 764 10164 796
rect 10196 764 10200 796
rect 10160 716 10200 764
rect 10160 684 10164 716
rect 10196 684 10200 716
rect 10160 636 10200 684
rect 10160 604 10164 636
rect 10196 604 10200 636
rect 10160 556 10200 604
rect 10160 524 10164 556
rect 10196 524 10200 556
rect 10160 476 10200 524
rect 10160 444 10164 476
rect 10196 444 10200 476
rect 10160 396 10200 444
rect 10160 364 10164 396
rect 10196 364 10200 396
rect 10160 316 10200 364
rect 10160 284 10164 316
rect 10196 284 10200 316
rect 10160 236 10200 284
rect 10160 204 10164 236
rect 10196 204 10200 236
rect 10160 156 10200 204
rect 10160 124 10164 156
rect 10196 124 10200 156
rect 10160 76 10200 124
rect 10160 44 10164 76
rect 10196 44 10200 76
rect 10160 -4 10200 44
rect 10160 -36 10164 -4
rect 10196 -36 10200 -4
rect 10160 -84 10200 -36
rect 10160 -116 10164 -84
rect 10196 -116 10200 -84
rect 10160 -164 10200 -116
rect 10160 -196 10164 -164
rect 10196 -196 10200 -164
rect 10160 -244 10200 -196
rect 10160 -276 10164 -244
rect 10196 -276 10200 -244
rect 10160 -324 10200 -276
rect 10160 -356 10164 -324
rect 10196 -356 10200 -324
rect 10160 -404 10200 -356
rect 10160 -436 10164 -404
rect 10196 -436 10200 -404
rect 10160 -484 10200 -436
rect 10160 -516 10164 -484
rect 10196 -516 10200 -484
rect 10160 -564 10200 -516
rect 10160 -596 10164 -564
rect 10196 -596 10200 -564
rect 10160 -644 10200 -596
rect 10160 -676 10164 -644
rect 10196 -676 10200 -644
rect 10160 -724 10200 -676
rect 10160 -756 10164 -724
rect 10196 -756 10200 -724
rect 10160 -804 10200 -756
rect 10160 -836 10164 -804
rect 10196 -836 10200 -804
rect 10160 -884 10200 -836
rect 10160 -916 10164 -884
rect 10196 -916 10200 -884
rect 10160 -964 10200 -916
rect 10160 -996 10164 -964
rect 10196 -996 10200 -964
rect 10160 -1044 10200 -996
rect 10160 -1076 10164 -1044
rect 10196 -1076 10200 -1044
rect 10160 -1124 10200 -1076
rect 10160 -1156 10164 -1124
rect 10196 -1156 10200 -1124
rect 10160 -1204 10200 -1156
rect 10160 -1236 10164 -1204
rect 10196 -1236 10200 -1204
rect 10160 -1284 10200 -1236
rect 10160 -1316 10164 -1284
rect 10196 -1316 10200 -1284
rect 10160 -1364 10200 -1316
rect 10160 -1396 10164 -1364
rect 10196 -1396 10200 -1364
rect 10160 -1444 10200 -1396
rect 10160 -1476 10164 -1444
rect 10196 -1476 10200 -1444
rect 10160 -1524 10200 -1476
rect 10160 -1556 10164 -1524
rect 10196 -1556 10200 -1524
rect 10160 -1604 10200 -1556
rect 10160 -1636 10164 -1604
rect 10196 -1636 10200 -1604
rect 10160 -1684 10200 -1636
rect 10160 -1716 10164 -1684
rect 10196 -1716 10200 -1684
rect 10160 -1764 10200 -1716
rect 10160 -1796 10164 -1764
rect 10196 -1796 10200 -1764
rect 10160 -1844 10200 -1796
rect 10160 -1876 10164 -1844
rect 10196 -1876 10200 -1844
rect 10160 -1924 10200 -1876
rect 10160 -1956 10164 -1924
rect 10196 -1956 10200 -1924
rect 10160 -2004 10200 -1956
rect 10160 -2036 10164 -2004
rect 10196 -2036 10200 -2004
rect 10160 -2084 10200 -2036
rect 10160 -2116 10164 -2084
rect 10196 -2116 10200 -2084
rect 10160 -2164 10200 -2116
rect 10160 -2196 10164 -2164
rect 10196 -2196 10200 -2164
rect 10160 -2244 10200 -2196
rect 10160 -2276 10164 -2244
rect 10196 -2276 10200 -2244
rect 10160 -2324 10200 -2276
rect 10160 -2356 10164 -2324
rect 10196 -2356 10200 -2324
rect 10160 -2404 10200 -2356
rect 10160 -2436 10164 -2404
rect 10196 -2436 10200 -2404
rect 10160 -2484 10200 -2436
rect 10160 -2516 10164 -2484
rect 10196 -2516 10200 -2484
rect 10160 -2564 10200 -2516
rect 10160 -2596 10164 -2564
rect 10196 -2596 10200 -2564
rect 10160 -2644 10200 -2596
rect 10160 -2676 10164 -2644
rect 10196 -2676 10200 -2644
rect 10160 -2724 10200 -2676
rect 10160 -2756 10164 -2724
rect 10196 -2756 10200 -2724
rect 10160 -2804 10200 -2756
rect 10160 -2836 10164 -2804
rect 10196 -2836 10200 -2804
rect 10160 -2884 10200 -2836
rect 10160 -2916 10164 -2884
rect 10196 -2916 10200 -2884
rect 10160 -2964 10200 -2916
rect 10160 -2996 10164 -2964
rect 10196 -2996 10200 -2964
rect 10160 -3044 10200 -2996
rect 10160 -3076 10164 -3044
rect 10196 -3076 10200 -3044
rect 10160 -3124 10200 -3076
rect 10160 -3156 10164 -3124
rect 10196 -3156 10200 -3124
rect 10160 -3204 10200 -3156
rect 10160 -3236 10164 -3204
rect 10196 -3236 10200 -3204
rect 10160 -3284 10200 -3236
rect 10160 -3316 10164 -3284
rect 10196 -3316 10200 -3284
rect 10160 -3364 10200 -3316
rect 10160 -3396 10164 -3364
rect 10196 -3396 10200 -3364
rect 10160 -3444 10200 -3396
rect 10160 -3476 10164 -3444
rect 10196 -3476 10200 -3444
rect 10160 -3524 10200 -3476
rect 10160 -3556 10164 -3524
rect 10196 -3556 10200 -3524
rect 10160 -3604 10200 -3556
rect 10160 -3636 10164 -3604
rect 10196 -3636 10200 -3604
rect 10160 -3684 10200 -3636
rect 10160 -3716 10164 -3684
rect 10196 -3716 10200 -3684
rect 10160 -3720 10200 -3716
rect 10240 1036 10280 1040
rect 10240 1004 10244 1036
rect 10276 1004 10280 1036
rect 10240 956 10280 1004
rect 10240 924 10244 956
rect 10276 924 10280 956
rect 10240 876 10280 924
rect 10240 844 10244 876
rect 10276 844 10280 876
rect 10240 796 10280 844
rect 10240 764 10244 796
rect 10276 764 10280 796
rect 10240 716 10280 764
rect 10240 684 10244 716
rect 10276 684 10280 716
rect 10240 636 10280 684
rect 10240 604 10244 636
rect 10276 604 10280 636
rect 10240 556 10280 604
rect 10240 524 10244 556
rect 10276 524 10280 556
rect 10240 476 10280 524
rect 10240 444 10244 476
rect 10276 444 10280 476
rect 10240 396 10280 444
rect 10240 364 10244 396
rect 10276 364 10280 396
rect 10240 316 10280 364
rect 10240 284 10244 316
rect 10276 284 10280 316
rect 10240 236 10280 284
rect 10240 204 10244 236
rect 10276 204 10280 236
rect 10240 156 10280 204
rect 10240 124 10244 156
rect 10276 124 10280 156
rect 10240 76 10280 124
rect 10240 44 10244 76
rect 10276 44 10280 76
rect 10240 -4 10280 44
rect 10240 -36 10244 -4
rect 10276 -36 10280 -4
rect 10240 -84 10280 -36
rect 10240 -116 10244 -84
rect 10276 -116 10280 -84
rect 10240 -164 10280 -116
rect 10240 -196 10244 -164
rect 10276 -196 10280 -164
rect 10240 -244 10280 -196
rect 10240 -276 10244 -244
rect 10276 -276 10280 -244
rect 10240 -324 10280 -276
rect 10240 -356 10244 -324
rect 10276 -356 10280 -324
rect 10240 -404 10280 -356
rect 10240 -436 10244 -404
rect 10276 -436 10280 -404
rect 10240 -484 10280 -436
rect 10240 -516 10244 -484
rect 10276 -516 10280 -484
rect 10240 -564 10280 -516
rect 10240 -596 10244 -564
rect 10276 -596 10280 -564
rect 10240 -644 10280 -596
rect 10240 -676 10244 -644
rect 10276 -676 10280 -644
rect 10240 -724 10280 -676
rect 10240 -756 10244 -724
rect 10276 -756 10280 -724
rect 10240 -804 10280 -756
rect 10240 -836 10244 -804
rect 10276 -836 10280 -804
rect 10240 -884 10280 -836
rect 10240 -916 10244 -884
rect 10276 -916 10280 -884
rect 10240 -964 10280 -916
rect 10240 -996 10244 -964
rect 10276 -996 10280 -964
rect 10240 -1044 10280 -996
rect 10240 -1076 10244 -1044
rect 10276 -1076 10280 -1044
rect 10240 -1124 10280 -1076
rect 10240 -1156 10244 -1124
rect 10276 -1156 10280 -1124
rect 10240 -1204 10280 -1156
rect 10240 -1236 10244 -1204
rect 10276 -1236 10280 -1204
rect 10240 -1284 10280 -1236
rect 10240 -1316 10244 -1284
rect 10276 -1316 10280 -1284
rect 10240 -1364 10280 -1316
rect 10240 -1396 10244 -1364
rect 10276 -1396 10280 -1364
rect 10240 -1444 10280 -1396
rect 10240 -1476 10244 -1444
rect 10276 -1476 10280 -1444
rect 10240 -1524 10280 -1476
rect 10240 -1556 10244 -1524
rect 10276 -1556 10280 -1524
rect 10240 -1604 10280 -1556
rect 10240 -1636 10244 -1604
rect 10276 -1636 10280 -1604
rect 10240 -1684 10280 -1636
rect 10240 -1716 10244 -1684
rect 10276 -1716 10280 -1684
rect 10240 -1764 10280 -1716
rect 10240 -1796 10244 -1764
rect 10276 -1796 10280 -1764
rect 10240 -1844 10280 -1796
rect 10240 -1876 10244 -1844
rect 10276 -1876 10280 -1844
rect 10240 -1924 10280 -1876
rect 10240 -1956 10244 -1924
rect 10276 -1956 10280 -1924
rect 10240 -2004 10280 -1956
rect 10240 -2036 10244 -2004
rect 10276 -2036 10280 -2004
rect 10240 -2084 10280 -2036
rect 10240 -2116 10244 -2084
rect 10276 -2116 10280 -2084
rect 10240 -2164 10280 -2116
rect 10240 -2196 10244 -2164
rect 10276 -2196 10280 -2164
rect 10240 -2244 10280 -2196
rect 10240 -2276 10244 -2244
rect 10276 -2276 10280 -2244
rect 10240 -2324 10280 -2276
rect 10240 -2356 10244 -2324
rect 10276 -2356 10280 -2324
rect 10240 -2404 10280 -2356
rect 10240 -2436 10244 -2404
rect 10276 -2436 10280 -2404
rect 10240 -2484 10280 -2436
rect 10240 -2516 10244 -2484
rect 10276 -2516 10280 -2484
rect 10240 -2564 10280 -2516
rect 10240 -2596 10244 -2564
rect 10276 -2596 10280 -2564
rect 10240 -2644 10280 -2596
rect 10240 -2676 10244 -2644
rect 10276 -2676 10280 -2644
rect 10240 -2724 10280 -2676
rect 10240 -2756 10244 -2724
rect 10276 -2756 10280 -2724
rect 10240 -2804 10280 -2756
rect 10240 -2836 10244 -2804
rect 10276 -2836 10280 -2804
rect 10240 -2884 10280 -2836
rect 10240 -2916 10244 -2884
rect 10276 -2916 10280 -2884
rect 10240 -2964 10280 -2916
rect 10240 -2996 10244 -2964
rect 10276 -2996 10280 -2964
rect 10240 -3044 10280 -2996
rect 10240 -3076 10244 -3044
rect 10276 -3076 10280 -3044
rect 10240 -3124 10280 -3076
rect 10240 -3156 10244 -3124
rect 10276 -3156 10280 -3124
rect 10240 -3204 10280 -3156
rect 10240 -3236 10244 -3204
rect 10276 -3236 10280 -3204
rect 10240 -3284 10280 -3236
rect 10240 -3316 10244 -3284
rect 10276 -3316 10280 -3284
rect 10240 -3364 10280 -3316
rect 10240 -3396 10244 -3364
rect 10276 -3396 10280 -3364
rect 10240 -3444 10280 -3396
rect 10240 -3476 10244 -3444
rect 10276 -3476 10280 -3444
rect 10240 -3524 10280 -3476
rect 10240 -3556 10244 -3524
rect 10276 -3556 10280 -3524
rect 10240 -3604 10280 -3556
rect 10240 -3636 10244 -3604
rect 10276 -3636 10280 -3604
rect 10240 -3684 10280 -3636
rect 10240 -3716 10244 -3684
rect 10276 -3716 10280 -3684
rect 10240 -3720 10280 -3716
rect 10320 1036 10360 1040
rect 10320 1004 10324 1036
rect 10356 1004 10360 1036
rect 10320 956 10360 1004
rect 10320 924 10324 956
rect 10356 924 10360 956
rect 10320 876 10360 924
rect 10320 844 10324 876
rect 10356 844 10360 876
rect 10320 796 10360 844
rect 10320 764 10324 796
rect 10356 764 10360 796
rect 10320 716 10360 764
rect 10320 684 10324 716
rect 10356 684 10360 716
rect 10320 636 10360 684
rect 10320 604 10324 636
rect 10356 604 10360 636
rect 10320 556 10360 604
rect 10320 524 10324 556
rect 10356 524 10360 556
rect 10320 476 10360 524
rect 10320 444 10324 476
rect 10356 444 10360 476
rect 10320 396 10360 444
rect 10320 364 10324 396
rect 10356 364 10360 396
rect 10320 316 10360 364
rect 10320 284 10324 316
rect 10356 284 10360 316
rect 10320 236 10360 284
rect 10320 204 10324 236
rect 10356 204 10360 236
rect 10320 156 10360 204
rect 10320 124 10324 156
rect 10356 124 10360 156
rect 10320 76 10360 124
rect 10320 44 10324 76
rect 10356 44 10360 76
rect 10320 -4 10360 44
rect 10320 -36 10324 -4
rect 10356 -36 10360 -4
rect 10320 -84 10360 -36
rect 10320 -116 10324 -84
rect 10356 -116 10360 -84
rect 10320 -164 10360 -116
rect 10320 -196 10324 -164
rect 10356 -196 10360 -164
rect 10320 -244 10360 -196
rect 10320 -276 10324 -244
rect 10356 -276 10360 -244
rect 10320 -324 10360 -276
rect 10320 -356 10324 -324
rect 10356 -356 10360 -324
rect 10320 -404 10360 -356
rect 10320 -436 10324 -404
rect 10356 -436 10360 -404
rect 10320 -484 10360 -436
rect 10320 -516 10324 -484
rect 10356 -516 10360 -484
rect 10320 -564 10360 -516
rect 10320 -596 10324 -564
rect 10356 -596 10360 -564
rect 10320 -644 10360 -596
rect 10320 -676 10324 -644
rect 10356 -676 10360 -644
rect 10320 -724 10360 -676
rect 10320 -756 10324 -724
rect 10356 -756 10360 -724
rect 10320 -804 10360 -756
rect 10320 -836 10324 -804
rect 10356 -836 10360 -804
rect 10320 -884 10360 -836
rect 10320 -916 10324 -884
rect 10356 -916 10360 -884
rect 10320 -964 10360 -916
rect 10320 -996 10324 -964
rect 10356 -996 10360 -964
rect 10320 -1044 10360 -996
rect 10320 -1076 10324 -1044
rect 10356 -1076 10360 -1044
rect 10320 -1124 10360 -1076
rect 10320 -1156 10324 -1124
rect 10356 -1156 10360 -1124
rect 10320 -1204 10360 -1156
rect 10320 -1236 10324 -1204
rect 10356 -1236 10360 -1204
rect 10320 -1284 10360 -1236
rect 10320 -1316 10324 -1284
rect 10356 -1316 10360 -1284
rect 10320 -1364 10360 -1316
rect 10320 -1396 10324 -1364
rect 10356 -1396 10360 -1364
rect 10320 -1444 10360 -1396
rect 10320 -1476 10324 -1444
rect 10356 -1476 10360 -1444
rect 10320 -1524 10360 -1476
rect 10320 -1556 10324 -1524
rect 10356 -1556 10360 -1524
rect 10320 -1604 10360 -1556
rect 10320 -1636 10324 -1604
rect 10356 -1636 10360 -1604
rect 10320 -1684 10360 -1636
rect 10320 -1716 10324 -1684
rect 10356 -1716 10360 -1684
rect 10320 -1764 10360 -1716
rect 10320 -1796 10324 -1764
rect 10356 -1796 10360 -1764
rect 10320 -1844 10360 -1796
rect 10320 -1876 10324 -1844
rect 10356 -1876 10360 -1844
rect 10320 -1924 10360 -1876
rect 10320 -1956 10324 -1924
rect 10356 -1956 10360 -1924
rect 10320 -2004 10360 -1956
rect 10320 -2036 10324 -2004
rect 10356 -2036 10360 -2004
rect 10320 -2084 10360 -2036
rect 10320 -2116 10324 -2084
rect 10356 -2116 10360 -2084
rect 10320 -2164 10360 -2116
rect 10320 -2196 10324 -2164
rect 10356 -2196 10360 -2164
rect 10320 -2244 10360 -2196
rect 10320 -2276 10324 -2244
rect 10356 -2276 10360 -2244
rect 10320 -2324 10360 -2276
rect 10320 -2356 10324 -2324
rect 10356 -2356 10360 -2324
rect 10320 -2404 10360 -2356
rect 10320 -2436 10324 -2404
rect 10356 -2436 10360 -2404
rect 10320 -2484 10360 -2436
rect 10320 -2516 10324 -2484
rect 10356 -2516 10360 -2484
rect 10320 -2564 10360 -2516
rect 10320 -2596 10324 -2564
rect 10356 -2596 10360 -2564
rect 10320 -2644 10360 -2596
rect 10320 -2676 10324 -2644
rect 10356 -2676 10360 -2644
rect 10320 -2724 10360 -2676
rect 10320 -2756 10324 -2724
rect 10356 -2756 10360 -2724
rect 10320 -2804 10360 -2756
rect 10320 -2836 10324 -2804
rect 10356 -2836 10360 -2804
rect 10320 -2884 10360 -2836
rect 10320 -2916 10324 -2884
rect 10356 -2916 10360 -2884
rect 10320 -2964 10360 -2916
rect 10320 -2996 10324 -2964
rect 10356 -2996 10360 -2964
rect 10320 -3044 10360 -2996
rect 10320 -3076 10324 -3044
rect 10356 -3076 10360 -3044
rect 10320 -3124 10360 -3076
rect 10320 -3156 10324 -3124
rect 10356 -3156 10360 -3124
rect 10320 -3204 10360 -3156
rect 10320 -3236 10324 -3204
rect 10356 -3236 10360 -3204
rect 10320 -3284 10360 -3236
rect 10320 -3316 10324 -3284
rect 10356 -3316 10360 -3284
rect 10320 -3364 10360 -3316
rect 10320 -3396 10324 -3364
rect 10356 -3396 10360 -3364
rect 10320 -3444 10360 -3396
rect 10320 -3476 10324 -3444
rect 10356 -3476 10360 -3444
rect 10320 -3524 10360 -3476
rect 10320 -3556 10324 -3524
rect 10356 -3556 10360 -3524
rect 10320 -3604 10360 -3556
rect 10320 -3636 10324 -3604
rect 10356 -3636 10360 -3604
rect 10320 -3684 10360 -3636
rect 10320 -3716 10324 -3684
rect 10356 -3716 10360 -3684
rect 10320 -3720 10360 -3716
rect 10400 1036 10440 1040
rect 10400 1004 10404 1036
rect 10436 1004 10440 1036
rect 10400 956 10440 1004
rect 10400 924 10404 956
rect 10436 924 10440 956
rect 10400 876 10440 924
rect 10400 844 10404 876
rect 10436 844 10440 876
rect 10400 796 10440 844
rect 10400 764 10404 796
rect 10436 764 10440 796
rect 10400 716 10440 764
rect 10400 684 10404 716
rect 10436 684 10440 716
rect 10400 636 10440 684
rect 10400 604 10404 636
rect 10436 604 10440 636
rect 10400 556 10440 604
rect 10400 524 10404 556
rect 10436 524 10440 556
rect 10400 476 10440 524
rect 10400 444 10404 476
rect 10436 444 10440 476
rect 10400 396 10440 444
rect 10400 364 10404 396
rect 10436 364 10440 396
rect 10400 316 10440 364
rect 10400 284 10404 316
rect 10436 284 10440 316
rect 10400 236 10440 284
rect 10400 204 10404 236
rect 10436 204 10440 236
rect 10400 156 10440 204
rect 10400 124 10404 156
rect 10436 124 10440 156
rect 10400 76 10440 124
rect 10400 44 10404 76
rect 10436 44 10440 76
rect 10400 -4 10440 44
rect 10400 -36 10404 -4
rect 10436 -36 10440 -4
rect 10400 -84 10440 -36
rect 10400 -116 10404 -84
rect 10436 -116 10440 -84
rect 10400 -164 10440 -116
rect 10400 -196 10404 -164
rect 10436 -196 10440 -164
rect 10400 -244 10440 -196
rect 10400 -276 10404 -244
rect 10436 -276 10440 -244
rect 10400 -324 10440 -276
rect 10400 -356 10404 -324
rect 10436 -356 10440 -324
rect 10400 -404 10440 -356
rect 10400 -436 10404 -404
rect 10436 -436 10440 -404
rect 10400 -484 10440 -436
rect 10400 -516 10404 -484
rect 10436 -516 10440 -484
rect 10400 -564 10440 -516
rect 10400 -596 10404 -564
rect 10436 -596 10440 -564
rect 10400 -644 10440 -596
rect 10400 -676 10404 -644
rect 10436 -676 10440 -644
rect 10400 -724 10440 -676
rect 10400 -756 10404 -724
rect 10436 -756 10440 -724
rect 10400 -804 10440 -756
rect 10400 -836 10404 -804
rect 10436 -836 10440 -804
rect 10400 -884 10440 -836
rect 10400 -916 10404 -884
rect 10436 -916 10440 -884
rect 10400 -964 10440 -916
rect 10400 -996 10404 -964
rect 10436 -996 10440 -964
rect 10400 -1044 10440 -996
rect 10400 -1076 10404 -1044
rect 10436 -1076 10440 -1044
rect 10400 -1124 10440 -1076
rect 10400 -1156 10404 -1124
rect 10436 -1156 10440 -1124
rect 10400 -1204 10440 -1156
rect 10400 -1236 10404 -1204
rect 10436 -1236 10440 -1204
rect 10400 -1284 10440 -1236
rect 10400 -1316 10404 -1284
rect 10436 -1316 10440 -1284
rect 10400 -1364 10440 -1316
rect 10400 -1396 10404 -1364
rect 10436 -1396 10440 -1364
rect 10400 -1444 10440 -1396
rect 10400 -1476 10404 -1444
rect 10436 -1476 10440 -1444
rect 10400 -1524 10440 -1476
rect 10400 -1556 10404 -1524
rect 10436 -1556 10440 -1524
rect 10400 -1604 10440 -1556
rect 10400 -1636 10404 -1604
rect 10436 -1636 10440 -1604
rect 10400 -1684 10440 -1636
rect 10400 -1716 10404 -1684
rect 10436 -1716 10440 -1684
rect 10400 -1764 10440 -1716
rect 10400 -1796 10404 -1764
rect 10436 -1796 10440 -1764
rect 10400 -1844 10440 -1796
rect 10400 -1876 10404 -1844
rect 10436 -1876 10440 -1844
rect 10400 -1924 10440 -1876
rect 10400 -1956 10404 -1924
rect 10436 -1956 10440 -1924
rect 10400 -2004 10440 -1956
rect 10400 -2036 10404 -2004
rect 10436 -2036 10440 -2004
rect 10400 -2084 10440 -2036
rect 10400 -2116 10404 -2084
rect 10436 -2116 10440 -2084
rect 10400 -2164 10440 -2116
rect 10400 -2196 10404 -2164
rect 10436 -2196 10440 -2164
rect 10400 -2244 10440 -2196
rect 10400 -2276 10404 -2244
rect 10436 -2276 10440 -2244
rect 10400 -2324 10440 -2276
rect 10400 -2356 10404 -2324
rect 10436 -2356 10440 -2324
rect 10400 -2404 10440 -2356
rect 10400 -2436 10404 -2404
rect 10436 -2436 10440 -2404
rect 10400 -2484 10440 -2436
rect 10400 -2516 10404 -2484
rect 10436 -2516 10440 -2484
rect 10400 -2564 10440 -2516
rect 10400 -2596 10404 -2564
rect 10436 -2596 10440 -2564
rect 10400 -2644 10440 -2596
rect 10400 -2676 10404 -2644
rect 10436 -2676 10440 -2644
rect 10400 -2724 10440 -2676
rect 10400 -2756 10404 -2724
rect 10436 -2756 10440 -2724
rect 10400 -2804 10440 -2756
rect 10400 -2836 10404 -2804
rect 10436 -2836 10440 -2804
rect 10400 -2884 10440 -2836
rect 10400 -2916 10404 -2884
rect 10436 -2916 10440 -2884
rect 10400 -2964 10440 -2916
rect 10400 -2996 10404 -2964
rect 10436 -2996 10440 -2964
rect 10400 -3044 10440 -2996
rect 10400 -3076 10404 -3044
rect 10436 -3076 10440 -3044
rect 10400 -3124 10440 -3076
rect 10400 -3156 10404 -3124
rect 10436 -3156 10440 -3124
rect 10400 -3204 10440 -3156
rect 10400 -3236 10404 -3204
rect 10436 -3236 10440 -3204
rect 10400 -3284 10440 -3236
rect 10400 -3316 10404 -3284
rect 10436 -3316 10440 -3284
rect 10400 -3364 10440 -3316
rect 10400 -3396 10404 -3364
rect 10436 -3396 10440 -3364
rect 10400 -3444 10440 -3396
rect 10400 -3476 10404 -3444
rect 10436 -3476 10440 -3444
rect 10400 -3524 10440 -3476
rect 10400 -3556 10404 -3524
rect 10436 -3556 10440 -3524
rect 10400 -3604 10440 -3556
rect 10400 -3636 10404 -3604
rect 10436 -3636 10440 -3604
rect 10400 -3684 10440 -3636
rect 10400 -3716 10404 -3684
rect 10436 -3716 10440 -3684
rect 10400 -3720 10440 -3716
rect 10480 1036 10520 1040
rect 10480 1004 10484 1036
rect 10516 1004 10520 1036
rect 10480 956 10520 1004
rect 10480 924 10484 956
rect 10516 924 10520 956
rect 10480 876 10520 924
rect 10480 844 10484 876
rect 10516 844 10520 876
rect 10480 796 10520 844
rect 10480 764 10484 796
rect 10516 764 10520 796
rect 10480 716 10520 764
rect 10480 684 10484 716
rect 10516 684 10520 716
rect 10480 636 10520 684
rect 10480 604 10484 636
rect 10516 604 10520 636
rect 10480 556 10520 604
rect 10480 524 10484 556
rect 10516 524 10520 556
rect 10480 476 10520 524
rect 10480 444 10484 476
rect 10516 444 10520 476
rect 10480 396 10520 444
rect 10480 364 10484 396
rect 10516 364 10520 396
rect 10480 316 10520 364
rect 10480 284 10484 316
rect 10516 284 10520 316
rect 10480 236 10520 284
rect 10480 204 10484 236
rect 10516 204 10520 236
rect 10480 156 10520 204
rect 10480 124 10484 156
rect 10516 124 10520 156
rect 10480 76 10520 124
rect 10480 44 10484 76
rect 10516 44 10520 76
rect 10480 -4 10520 44
rect 10480 -36 10484 -4
rect 10516 -36 10520 -4
rect 10480 -84 10520 -36
rect 10480 -116 10484 -84
rect 10516 -116 10520 -84
rect 10480 -164 10520 -116
rect 10480 -196 10484 -164
rect 10516 -196 10520 -164
rect 10480 -244 10520 -196
rect 10480 -276 10484 -244
rect 10516 -276 10520 -244
rect 10480 -324 10520 -276
rect 10480 -356 10484 -324
rect 10516 -356 10520 -324
rect 10480 -404 10520 -356
rect 10480 -436 10484 -404
rect 10516 -436 10520 -404
rect 10480 -484 10520 -436
rect 10480 -516 10484 -484
rect 10516 -516 10520 -484
rect 10480 -564 10520 -516
rect 10480 -596 10484 -564
rect 10516 -596 10520 -564
rect 10480 -644 10520 -596
rect 10480 -676 10484 -644
rect 10516 -676 10520 -644
rect 10480 -724 10520 -676
rect 10480 -756 10484 -724
rect 10516 -756 10520 -724
rect 10480 -804 10520 -756
rect 10480 -836 10484 -804
rect 10516 -836 10520 -804
rect 10480 -884 10520 -836
rect 10480 -916 10484 -884
rect 10516 -916 10520 -884
rect 10480 -964 10520 -916
rect 10480 -996 10484 -964
rect 10516 -996 10520 -964
rect 10480 -1044 10520 -996
rect 10480 -1076 10484 -1044
rect 10516 -1076 10520 -1044
rect 10480 -1124 10520 -1076
rect 10480 -1156 10484 -1124
rect 10516 -1156 10520 -1124
rect 10480 -1204 10520 -1156
rect 10480 -1236 10484 -1204
rect 10516 -1236 10520 -1204
rect 10480 -1284 10520 -1236
rect 10480 -1316 10484 -1284
rect 10516 -1316 10520 -1284
rect 10480 -1364 10520 -1316
rect 10480 -1396 10484 -1364
rect 10516 -1396 10520 -1364
rect 10480 -1444 10520 -1396
rect 10480 -1476 10484 -1444
rect 10516 -1476 10520 -1444
rect 10480 -1524 10520 -1476
rect 10480 -1556 10484 -1524
rect 10516 -1556 10520 -1524
rect 10480 -1604 10520 -1556
rect 10480 -1636 10484 -1604
rect 10516 -1636 10520 -1604
rect 10480 -1684 10520 -1636
rect 10480 -1716 10484 -1684
rect 10516 -1716 10520 -1684
rect 10480 -1764 10520 -1716
rect 10480 -1796 10484 -1764
rect 10516 -1796 10520 -1764
rect 10480 -1844 10520 -1796
rect 10480 -1876 10484 -1844
rect 10516 -1876 10520 -1844
rect 10480 -1924 10520 -1876
rect 10480 -1956 10484 -1924
rect 10516 -1956 10520 -1924
rect 10480 -2004 10520 -1956
rect 10480 -2036 10484 -2004
rect 10516 -2036 10520 -2004
rect 10480 -2084 10520 -2036
rect 10480 -2116 10484 -2084
rect 10516 -2116 10520 -2084
rect 10480 -2164 10520 -2116
rect 10480 -2196 10484 -2164
rect 10516 -2196 10520 -2164
rect 10480 -2244 10520 -2196
rect 10480 -2276 10484 -2244
rect 10516 -2276 10520 -2244
rect 10480 -2324 10520 -2276
rect 10480 -2356 10484 -2324
rect 10516 -2356 10520 -2324
rect 10480 -2404 10520 -2356
rect 10480 -2436 10484 -2404
rect 10516 -2436 10520 -2404
rect 10480 -2484 10520 -2436
rect 10480 -2516 10484 -2484
rect 10516 -2516 10520 -2484
rect 10480 -2564 10520 -2516
rect 10480 -2596 10484 -2564
rect 10516 -2596 10520 -2564
rect 10480 -2644 10520 -2596
rect 10480 -2676 10484 -2644
rect 10516 -2676 10520 -2644
rect 10480 -2724 10520 -2676
rect 10480 -2756 10484 -2724
rect 10516 -2756 10520 -2724
rect 10480 -2804 10520 -2756
rect 10480 -2836 10484 -2804
rect 10516 -2836 10520 -2804
rect 10480 -2884 10520 -2836
rect 10480 -2916 10484 -2884
rect 10516 -2916 10520 -2884
rect 10480 -2964 10520 -2916
rect 10480 -2996 10484 -2964
rect 10516 -2996 10520 -2964
rect 10480 -3044 10520 -2996
rect 10480 -3076 10484 -3044
rect 10516 -3076 10520 -3044
rect 10480 -3124 10520 -3076
rect 10480 -3156 10484 -3124
rect 10516 -3156 10520 -3124
rect 10480 -3204 10520 -3156
rect 10480 -3236 10484 -3204
rect 10516 -3236 10520 -3204
rect 10480 -3284 10520 -3236
rect 10480 -3316 10484 -3284
rect 10516 -3316 10520 -3284
rect 10480 -3364 10520 -3316
rect 10480 -3396 10484 -3364
rect 10516 -3396 10520 -3364
rect 10480 -3444 10520 -3396
rect 10480 -3476 10484 -3444
rect 10516 -3476 10520 -3444
rect 10480 -3524 10520 -3476
rect 10480 -3556 10484 -3524
rect 10516 -3556 10520 -3524
rect 10480 -3604 10520 -3556
rect 10480 -3636 10484 -3604
rect 10516 -3636 10520 -3604
rect 10480 -3684 10520 -3636
rect 10480 -3716 10484 -3684
rect 10516 -3716 10520 -3684
rect 10480 -3720 10520 -3716
rect 10560 -164 10600 1040
rect 10560 -196 10564 -164
rect 10596 -196 10600 -164
rect 10560 -244 10600 -196
rect 10560 -276 10564 -244
rect 10596 -276 10600 -244
rect 10560 -324 10600 -276
rect 10560 -356 10564 -324
rect 10596 -356 10600 -324
rect 10560 -404 10600 -356
rect 10560 -436 10564 -404
rect 10596 -436 10600 -404
rect 10560 -484 10600 -436
rect 10560 -516 10564 -484
rect 10596 -516 10600 -484
rect 10560 -564 10600 -516
rect 10560 -596 10564 -564
rect 10596 -596 10600 -564
rect 10560 -644 10600 -596
rect 10560 -676 10564 -644
rect 10596 -676 10600 -644
rect 10560 -724 10600 -676
rect 10560 -756 10564 -724
rect 10596 -756 10600 -724
rect 10560 -804 10600 -756
rect 10560 -836 10564 -804
rect 10596 -836 10600 -804
rect 10560 -884 10600 -836
rect 10560 -916 10564 -884
rect 10596 -916 10600 -884
rect 10560 -964 10600 -916
rect 10560 -996 10564 -964
rect 10596 -996 10600 -964
rect 10560 -1044 10600 -996
rect 10560 -1076 10564 -1044
rect 10596 -1076 10600 -1044
rect 10560 -1124 10600 -1076
rect 10560 -1156 10564 -1124
rect 10596 -1156 10600 -1124
rect 10560 -1204 10600 -1156
rect 10560 -1236 10564 -1204
rect 10596 -1236 10600 -1204
rect 10560 -1284 10600 -1236
rect 10560 -1316 10564 -1284
rect 10596 -1316 10600 -1284
rect 10560 -1364 10600 -1316
rect 10560 -1396 10564 -1364
rect 10596 -1396 10600 -1364
rect 10560 -1444 10600 -1396
rect 10560 -1476 10564 -1444
rect 10596 -1476 10600 -1444
rect 10560 -1524 10600 -1476
rect 10560 -1556 10564 -1524
rect 10596 -1556 10600 -1524
rect 10560 -1604 10600 -1556
rect 10560 -1636 10564 -1604
rect 10596 -1636 10600 -1604
rect 10560 -1684 10600 -1636
rect 10560 -1716 10564 -1684
rect 10596 -1716 10600 -1684
rect 10560 -1764 10600 -1716
rect 10560 -1796 10564 -1764
rect 10596 -1796 10600 -1764
rect 10560 -1844 10600 -1796
rect 10560 -1876 10564 -1844
rect 10596 -1876 10600 -1844
rect 10560 -1924 10600 -1876
rect 10560 -1956 10564 -1924
rect 10596 -1956 10600 -1924
rect 10560 -2004 10600 -1956
rect 10560 -2036 10564 -2004
rect 10596 -2036 10600 -2004
rect 10560 -2084 10600 -2036
rect 10560 -2116 10564 -2084
rect 10596 -2116 10600 -2084
rect 10560 -2164 10600 -2116
rect 10560 -2196 10564 -2164
rect 10596 -2196 10600 -2164
rect 10560 -2244 10600 -2196
rect 10560 -2276 10564 -2244
rect 10596 -2276 10600 -2244
rect 10560 -2324 10600 -2276
rect 10560 -2356 10564 -2324
rect 10596 -2356 10600 -2324
rect 10560 -2404 10600 -2356
rect 10560 -2436 10564 -2404
rect 10596 -2436 10600 -2404
rect 10560 -2484 10600 -2436
rect 10560 -2516 10564 -2484
rect 10596 -2516 10600 -2484
rect 10560 -3720 10600 -2516
rect 10640 1036 10680 1040
rect 10640 1004 10644 1036
rect 10676 1004 10680 1036
rect 10640 956 10680 1004
rect 10640 924 10644 956
rect 10676 924 10680 956
rect 10640 876 10680 924
rect 10640 844 10644 876
rect 10676 844 10680 876
rect 10640 796 10680 844
rect 10640 764 10644 796
rect 10676 764 10680 796
rect 10640 716 10680 764
rect 10640 684 10644 716
rect 10676 684 10680 716
rect 10640 636 10680 684
rect 10640 604 10644 636
rect 10676 604 10680 636
rect 10640 556 10680 604
rect 10640 524 10644 556
rect 10676 524 10680 556
rect 10640 476 10680 524
rect 10640 444 10644 476
rect 10676 444 10680 476
rect 10640 396 10680 444
rect 10640 364 10644 396
rect 10676 364 10680 396
rect 10640 316 10680 364
rect 10640 284 10644 316
rect 10676 284 10680 316
rect 10640 236 10680 284
rect 10640 204 10644 236
rect 10676 204 10680 236
rect 10640 156 10680 204
rect 10640 124 10644 156
rect 10676 124 10680 156
rect 10640 76 10680 124
rect 10640 44 10644 76
rect 10676 44 10680 76
rect 10640 -4 10680 44
rect 10640 -36 10644 -4
rect 10676 -36 10680 -4
rect 10640 -84 10680 -36
rect 10640 -116 10644 -84
rect 10676 -116 10680 -84
rect 10640 -164 10680 -116
rect 10640 -196 10644 -164
rect 10676 -196 10680 -164
rect 10640 -244 10680 -196
rect 10640 -276 10644 -244
rect 10676 -276 10680 -244
rect 10640 -324 10680 -276
rect 10640 -356 10644 -324
rect 10676 -356 10680 -324
rect 10640 -404 10680 -356
rect 10640 -436 10644 -404
rect 10676 -436 10680 -404
rect 10640 -484 10680 -436
rect 10640 -516 10644 -484
rect 10676 -516 10680 -484
rect 10640 -564 10680 -516
rect 10640 -596 10644 -564
rect 10676 -596 10680 -564
rect 10640 -644 10680 -596
rect 10640 -676 10644 -644
rect 10676 -676 10680 -644
rect 10640 -724 10680 -676
rect 10640 -756 10644 -724
rect 10676 -756 10680 -724
rect 10640 -804 10680 -756
rect 10640 -836 10644 -804
rect 10676 -836 10680 -804
rect 10640 -884 10680 -836
rect 10640 -916 10644 -884
rect 10676 -916 10680 -884
rect 10640 -964 10680 -916
rect 10640 -996 10644 -964
rect 10676 -996 10680 -964
rect 10640 -1044 10680 -996
rect 10640 -1076 10644 -1044
rect 10676 -1076 10680 -1044
rect 10640 -1124 10680 -1076
rect 10640 -1156 10644 -1124
rect 10676 -1156 10680 -1124
rect 10640 -1204 10680 -1156
rect 10640 -1236 10644 -1204
rect 10676 -1236 10680 -1204
rect 10640 -1284 10680 -1236
rect 10640 -1316 10644 -1284
rect 10676 -1316 10680 -1284
rect 10640 -1364 10680 -1316
rect 10640 -1396 10644 -1364
rect 10676 -1396 10680 -1364
rect 10640 -1444 10680 -1396
rect 10640 -1476 10644 -1444
rect 10676 -1476 10680 -1444
rect 10640 -1524 10680 -1476
rect 10640 -1556 10644 -1524
rect 10676 -1556 10680 -1524
rect 10640 -1604 10680 -1556
rect 10640 -1636 10644 -1604
rect 10676 -1636 10680 -1604
rect 10640 -1684 10680 -1636
rect 10640 -1716 10644 -1684
rect 10676 -1716 10680 -1684
rect 10640 -1764 10680 -1716
rect 10640 -1796 10644 -1764
rect 10676 -1796 10680 -1764
rect 10640 -1844 10680 -1796
rect 10640 -1876 10644 -1844
rect 10676 -1876 10680 -1844
rect 10640 -1924 10680 -1876
rect 10640 -1956 10644 -1924
rect 10676 -1956 10680 -1924
rect 10640 -2004 10680 -1956
rect 10640 -2036 10644 -2004
rect 10676 -2036 10680 -2004
rect 10640 -2084 10680 -2036
rect 10640 -2116 10644 -2084
rect 10676 -2116 10680 -2084
rect 10640 -2164 10680 -2116
rect 10640 -2196 10644 -2164
rect 10676 -2196 10680 -2164
rect 10640 -2244 10680 -2196
rect 10640 -2276 10644 -2244
rect 10676 -2276 10680 -2244
rect 10640 -2324 10680 -2276
rect 10640 -2356 10644 -2324
rect 10676 -2356 10680 -2324
rect 10640 -2404 10680 -2356
rect 10640 -2436 10644 -2404
rect 10676 -2436 10680 -2404
rect 10640 -2484 10680 -2436
rect 10640 -2516 10644 -2484
rect 10676 -2516 10680 -2484
rect 10640 -2564 10680 -2516
rect 10640 -2596 10644 -2564
rect 10676 -2596 10680 -2564
rect 10640 -2644 10680 -2596
rect 10640 -2676 10644 -2644
rect 10676 -2676 10680 -2644
rect 10640 -2724 10680 -2676
rect 10640 -2756 10644 -2724
rect 10676 -2756 10680 -2724
rect 10640 -2804 10680 -2756
rect 10640 -2836 10644 -2804
rect 10676 -2836 10680 -2804
rect 10640 -2884 10680 -2836
rect 10640 -2916 10644 -2884
rect 10676 -2916 10680 -2884
rect 10640 -2964 10680 -2916
rect 10640 -2996 10644 -2964
rect 10676 -2996 10680 -2964
rect 10640 -3044 10680 -2996
rect 10640 -3076 10644 -3044
rect 10676 -3076 10680 -3044
rect 10640 -3124 10680 -3076
rect 10640 -3156 10644 -3124
rect 10676 -3156 10680 -3124
rect 10640 -3204 10680 -3156
rect 10640 -3236 10644 -3204
rect 10676 -3236 10680 -3204
rect 10640 -3284 10680 -3236
rect 10640 -3316 10644 -3284
rect 10676 -3316 10680 -3284
rect 10640 -3364 10680 -3316
rect 10640 -3396 10644 -3364
rect 10676 -3396 10680 -3364
rect 10640 -3444 10680 -3396
rect 10640 -3476 10644 -3444
rect 10676 -3476 10680 -3444
rect 10640 -3524 10680 -3476
rect 10640 -3556 10644 -3524
rect 10676 -3556 10680 -3524
rect 10640 -3604 10680 -3556
rect 10640 -3636 10644 -3604
rect 10676 -3636 10680 -3604
rect 10640 -3684 10680 -3636
rect 10640 -3716 10644 -3684
rect 10676 -3716 10680 -3684
rect 10640 -3720 10680 -3716
rect 10720 155 10760 1080
rect 10720 125 10725 155
rect 10755 125 10760 155
rect 10720 -405 10760 125
rect 10720 -435 10725 -405
rect 10755 -435 10760 -405
rect 10720 -2245 10760 -435
rect 10720 -2275 10725 -2245
rect 10755 -2275 10760 -2245
rect 10720 -2805 10760 -2275
rect 10720 -2835 10725 -2805
rect 10755 -2835 10760 -2805
rect 10720 -3720 10760 -2835
rect 10800 1036 10840 1040
rect 10800 1004 10804 1036
rect 10836 1004 10840 1036
rect 10800 956 10840 1004
rect 10800 924 10804 956
rect 10836 924 10840 956
rect 10800 876 10840 924
rect 10800 844 10804 876
rect 10836 844 10840 876
rect 10800 796 10840 844
rect 10800 764 10804 796
rect 10836 764 10840 796
rect 10800 716 10840 764
rect 10800 684 10804 716
rect 10836 684 10840 716
rect 10800 636 10840 684
rect 10800 604 10804 636
rect 10836 604 10840 636
rect 10800 556 10840 604
rect 10800 524 10804 556
rect 10836 524 10840 556
rect 10800 476 10840 524
rect 10800 444 10804 476
rect 10836 444 10840 476
rect 10800 396 10840 444
rect 10800 364 10804 396
rect 10836 364 10840 396
rect 10800 316 10840 364
rect 10800 284 10804 316
rect 10836 284 10840 316
rect 10800 236 10840 284
rect 10800 204 10804 236
rect 10836 204 10840 236
rect 10800 156 10840 204
rect 10800 124 10804 156
rect 10836 124 10840 156
rect 10800 76 10840 124
rect 10800 44 10804 76
rect 10836 44 10840 76
rect 10800 -4 10840 44
rect 10800 -36 10804 -4
rect 10836 -36 10840 -4
rect 10800 -84 10840 -36
rect 10800 -116 10804 -84
rect 10836 -116 10840 -84
rect 10800 -164 10840 -116
rect 10800 -196 10804 -164
rect 10836 -196 10840 -164
rect 10800 -244 10840 -196
rect 10800 -276 10804 -244
rect 10836 -276 10840 -244
rect 10800 -324 10840 -276
rect 10800 -356 10804 -324
rect 10836 -356 10840 -324
rect 10800 -404 10840 -356
rect 10800 -436 10804 -404
rect 10836 -436 10840 -404
rect 10800 -484 10840 -436
rect 10800 -516 10804 -484
rect 10836 -516 10840 -484
rect 10800 -564 10840 -516
rect 10800 -596 10804 -564
rect 10836 -596 10840 -564
rect 10800 -644 10840 -596
rect 10800 -676 10804 -644
rect 10836 -676 10840 -644
rect 10800 -724 10840 -676
rect 10800 -756 10804 -724
rect 10836 -756 10840 -724
rect 10800 -804 10840 -756
rect 10800 -836 10804 -804
rect 10836 -836 10840 -804
rect 10800 -884 10840 -836
rect 10800 -916 10804 -884
rect 10836 -916 10840 -884
rect 10800 -964 10840 -916
rect 10800 -996 10804 -964
rect 10836 -996 10840 -964
rect 10800 -1044 10840 -996
rect 10800 -1076 10804 -1044
rect 10836 -1076 10840 -1044
rect 10800 -1124 10840 -1076
rect 10800 -1156 10804 -1124
rect 10836 -1156 10840 -1124
rect 10800 -1204 10840 -1156
rect 10800 -1236 10804 -1204
rect 10836 -1236 10840 -1204
rect 10800 -1284 10840 -1236
rect 10800 -1316 10804 -1284
rect 10836 -1316 10840 -1284
rect 10800 -1364 10840 -1316
rect 10800 -1396 10804 -1364
rect 10836 -1396 10840 -1364
rect 10800 -1444 10840 -1396
rect 10800 -1476 10804 -1444
rect 10836 -1476 10840 -1444
rect 10800 -1524 10840 -1476
rect 10800 -1556 10804 -1524
rect 10836 -1556 10840 -1524
rect 10800 -1604 10840 -1556
rect 10800 -1636 10804 -1604
rect 10836 -1636 10840 -1604
rect 10800 -1684 10840 -1636
rect 10800 -1716 10804 -1684
rect 10836 -1716 10840 -1684
rect 10800 -1764 10840 -1716
rect 10800 -1796 10804 -1764
rect 10836 -1796 10840 -1764
rect 10800 -1844 10840 -1796
rect 10800 -1876 10804 -1844
rect 10836 -1876 10840 -1844
rect 10800 -1924 10840 -1876
rect 10800 -1956 10804 -1924
rect 10836 -1956 10840 -1924
rect 10800 -2004 10840 -1956
rect 10800 -2036 10804 -2004
rect 10836 -2036 10840 -2004
rect 10800 -2084 10840 -2036
rect 10800 -2116 10804 -2084
rect 10836 -2116 10840 -2084
rect 10800 -2164 10840 -2116
rect 10800 -2196 10804 -2164
rect 10836 -2196 10840 -2164
rect 10800 -2244 10840 -2196
rect 10800 -2276 10804 -2244
rect 10836 -2276 10840 -2244
rect 10800 -2324 10840 -2276
rect 10800 -2356 10804 -2324
rect 10836 -2356 10840 -2324
rect 10800 -2404 10840 -2356
rect 10800 -2436 10804 -2404
rect 10836 -2436 10840 -2404
rect 10800 -2484 10840 -2436
rect 10800 -2516 10804 -2484
rect 10836 -2516 10840 -2484
rect 10800 -2564 10840 -2516
rect 10800 -2596 10804 -2564
rect 10836 -2596 10840 -2564
rect 10800 -2644 10840 -2596
rect 10800 -2676 10804 -2644
rect 10836 -2676 10840 -2644
rect 10800 -2724 10840 -2676
rect 10800 -2756 10804 -2724
rect 10836 -2756 10840 -2724
rect 10800 -2804 10840 -2756
rect 10800 -2836 10804 -2804
rect 10836 -2836 10840 -2804
rect 10800 -2884 10840 -2836
rect 10800 -2916 10804 -2884
rect 10836 -2916 10840 -2884
rect 10800 -2964 10840 -2916
rect 10800 -2996 10804 -2964
rect 10836 -2996 10840 -2964
rect 10800 -3044 10840 -2996
rect 10800 -3076 10804 -3044
rect 10836 -3076 10840 -3044
rect 10800 -3124 10840 -3076
rect 10800 -3156 10804 -3124
rect 10836 -3156 10840 -3124
rect 10800 -3204 10840 -3156
rect 10800 -3236 10804 -3204
rect 10836 -3236 10840 -3204
rect 10800 -3284 10840 -3236
rect 10800 -3316 10804 -3284
rect 10836 -3316 10840 -3284
rect 10800 -3364 10840 -3316
rect 10800 -3396 10804 -3364
rect 10836 -3396 10840 -3364
rect 10800 -3444 10840 -3396
rect 10800 -3476 10804 -3444
rect 10836 -3476 10840 -3444
rect 10800 -3524 10840 -3476
rect 10800 -3556 10804 -3524
rect 10836 -3556 10840 -3524
rect 10800 -3604 10840 -3556
rect 10800 -3636 10804 -3604
rect 10836 -3636 10840 -3604
rect 10800 -3684 10840 -3636
rect 10800 -3716 10804 -3684
rect 10836 -3716 10840 -3684
rect 10800 -3720 10840 -3716
rect 10880 315 10920 1080
rect 10880 285 10885 315
rect 10915 285 10920 315
rect 10880 -565 10920 285
rect 10880 -595 10885 -565
rect 10915 -595 10920 -565
rect 10880 -2085 10920 -595
rect 10880 -2115 10885 -2085
rect 10915 -2115 10920 -2085
rect 10880 -2965 10920 -2115
rect 10880 -2995 10885 -2965
rect 10915 -2995 10920 -2965
rect 10880 -3720 10920 -2995
rect 10960 1036 11000 1080
rect 10960 1004 10964 1036
rect 10996 1004 11000 1036
rect 10960 956 11000 1004
rect 10960 924 10964 956
rect 10996 924 11000 956
rect 10960 876 11000 924
rect 10960 844 10964 876
rect 10996 844 11000 876
rect 10960 796 11000 844
rect 10960 764 10964 796
rect 10996 764 11000 796
rect 10960 716 11000 764
rect 10960 684 10964 716
rect 10996 684 11000 716
rect 10960 636 11000 684
rect 10960 604 10964 636
rect 10996 604 11000 636
rect 10960 556 11000 604
rect 10960 524 10964 556
rect 10996 524 11000 556
rect 10960 476 11000 524
rect 10960 444 10964 476
rect 10996 444 11000 476
rect 10960 396 11000 444
rect 10960 364 10964 396
rect 10996 364 11000 396
rect 10960 316 11000 364
rect 10960 284 10964 316
rect 10996 284 11000 316
rect 10960 236 11000 284
rect 10960 204 10964 236
rect 10996 204 11000 236
rect 10960 156 11000 204
rect 10960 124 10964 156
rect 10996 124 11000 156
rect 10960 76 11000 124
rect 10960 44 10964 76
rect 10996 44 11000 76
rect 10960 -4 11000 44
rect 10960 -36 10964 -4
rect 10996 -36 11000 -4
rect 10960 -84 11000 -36
rect 10960 -116 10964 -84
rect 10996 -116 11000 -84
rect 10960 -164 11000 -116
rect 10960 -196 10964 -164
rect 10996 -196 11000 -164
rect 10960 -244 11000 -196
rect 10960 -276 10964 -244
rect 10996 -276 11000 -244
rect 10960 -324 11000 -276
rect 10960 -356 10964 -324
rect 10996 -356 11000 -324
rect 10960 -404 11000 -356
rect 10960 -436 10964 -404
rect 10996 -436 11000 -404
rect 10960 -484 11000 -436
rect 10960 -516 10964 -484
rect 10996 -516 11000 -484
rect 10960 -564 11000 -516
rect 10960 -596 10964 -564
rect 10996 -596 11000 -564
rect 10960 -644 11000 -596
rect 10960 -676 10964 -644
rect 10996 -676 11000 -644
rect 10960 -724 11000 -676
rect 10960 -756 10964 -724
rect 10996 -756 11000 -724
rect 10960 -804 11000 -756
rect 10960 -836 10964 -804
rect 10996 -836 11000 -804
rect 10960 -884 11000 -836
rect 10960 -916 10964 -884
rect 10996 -916 11000 -884
rect 10960 -964 11000 -916
rect 10960 -996 10964 -964
rect 10996 -996 11000 -964
rect 10960 -1044 11000 -996
rect 10960 -1076 10964 -1044
rect 10996 -1076 11000 -1044
rect 10960 -1124 11000 -1076
rect 10960 -1156 10964 -1124
rect 10996 -1156 11000 -1124
rect 10960 -1204 11000 -1156
rect 10960 -1236 10964 -1204
rect 10996 -1236 11000 -1204
rect 10960 -1284 11000 -1236
rect 10960 -1316 10964 -1284
rect 10996 -1316 11000 -1284
rect 10960 -1364 11000 -1316
rect 10960 -1396 10964 -1364
rect 10996 -1396 11000 -1364
rect 10960 -1444 11000 -1396
rect 10960 -1476 10964 -1444
rect 10996 -1476 11000 -1444
rect 10960 -1524 11000 -1476
rect 10960 -1556 10964 -1524
rect 10996 -1556 11000 -1524
rect 10960 -1604 11000 -1556
rect 10960 -1636 10964 -1604
rect 10996 -1636 11000 -1604
rect 10960 -1684 11000 -1636
rect 10960 -1716 10964 -1684
rect 10996 -1716 11000 -1684
rect 10960 -1764 11000 -1716
rect 10960 -1796 10964 -1764
rect 10996 -1796 11000 -1764
rect 10960 -1844 11000 -1796
rect 10960 -1876 10964 -1844
rect 10996 -1876 11000 -1844
rect 10960 -1924 11000 -1876
rect 10960 -1956 10964 -1924
rect 10996 -1956 11000 -1924
rect 10960 -2004 11000 -1956
rect 10960 -2036 10964 -2004
rect 10996 -2036 11000 -2004
rect 10960 -2084 11000 -2036
rect 10960 -2116 10964 -2084
rect 10996 -2116 11000 -2084
rect 10960 -2164 11000 -2116
rect 10960 -2196 10964 -2164
rect 10996 -2196 11000 -2164
rect 10960 -2244 11000 -2196
rect 10960 -2276 10964 -2244
rect 10996 -2276 11000 -2244
rect 10960 -2324 11000 -2276
rect 10960 -2356 10964 -2324
rect 10996 -2356 11000 -2324
rect 10960 -2404 11000 -2356
rect 10960 -2436 10964 -2404
rect 10996 -2436 11000 -2404
rect 10960 -2484 11000 -2436
rect 10960 -2516 10964 -2484
rect 10996 -2516 11000 -2484
rect 10960 -2564 11000 -2516
rect 10960 -2596 10964 -2564
rect 10996 -2596 11000 -2564
rect 10960 -2644 11000 -2596
rect 10960 -2676 10964 -2644
rect 10996 -2676 11000 -2644
rect 10960 -2724 11000 -2676
rect 10960 -2756 10964 -2724
rect 10996 -2756 11000 -2724
rect 10960 -2804 11000 -2756
rect 10960 -2836 10964 -2804
rect 10996 -2836 11000 -2804
rect 10960 -2884 11000 -2836
rect 10960 -2916 10964 -2884
rect 10996 -2916 11000 -2884
rect 10960 -2964 11000 -2916
rect 10960 -2996 10964 -2964
rect 10996 -2996 11000 -2964
rect 10960 -3044 11000 -2996
rect 10960 -3076 10964 -3044
rect 10996 -3076 11000 -3044
rect 10960 -3124 11000 -3076
rect 10960 -3156 10964 -3124
rect 10996 -3156 11000 -3124
rect 10960 -3204 11000 -3156
rect 10960 -3236 10964 -3204
rect 10996 -3236 11000 -3204
rect 10960 -3284 11000 -3236
rect 10960 -3316 10964 -3284
rect 10996 -3316 11000 -3284
rect 10960 -3364 11000 -3316
rect 10960 -3396 10964 -3364
rect 10996 -3396 11000 -3364
rect 10960 -3444 11000 -3396
rect 10960 -3476 10964 -3444
rect 10996 -3476 11000 -3444
rect 10960 -3524 11000 -3476
rect 10960 -3556 10964 -3524
rect 10996 -3556 11000 -3524
rect 10960 -3604 11000 -3556
rect 10960 -3636 10964 -3604
rect 10996 -3636 11000 -3604
rect 10960 -3684 11000 -3636
rect 10960 -3716 10964 -3684
rect 10996 -3716 11000 -3684
rect 10960 -3720 11000 -3716
<< via3 >>
rect -716 1035 -684 1036
rect -716 1005 -715 1035
rect -715 1005 -685 1035
rect -685 1005 -684 1035
rect -716 1004 -684 1005
rect -716 955 -684 956
rect -716 925 -715 955
rect -715 925 -685 955
rect -685 925 -684 955
rect -716 924 -684 925
rect -716 875 -684 876
rect -716 845 -715 875
rect -715 845 -685 875
rect -685 845 -684 875
rect -716 844 -684 845
rect -716 764 -684 796
rect -716 684 -684 716
rect -716 635 -684 636
rect -716 605 -715 635
rect -715 605 -685 635
rect -685 605 -684 635
rect -716 604 -684 605
rect -716 555 -684 556
rect -716 525 -715 555
rect -715 525 -685 555
rect -685 525 -684 555
rect -716 524 -684 525
rect -716 475 -684 476
rect -716 445 -715 475
rect -715 445 -685 475
rect -685 445 -684 475
rect -716 444 -684 445
rect -716 395 -684 396
rect -716 365 -715 395
rect -715 365 -685 395
rect -685 365 -684 395
rect -716 364 -684 365
rect -716 315 -684 316
rect -716 285 -715 315
rect -715 285 -685 315
rect -685 285 -684 315
rect -716 284 -684 285
rect -716 235 -684 236
rect -716 205 -715 235
rect -715 205 -685 235
rect -685 205 -684 235
rect -716 204 -684 205
rect -716 155 -684 156
rect -716 125 -715 155
rect -715 125 -685 155
rect -685 125 -684 155
rect -716 124 -684 125
rect -716 75 -684 76
rect -716 45 -715 75
rect -715 45 -685 75
rect -685 45 -684 75
rect -716 44 -684 45
rect -716 -5 -684 -4
rect -716 -35 -715 -5
rect -715 -35 -685 -5
rect -685 -35 -684 -5
rect -716 -36 -684 -35
rect -716 -85 -684 -84
rect -716 -115 -715 -85
rect -715 -115 -685 -85
rect -685 -115 -684 -85
rect -716 -116 -684 -115
rect -716 -165 -684 -164
rect -716 -195 -715 -165
rect -715 -195 -685 -165
rect -685 -195 -684 -165
rect -716 -196 -684 -195
rect -716 -245 -684 -244
rect -716 -275 -715 -245
rect -715 -275 -685 -245
rect -685 -275 -684 -245
rect -716 -276 -684 -275
rect -716 -325 -684 -324
rect -716 -355 -715 -325
rect -715 -355 -685 -325
rect -685 -355 -684 -325
rect -716 -356 -684 -355
rect -716 -405 -684 -404
rect -716 -435 -715 -405
rect -715 -435 -685 -405
rect -685 -435 -684 -405
rect -716 -436 -684 -435
rect -716 -485 -684 -484
rect -716 -515 -715 -485
rect -715 -515 -685 -485
rect -685 -515 -684 -485
rect -716 -516 -684 -515
rect -716 -565 -684 -564
rect -716 -595 -715 -565
rect -715 -595 -685 -565
rect -685 -595 -684 -565
rect -716 -596 -684 -595
rect -716 -645 -684 -644
rect -716 -675 -715 -645
rect -715 -675 -685 -645
rect -685 -675 -684 -645
rect -716 -676 -684 -675
rect -716 -725 -684 -724
rect -716 -755 -715 -725
rect -715 -755 -685 -725
rect -685 -755 -684 -725
rect -716 -756 -684 -755
rect -716 -805 -684 -804
rect -716 -835 -715 -805
rect -715 -835 -685 -805
rect -685 -835 -684 -805
rect -716 -836 -684 -835
rect -716 -885 -684 -884
rect -716 -915 -715 -885
rect -715 -915 -685 -885
rect -685 -915 -684 -885
rect -716 -916 -684 -915
rect -716 -996 -684 -964
rect -716 -1076 -684 -1044
rect -716 -1125 -684 -1124
rect -716 -1155 -715 -1125
rect -715 -1155 -685 -1125
rect -685 -1155 -684 -1125
rect -716 -1156 -684 -1155
rect -716 -1205 -684 -1204
rect -716 -1235 -715 -1205
rect -715 -1235 -685 -1205
rect -685 -1235 -684 -1205
rect -716 -1236 -684 -1235
rect -716 -1285 -684 -1284
rect -716 -1315 -715 -1285
rect -715 -1315 -685 -1285
rect -685 -1315 -684 -1285
rect -716 -1316 -684 -1315
rect -716 -1365 -684 -1364
rect -716 -1395 -715 -1365
rect -715 -1395 -685 -1365
rect -685 -1395 -684 -1365
rect -716 -1396 -684 -1395
rect -716 -1445 -684 -1444
rect -716 -1475 -715 -1445
rect -715 -1475 -685 -1445
rect -685 -1475 -684 -1445
rect -716 -1476 -684 -1475
rect -716 -1525 -684 -1524
rect -716 -1555 -715 -1525
rect -715 -1555 -685 -1525
rect -685 -1555 -684 -1525
rect -716 -1556 -684 -1555
rect -716 -1636 -684 -1604
rect -716 -1716 -684 -1684
rect -716 -1765 -684 -1764
rect -716 -1795 -715 -1765
rect -715 -1795 -685 -1765
rect -685 -1795 -684 -1765
rect -716 -1796 -684 -1795
rect -716 -1845 -684 -1844
rect -716 -1875 -715 -1845
rect -715 -1875 -685 -1845
rect -685 -1875 -684 -1845
rect -716 -1876 -684 -1875
rect -716 -1925 -684 -1924
rect -716 -1955 -715 -1925
rect -715 -1955 -685 -1925
rect -685 -1955 -684 -1925
rect -716 -1956 -684 -1955
rect -716 -2005 -684 -2004
rect -716 -2035 -715 -2005
rect -715 -2035 -685 -2005
rect -685 -2035 -684 -2005
rect -716 -2036 -684 -2035
rect -716 -2085 -684 -2084
rect -716 -2115 -715 -2085
rect -715 -2115 -685 -2085
rect -685 -2115 -684 -2085
rect -716 -2116 -684 -2115
rect -716 -2165 -684 -2164
rect -716 -2195 -715 -2165
rect -715 -2195 -685 -2165
rect -685 -2195 -684 -2165
rect -716 -2196 -684 -2195
rect -716 -2245 -684 -2244
rect -716 -2275 -715 -2245
rect -715 -2275 -685 -2245
rect -685 -2275 -684 -2245
rect -716 -2276 -684 -2275
rect -716 -2325 -684 -2324
rect -716 -2355 -715 -2325
rect -715 -2355 -685 -2325
rect -685 -2355 -684 -2325
rect -716 -2356 -684 -2355
rect -716 -2405 -684 -2404
rect -716 -2435 -715 -2405
rect -715 -2435 -685 -2405
rect -685 -2435 -684 -2405
rect -716 -2436 -684 -2435
rect -716 -2485 -684 -2484
rect -716 -2515 -715 -2485
rect -715 -2515 -685 -2485
rect -685 -2515 -684 -2485
rect -716 -2516 -684 -2515
rect -716 -2565 -684 -2564
rect -716 -2595 -715 -2565
rect -715 -2595 -685 -2565
rect -685 -2595 -684 -2565
rect -716 -2596 -684 -2595
rect -716 -2645 -684 -2644
rect -716 -2675 -715 -2645
rect -715 -2675 -685 -2645
rect -685 -2675 -684 -2645
rect -716 -2676 -684 -2675
rect -716 -2725 -684 -2724
rect -716 -2755 -715 -2725
rect -715 -2755 -685 -2725
rect -685 -2755 -684 -2725
rect -716 -2756 -684 -2755
rect -716 -2805 -684 -2804
rect -716 -2835 -715 -2805
rect -715 -2835 -685 -2805
rect -685 -2835 -684 -2805
rect -716 -2836 -684 -2835
rect -716 -2885 -684 -2884
rect -716 -2915 -715 -2885
rect -715 -2915 -685 -2885
rect -685 -2915 -684 -2885
rect -716 -2916 -684 -2915
rect -716 -2965 -684 -2964
rect -716 -2995 -715 -2965
rect -715 -2995 -685 -2965
rect -685 -2995 -684 -2965
rect -716 -2996 -684 -2995
rect -716 -3045 -684 -3044
rect -716 -3075 -715 -3045
rect -715 -3075 -685 -3045
rect -685 -3075 -684 -3045
rect -716 -3076 -684 -3075
rect -716 -3125 -684 -3124
rect -716 -3155 -715 -3125
rect -715 -3155 -685 -3125
rect -685 -3155 -684 -3125
rect -716 -3156 -684 -3155
rect -716 -3205 -684 -3204
rect -716 -3235 -715 -3205
rect -715 -3235 -685 -3205
rect -685 -3235 -684 -3205
rect -716 -3236 -684 -3235
rect -716 -3285 -684 -3284
rect -716 -3315 -715 -3285
rect -715 -3315 -685 -3285
rect -685 -3315 -684 -3285
rect -716 -3316 -684 -3315
rect -716 -3396 -684 -3364
rect -716 -3476 -684 -3444
rect -716 -3525 -684 -3524
rect -716 -3555 -715 -3525
rect -715 -3555 -685 -3525
rect -685 -3555 -684 -3525
rect -716 -3556 -684 -3555
rect -716 -3605 -684 -3604
rect -716 -3635 -715 -3605
rect -715 -3635 -685 -3605
rect -685 -3635 -684 -3605
rect -716 -3636 -684 -3635
rect -716 -3685 -684 -3684
rect -716 -3715 -715 -3685
rect -715 -3715 -685 -3685
rect -685 -3715 -684 -3685
rect -716 -3716 -684 -3715
rect -556 1035 -524 1036
rect -556 1005 -555 1035
rect -555 1005 -525 1035
rect -525 1005 -524 1035
rect -556 1004 -524 1005
rect -556 955 -524 956
rect -556 925 -555 955
rect -555 925 -525 955
rect -525 925 -524 955
rect -556 924 -524 925
rect -556 875 -524 876
rect -556 845 -555 875
rect -555 845 -525 875
rect -525 845 -524 875
rect -556 844 -524 845
rect -556 764 -524 796
rect -556 684 -524 716
rect -556 635 -524 636
rect -556 605 -555 635
rect -555 605 -525 635
rect -525 605 -524 635
rect -556 604 -524 605
rect -556 555 -524 556
rect -556 525 -555 555
rect -555 525 -525 555
rect -525 525 -524 555
rect -556 524 -524 525
rect -556 475 -524 476
rect -556 445 -555 475
rect -555 445 -525 475
rect -525 445 -524 475
rect -556 444 -524 445
rect -556 395 -524 396
rect -556 365 -555 395
rect -555 365 -525 395
rect -525 365 -524 395
rect -556 364 -524 365
rect -556 315 -524 316
rect -556 285 -555 315
rect -555 285 -525 315
rect -525 285 -524 315
rect -556 284 -524 285
rect -556 235 -524 236
rect -556 205 -555 235
rect -555 205 -525 235
rect -525 205 -524 235
rect -556 204 -524 205
rect -556 155 -524 156
rect -556 125 -555 155
rect -555 125 -525 155
rect -525 125 -524 155
rect -556 124 -524 125
rect -556 75 -524 76
rect -556 45 -555 75
rect -555 45 -525 75
rect -525 45 -524 75
rect -556 44 -524 45
rect -556 -5 -524 -4
rect -556 -35 -555 -5
rect -555 -35 -525 -5
rect -525 -35 -524 -5
rect -556 -36 -524 -35
rect -556 -85 -524 -84
rect -556 -115 -555 -85
rect -555 -115 -525 -85
rect -525 -115 -524 -85
rect -556 -116 -524 -115
rect -556 -165 -524 -164
rect -556 -195 -555 -165
rect -555 -195 -525 -165
rect -525 -195 -524 -165
rect -556 -196 -524 -195
rect -556 -245 -524 -244
rect -556 -275 -555 -245
rect -555 -275 -525 -245
rect -525 -275 -524 -245
rect -556 -276 -524 -275
rect -556 -325 -524 -324
rect -556 -355 -555 -325
rect -555 -355 -525 -325
rect -525 -355 -524 -325
rect -556 -356 -524 -355
rect -556 -405 -524 -404
rect -556 -435 -555 -405
rect -555 -435 -525 -405
rect -525 -435 -524 -405
rect -556 -436 -524 -435
rect -556 -485 -524 -484
rect -556 -515 -555 -485
rect -555 -515 -525 -485
rect -525 -515 -524 -485
rect -556 -516 -524 -515
rect -556 -565 -524 -564
rect -556 -595 -555 -565
rect -555 -595 -525 -565
rect -525 -595 -524 -565
rect -556 -596 -524 -595
rect -556 -645 -524 -644
rect -556 -675 -555 -645
rect -555 -675 -525 -645
rect -525 -675 -524 -645
rect -556 -676 -524 -675
rect -556 -725 -524 -724
rect -556 -755 -555 -725
rect -555 -755 -525 -725
rect -525 -755 -524 -725
rect -556 -756 -524 -755
rect -556 -805 -524 -804
rect -556 -835 -555 -805
rect -555 -835 -525 -805
rect -525 -835 -524 -805
rect -556 -836 -524 -835
rect -556 -885 -524 -884
rect -556 -915 -555 -885
rect -555 -915 -525 -885
rect -525 -915 -524 -885
rect -556 -916 -524 -915
rect -556 -996 -524 -964
rect -556 -1076 -524 -1044
rect -556 -1125 -524 -1124
rect -556 -1155 -555 -1125
rect -555 -1155 -525 -1125
rect -525 -1155 -524 -1125
rect -556 -1156 -524 -1155
rect -556 -1205 -524 -1204
rect -556 -1235 -555 -1205
rect -555 -1235 -525 -1205
rect -525 -1235 -524 -1205
rect -556 -1236 -524 -1235
rect -556 -1285 -524 -1284
rect -556 -1315 -555 -1285
rect -555 -1315 -525 -1285
rect -525 -1315 -524 -1285
rect -556 -1316 -524 -1315
rect -556 -1365 -524 -1364
rect -556 -1395 -555 -1365
rect -555 -1395 -525 -1365
rect -525 -1395 -524 -1365
rect -556 -1396 -524 -1395
rect -556 -1445 -524 -1444
rect -556 -1475 -555 -1445
rect -555 -1475 -525 -1445
rect -525 -1475 -524 -1445
rect -556 -1476 -524 -1475
rect -556 -1525 -524 -1524
rect -556 -1555 -555 -1525
rect -555 -1555 -525 -1525
rect -525 -1555 -524 -1525
rect -556 -1556 -524 -1555
rect -556 -1636 -524 -1604
rect -556 -1716 -524 -1684
rect -556 -1765 -524 -1764
rect -556 -1795 -555 -1765
rect -555 -1795 -525 -1765
rect -525 -1795 -524 -1765
rect -556 -1796 -524 -1795
rect -556 -1845 -524 -1844
rect -556 -1875 -555 -1845
rect -555 -1875 -525 -1845
rect -525 -1875 -524 -1845
rect -556 -1876 -524 -1875
rect -556 -1925 -524 -1924
rect -556 -1955 -555 -1925
rect -555 -1955 -525 -1925
rect -525 -1955 -524 -1925
rect -556 -1956 -524 -1955
rect -556 -2005 -524 -2004
rect -556 -2035 -555 -2005
rect -555 -2035 -525 -2005
rect -525 -2035 -524 -2005
rect -556 -2036 -524 -2035
rect -556 -2085 -524 -2084
rect -556 -2115 -555 -2085
rect -555 -2115 -525 -2085
rect -525 -2115 -524 -2085
rect -556 -2116 -524 -2115
rect -556 -2165 -524 -2164
rect -556 -2195 -555 -2165
rect -555 -2195 -525 -2165
rect -525 -2195 -524 -2165
rect -556 -2196 -524 -2195
rect -556 -2245 -524 -2244
rect -556 -2275 -555 -2245
rect -555 -2275 -525 -2245
rect -525 -2275 -524 -2245
rect -556 -2276 -524 -2275
rect -556 -2325 -524 -2324
rect -556 -2355 -555 -2325
rect -555 -2355 -525 -2325
rect -525 -2355 -524 -2325
rect -556 -2356 -524 -2355
rect -556 -2405 -524 -2404
rect -556 -2435 -555 -2405
rect -555 -2435 -525 -2405
rect -525 -2435 -524 -2405
rect -556 -2436 -524 -2435
rect -556 -2485 -524 -2484
rect -556 -2515 -555 -2485
rect -555 -2515 -525 -2485
rect -525 -2515 -524 -2485
rect -556 -2516 -524 -2515
rect -556 -2565 -524 -2564
rect -556 -2595 -555 -2565
rect -555 -2595 -525 -2565
rect -525 -2595 -524 -2565
rect -556 -2596 -524 -2595
rect -556 -2645 -524 -2644
rect -556 -2675 -555 -2645
rect -555 -2675 -525 -2645
rect -525 -2675 -524 -2645
rect -556 -2676 -524 -2675
rect -556 -2725 -524 -2724
rect -556 -2755 -555 -2725
rect -555 -2755 -525 -2725
rect -525 -2755 -524 -2725
rect -556 -2756 -524 -2755
rect -556 -2805 -524 -2804
rect -556 -2835 -555 -2805
rect -555 -2835 -525 -2805
rect -525 -2835 -524 -2805
rect -556 -2836 -524 -2835
rect -556 -2885 -524 -2884
rect -556 -2915 -555 -2885
rect -555 -2915 -525 -2885
rect -525 -2915 -524 -2885
rect -556 -2916 -524 -2915
rect -556 -2965 -524 -2964
rect -556 -2995 -555 -2965
rect -555 -2995 -525 -2965
rect -525 -2995 -524 -2965
rect -556 -2996 -524 -2995
rect -556 -3045 -524 -3044
rect -556 -3075 -555 -3045
rect -555 -3075 -525 -3045
rect -525 -3075 -524 -3045
rect -556 -3076 -524 -3075
rect -556 -3125 -524 -3124
rect -556 -3155 -555 -3125
rect -555 -3155 -525 -3125
rect -525 -3155 -524 -3125
rect -556 -3156 -524 -3155
rect -556 -3205 -524 -3204
rect -556 -3235 -555 -3205
rect -555 -3235 -525 -3205
rect -525 -3235 -524 -3205
rect -556 -3236 -524 -3235
rect -556 -3285 -524 -3284
rect -556 -3315 -555 -3285
rect -555 -3315 -525 -3285
rect -525 -3315 -524 -3285
rect -556 -3316 -524 -3315
rect -556 -3396 -524 -3364
rect -556 -3476 -524 -3444
rect -556 -3525 -524 -3524
rect -556 -3555 -555 -3525
rect -555 -3555 -525 -3525
rect -525 -3555 -524 -3525
rect -556 -3556 -524 -3555
rect -556 -3605 -524 -3604
rect -556 -3635 -555 -3605
rect -555 -3635 -525 -3605
rect -525 -3635 -524 -3605
rect -556 -3636 -524 -3635
rect -556 -3685 -524 -3684
rect -556 -3715 -555 -3685
rect -555 -3715 -525 -3685
rect -525 -3715 -524 -3685
rect -556 -3716 -524 -3715
rect -396 1035 -364 1036
rect -396 1005 -395 1035
rect -395 1005 -365 1035
rect -365 1005 -364 1035
rect -396 1004 -364 1005
rect -396 955 -364 956
rect -396 925 -395 955
rect -395 925 -365 955
rect -365 925 -364 955
rect -396 924 -364 925
rect -396 875 -364 876
rect -396 845 -395 875
rect -395 845 -365 875
rect -365 845 -364 875
rect -396 844 -364 845
rect -396 764 -364 796
rect -396 684 -364 716
rect -396 635 -364 636
rect -396 605 -395 635
rect -395 605 -365 635
rect -365 605 -364 635
rect -396 604 -364 605
rect -396 555 -364 556
rect -396 525 -395 555
rect -395 525 -365 555
rect -365 525 -364 555
rect -396 524 -364 525
rect -396 444 -364 476
rect -396 395 -364 396
rect -396 365 -395 395
rect -395 365 -365 395
rect -365 365 -364 395
rect -396 364 -364 365
rect -396 315 -364 316
rect -396 285 -395 315
rect -395 285 -365 315
rect -365 285 -364 315
rect -396 284 -364 285
rect -396 235 -364 236
rect -396 205 -395 235
rect -395 205 -365 235
rect -365 205 -364 235
rect -396 204 -364 205
rect -396 155 -364 156
rect -396 125 -395 155
rect -395 125 -365 155
rect -365 125 -364 155
rect -396 124 -364 125
rect -396 75 -364 76
rect -396 45 -395 75
rect -395 45 -365 75
rect -365 45 -364 75
rect -396 44 -364 45
rect -396 -5 -364 -4
rect -396 -35 -395 -5
rect -395 -35 -365 -5
rect -365 -35 -364 -5
rect -396 -36 -364 -35
rect -396 -85 -364 -84
rect -396 -115 -395 -85
rect -395 -115 -365 -85
rect -365 -115 -364 -85
rect -396 -116 -364 -115
rect -396 -165 -364 -164
rect -396 -195 -395 -165
rect -395 -195 -365 -165
rect -365 -195 -364 -165
rect -396 -196 -364 -195
rect -396 -245 -364 -244
rect -396 -275 -395 -245
rect -395 -275 -365 -245
rect -365 -275 -364 -245
rect -396 -276 -364 -275
rect -396 -325 -364 -324
rect -396 -355 -395 -325
rect -395 -355 -365 -325
rect -365 -355 -364 -325
rect -396 -356 -364 -355
rect -396 -405 -364 -404
rect -396 -435 -395 -405
rect -395 -435 -365 -405
rect -365 -435 -364 -405
rect -396 -436 -364 -435
rect -396 -485 -364 -484
rect -396 -515 -395 -485
rect -395 -515 -365 -485
rect -365 -515 -364 -485
rect -396 -516 -364 -515
rect -396 -565 -364 -564
rect -396 -595 -395 -565
rect -395 -595 -365 -565
rect -365 -595 -364 -565
rect -396 -596 -364 -595
rect -396 -645 -364 -644
rect -396 -675 -395 -645
rect -395 -675 -365 -645
rect -365 -675 -364 -645
rect -396 -676 -364 -675
rect -396 -756 -364 -724
rect -396 -805 -364 -804
rect -396 -835 -395 -805
rect -395 -835 -365 -805
rect -365 -835 -364 -805
rect -396 -836 -364 -835
rect -396 -885 -364 -884
rect -396 -915 -395 -885
rect -395 -915 -365 -885
rect -365 -915 -364 -885
rect -396 -916 -364 -915
rect -396 -996 -364 -964
rect -396 -1076 -364 -1044
rect -396 -1125 -364 -1124
rect -396 -1155 -395 -1125
rect -395 -1155 -365 -1125
rect -365 -1155 -364 -1125
rect -396 -1156 -364 -1155
rect -396 -1205 -364 -1204
rect -396 -1235 -395 -1205
rect -395 -1235 -365 -1205
rect -365 -1235 -364 -1205
rect -396 -1236 -364 -1235
rect -396 -1285 -364 -1284
rect -396 -1315 -395 -1285
rect -395 -1315 -365 -1285
rect -365 -1315 -364 -1285
rect -396 -1316 -364 -1315
rect -396 -1365 -364 -1364
rect -396 -1395 -395 -1365
rect -395 -1395 -365 -1365
rect -365 -1395 -364 -1365
rect -396 -1396 -364 -1395
rect -396 -1445 -364 -1444
rect -396 -1475 -395 -1445
rect -395 -1475 -365 -1445
rect -365 -1475 -364 -1445
rect -396 -1476 -364 -1475
rect -396 -1525 -364 -1524
rect -396 -1555 -395 -1525
rect -395 -1555 -365 -1525
rect -365 -1555 -364 -1525
rect -396 -1556 -364 -1555
rect -396 -1636 -364 -1604
rect -396 -1716 -364 -1684
rect -396 -1765 -364 -1764
rect -396 -1795 -395 -1765
rect -395 -1795 -365 -1765
rect -365 -1795 -364 -1765
rect -396 -1796 -364 -1795
rect -396 -1845 -364 -1844
rect -396 -1875 -395 -1845
rect -395 -1875 -365 -1845
rect -365 -1875 -364 -1845
rect -396 -1876 -364 -1875
rect -396 -1956 -364 -1924
rect -396 -2005 -364 -2004
rect -396 -2035 -395 -2005
rect -395 -2035 -365 -2005
rect -365 -2035 -364 -2005
rect -396 -2036 -364 -2035
rect -396 -2085 -364 -2084
rect -396 -2115 -395 -2085
rect -395 -2115 -365 -2085
rect -365 -2115 -364 -2085
rect -396 -2116 -364 -2115
rect -396 -2165 -364 -2164
rect -396 -2195 -395 -2165
rect -395 -2195 -365 -2165
rect -365 -2195 -364 -2165
rect -396 -2196 -364 -2195
rect -396 -2245 -364 -2244
rect -396 -2275 -395 -2245
rect -395 -2275 -365 -2245
rect -365 -2275 -364 -2245
rect -396 -2276 -364 -2275
rect -396 -2325 -364 -2324
rect -396 -2355 -395 -2325
rect -395 -2355 -365 -2325
rect -365 -2355 -364 -2325
rect -396 -2356 -364 -2355
rect -396 -2405 -364 -2404
rect -396 -2435 -395 -2405
rect -395 -2435 -365 -2405
rect -365 -2435 -364 -2405
rect -396 -2436 -364 -2435
rect -396 -2485 -364 -2484
rect -396 -2515 -395 -2485
rect -395 -2515 -365 -2485
rect -365 -2515 -364 -2485
rect -396 -2516 -364 -2515
rect -396 -2565 -364 -2564
rect -396 -2595 -395 -2565
rect -395 -2595 -365 -2565
rect -365 -2595 -364 -2565
rect -396 -2596 -364 -2595
rect -396 -2645 -364 -2644
rect -396 -2675 -395 -2645
rect -395 -2675 -365 -2645
rect -365 -2675 -364 -2645
rect -396 -2676 -364 -2675
rect -396 -2725 -364 -2724
rect -396 -2755 -395 -2725
rect -395 -2755 -365 -2725
rect -365 -2755 -364 -2725
rect -396 -2756 -364 -2755
rect -396 -2805 -364 -2804
rect -396 -2835 -395 -2805
rect -395 -2835 -365 -2805
rect -365 -2835 -364 -2805
rect -396 -2836 -364 -2835
rect -396 -2885 -364 -2884
rect -396 -2915 -395 -2885
rect -395 -2915 -365 -2885
rect -365 -2915 -364 -2885
rect -396 -2916 -364 -2915
rect -396 -2965 -364 -2964
rect -396 -2995 -395 -2965
rect -395 -2995 -365 -2965
rect -365 -2995 -364 -2965
rect -396 -2996 -364 -2995
rect -396 -3045 -364 -3044
rect -396 -3075 -395 -3045
rect -395 -3075 -365 -3045
rect -365 -3075 -364 -3045
rect -396 -3076 -364 -3075
rect -396 -3156 -364 -3124
rect -396 -3205 -364 -3204
rect -396 -3235 -395 -3205
rect -395 -3235 -365 -3205
rect -365 -3235 -364 -3205
rect -396 -3236 -364 -3235
rect -396 -3285 -364 -3284
rect -396 -3315 -395 -3285
rect -395 -3315 -365 -3285
rect -365 -3315 -364 -3285
rect -396 -3316 -364 -3315
rect -396 -3396 -364 -3364
rect -396 -3476 -364 -3444
rect -396 -3525 -364 -3524
rect -396 -3555 -395 -3525
rect -395 -3555 -365 -3525
rect -365 -3555 -364 -3525
rect -396 -3556 -364 -3555
rect -396 -3605 -364 -3604
rect -396 -3635 -395 -3605
rect -395 -3635 -365 -3605
rect -365 -3635 -364 -3605
rect -396 -3636 -364 -3635
rect -396 -3685 -364 -3684
rect -396 -3715 -395 -3685
rect -395 -3715 -365 -3685
rect -365 -3715 -364 -3685
rect -396 -3716 -364 -3715
rect -316 1035 -284 1036
rect -316 1005 -315 1035
rect -315 1005 -285 1035
rect -285 1005 -284 1035
rect -316 1004 -284 1005
rect -316 955 -284 956
rect -316 925 -315 955
rect -315 925 -285 955
rect -285 925 -284 955
rect -316 924 -284 925
rect -316 875 -284 876
rect -316 845 -315 875
rect -315 845 -285 875
rect -285 845 -284 875
rect -316 844 -284 845
rect -316 764 -284 796
rect -316 684 -284 716
rect -316 635 -284 636
rect -316 605 -315 635
rect -315 605 -285 635
rect -285 605 -284 635
rect -316 604 -284 605
rect -316 555 -284 556
rect -316 525 -315 555
rect -315 525 -285 555
rect -285 525 -284 555
rect -316 524 -284 525
rect -316 444 -284 476
rect -316 395 -284 396
rect -316 365 -315 395
rect -315 365 -285 395
rect -285 365 -284 395
rect -316 364 -284 365
rect -316 284 -284 316
rect -316 235 -284 236
rect -316 205 -315 235
rect -315 205 -285 235
rect -285 205 -284 235
rect -316 204 -284 205
rect -316 124 -284 156
rect -316 75 -284 76
rect -316 45 -315 75
rect -315 45 -285 75
rect -285 45 -284 75
rect -316 44 -284 45
rect -316 -5 -284 -4
rect -316 -35 -315 -5
rect -315 -35 -285 -5
rect -285 -35 -284 -5
rect -316 -36 -284 -35
rect -316 -85 -284 -84
rect -316 -115 -315 -85
rect -315 -115 -285 -85
rect -285 -115 -284 -85
rect -316 -116 -284 -115
rect -316 -2565 -284 -2564
rect -316 -2595 -315 -2565
rect -315 -2595 -285 -2565
rect -285 -2595 -284 -2565
rect -316 -2596 -284 -2595
rect -316 -2645 -284 -2644
rect -316 -2675 -315 -2645
rect -315 -2675 -285 -2645
rect -285 -2675 -284 -2645
rect -316 -2676 -284 -2675
rect -316 -2725 -284 -2724
rect -316 -2755 -315 -2725
rect -315 -2755 -285 -2725
rect -285 -2755 -284 -2725
rect -316 -2756 -284 -2755
rect -316 -2836 -284 -2804
rect -316 -2885 -284 -2884
rect -316 -2915 -315 -2885
rect -315 -2915 -285 -2885
rect -285 -2915 -284 -2885
rect -316 -2916 -284 -2915
rect -316 -2996 -284 -2964
rect -316 -3045 -284 -3044
rect -316 -3075 -315 -3045
rect -315 -3075 -285 -3045
rect -285 -3075 -284 -3045
rect -316 -3076 -284 -3075
rect -316 -3156 -284 -3124
rect -316 -3205 -284 -3204
rect -316 -3235 -315 -3205
rect -315 -3235 -285 -3205
rect -285 -3235 -284 -3205
rect -316 -3236 -284 -3235
rect -316 -3285 -284 -3284
rect -316 -3315 -315 -3285
rect -315 -3315 -285 -3285
rect -285 -3315 -284 -3285
rect -316 -3316 -284 -3315
rect -316 -3396 -284 -3364
rect -316 -3476 -284 -3444
rect -316 -3525 -284 -3524
rect -316 -3555 -315 -3525
rect -315 -3555 -285 -3525
rect -285 -3555 -284 -3525
rect -316 -3556 -284 -3555
rect -316 -3605 -284 -3604
rect -316 -3635 -315 -3605
rect -315 -3635 -285 -3605
rect -285 -3635 -284 -3605
rect -316 -3636 -284 -3635
rect -316 -3685 -284 -3684
rect -316 -3715 -315 -3685
rect -315 -3715 -285 -3685
rect -285 -3715 -284 -3685
rect -316 -3716 -284 -3715
rect -236 1035 -204 1036
rect -236 1005 -235 1035
rect -235 1005 -205 1035
rect -205 1005 -204 1035
rect -236 1004 -204 1005
rect -236 955 -204 956
rect -236 925 -235 955
rect -235 925 -205 955
rect -205 925 -204 955
rect -236 924 -204 925
rect -236 875 -204 876
rect -236 845 -235 875
rect -235 845 -205 875
rect -205 845 -204 875
rect -236 844 -204 845
rect -236 764 -204 796
rect -236 684 -204 716
rect -236 635 -204 636
rect -236 605 -235 635
rect -235 605 -205 635
rect -205 605 -204 635
rect -236 604 -204 605
rect -236 555 -204 556
rect -236 525 -235 555
rect -235 525 -205 555
rect -205 525 -204 555
rect -236 524 -204 525
rect -236 444 -204 476
rect -236 395 -204 396
rect -236 365 -235 395
rect -235 365 -205 395
rect -205 365 -204 395
rect -236 364 -204 365
rect -236 284 -204 316
rect -236 235 -204 236
rect -236 205 -235 235
rect -235 205 -205 235
rect -205 205 -204 235
rect -236 204 -204 205
rect -236 124 -204 156
rect -236 75 -204 76
rect -236 45 -235 75
rect -235 45 -205 75
rect -205 45 -204 75
rect -236 44 -204 45
rect -236 -5 -204 -4
rect -236 -35 -235 -5
rect -235 -35 -205 -5
rect -205 -35 -204 -5
rect -236 -36 -204 -35
rect -236 -85 -204 -84
rect -236 -115 -235 -85
rect -235 -115 -205 -85
rect -205 -115 -204 -85
rect -236 -116 -204 -115
rect -236 -165 -204 -164
rect -236 -195 -235 -165
rect -235 -195 -205 -165
rect -205 -195 -204 -165
rect -236 -196 -204 -195
rect -236 -245 -204 -244
rect -236 -275 -235 -245
rect -235 -275 -205 -245
rect -205 -275 -204 -245
rect -236 -276 -204 -275
rect -236 -325 -204 -324
rect -236 -355 -235 -325
rect -235 -355 -205 -325
rect -205 -355 -204 -325
rect -236 -356 -204 -355
rect -236 -436 -204 -404
rect -236 -485 -204 -484
rect -236 -515 -235 -485
rect -235 -515 -205 -485
rect -205 -515 -204 -485
rect -236 -516 -204 -515
rect -236 -596 -204 -564
rect -236 -645 -204 -644
rect -236 -675 -235 -645
rect -235 -675 -205 -645
rect -205 -675 -204 -645
rect -236 -676 -204 -675
rect -236 -756 -204 -724
rect -236 -805 -204 -804
rect -236 -835 -235 -805
rect -235 -835 -205 -805
rect -205 -835 -204 -805
rect -236 -836 -204 -835
rect -236 -885 -204 -884
rect -236 -915 -235 -885
rect -235 -915 -205 -885
rect -205 -915 -204 -885
rect -236 -916 -204 -915
rect -236 -996 -204 -964
rect -236 -1076 -204 -1044
rect -236 -1125 -204 -1124
rect -236 -1155 -235 -1125
rect -235 -1155 -205 -1125
rect -205 -1155 -204 -1125
rect -236 -1156 -204 -1155
rect -236 -1205 -204 -1204
rect -236 -1235 -235 -1205
rect -235 -1235 -205 -1205
rect -205 -1235 -204 -1205
rect -236 -1236 -204 -1235
rect -236 -1285 -204 -1284
rect -236 -1315 -235 -1285
rect -235 -1315 -205 -1285
rect -205 -1315 -204 -1285
rect -236 -1316 -204 -1315
rect -236 -1365 -204 -1364
rect -236 -1395 -235 -1365
rect -235 -1395 -205 -1365
rect -205 -1395 -204 -1365
rect -236 -1396 -204 -1395
rect -236 -1445 -204 -1444
rect -236 -1475 -235 -1445
rect -235 -1475 -205 -1445
rect -205 -1475 -204 -1445
rect -236 -1476 -204 -1475
rect -236 -1525 -204 -1524
rect -236 -1555 -235 -1525
rect -235 -1555 -205 -1525
rect -205 -1555 -204 -1525
rect -236 -1556 -204 -1555
rect -236 -1636 -204 -1604
rect -236 -1716 -204 -1684
rect -236 -1765 -204 -1764
rect -236 -1795 -235 -1765
rect -235 -1795 -205 -1765
rect -205 -1795 -204 -1765
rect -236 -1796 -204 -1795
rect -236 -1845 -204 -1844
rect -236 -1875 -235 -1845
rect -235 -1875 -205 -1845
rect -205 -1875 -204 -1845
rect -236 -1876 -204 -1875
rect -236 -1956 -204 -1924
rect -236 -2005 -204 -2004
rect -236 -2035 -235 -2005
rect -235 -2035 -205 -2005
rect -205 -2035 -204 -2005
rect -236 -2036 -204 -2035
rect -236 -2116 -204 -2084
rect -236 -2165 -204 -2164
rect -236 -2195 -235 -2165
rect -235 -2195 -205 -2165
rect -205 -2195 -204 -2165
rect -236 -2196 -204 -2195
rect -236 -2276 -204 -2244
rect -236 -2325 -204 -2324
rect -236 -2355 -235 -2325
rect -235 -2355 -205 -2325
rect -205 -2355 -204 -2325
rect -236 -2356 -204 -2355
rect -236 -2405 -204 -2404
rect -236 -2435 -235 -2405
rect -235 -2435 -205 -2405
rect -205 -2435 -204 -2405
rect -236 -2436 -204 -2435
rect -236 -2485 -204 -2484
rect -236 -2515 -235 -2485
rect -235 -2515 -205 -2485
rect -205 -2515 -204 -2485
rect -236 -2516 -204 -2515
rect -236 -2565 -204 -2564
rect -236 -2595 -235 -2565
rect -235 -2595 -205 -2565
rect -205 -2595 -204 -2565
rect -236 -2596 -204 -2595
rect -236 -2645 -204 -2644
rect -236 -2675 -235 -2645
rect -235 -2675 -205 -2645
rect -205 -2675 -204 -2645
rect -236 -2676 -204 -2675
rect -236 -2725 -204 -2724
rect -236 -2755 -235 -2725
rect -235 -2755 -205 -2725
rect -205 -2755 -204 -2725
rect -236 -2756 -204 -2755
rect -236 -2836 -204 -2804
rect -236 -2885 -204 -2884
rect -236 -2915 -235 -2885
rect -235 -2915 -205 -2885
rect -205 -2915 -204 -2885
rect -236 -2916 -204 -2915
rect -236 -2996 -204 -2964
rect -236 -3045 -204 -3044
rect -236 -3075 -235 -3045
rect -235 -3075 -205 -3045
rect -205 -3075 -204 -3045
rect -236 -3076 -204 -3075
rect -236 -3156 -204 -3124
rect -236 -3205 -204 -3204
rect -236 -3235 -235 -3205
rect -235 -3235 -205 -3205
rect -205 -3235 -204 -3205
rect -236 -3236 -204 -3235
rect -236 -3285 -204 -3284
rect -236 -3315 -235 -3285
rect -235 -3315 -205 -3285
rect -205 -3315 -204 -3285
rect -236 -3316 -204 -3315
rect -236 -3396 -204 -3364
rect -236 -3476 -204 -3444
rect -236 -3525 -204 -3524
rect -236 -3555 -235 -3525
rect -235 -3555 -205 -3525
rect -205 -3555 -204 -3525
rect -236 -3556 -204 -3555
rect -236 -3605 -204 -3604
rect -236 -3635 -235 -3605
rect -235 -3635 -205 -3605
rect -205 -3635 -204 -3605
rect -236 -3636 -204 -3635
rect -236 -3685 -204 -3684
rect -236 -3715 -235 -3685
rect -235 -3715 -205 -3685
rect -205 -3715 -204 -3685
rect -236 -3716 -204 -3715
rect -156 1035 -124 1036
rect -156 1005 -155 1035
rect -155 1005 -125 1035
rect -125 1005 -124 1035
rect -156 1004 -124 1005
rect -156 955 -124 956
rect -156 925 -155 955
rect -155 925 -125 955
rect -125 925 -124 955
rect -156 924 -124 925
rect -156 875 -124 876
rect -156 845 -155 875
rect -155 845 -125 875
rect -125 845 -124 875
rect -156 844 -124 845
rect -156 764 -124 796
rect -156 684 -124 716
rect -156 635 -124 636
rect -156 605 -155 635
rect -155 605 -125 635
rect -125 605 -124 635
rect -156 604 -124 605
rect -156 555 -124 556
rect -156 525 -155 555
rect -155 525 -125 555
rect -125 525 -124 555
rect -156 524 -124 525
rect -156 444 -124 476
rect -156 395 -124 396
rect -156 365 -155 395
rect -155 365 -125 395
rect -125 365 -124 395
rect -156 364 -124 365
rect -156 284 -124 316
rect -156 235 -124 236
rect -156 205 -155 235
rect -155 205 -125 235
rect -125 205 -124 235
rect -156 204 -124 205
rect -156 124 -124 156
rect -156 75 -124 76
rect -156 45 -155 75
rect -155 45 -125 75
rect -125 45 -124 75
rect -156 44 -124 45
rect -156 -5 -124 -4
rect -156 -35 -155 -5
rect -155 -35 -125 -5
rect -125 -35 -124 -5
rect -156 -36 -124 -35
rect -156 -85 -124 -84
rect -156 -115 -155 -85
rect -155 -115 -125 -85
rect -125 -115 -124 -85
rect -156 -116 -124 -115
rect -156 -165 -124 -164
rect -156 -195 -155 -165
rect -155 -195 -125 -165
rect -125 -195 -124 -165
rect -156 -196 -124 -195
rect -156 -245 -124 -244
rect -156 -275 -155 -245
rect -155 -275 -125 -245
rect -125 -275 -124 -245
rect -156 -276 -124 -275
rect -156 -325 -124 -324
rect -156 -355 -155 -325
rect -155 -355 -125 -325
rect -125 -355 -124 -325
rect -156 -356 -124 -355
rect -156 -436 -124 -404
rect -156 -485 -124 -484
rect -156 -515 -155 -485
rect -155 -515 -125 -485
rect -125 -515 -124 -485
rect -156 -516 -124 -515
rect -156 -596 -124 -564
rect -156 -645 -124 -644
rect -156 -675 -155 -645
rect -155 -675 -125 -645
rect -125 -675 -124 -645
rect -156 -676 -124 -675
rect -156 -756 -124 -724
rect -156 -805 -124 -804
rect -156 -835 -155 -805
rect -155 -835 -125 -805
rect -125 -835 -124 -805
rect -156 -836 -124 -835
rect -156 -885 -124 -884
rect -156 -915 -155 -885
rect -155 -915 -125 -885
rect -125 -915 -124 -885
rect -156 -916 -124 -915
rect -156 -996 -124 -964
rect -156 -1076 -124 -1044
rect -156 -1125 -124 -1124
rect -156 -1155 -155 -1125
rect -155 -1155 -125 -1125
rect -125 -1155 -124 -1125
rect -156 -1156 -124 -1155
rect -156 -1205 -124 -1204
rect -156 -1235 -155 -1205
rect -155 -1235 -125 -1205
rect -125 -1235 -124 -1205
rect -156 -1236 -124 -1235
rect -156 -1285 -124 -1284
rect -156 -1315 -155 -1285
rect -155 -1315 -125 -1285
rect -125 -1315 -124 -1285
rect -156 -1316 -124 -1315
rect -156 -1365 -124 -1364
rect -156 -1395 -155 -1365
rect -155 -1395 -125 -1365
rect -125 -1395 -124 -1365
rect -156 -1396 -124 -1395
rect -156 -1445 -124 -1444
rect -156 -1475 -155 -1445
rect -155 -1475 -125 -1445
rect -125 -1475 -124 -1445
rect -156 -1476 -124 -1475
rect -156 -1525 -124 -1524
rect -156 -1555 -155 -1525
rect -155 -1555 -125 -1525
rect -125 -1555 -124 -1525
rect -156 -1556 -124 -1555
rect -156 -1636 -124 -1604
rect -156 -1716 -124 -1684
rect -156 -1765 -124 -1764
rect -156 -1795 -155 -1765
rect -155 -1795 -125 -1765
rect -125 -1795 -124 -1765
rect -156 -1796 -124 -1795
rect -156 -1845 -124 -1844
rect -156 -1875 -155 -1845
rect -155 -1875 -125 -1845
rect -125 -1875 -124 -1845
rect -156 -1876 -124 -1875
rect -156 -1956 -124 -1924
rect -156 -2005 -124 -2004
rect -156 -2035 -155 -2005
rect -155 -2035 -125 -2005
rect -125 -2035 -124 -2005
rect -156 -2036 -124 -2035
rect -156 -2116 -124 -2084
rect -156 -2165 -124 -2164
rect -156 -2195 -155 -2165
rect -155 -2195 -125 -2165
rect -125 -2195 -124 -2165
rect -156 -2196 -124 -2195
rect -156 -2276 -124 -2244
rect -156 -2325 -124 -2324
rect -156 -2355 -155 -2325
rect -155 -2355 -125 -2325
rect -125 -2355 -124 -2325
rect -156 -2356 -124 -2355
rect -156 -2405 -124 -2404
rect -156 -2435 -155 -2405
rect -155 -2435 -125 -2405
rect -125 -2435 -124 -2405
rect -156 -2436 -124 -2435
rect -156 -2485 -124 -2484
rect -156 -2515 -155 -2485
rect -155 -2515 -125 -2485
rect -125 -2515 -124 -2485
rect -156 -2516 -124 -2515
rect -156 -2565 -124 -2564
rect -156 -2595 -155 -2565
rect -155 -2595 -125 -2565
rect -125 -2595 -124 -2565
rect -156 -2596 -124 -2595
rect -156 -2645 -124 -2644
rect -156 -2675 -155 -2645
rect -155 -2675 -125 -2645
rect -125 -2675 -124 -2645
rect -156 -2676 -124 -2675
rect -156 -2725 -124 -2724
rect -156 -2755 -155 -2725
rect -155 -2755 -125 -2725
rect -125 -2755 -124 -2725
rect -156 -2756 -124 -2755
rect -156 -2836 -124 -2804
rect -156 -2885 -124 -2884
rect -156 -2915 -155 -2885
rect -155 -2915 -125 -2885
rect -125 -2915 -124 -2885
rect -156 -2916 -124 -2915
rect -156 -2996 -124 -2964
rect -156 -3045 -124 -3044
rect -156 -3075 -155 -3045
rect -155 -3075 -125 -3045
rect -125 -3075 -124 -3045
rect -156 -3076 -124 -3075
rect -156 -3156 -124 -3124
rect -156 -3205 -124 -3204
rect -156 -3235 -155 -3205
rect -155 -3235 -125 -3205
rect -125 -3235 -124 -3205
rect -156 -3236 -124 -3235
rect -156 -3285 -124 -3284
rect -156 -3315 -155 -3285
rect -155 -3315 -125 -3285
rect -125 -3315 -124 -3285
rect -156 -3316 -124 -3315
rect -156 -3396 -124 -3364
rect -156 -3476 -124 -3444
rect -156 -3525 -124 -3524
rect -156 -3555 -155 -3525
rect -155 -3555 -125 -3525
rect -125 -3555 -124 -3525
rect -156 -3556 -124 -3555
rect -156 -3605 -124 -3604
rect -156 -3635 -155 -3605
rect -155 -3635 -125 -3605
rect -125 -3635 -124 -3605
rect -156 -3636 -124 -3635
rect -156 -3685 -124 -3684
rect -156 -3715 -155 -3685
rect -155 -3715 -125 -3685
rect -125 -3715 -124 -3685
rect -156 -3716 -124 -3715
rect -76 1035 -44 1036
rect -76 1005 -75 1035
rect -75 1005 -45 1035
rect -45 1005 -44 1035
rect -76 1004 -44 1005
rect -76 955 -44 956
rect -76 925 -75 955
rect -75 925 -45 955
rect -45 925 -44 955
rect -76 924 -44 925
rect -76 875 -44 876
rect -76 845 -75 875
rect -75 845 -45 875
rect -45 845 -44 875
rect -76 844 -44 845
rect -76 764 -44 796
rect -76 684 -44 716
rect -76 635 -44 636
rect -76 605 -75 635
rect -75 605 -45 635
rect -45 605 -44 635
rect -76 604 -44 605
rect -76 555 -44 556
rect -76 525 -75 555
rect -75 525 -45 555
rect -45 525 -44 555
rect -76 524 -44 525
rect -76 444 -44 476
rect -76 395 -44 396
rect -76 365 -75 395
rect -75 365 -45 395
rect -45 365 -44 395
rect -76 364 -44 365
rect -76 284 -44 316
rect -76 235 -44 236
rect -76 205 -75 235
rect -75 205 -45 235
rect -45 205 -44 235
rect -76 204 -44 205
rect -76 124 -44 156
rect -76 75 -44 76
rect -76 45 -75 75
rect -75 45 -45 75
rect -45 45 -44 75
rect -76 44 -44 45
rect -76 -5 -44 -4
rect -76 -35 -75 -5
rect -75 -35 -45 -5
rect -45 -35 -44 -5
rect -76 -36 -44 -35
rect -76 -85 -44 -84
rect -76 -115 -75 -85
rect -75 -115 -45 -85
rect -45 -115 -44 -85
rect -76 -116 -44 -115
rect -76 -165 -44 -164
rect -76 -195 -75 -165
rect -75 -195 -45 -165
rect -45 -195 -44 -165
rect -76 -196 -44 -195
rect -76 -245 -44 -244
rect -76 -275 -75 -245
rect -75 -275 -45 -245
rect -45 -275 -44 -245
rect -76 -276 -44 -275
rect -76 -325 -44 -324
rect -76 -355 -75 -325
rect -75 -355 -45 -325
rect -45 -355 -44 -325
rect -76 -356 -44 -355
rect -76 -436 -44 -404
rect -76 -485 -44 -484
rect -76 -515 -75 -485
rect -75 -515 -45 -485
rect -45 -515 -44 -485
rect -76 -516 -44 -515
rect -76 -596 -44 -564
rect -76 -645 -44 -644
rect -76 -675 -75 -645
rect -75 -675 -45 -645
rect -45 -675 -44 -645
rect -76 -676 -44 -675
rect -76 -756 -44 -724
rect -76 -805 -44 -804
rect -76 -835 -75 -805
rect -75 -835 -45 -805
rect -45 -835 -44 -805
rect -76 -836 -44 -835
rect -76 -885 -44 -884
rect -76 -915 -75 -885
rect -75 -915 -45 -885
rect -45 -915 -44 -885
rect -76 -916 -44 -915
rect -76 -996 -44 -964
rect -76 -1076 -44 -1044
rect -76 -1125 -44 -1124
rect -76 -1155 -75 -1125
rect -75 -1155 -45 -1125
rect -45 -1155 -44 -1125
rect -76 -1156 -44 -1155
rect -76 -1205 -44 -1204
rect -76 -1235 -75 -1205
rect -75 -1235 -45 -1205
rect -45 -1235 -44 -1205
rect -76 -1236 -44 -1235
rect -76 -1285 -44 -1284
rect -76 -1315 -75 -1285
rect -75 -1315 -45 -1285
rect -45 -1315 -44 -1285
rect -76 -1316 -44 -1315
rect -76 -1365 -44 -1364
rect -76 -1395 -75 -1365
rect -75 -1395 -45 -1365
rect -45 -1395 -44 -1365
rect -76 -1396 -44 -1395
rect -76 -1445 -44 -1444
rect -76 -1475 -75 -1445
rect -75 -1475 -45 -1445
rect -45 -1475 -44 -1445
rect -76 -1476 -44 -1475
rect -76 -1525 -44 -1524
rect -76 -1555 -75 -1525
rect -75 -1555 -45 -1525
rect -45 -1555 -44 -1525
rect -76 -1556 -44 -1555
rect -76 -1636 -44 -1604
rect -76 -1716 -44 -1684
rect -76 -1765 -44 -1764
rect -76 -1795 -75 -1765
rect -75 -1795 -45 -1765
rect -45 -1795 -44 -1765
rect -76 -1796 -44 -1795
rect -76 -1845 -44 -1844
rect -76 -1875 -75 -1845
rect -75 -1875 -45 -1845
rect -45 -1875 -44 -1845
rect -76 -1876 -44 -1875
rect -76 -1956 -44 -1924
rect -76 -2005 -44 -2004
rect -76 -2035 -75 -2005
rect -75 -2035 -45 -2005
rect -45 -2035 -44 -2005
rect -76 -2036 -44 -2035
rect -76 -2116 -44 -2084
rect -76 -2165 -44 -2164
rect -76 -2195 -75 -2165
rect -75 -2195 -45 -2165
rect -45 -2195 -44 -2165
rect -76 -2196 -44 -2195
rect -76 -2276 -44 -2244
rect -76 -2325 -44 -2324
rect -76 -2355 -75 -2325
rect -75 -2355 -45 -2325
rect -45 -2355 -44 -2325
rect -76 -2356 -44 -2355
rect -76 -2405 -44 -2404
rect -76 -2435 -75 -2405
rect -75 -2435 -45 -2405
rect -45 -2435 -44 -2405
rect -76 -2436 -44 -2435
rect -76 -2485 -44 -2484
rect -76 -2515 -75 -2485
rect -75 -2515 -45 -2485
rect -45 -2515 -44 -2485
rect -76 -2516 -44 -2515
rect -76 -2565 -44 -2564
rect -76 -2595 -75 -2565
rect -75 -2595 -45 -2565
rect -45 -2595 -44 -2565
rect -76 -2596 -44 -2595
rect -76 -2645 -44 -2644
rect -76 -2675 -75 -2645
rect -75 -2675 -45 -2645
rect -45 -2675 -44 -2645
rect -76 -2676 -44 -2675
rect -76 -2725 -44 -2724
rect -76 -2755 -75 -2725
rect -75 -2755 -45 -2725
rect -45 -2755 -44 -2725
rect -76 -2756 -44 -2755
rect -76 -2836 -44 -2804
rect -76 -2885 -44 -2884
rect -76 -2915 -75 -2885
rect -75 -2915 -45 -2885
rect -45 -2915 -44 -2885
rect -76 -2916 -44 -2915
rect -76 -2996 -44 -2964
rect -76 -3045 -44 -3044
rect -76 -3075 -75 -3045
rect -75 -3075 -45 -3045
rect -45 -3075 -44 -3045
rect -76 -3076 -44 -3075
rect -76 -3156 -44 -3124
rect -76 -3205 -44 -3204
rect -76 -3235 -75 -3205
rect -75 -3235 -45 -3205
rect -45 -3235 -44 -3205
rect -76 -3236 -44 -3235
rect -76 -3285 -44 -3284
rect -76 -3315 -75 -3285
rect -75 -3315 -45 -3285
rect -45 -3315 -44 -3285
rect -76 -3316 -44 -3315
rect -76 -3396 -44 -3364
rect -76 -3476 -44 -3444
rect -76 -3525 -44 -3524
rect -76 -3555 -75 -3525
rect -75 -3555 -45 -3525
rect -45 -3555 -44 -3525
rect -76 -3556 -44 -3555
rect -76 -3605 -44 -3604
rect -76 -3635 -75 -3605
rect -75 -3635 -45 -3605
rect -45 -3635 -44 -3605
rect -76 -3636 -44 -3635
rect -76 -3685 -44 -3684
rect -76 -3715 -75 -3685
rect -75 -3715 -45 -3685
rect -45 -3715 -44 -3685
rect -76 -3716 -44 -3715
rect 4 1035 36 1036
rect 4 1005 5 1035
rect 5 1005 35 1035
rect 35 1005 36 1035
rect 4 1004 36 1005
rect 4 955 36 956
rect 4 925 5 955
rect 5 925 35 955
rect 35 925 36 955
rect 4 924 36 925
rect 4 875 36 876
rect 4 845 5 875
rect 5 845 35 875
rect 35 845 36 875
rect 4 844 36 845
rect 4 764 36 796
rect 4 684 36 716
rect 4 635 36 636
rect 4 605 5 635
rect 5 605 35 635
rect 35 605 36 635
rect 4 604 36 605
rect 4 555 36 556
rect 4 525 5 555
rect 5 525 35 555
rect 35 525 36 555
rect 4 524 36 525
rect 4 444 36 476
rect 4 395 36 396
rect 4 365 5 395
rect 5 365 35 395
rect 35 365 36 395
rect 4 364 36 365
rect 4 284 36 316
rect 4 235 36 236
rect 4 205 5 235
rect 5 205 35 235
rect 35 205 36 235
rect 4 204 36 205
rect 4 124 36 156
rect 4 75 36 76
rect 4 45 5 75
rect 5 45 35 75
rect 35 45 36 75
rect 4 44 36 45
rect 4 -5 36 -4
rect 4 -35 5 -5
rect 5 -35 35 -5
rect 35 -35 36 -5
rect 4 -36 36 -35
rect 4 -85 36 -84
rect 4 -115 5 -85
rect 5 -115 35 -85
rect 35 -115 36 -85
rect 4 -116 36 -115
rect 4 -165 36 -164
rect 4 -195 5 -165
rect 5 -195 35 -165
rect 35 -195 36 -165
rect 4 -196 36 -195
rect 4 -245 36 -244
rect 4 -275 5 -245
rect 5 -275 35 -245
rect 35 -275 36 -245
rect 4 -276 36 -275
rect 4 -325 36 -324
rect 4 -355 5 -325
rect 5 -355 35 -325
rect 35 -355 36 -325
rect 4 -356 36 -355
rect 4 -436 36 -404
rect 4 -485 36 -484
rect 4 -515 5 -485
rect 5 -515 35 -485
rect 35 -515 36 -485
rect 4 -516 36 -515
rect 4 -596 36 -564
rect 4 -645 36 -644
rect 4 -675 5 -645
rect 5 -675 35 -645
rect 35 -675 36 -645
rect 4 -676 36 -675
rect 4 -756 36 -724
rect 4 -805 36 -804
rect 4 -835 5 -805
rect 5 -835 35 -805
rect 35 -835 36 -805
rect 4 -836 36 -835
rect 4 -885 36 -884
rect 4 -915 5 -885
rect 5 -915 35 -885
rect 35 -915 36 -885
rect 4 -916 36 -915
rect 4 -996 36 -964
rect 4 -1076 36 -1044
rect 4 -1125 36 -1124
rect 4 -1155 5 -1125
rect 5 -1155 35 -1125
rect 35 -1155 36 -1125
rect 4 -1156 36 -1155
rect 4 -1205 36 -1204
rect 4 -1235 5 -1205
rect 5 -1235 35 -1205
rect 35 -1235 36 -1205
rect 4 -1236 36 -1235
rect 4 -1285 36 -1284
rect 4 -1315 5 -1285
rect 5 -1315 35 -1285
rect 35 -1315 36 -1285
rect 4 -1316 36 -1315
rect 4 -1365 36 -1364
rect 4 -1395 5 -1365
rect 5 -1395 35 -1365
rect 35 -1395 36 -1365
rect 4 -1396 36 -1395
rect 4 -1445 36 -1444
rect 4 -1475 5 -1445
rect 5 -1475 35 -1445
rect 35 -1475 36 -1445
rect 4 -1476 36 -1475
rect 4 -1525 36 -1524
rect 4 -1555 5 -1525
rect 5 -1555 35 -1525
rect 35 -1555 36 -1525
rect 4 -1556 36 -1555
rect 4 -1636 36 -1604
rect 4 -1716 36 -1684
rect 4 -1765 36 -1764
rect 4 -1795 5 -1765
rect 5 -1795 35 -1765
rect 35 -1795 36 -1765
rect 4 -1796 36 -1795
rect 4 -1845 36 -1844
rect 4 -1875 5 -1845
rect 5 -1875 35 -1845
rect 35 -1875 36 -1845
rect 4 -1876 36 -1875
rect 4 -1956 36 -1924
rect 4 -2005 36 -2004
rect 4 -2035 5 -2005
rect 5 -2035 35 -2005
rect 35 -2035 36 -2005
rect 4 -2036 36 -2035
rect 4 -2116 36 -2084
rect 4 -2165 36 -2164
rect 4 -2195 5 -2165
rect 5 -2195 35 -2165
rect 35 -2195 36 -2165
rect 4 -2196 36 -2195
rect 4 -2276 36 -2244
rect 4 -2325 36 -2324
rect 4 -2355 5 -2325
rect 5 -2355 35 -2325
rect 35 -2355 36 -2325
rect 4 -2356 36 -2355
rect 4 -2405 36 -2404
rect 4 -2435 5 -2405
rect 5 -2435 35 -2405
rect 35 -2435 36 -2405
rect 4 -2436 36 -2435
rect 4 -2485 36 -2484
rect 4 -2515 5 -2485
rect 5 -2515 35 -2485
rect 35 -2515 36 -2485
rect 4 -2516 36 -2515
rect 4 -2565 36 -2564
rect 4 -2595 5 -2565
rect 5 -2595 35 -2565
rect 35 -2595 36 -2565
rect 4 -2596 36 -2595
rect 4 -2645 36 -2644
rect 4 -2675 5 -2645
rect 5 -2675 35 -2645
rect 35 -2675 36 -2645
rect 4 -2676 36 -2675
rect 4 -2725 36 -2724
rect 4 -2755 5 -2725
rect 5 -2755 35 -2725
rect 35 -2755 36 -2725
rect 4 -2756 36 -2755
rect 4 -2836 36 -2804
rect 4 -2885 36 -2884
rect 4 -2915 5 -2885
rect 5 -2915 35 -2885
rect 35 -2915 36 -2885
rect 4 -2916 36 -2915
rect 4 -2996 36 -2964
rect 4 -3045 36 -3044
rect 4 -3075 5 -3045
rect 5 -3075 35 -3045
rect 35 -3075 36 -3045
rect 4 -3076 36 -3075
rect 4 -3156 36 -3124
rect 4 -3205 36 -3204
rect 4 -3235 5 -3205
rect 5 -3235 35 -3205
rect 35 -3235 36 -3205
rect 4 -3236 36 -3235
rect 4 -3285 36 -3284
rect 4 -3315 5 -3285
rect 5 -3315 35 -3285
rect 35 -3315 36 -3285
rect 4 -3316 36 -3315
rect 4 -3396 36 -3364
rect 4 -3476 36 -3444
rect 4 -3525 36 -3524
rect 4 -3555 5 -3525
rect 5 -3555 35 -3525
rect 35 -3555 36 -3525
rect 4 -3556 36 -3555
rect 4 -3605 36 -3604
rect 4 -3635 5 -3605
rect 5 -3635 35 -3605
rect 35 -3635 36 -3605
rect 4 -3636 36 -3635
rect 4 -3685 36 -3684
rect 4 -3715 5 -3685
rect 5 -3715 35 -3685
rect 35 -3715 36 -3685
rect 4 -3716 36 -3715
rect 84 1035 116 1036
rect 84 1005 85 1035
rect 85 1005 115 1035
rect 115 1005 116 1035
rect 84 1004 116 1005
rect 84 955 116 956
rect 84 925 85 955
rect 85 925 115 955
rect 115 925 116 955
rect 84 924 116 925
rect 84 875 116 876
rect 84 845 85 875
rect 85 845 115 875
rect 115 845 116 875
rect 84 844 116 845
rect 84 764 116 796
rect 84 684 116 716
rect 84 635 116 636
rect 84 605 85 635
rect 85 605 115 635
rect 115 605 116 635
rect 84 604 116 605
rect 84 555 116 556
rect 84 525 85 555
rect 85 525 115 555
rect 115 525 116 555
rect 84 524 116 525
rect 84 444 116 476
rect 84 395 116 396
rect 84 365 85 395
rect 85 365 115 395
rect 115 365 116 395
rect 84 364 116 365
rect 84 284 116 316
rect 84 235 116 236
rect 84 205 85 235
rect 85 205 115 235
rect 115 205 116 235
rect 84 204 116 205
rect 84 124 116 156
rect 84 75 116 76
rect 84 45 85 75
rect 85 45 115 75
rect 115 45 116 75
rect 84 44 116 45
rect 84 -5 116 -4
rect 84 -35 85 -5
rect 85 -35 115 -5
rect 115 -35 116 -5
rect 84 -36 116 -35
rect 84 -85 116 -84
rect 84 -115 85 -85
rect 85 -115 115 -85
rect 115 -115 116 -85
rect 84 -116 116 -115
rect 84 -165 116 -164
rect 84 -195 85 -165
rect 85 -195 115 -165
rect 115 -195 116 -165
rect 84 -196 116 -195
rect 84 -245 116 -244
rect 84 -275 85 -245
rect 85 -275 115 -245
rect 115 -275 116 -245
rect 84 -276 116 -275
rect 84 -325 116 -324
rect 84 -355 85 -325
rect 85 -355 115 -325
rect 115 -355 116 -325
rect 84 -356 116 -355
rect 84 -436 116 -404
rect 84 -485 116 -484
rect 84 -515 85 -485
rect 85 -515 115 -485
rect 115 -515 116 -485
rect 84 -516 116 -515
rect 84 -596 116 -564
rect 84 -645 116 -644
rect 84 -675 85 -645
rect 85 -675 115 -645
rect 115 -675 116 -645
rect 84 -676 116 -675
rect 84 -756 116 -724
rect 84 -805 116 -804
rect 84 -835 85 -805
rect 85 -835 115 -805
rect 115 -835 116 -805
rect 84 -836 116 -835
rect 84 -885 116 -884
rect 84 -915 85 -885
rect 85 -915 115 -885
rect 115 -915 116 -885
rect 84 -916 116 -915
rect 84 -996 116 -964
rect 84 -1076 116 -1044
rect 84 -1125 116 -1124
rect 84 -1155 85 -1125
rect 85 -1155 115 -1125
rect 115 -1155 116 -1125
rect 84 -1156 116 -1155
rect 84 -1205 116 -1204
rect 84 -1235 85 -1205
rect 85 -1235 115 -1205
rect 115 -1235 116 -1205
rect 84 -1236 116 -1235
rect 84 -1285 116 -1284
rect 84 -1315 85 -1285
rect 85 -1315 115 -1285
rect 115 -1315 116 -1285
rect 84 -1316 116 -1315
rect 84 -1365 116 -1364
rect 84 -1395 85 -1365
rect 85 -1395 115 -1365
rect 115 -1395 116 -1365
rect 84 -1396 116 -1395
rect 84 -1445 116 -1444
rect 84 -1475 85 -1445
rect 85 -1475 115 -1445
rect 115 -1475 116 -1445
rect 84 -1476 116 -1475
rect 84 -1525 116 -1524
rect 84 -1555 85 -1525
rect 85 -1555 115 -1525
rect 115 -1555 116 -1525
rect 84 -1556 116 -1555
rect 84 -1636 116 -1604
rect 84 -1716 116 -1684
rect 84 -1765 116 -1764
rect 84 -1795 85 -1765
rect 85 -1795 115 -1765
rect 115 -1795 116 -1765
rect 84 -1796 116 -1795
rect 84 -1845 116 -1844
rect 84 -1875 85 -1845
rect 85 -1875 115 -1845
rect 115 -1875 116 -1845
rect 84 -1876 116 -1875
rect 84 -1956 116 -1924
rect 84 -2005 116 -2004
rect 84 -2035 85 -2005
rect 85 -2035 115 -2005
rect 115 -2035 116 -2005
rect 84 -2036 116 -2035
rect 84 -2116 116 -2084
rect 84 -2165 116 -2164
rect 84 -2195 85 -2165
rect 85 -2195 115 -2165
rect 115 -2195 116 -2165
rect 84 -2196 116 -2195
rect 84 -2276 116 -2244
rect 84 -2325 116 -2324
rect 84 -2355 85 -2325
rect 85 -2355 115 -2325
rect 115 -2355 116 -2325
rect 84 -2356 116 -2355
rect 84 -2405 116 -2404
rect 84 -2435 85 -2405
rect 85 -2435 115 -2405
rect 115 -2435 116 -2405
rect 84 -2436 116 -2435
rect 84 -2485 116 -2484
rect 84 -2515 85 -2485
rect 85 -2515 115 -2485
rect 115 -2515 116 -2485
rect 84 -2516 116 -2515
rect 84 -2565 116 -2564
rect 84 -2595 85 -2565
rect 85 -2595 115 -2565
rect 115 -2595 116 -2565
rect 84 -2596 116 -2595
rect 84 -2645 116 -2644
rect 84 -2675 85 -2645
rect 85 -2675 115 -2645
rect 115 -2675 116 -2645
rect 84 -2676 116 -2675
rect 84 -2725 116 -2724
rect 84 -2755 85 -2725
rect 85 -2755 115 -2725
rect 115 -2755 116 -2725
rect 84 -2756 116 -2755
rect 84 -2836 116 -2804
rect 84 -2885 116 -2884
rect 84 -2915 85 -2885
rect 85 -2915 115 -2885
rect 115 -2915 116 -2885
rect 84 -2916 116 -2915
rect 84 -2996 116 -2964
rect 84 -3045 116 -3044
rect 84 -3075 85 -3045
rect 85 -3075 115 -3045
rect 115 -3075 116 -3045
rect 84 -3076 116 -3075
rect 84 -3156 116 -3124
rect 84 -3205 116 -3204
rect 84 -3235 85 -3205
rect 85 -3235 115 -3205
rect 115 -3235 116 -3205
rect 84 -3236 116 -3235
rect 84 -3285 116 -3284
rect 84 -3315 85 -3285
rect 85 -3315 115 -3285
rect 115 -3315 116 -3285
rect 84 -3316 116 -3315
rect 84 -3396 116 -3364
rect 84 -3476 116 -3444
rect 84 -3525 116 -3524
rect 84 -3555 85 -3525
rect 85 -3555 115 -3525
rect 115 -3555 116 -3525
rect 84 -3556 116 -3555
rect 84 -3605 116 -3604
rect 84 -3635 85 -3605
rect 85 -3635 115 -3605
rect 115 -3635 116 -3605
rect 84 -3636 116 -3635
rect 84 -3685 116 -3684
rect 84 -3715 85 -3685
rect 85 -3715 115 -3685
rect 115 -3715 116 -3685
rect 84 -3716 116 -3715
rect 164 1035 196 1036
rect 164 1005 165 1035
rect 165 1005 195 1035
rect 195 1005 196 1035
rect 164 1004 196 1005
rect 164 955 196 956
rect 164 925 165 955
rect 165 925 195 955
rect 195 925 196 955
rect 164 924 196 925
rect 164 875 196 876
rect 164 845 165 875
rect 165 845 195 875
rect 195 845 196 875
rect 164 844 196 845
rect 164 764 196 796
rect 164 684 196 716
rect 164 635 196 636
rect 164 605 165 635
rect 165 605 195 635
rect 195 605 196 635
rect 164 604 196 605
rect 164 555 196 556
rect 164 525 165 555
rect 165 525 195 555
rect 195 525 196 555
rect 164 524 196 525
rect 164 444 196 476
rect 164 395 196 396
rect 164 365 165 395
rect 165 365 195 395
rect 195 365 196 395
rect 164 364 196 365
rect 164 284 196 316
rect 164 235 196 236
rect 164 205 165 235
rect 165 205 195 235
rect 195 205 196 235
rect 164 204 196 205
rect 164 124 196 156
rect 164 75 196 76
rect 164 45 165 75
rect 165 45 195 75
rect 195 45 196 75
rect 164 44 196 45
rect 164 -5 196 -4
rect 164 -35 165 -5
rect 165 -35 195 -5
rect 195 -35 196 -5
rect 164 -36 196 -35
rect 164 -85 196 -84
rect 164 -115 165 -85
rect 165 -115 195 -85
rect 195 -115 196 -85
rect 164 -116 196 -115
rect 164 -165 196 -164
rect 164 -195 165 -165
rect 165 -195 195 -165
rect 195 -195 196 -165
rect 164 -196 196 -195
rect 164 -245 196 -244
rect 164 -275 165 -245
rect 165 -275 195 -245
rect 195 -275 196 -245
rect 164 -276 196 -275
rect 164 -325 196 -324
rect 164 -355 165 -325
rect 165 -355 195 -325
rect 195 -355 196 -325
rect 164 -356 196 -355
rect 164 -436 196 -404
rect 164 -485 196 -484
rect 164 -515 165 -485
rect 165 -515 195 -485
rect 195 -515 196 -485
rect 164 -516 196 -515
rect 164 -596 196 -564
rect 164 -645 196 -644
rect 164 -675 165 -645
rect 165 -675 195 -645
rect 195 -675 196 -645
rect 164 -676 196 -675
rect 164 -756 196 -724
rect 164 -805 196 -804
rect 164 -835 165 -805
rect 165 -835 195 -805
rect 195 -835 196 -805
rect 164 -836 196 -835
rect 164 -885 196 -884
rect 164 -915 165 -885
rect 165 -915 195 -885
rect 195 -915 196 -885
rect 164 -916 196 -915
rect 164 -996 196 -964
rect 164 -1076 196 -1044
rect 164 -1125 196 -1124
rect 164 -1155 165 -1125
rect 165 -1155 195 -1125
rect 195 -1155 196 -1125
rect 164 -1156 196 -1155
rect 164 -1205 196 -1204
rect 164 -1235 165 -1205
rect 165 -1235 195 -1205
rect 195 -1235 196 -1205
rect 164 -1236 196 -1235
rect 164 -1285 196 -1284
rect 164 -1315 165 -1285
rect 165 -1315 195 -1285
rect 195 -1315 196 -1285
rect 164 -1316 196 -1315
rect 164 -1365 196 -1364
rect 164 -1395 165 -1365
rect 165 -1395 195 -1365
rect 195 -1395 196 -1365
rect 164 -1396 196 -1395
rect 164 -1445 196 -1444
rect 164 -1475 165 -1445
rect 165 -1475 195 -1445
rect 195 -1475 196 -1445
rect 164 -1476 196 -1475
rect 164 -1525 196 -1524
rect 164 -1555 165 -1525
rect 165 -1555 195 -1525
rect 195 -1555 196 -1525
rect 164 -1556 196 -1555
rect 164 -1636 196 -1604
rect 164 -1716 196 -1684
rect 164 -1765 196 -1764
rect 164 -1795 165 -1765
rect 165 -1795 195 -1765
rect 195 -1795 196 -1765
rect 164 -1796 196 -1795
rect 164 -1845 196 -1844
rect 164 -1875 165 -1845
rect 165 -1875 195 -1845
rect 195 -1875 196 -1845
rect 164 -1876 196 -1875
rect 164 -1956 196 -1924
rect 164 -2005 196 -2004
rect 164 -2035 165 -2005
rect 165 -2035 195 -2005
rect 195 -2035 196 -2005
rect 164 -2036 196 -2035
rect 164 -2116 196 -2084
rect 164 -2165 196 -2164
rect 164 -2195 165 -2165
rect 165 -2195 195 -2165
rect 195 -2195 196 -2165
rect 164 -2196 196 -2195
rect 164 -2276 196 -2244
rect 164 -2325 196 -2324
rect 164 -2355 165 -2325
rect 165 -2355 195 -2325
rect 195 -2355 196 -2325
rect 164 -2356 196 -2355
rect 164 -2405 196 -2404
rect 164 -2435 165 -2405
rect 165 -2435 195 -2405
rect 195 -2435 196 -2405
rect 164 -2436 196 -2435
rect 164 -2485 196 -2484
rect 164 -2515 165 -2485
rect 165 -2515 195 -2485
rect 195 -2515 196 -2485
rect 164 -2516 196 -2515
rect 164 -2565 196 -2564
rect 164 -2595 165 -2565
rect 165 -2595 195 -2565
rect 195 -2595 196 -2565
rect 164 -2596 196 -2595
rect 164 -2645 196 -2644
rect 164 -2675 165 -2645
rect 165 -2675 195 -2645
rect 195 -2675 196 -2645
rect 164 -2676 196 -2675
rect 164 -2725 196 -2724
rect 164 -2755 165 -2725
rect 165 -2755 195 -2725
rect 195 -2755 196 -2725
rect 164 -2756 196 -2755
rect 164 -2836 196 -2804
rect 164 -2885 196 -2884
rect 164 -2915 165 -2885
rect 165 -2915 195 -2885
rect 195 -2915 196 -2885
rect 164 -2916 196 -2915
rect 164 -2996 196 -2964
rect 164 -3045 196 -3044
rect 164 -3075 165 -3045
rect 165 -3075 195 -3045
rect 195 -3075 196 -3045
rect 164 -3076 196 -3075
rect 164 -3156 196 -3124
rect 164 -3205 196 -3204
rect 164 -3235 165 -3205
rect 165 -3235 195 -3205
rect 195 -3235 196 -3205
rect 164 -3236 196 -3235
rect 164 -3285 196 -3284
rect 164 -3315 165 -3285
rect 165 -3315 195 -3285
rect 195 -3315 196 -3285
rect 164 -3316 196 -3315
rect 164 -3396 196 -3364
rect 164 -3476 196 -3444
rect 164 -3525 196 -3524
rect 164 -3555 165 -3525
rect 165 -3555 195 -3525
rect 195 -3555 196 -3525
rect 164 -3556 196 -3555
rect 164 -3605 196 -3604
rect 164 -3635 165 -3605
rect 165 -3635 195 -3605
rect 195 -3635 196 -3605
rect 164 -3636 196 -3635
rect 164 -3685 196 -3684
rect 164 -3715 165 -3685
rect 165 -3715 195 -3685
rect 195 -3715 196 -3685
rect 164 -3716 196 -3715
rect 244 1035 276 1036
rect 244 1005 245 1035
rect 245 1005 275 1035
rect 275 1005 276 1035
rect 244 1004 276 1005
rect 244 955 276 956
rect 244 925 245 955
rect 245 925 275 955
rect 275 925 276 955
rect 244 924 276 925
rect 244 875 276 876
rect 244 845 245 875
rect 245 845 275 875
rect 275 845 276 875
rect 244 844 276 845
rect 244 764 276 796
rect 244 684 276 716
rect 244 635 276 636
rect 244 605 245 635
rect 245 605 275 635
rect 275 605 276 635
rect 244 604 276 605
rect 244 555 276 556
rect 244 525 245 555
rect 245 525 275 555
rect 275 525 276 555
rect 244 524 276 525
rect 244 444 276 476
rect 244 395 276 396
rect 244 365 245 395
rect 245 365 275 395
rect 275 365 276 395
rect 244 364 276 365
rect 244 284 276 316
rect 244 235 276 236
rect 244 205 245 235
rect 245 205 275 235
rect 275 205 276 235
rect 244 204 276 205
rect 244 124 276 156
rect 244 75 276 76
rect 244 45 245 75
rect 245 45 275 75
rect 275 45 276 75
rect 244 44 276 45
rect 244 -5 276 -4
rect 244 -35 245 -5
rect 245 -35 275 -5
rect 275 -35 276 -5
rect 244 -36 276 -35
rect 244 -85 276 -84
rect 244 -115 245 -85
rect 245 -115 275 -85
rect 275 -115 276 -85
rect 244 -116 276 -115
rect 244 -165 276 -164
rect 244 -195 245 -165
rect 245 -195 275 -165
rect 275 -195 276 -165
rect 244 -196 276 -195
rect 244 -245 276 -244
rect 244 -275 245 -245
rect 245 -275 275 -245
rect 275 -275 276 -245
rect 244 -276 276 -275
rect 244 -325 276 -324
rect 244 -355 245 -325
rect 245 -355 275 -325
rect 275 -355 276 -325
rect 244 -356 276 -355
rect 244 -436 276 -404
rect 244 -485 276 -484
rect 244 -515 245 -485
rect 245 -515 275 -485
rect 275 -515 276 -485
rect 244 -516 276 -515
rect 244 -596 276 -564
rect 244 -645 276 -644
rect 244 -675 245 -645
rect 245 -675 275 -645
rect 275 -675 276 -645
rect 244 -676 276 -675
rect 244 -756 276 -724
rect 244 -805 276 -804
rect 244 -835 245 -805
rect 245 -835 275 -805
rect 275 -835 276 -805
rect 244 -836 276 -835
rect 244 -885 276 -884
rect 244 -915 245 -885
rect 245 -915 275 -885
rect 275 -915 276 -885
rect 244 -916 276 -915
rect 244 -996 276 -964
rect 244 -1076 276 -1044
rect 244 -1125 276 -1124
rect 244 -1155 245 -1125
rect 245 -1155 275 -1125
rect 275 -1155 276 -1125
rect 244 -1156 276 -1155
rect 244 -1205 276 -1204
rect 244 -1235 245 -1205
rect 245 -1235 275 -1205
rect 275 -1235 276 -1205
rect 244 -1236 276 -1235
rect 244 -1285 276 -1284
rect 244 -1315 245 -1285
rect 245 -1315 275 -1285
rect 275 -1315 276 -1285
rect 244 -1316 276 -1315
rect 244 -1365 276 -1364
rect 244 -1395 245 -1365
rect 245 -1395 275 -1365
rect 275 -1395 276 -1365
rect 244 -1396 276 -1395
rect 244 -1445 276 -1444
rect 244 -1475 245 -1445
rect 245 -1475 275 -1445
rect 275 -1475 276 -1445
rect 244 -1476 276 -1475
rect 244 -1525 276 -1524
rect 244 -1555 245 -1525
rect 245 -1555 275 -1525
rect 275 -1555 276 -1525
rect 244 -1556 276 -1555
rect 244 -1636 276 -1604
rect 244 -1716 276 -1684
rect 244 -1765 276 -1764
rect 244 -1795 245 -1765
rect 245 -1795 275 -1765
rect 275 -1795 276 -1765
rect 244 -1796 276 -1795
rect 244 -1845 276 -1844
rect 244 -1875 245 -1845
rect 245 -1875 275 -1845
rect 275 -1875 276 -1845
rect 244 -1876 276 -1875
rect 244 -1956 276 -1924
rect 244 -2005 276 -2004
rect 244 -2035 245 -2005
rect 245 -2035 275 -2005
rect 275 -2035 276 -2005
rect 244 -2036 276 -2035
rect 244 -2116 276 -2084
rect 244 -2165 276 -2164
rect 244 -2195 245 -2165
rect 245 -2195 275 -2165
rect 275 -2195 276 -2165
rect 244 -2196 276 -2195
rect 244 -2276 276 -2244
rect 244 -2325 276 -2324
rect 244 -2355 245 -2325
rect 245 -2355 275 -2325
rect 275 -2355 276 -2325
rect 244 -2356 276 -2355
rect 244 -2405 276 -2404
rect 244 -2435 245 -2405
rect 245 -2435 275 -2405
rect 275 -2435 276 -2405
rect 244 -2436 276 -2435
rect 244 -2485 276 -2484
rect 244 -2515 245 -2485
rect 245 -2515 275 -2485
rect 275 -2515 276 -2485
rect 244 -2516 276 -2515
rect 244 -2565 276 -2564
rect 244 -2595 245 -2565
rect 245 -2595 275 -2565
rect 275 -2595 276 -2565
rect 244 -2596 276 -2595
rect 244 -2645 276 -2644
rect 244 -2675 245 -2645
rect 245 -2675 275 -2645
rect 275 -2675 276 -2645
rect 244 -2676 276 -2675
rect 244 -2725 276 -2724
rect 244 -2755 245 -2725
rect 245 -2755 275 -2725
rect 275 -2755 276 -2725
rect 244 -2756 276 -2755
rect 244 -2836 276 -2804
rect 244 -2885 276 -2884
rect 244 -2915 245 -2885
rect 245 -2915 275 -2885
rect 275 -2915 276 -2885
rect 244 -2916 276 -2915
rect 244 -2996 276 -2964
rect 244 -3045 276 -3044
rect 244 -3075 245 -3045
rect 245 -3075 275 -3045
rect 275 -3075 276 -3045
rect 244 -3076 276 -3075
rect 244 -3156 276 -3124
rect 244 -3205 276 -3204
rect 244 -3235 245 -3205
rect 245 -3235 275 -3205
rect 275 -3235 276 -3205
rect 244 -3236 276 -3235
rect 244 -3285 276 -3284
rect 244 -3315 245 -3285
rect 245 -3315 275 -3285
rect 275 -3315 276 -3285
rect 244 -3316 276 -3315
rect 244 -3396 276 -3364
rect 244 -3476 276 -3444
rect 244 -3525 276 -3524
rect 244 -3555 245 -3525
rect 245 -3555 275 -3525
rect 275 -3555 276 -3525
rect 244 -3556 276 -3555
rect 244 -3605 276 -3604
rect 244 -3635 245 -3605
rect 245 -3635 275 -3605
rect 275 -3635 276 -3605
rect 244 -3636 276 -3635
rect 244 -3685 276 -3684
rect 244 -3715 245 -3685
rect 245 -3715 275 -3685
rect 275 -3715 276 -3685
rect 244 -3716 276 -3715
rect 324 1035 356 1036
rect 324 1005 325 1035
rect 325 1005 355 1035
rect 355 1005 356 1035
rect 324 1004 356 1005
rect 324 955 356 956
rect 324 925 325 955
rect 325 925 355 955
rect 355 925 356 955
rect 324 924 356 925
rect 324 875 356 876
rect 324 845 325 875
rect 325 845 355 875
rect 355 845 356 875
rect 324 844 356 845
rect 324 764 356 796
rect 324 684 356 716
rect 324 635 356 636
rect 324 605 325 635
rect 325 605 355 635
rect 355 605 356 635
rect 324 604 356 605
rect 324 555 356 556
rect 324 525 325 555
rect 325 525 355 555
rect 355 525 356 555
rect 324 524 356 525
rect 324 444 356 476
rect 324 395 356 396
rect 324 365 325 395
rect 325 365 355 395
rect 355 365 356 395
rect 324 364 356 365
rect 324 284 356 316
rect 324 235 356 236
rect 324 205 325 235
rect 325 205 355 235
rect 355 205 356 235
rect 324 204 356 205
rect 324 124 356 156
rect 324 75 356 76
rect 324 45 325 75
rect 325 45 355 75
rect 355 45 356 75
rect 324 44 356 45
rect 324 -5 356 -4
rect 324 -35 325 -5
rect 325 -35 355 -5
rect 355 -35 356 -5
rect 324 -36 356 -35
rect 324 -85 356 -84
rect 324 -115 325 -85
rect 325 -115 355 -85
rect 355 -115 356 -85
rect 324 -116 356 -115
rect 324 -165 356 -164
rect 324 -195 325 -165
rect 325 -195 355 -165
rect 355 -195 356 -165
rect 324 -196 356 -195
rect 324 -245 356 -244
rect 324 -275 325 -245
rect 325 -275 355 -245
rect 355 -275 356 -245
rect 324 -276 356 -275
rect 324 -325 356 -324
rect 324 -355 325 -325
rect 325 -355 355 -325
rect 355 -355 356 -325
rect 324 -356 356 -355
rect 324 -436 356 -404
rect 324 -485 356 -484
rect 324 -515 325 -485
rect 325 -515 355 -485
rect 355 -515 356 -485
rect 324 -516 356 -515
rect 324 -596 356 -564
rect 324 -645 356 -644
rect 324 -675 325 -645
rect 325 -675 355 -645
rect 355 -675 356 -645
rect 324 -676 356 -675
rect 324 -756 356 -724
rect 324 -805 356 -804
rect 324 -835 325 -805
rect 325 -835 355 -805
rect 355 -835 356 -805
rect 324 -836 356 -835
rect 324 -885 356 -884
rect 324 -915 325 -885
rect 325 -915 355 -885
rect 355 -915 356 -885
rect 324 -916 356 -915
rect 324 -996 356 -964
rect 324 -1076 356 -1044
rect 324 -1125 356 -1124
rect 324 -1155 325 -1125
rect 325 -1155 355 -1125
rect 355 -1155 356 -1125
rect 324 -1156 356 -1155
rect 324 -1205 356 -1204
rect 324 -1235 325 -1205
rect 325 -1235 355 -1205
rect 355 -1235 356 -1205
rect 324 -1236 356 -1235
rect 324 -1285 356 -1284
rect 324 -1315 325 -1285
rect 325 -1315 355 -1285
rect 355 -1315 356 -1285
rect 324 -1316 356 -1315
rect 324 -1365 356 -1364
rect 324 -1395 325 -1365
rect 325 -1395 355 -1365
rect 355 -1395 356 -1365
rect 324 -1396 356 -1395
rect 324 -1445 356 -1444
rect 324 -1475 325 -1445
rect 325 -1475 355 -1445
rect 355 -1475 356 -1445
rect 324 -1476 356 -1475
rect 324 -1525 356 -1524
rect 324 -1555 325 -1525
rect 325 -1555 355 -1525
rect 355 -1555 356 -1525
rect 324 -1556 356 -1555
rect 324 -1636 356 -1604
rect 324 -1716 356 -1684
rect 324 -1765 356 -1764
rect 324 -1795 325 -1765
rect 325 -1795 355 -1765
rect 355 -1795 356 -1765
rect 324 -1796 356 -1795
rect 324 -1845 356 -1844
rect 324 -1875 325 -1845
rect 325 -1875 355 -1845
rect 355 -1875 356 -1845
rect 324 -1876 356 -1875
rect 324 -1956 356 -1924
rect 324 -2005 356 -2004
rect 324 -2035 325 -2005
rect 325 -2035 355 -2005
rect 355 -2035 356 -2005
rect 324 -2036 356 -2035
rect 324 -2116 356 -2084
rect 324 -2165 356 -2164
rect 324 -2195 325 -2165
rect 325 -2195 355 -2165
rect 355 -2195 356 -2165
rect 324 -2196 356 -2195
rect 324 -2276 356 -2244
rect 324 -2325 356 -2324
rect 324 -2355 325 -2325
rect 325 -2355 355 -2325
rect 355 -2355 356 -2325
rect 324 -2356 356 -2355
rect 324 -2405 356 -2404
rect 324 -2435 325 -2405
rect 325 -2435 355 -2405
rect 355 -2435 356 -2405
rect 324 -2436 356 -2435
rect 324 -2485 356 -2484
rect 324 -2515 325 -2485
rect 325 -2515 355 -2485
rect 355 -2515 356 -2485
rect 324 -2516 356 -2515
rect 324 -2565 356 -2564
rect 324 -2595 325 -2565
rect 325 -2595 355 -2565
rect 355 -2595 356 -2565
rect 324 -2596 356 -2595
rect 324 -2645 356 -2644
rect 324 -2675 325 -2645
rect 325 -2675 355 -2645
rect 355 -2675 356 -2645
rect 324 -2676 356 -2675
rect 324 -2725 356 -2724
rect 324 -2755 325 -2725
rect 325 -2755 355 -2725
rect 355 -2755 356 -2725
rect 324 -2756 356 -2755
rect 324 -2836 356 -2804
rect 324 -2885 356 -2884
rect 324 -2915 325 -2885
rect 325 -2915 355 -2885
rect 355 -2915 356 -2885
rect 324 -2916 356 -2915
rect 324 -2996 356 -2964
rect 324 -3045 356 -3044
rect 324 -3075 325 -3045
rect 325 -3075 355 -3045
rect 355 -3075 356 -3045
rect 324 -3076 356 -3075
rect 324 -3156 356 -3124
rect 324 -3205 356 -3204
rect 324 -3235 325 -3205
rect 325 -3235 355 -3205
rect 355 -3235 356 -3205
rect 324 -3236 356 -3235
rect 324 -3285 356 -3284
rect 324 -3315 325 -3285
rect 325 -3315 355 -3285
rect 355 -3315 356 -3285
rect 324 -3316 356 -3315
rect 324 -3396 356 -3364
rect 324 -3476 356 -3444
rect 324 -3525 356 -3524
rect 324 -3555 325 -3525
rect 325 -3555 355 -3525
rect 355 -3555 356 -3525
rect 324 -3556 356 -3555
rect 324 -3605 356 -3604
rect 324 -3635 325 -3605
rect 325 -3635 355 -3605
rect 355 -3635 356 -3605
rect 324 -3636 356 -3635
rect 324 -3685 356 -3684
rect 324 -3715 325 -3685
rect 325 -3715 355 -3685
rect 355 -3715 356 -3685
rect 324 -3716 356 -3715
rect 404 1035 436 1036
rect 404 1005 405 1035
rect 405 1005 435 1035
rect 435 1005 436 1035
rect 404 1004 436 1005
rect 404 955 436 956
rect 404 925 405 955
rect 405 925 435 955
rect 435 925 436 955
rect 404 924 436 925
rect 404 875 436 876
rect 404 845 405 875
rect 405 845 435 875
rect 435 845 436 875
rect 404 844 436 845
rect 404 764 436 796
rect 404 684 436 716
rect 404 635 436 636
rect 404 605 405 635
rect 405 605 435 635
rect 435 605 436 635
rect 404 604 436 605
rect 404 555 436 556
rect 404 525 405 555
rect 405 525 435 555
rect 435 525 436 555
rect 404 524 436 525
rect 404 444 436 476
rect 404 395 436 396
rect 404 365 405 395
rect 405 365 435 395
rect 435 365 436 395
rect 404 364 436 365
rect 404 284 436 316
rect 404 235 436 236
rect 404 205 405 235
rect 405 205 435 235
rect 435 205 436 235
rect 404 204 436 205
rect 404 124 436 156
rect 404 75 436 76
rect 404 45 405 75
rect 405 45 435 75
rect 435 45 436 75
rect 404 44 436 45
rect 404 -5 436 -4
rect 404 -35 405 -5
rect 405 -35 435 -5
rect 435 -35 436 -5
rect 404 -36 436 -35
rect 404 -85 436 -84
rect 404 -115 405 -85
rect 405 -115 435 -85
rect 435 -115 436 -85
rect 404 -116 436 -115
rect 404 -165 436 -164
rect 404 -195 405 -165
rect 405 -195 435 -165
rect 435 -195 436 -165
rect 404 -196 436 -195
rect 404 -245 436 -244
rect 404 -275 405 -245
rect 405 -275 435 -245
rect 435 -275 436 -245
rect 404 -276 436 -275
rect 404 -325 436 -324
rect 404 -355 405 -325
rect 405 -355 435 -325
rect 435 -355 436 -325
rect 404 -356 436 -355
rect 404 -436 436 -404
rect 404 -485 436 -484
rect 404 -515 405 -485
rect 405 -515 435 -485
rect 435 -515 436 -485
rect 404 -516 436 -515
rect 404 -596 436 -564
rect 404 -645 436 -644
rect 404 -675 405 -645
rect 405 -675 435 -645
rect 435 -675 436 -645
rect 404 -676 436 -675
rect 404 -756 436 -724
rect 404 -805 436 -804
rect 404 -835 405 -805
rect 405 -835 435 -805
rect 435 -835 436 -805
rect 404 -836 436 -835
rect 404 -885 436 -884
rect 404 -915 405 -885
rect 405 -915 435 -885
rect 435 -915 436 -885
rect 404 -916 436 -915
rect 404 -996 436 -964
rect 404 -1076 436 -1044
rect 404 -1125 436 -1124
rect 404 -1155 405 -1125
rect 405 -1155 435 -1125
rect 435 -1155 436 -1125
rect 404 -1156 436 -1155
rect 404 -1205 436 -1204
rect 404 -1235 405 -1205
rect 405 -1235 435 -1205
rect 435 -1235 436 -1205
rect 404 -1236 436 -1235
rect 404 -1285 436 -1284
rect 404 -1315 405 -1285
rect 405 -1315 435 -1285
rect 435 -1315 436 -1285
rect 404 -1316 436 -1315
rect 404 -1365 436 -1364
rect 404 -1395 405 -1365
rect 405 -1395 435 -1365
rect 435 -1395 436 -1365
rect 404 -1396 436 -1395
rect 404 -1445 436 -1444
rect 404 -1475 405 -1445
rect 405 -1475 435 -1445
rect 435 -1475 436 -1445
rect 404 -1476 436 -1475
rect 404 -1525 436 -1524
rect 404 -1555 405 -1525
rect 405 -1555 435 -1525
rect 435 -1555 436 -1525
rect 404 -1556 436 -1555
rect 404 -1636 436 -1604
rect 404 -1716 436 -1684
rect 404 -1765 436 -1764
rect 404 -1795 405 -1765
rect 405 -1795 435 -1765
rect 435 -1795 436 -1765
rect 404 -1796 436 -1795
rect 404 -1845 436 -1844
rect 404 -1875 405 -1845
rect 405 -1875 435 -1845
rect 435 -1875 436 -1845
rect 404 -1876 436 -1875
rect 404 -1956 436 -1924
rect 404 -2005 436 -2004
rect 404 -2035 405 -2005
rect 405 -2035 435 -2005
rect 435 -2035 436 -2005
rect 404 -2036 436 -2035
rect 404 -2116 436 -2084
rect 404 -2165 436 -2164
rect 404 -2195 405 -2165
rect 405 -2195 435 -2165
rect 435 -2195 436 -2165
rect 404 -2196 436 -2195
rect 404 -2276 436 -2244
rect 404 -2325 436 -2324
rect 404 -2355 405 -2325
rect 405 -2355 435 -2325
rect 435 -2355 436 -2325
rect 404 -2356 436 -2355
rect 404 -2405 436 -2404
rect 404 -2435 405 -2405
rect 405 -2435 435 -2405
rect 435 -2435 436 -2405
rect 404 -2436 436 -2435
rect 404 -2485 436 -2484
rect 404 -2515 405 -2485
rect 405 -2515 435 -2485
rect 435 -2515 436 -2485
rect 404 -2516 436 -2515
rect 404 -2565 436 -2564
rect 404 -2595 405 -2565
rect 405 -2595 435 -2565
rect 435 -2595 436 -2565
rect 404 -2596 436 -2595
rect 404 -2645 436 -2644
rect 404 -2675 405 -2645
rect 405 -2675 435 -2645
rect 435 -2675 436 -2645
rect 404 -2676 436 -2675
rect 404 -2725 436 -2724
rect 404 -2755 405 -2725
rect 405 -2755 435 -2725
rect 435 -2755 436 -2725
rect 404 -2756 436 -2755
rect 404 -2836 436 -2804
rect 404 -2885 436 -2884
rect 404 -2915 405 -2885
rect 405 -2915 435 -2885
rect 435 -2915 436 -2885
rect 404 -2916 436 -2915
rect 404 -2996 436 -2964
rect 404 -3045 436 -3044
rect 404 -3075 405 -3045
rect 405 -3075 435 -3045
rect 435 -3075 436 -3045
rect 404 -3076 436 -3075
rect 404 -3156 436 -3124
rect 404 -3205 436 -3204
rect 404 -3235 405 -3205
rect 405 -3235 435 -3205
rect 435 -3235 436 -3205
rect 404 -3236 436 -3235
rect 404 -3285 436 -3284
rect 404 -3315 405 -3285
rect 405 -3315 435 -3285
rect 435 -3315 436 -3285
rect 404 -3316 436 -3315
rect 404 -3396 436 -3364
rect 404 -3476 436 -3444
rect 404 -3525 436 -3524
rect 404 -3555 405 -3525
rect 405 -3555 435 -3525
rect 435 -3555 436 -3525
rect 404 -3556 436 -3555
rect 404 -3605 436 -3604
rect 404 -3635 405 -3605
rect 405 -3635 435 -3605
rect 435 -3635 436 -3605
rect 404 -3636 436 -3635
rect 404 -3685 436 -3684
rect 404 -3715 405 -3685
rect 405 -3715 435 -3685
rect 435 -3715 436 -3685
rect 404 -3716 436 -3715
rect 484 1035 516 1036
rect 484 1005 485 1035
rect 485 1005 515 1035
rect 515 1005 516 1035
rect 484 1004 516 1005
rect 484 955 516 956
rect 484 925 485 955
rect 485 925 515 955
rect 515 925 516 955
rect 484 924 516 925
rect 484 875 516 876
rect 484 845 485 875
rect 485 845 515 875
rect 515 845 516 875
rect 484 844 516 845
rect 484 764 516 796
rect 484 684 516 716
rect 484 635 516 636
rect 484 605 485 635
rect 485 605 515 635
rect 515 605 516 635
rect 484 604 516 605
rect 484 555 516 556
rect 484 525 485 555
rect 485 525 515 555
rect 515 525 516 555
rect 484 524 516 525
rect 484 444 516 476
rect 484 395 516 396
rect 484 365 485 395
rect 485 365 515 395
rect 515 365 516 395
rect 484 364 516 365
rect 484 284 516 316
rect 484 235 516 236
rect 484 205 485 235
rect 485 205 515 235
rect 515 205 516 235
rect 484 204 516 205
rect 484 124 516 156
rect 484 75 516 76
rect 484 45 485 75
rect 485 45 515 75
rect 515 45 516 75
rect 484 44 516 45
rect 484 -5 516 -4
rect 484 -35 485 -5
rect 485 -35 515 -5
rect 515 -35 516 -5
rect 484 -36 516 -35
rect 484 -85 516 -84
rect 484 -115 485 -85
rect 485 -115 515 -85
rect 515 -115 516 -85
rect 484 -116 516 -115
rect 484 -165 516 -164
rect 484 -195 485 -165
rect 485 -195 515 -165
rect 515 -195 516 -165
rect 484 -196 516 -195
rect 484 -245 516 -244
rect 484 -275 485 -245
rect 485 -275 515 -245
rect 515 -275 516 -245
rect 484 -276 516 -275
rect 484 -325 516 -324
rect 484 -355 485 -325
rect 485 -355 515 -325
rect 515 -355 516 -325
rect 484 -356 516 -355
rect 484 -436 516 -404
rect 484 -485 516 -484
rect 484 -515 485 -485
rect 485 -515 515 -485
rect 515 -515 516 -485
rect 484 -516 516 -515
rect 484 -596 516 -564
rect 484 -645 516 -644
rect 484 -675 485 -645
rect 485 -675 515 -645
rect 515 -675 516 -645
rect 484 -676 516 -675
rect 484 -756 516 -724
rect 484 -805 516 -804
rect 484 -835 485 -805
rect 485 -835 515 -805
rect 515 -835 516 -805
rect 484 -836 516 -835
rect 484 -885 516 -884
rect 484 -915 485 -885
rect 485 -915 515 -885
rect 515 -915 516 -885
rect 484 -916 516 -915
rect 484 -996 516 -964
rect 484 -1076 516 -1044
rect 484 -1125 516 -1124
rect 484 -1155 485 -1125
rect 485 -1155 515 -1125
rect 515 -1155 516 -1125
rect 484 -1156 516 -1155
rect 484 -1205 516 -1204
rect 484 -1235 485 -1205
rect 485 -1235 515 -1205
rect 515 -1235 516 -1205
rect 484 -1236 516 -1235
rect 484 -1285 516 -1284
rect 484 -1315 485 -1285
rect 485 -1315 515 -1285
rect 515 -1315 516 -1285
rect 484 -1316 516 -1315
rect 484 -1365 516 -1364
rect 484 -1395 485 -1365
rect 485 -1395 515 -1365
rect 515 -1395 516 -1365
rect 484 -1396 516 -1395
rect 484 -1445 516 -1444
rect 484 -1475 485 -1445
rect 485 -1475 515 -1445
rect 515 -1475 516 -1445
rect 484 -1476 516 -1475
rect 484 -1525 516 -1524
rect 484 -1555 485 -1525
rect 485 -1555 515 -1525
rect 515 -1555 516 -1525
rect 484 -1556 516 -1555
rect 484 -1636 516 -1604
rect 484 -1716 516 -1684
rect 484 -1765 516 -1764
rect 484 -1795 485 -1765
rect 485 -1795 515 -1765
rect 515 -1795 516 -1765
rect 484 -1796 516 -1795
rect 484 -1845 516 -1844
rect 484 -1875 485 -1845
rect 485 -1875 515 -1845
rect 515 -1875 516 -1845
rect 484 -1876 516 -1875
rect 484 -1956 516 -1924
rect 484 -2005 516 -2004
rect 484 -2035 485 -2005
rect 485 -2035 515 -2005
rect 515 -2035 516 -2005
rect 484 -2036 516 -2035
rect 484 -2116 516 -2084
rect 484 -2165 516 -2164
rect 484 -2195 485 -2165
rect 485 -2195 515 -2165
rect 515 -2195 516 -2165
rect 484 -2196 516 -2195
rect 484 -2276 516 -2244
rect 484 -2325 516 -2324
rect 484 -2355 485 -2325
rect 485 -2355 515 -2325
rect 515 -2355 516 -2325
rect 484 -2356 516 -2355
rect 484 -2405 516 -2404
rect 484 -2435 485 -2405
rect 485 -2435 515 -2405
rect 515 -2435 516 -2405
rect 484 -2436 516 -2435
rect 484 -2485 516 -2484
rect 484 -2515 485 -2485
rect 485 -2515 515 -2485
rect 515 -2515 516 -2485
rect 484 -2516 516 -2515
rect 484 -2565 516 -2564
rect 484 -2595 485 -2565
rect 485 -2595 515 -2565
rect 515 -2595 516 -2565
rect 484 -2596 516 -2595
rect 484 -2645 516 -2644
rect 484 -2675 485 -2645
rect 485 -2675 515 -2645
rect 515 -2675 516 -2645
rect 484 -2676 516 -2675
rect 484 -2725 516 -2724
rect 484 -2755 485 -2725
rect 485 -2755 515 -2725
rect 515 -2755 516 -2725
rect 484 -2756 516 -2755
rect 484 -2836 516 -2804
rect 484 -2885 516 -2884
rect 484 -2915 485 -2885
rect 485 -2915 515 -2885
rect 515 -2915 516 -2885
rect 484 -2916 516 -2915
rect 484 -2996 516 -2964
rect 484 -3045 516 -3044
rect 484 -3075 485 -3045
rect 485 -3075 515 -3045
rect 515 -3075 516 -3045
rect 484 -3076 516 -3075
rect 484 -3156 516 -3124
rect 484 -3205 516 -3204
rect 484 -3235 485 -3205
rect 485 -3235 515 -3205
rect 515 -3235 516 -3205
rect 484 -3236 516 -3235
rect 484 -3285 516 -3284
rect 484 -3315 485 -3285
rect 485 -3315 515 -3285
rect 515 -3315 516 -3285
rect 484 -3316 516 -3315
rect 484 -3396 516 -3364
rect 484 -3476 516 -3444
rect 484 -3525 516 -3524
rect 484 -3555 485 -3525
rect 485 -3555 515 -3525
rect 515 -3555 516 -3525
rect 484 -3556 516 -3555
rect 484 -3605 516 -3604
rect 484 -3635 485 -3605
rect 485 -3635 515 -3605
rect 515 -3635 516 -3605
rect 484 -3636 516 -3635
rect 484 -3685 516 -3684
rect 484 -3715 485 -3685
rect 485 -3715 515 -3685
rect 515 -3715 516 -3685
rect 484 -3716 516 -3715
rect 564 1035 596 1036
rect 564 1005 565 1035
rect 565 1005 595 1035
rect 595 1005 596 1035
rect 564 1004 596 1005
rect 564 955 596 956
rect 564 925 565 955
rect 565 925 595 955
rect 595 925 596 955
rect 564 924 596 925
rect 564 875 596 876
rect 564 845 565 875
rect 565 845 595 875
rect 595 845 596 875
rect 564 844 596 845
rect 564 764 596 796
rect 564 684 596 716
rect 564 635 596 636
rect 564 605 565 635
rect 565 605 595 635
rect 595 605 596 635
rect 564 604 596 605
rect 564 555 596 556
rect 564 525 565 555
rect 565 525 595 555
rect 595 525 596 555
rect 564 524 596 525
rect 564 444 596 476
rect 564 395 596 396
rect 564 365 565 395
rect 565 365 595 395
rect 595 365 596 395
rect 564 364 596 365
rect 564 284 596 316
rect 564 235 596 236
rect 564 205 565 235
rect 565 205 595 235
rect 595 205 596 235
rect 564 204 596 205
rect 564 124 596 156
rect 564 75 596 76
rect 564 45 565 75
rect 565 45 595 75
rect 595 45 596 75
rect 564 44 596 45
rect 564 -5 596 -4
rect 564 -35 565 -5
rect 565 -35 595 -5
rect 595 -35 596 -5
rect 564 -36 596 -35
rect 564 -85 596 -84
rect 564 -115 565 -85
rect 565 -115 595 -85
rect 595 -115 596 -85
rect 564 -116 596 -115
rect 564 -165 596 -164
rect 564 -195 565 -165
rect 565 -195 595 -165
rect 595 -195 596 -165
rect 564 -196 596 -195
rect 564 -245 596 -244
rect 564 -275 565 -245
rect 565 -275 595 -245
rect 595 -275 596 -245
rect 564 -276 596 -275
rect 564 -325 596 -324
rect 564 -355 565 -325
rect 565 -355 595 -325
rect 595 -355 596 -325
rect 564 -356 596 -355
rect 564 -436 596 -404
rect 564 -485 596 -484
rect 564 -515 565 -485
rect 565 -515 595 -485
rect 595 -515 596 -485
rect 564 -516 596 -515
rect 564 -596 596 -564
rect 564 -645 596 -644
rect 564 -675 565 -645
rect 565 -675 595 -645
rect 595 -675 596 -645
rect 564 -676 596 -675
rect 564 -756 596 -724
rect 564 -805 596 -804
rect 564 -835 565 -805
rect 565 -835 595 -805
rect 595 -835 596 -805
rect 564 -836 596 -835
rect 564 -885 596 -884
rect 564 -915 565 -885
rect 565 -915 595 -885
rect 595 -915 596 -885
rect 564 -916 596 -915
rect 564 -996 596 -964
rect 564 -1076 596 -1044
rect 564 -1125 596 -1124
rect 564 -1155 565 -1125
rect 565 -1155 595 -1125
rect 595 -1155 596 -1125
rect 564 -1156 596 -1155
rect 564 -1205 596 -1204
rect 564 -1235 565 -1205
rect 565 -1235 595 -1205
rect 595 -1235 596 -1205
rect 564 -1236 596 -1235
rect 564 -1285 596 -1284
rect 564 -1315 565 -1285
rect 565 -1315 595 -1285
rect 595 -1315 596 -1285
rect 564 -1316 596 -1315
rect 564 -1365 596 -1364
rect 564 -1395 565 -1365
rect 565 -1395 595 -1365
rect 595 -1395 596 -1365
rect 564 -1396 596 -1395
rect 564 -1445 596 -1444
rect 564 -1475 565 -1445
rect 565 -1475 595 -1445
rect 595 -1475 596 -1445
rect 564 -1476 596 -1475
rect 564 -1525 596 -1524
rect 564 -1555 565 -1525
rect 565 -1555 595 -1525
rect 595 -1555 596 -1525
rect 564 -1556 596 -1555
rect 564 -1636 596 -1604
rect 564 -1716 596 -1684
rect 564 -1765 596 -1764
rect 564 -1795 565 -1765
rect 565 -1795 595 -1765
rect 595 -1795 596 -1765
rect 564 -1796 596 -1795
rect 564 -1845 596 -1844
rect 564 -1875 565 -1845
rect 565 -1875 595 -1845
rect 595 -1875 596 -1845
rect 564 -1876 596 -1875
rect 564 -1956 596 -1924
rect 564 -2005 596 -2004
rect 564 -2035 565 -2005
rect 565 -2035 595 -2005
rect 595 -2035 596 -2005
rect 564 -2036 596 -2035
rect 564 -2116 596 -2084
rect 564 -2165 596 -2164
rect 564 -2195 565 -2165
rect 565 -2195 595 -2165
rect 595 -2195 596 -2165
rect 564 -2196 596 -2195
rect 564 -2276 596 -2244
rect 564 -2325 596 -2324
rect 564 -2355 565 -2325
rect 565 -2355 595 -2325
rect 595 -2355 596 -2325
rect 564 -2356 596 -2355
rect 564 -2405 596 -2404
rect 564 -2435 565 -2405
rect 565 -2435 595 -2405
rect 595 -2435 596 -2405
rect 564 -2436 596 -2435
rect 564 -2485 596 -2484
rect 564 -2515 565 -2485
rect 565 -2515 595 -2485
rect 595 -2515 596 -2485
rect 564 -2516 596 -2515
rect 564 -2565 596 -2564
rect 564 -2595 565 -2565
rect 565 -2595 595 -2565
rect 595 -2595 596 -2565
rect 564 -2596 596 -2595
rect 564 -2645 596 -2644
rect 564 -2675 565 -2645
rect 565 -2675 595 -2645
rect 595 -2675 596 -2645
rect 564 -2676 596 -2675
rect 564 -2725 596 -2724
rect 564 -2755 565 -2725
rect 565 -2755 595 -2725
rect 595 -2755 596 -2725
rect 564 -2756 596 -2755
rect 564 -2836 596 -2804
rect 564 -2885 596 -2884
rect 564 -2915 565 -2885
rect 565 -2915 595 -2885
rect 595 -2915 596 -2885
rect 564 -2916 596 -2915
rect 564 -2996 596 -2964
rect 564 -3045 596 -3044
rect 564 -3075 565 -3045
rect 565 -3075 595 -3045
rect 595 -3075 596 -3045
rect 564 -3076 596 -3075
rect 564 -3156 596 -3124
rect 564 -3205 596 -3204
rect 564 -3235 565 -3205
rect 565 -3235 595 -3205
rect 595 -3235 596 -3205
rect 564 -3236 596 -3235
rect 564 -3285 596 -3284
rect 564 -3315 565 -3285
rect 565 -3315 595 -3285
rect 595 -3315 596 -3285
rect 564 -3316 596 -3315
rect 564 -3396 596 -3364
rect 564 -3476 596 -3444
rect 564 -3525 596 -3524
rect 564 -3555 565 -3525
rect 565 -3555 595 -3525
rect 595 -3555 596 -3525
rect 564 -3556 596 -3555
rect 564 -3605 596 -3604
rect 564 -3635 565 -3605
rect 565 -3635 595 -3605
rect 595 -3635 596 -3605
rect 564 -3636 596 -3635
rect 564 -3685 596 -3684
rect 564 -3715 565 -3685
rect 565 -3715 595 -3685
rect 595 -3715 596 -3685
rect 564 -3716 596 -3715
rect 644 1035 676 1036
rect 644 1005 645 1035
rect 645 1005 675 1035
rect 675 1005 676 1035
rect 644 1004 676 1005
rect 644 955 676 956
rect 644 925 645 955
rect 645 925 675 955
rect 675 925 676 955
rect 644 924 676 925
rect 644 875 676 876
rect 644 845 645 875
rect 645 845 675 875
rect 675 845 676 875
rect 644 844 676 845
rect 644 764 676 796
rect 644 684 676 716
rect 644 635 676 636
rect 644 605 645 635
rect 645 605 675 635
rect 675 605 676 635
rect 644 604 676 605
rect 644 555 676 556
rect 644 525 645 555
rect 645 525 675 555
rect 675 525 676 555
rect 644 524 676 525
rect 644 444 676 476
rect 644 395 676 396
rect 644 365 645 395
rect 645 365 675 395
rect 675 365 676 395
rect 644 364 676 365
rect 644 284 676 316
rect 644 235 676 236
rect 644 205 645 235
rect 645 205 675 235
rect 675 205 676 235
rect 644 204 676 205
rect 644 124 676 156
rect 644 75 676 76
rect 644 45 645 75
rect 645 45 675 75
rect 675 45 676 75
rect 644 44 676 45
rect 644 -5 676 -4
rect 644 -35 645 -5
rect 645 -35 675 -5
rect 675 -35 676 -5
rect 644 -36 676 -35
rect 644 -85 676 -84
rect 644 -115 645 -85
rect 645 -115 675 -85
rect 675 -115 676 -85
rect 644 -116 676 -115
rect 644 -165 676 -164
rect 644 -195 645 -165
rect 645 -195 675 -165
rect 675 -195 676 -165
rect 644 -196 676 -195
rect 644 -245 676 -244
rect 644 -275 645 -245
rect 645 -275 675 -245
rect 675 -275 676 -245
rect 644 -276 676 -275
rect 644 -325 676 -324
rect 644 -355 645 -325
rect 645 -355 675 -325
rect 675 -355 676 -325
rect 644 -356 676 -355
rect 644 -436 676 -404
rect 644 -485 676 -484
rect 644 -515 645 -485
rect 645 -515 675 -485
rect 675 -515 676 -485
rect 644 -516 676 -515
rect 644 -596 676 -564
rect 644 -645 676 -644
rect 644 -675 645 -645
rect 645 -675 675 -645
rect 675 -675 676 -645
rect 644 -676 676 -675
rect 644 -756 676 -724
rect 644 -805 676 -804
rect 644 -835 645 -805
rect 645 -835 675 -805
rect 675 -835 676 -805
rect 644 -836 676 -835
rect 644 -885 676 -884
rect 644 -915 645 -885
rect 645 -915 675 -885
rect 675 -915 676 -885
rect 644 -916 676 -915
rect 644 -996 676 -964
rect 644 -1076 676 -1044
rect 644 -1125 676 -1124
rect 644 -1155 645 -1125
rect 645 -1155 675 -1125
rect 675 -1155 676 -1125
rect 644 -1156 676 -1155
rect 644 -1205 676 -1204
rect 644 -1235 645 -1205
rect 645 -1235 675 -1205
rect 675 -1235 676 -1205
rect 644 -1236 676 -1235
rect 644 -1285 676 -1284
rect 644 -1315 645 -1285
rect 645 -1315 675 -1285
rect 675 -1315 676 -1285
rect 644 -1316 676 -1315
rect 644 -1365 676 -1364
rect 644 -1395 645 -1365
rect 645 -1395 675 -1365
rect 675 -1395 676 -1365
rect 644 -1396 676 -1395
rect 644 -1445 676 -1444
rect 644 -1475 645 -1445
rect 645 -1475 675 -1445
rect 675 -1475 676 -1445
rect 644 -1476 676 -1475
rect 644 -1525 676 -1524
rect 644 -1555 645 -1525
rect 645 -1555 675 -1525
rect 675 -1555 676 -1525
rect 644 -1556 676 -1555
rect 644 -1636 676 -1604
rect 644 -1716 676 -1684
rect 644 -1765 676 -1764
rect 644 -1795 645 -1765
rect 645 -1795 675 -1765
rect 675 -1795 676 -1765
rect 644 -1796 676 -1795
rect 644 -1845 676 -1844
rect 644 -1875 645 -1845
rect 645 -1875 675 -1845
rect 675 -1875 676 -1845
rect 644 -1876 676 -1875
rect 644 -1956 676 -1924
rect 644 -2005 676 -2004
rect 644 -2035 645 -2005
rect 645 -2035 675 -2005
rect 675 -2035 676 -2005
rect 644 -2036 676 -2035
rect 644 -2116 676 -2084
rect 644 -2165 676 -2164
rect 644 -2195 645 -2165
rect 645 -2195 675 -2165
rect 675 -2195 676 -2165
rect 644 -2196 676 -2195
rect 644 -2276 676 -2244
rect 644 -2325 676 -2324
rect 644 -2355 645 -2325
rect 645 -2355 675 -2325
rect 675 -2355 676 -2325
rect 644 -2356 676 -2355
rect 644 -2405 676 -2404
rect 644 -2435 645 -2405
rect 645 -2435 675 -2405
rect 675 -2435 676 -2405
rect 644 -2436 676 -2435
rect 644 -2485 676 -2484
rect 644 -2515 645 -2485
rect 645 -2515 675 -2485
rect 675 -2515 676 -2485
rect 644 -2516 676 -2515
rect 644 -2565 676 -2564
rect 644 -2595 645 -2565
rect 645 -2595 675 -2565
rect 675 -2595 676 -2565
rect 644 -2596 676 -2595
rect 644 -2645 676 -2644
rect 644 -2675 645 -2645
rect 645 -2675 675 -2645
rect 675 -2675 676 -2645
rect 644 -2676 676 -2675
rect 644 -2725 676 -2724
rect 644 -2755 645 -2725
rect 645 -2755 675 -2725
rect 675 -2755 676 -2725
rect 644 -2756 676 -2755
rect 644 -2836 676 -2804
rect 644 -2885 676 -2884
rect 644 -2915 645 -2885
rect 645 -2915 675 -2885
rect 675 -2915 676 -2885
rect 644 -2916 676 -2915
rect 644 -2996 676 -2964
rect 644 -3045 676 -3044
rect 644 -3075 645 -3045
rect 645 -3075 675 -3045
rect 675 -3075 676 -3045
rect 644 -3076 676 -3075
rect 644 -3156 676 -3124
rect 644 -3205 676 -3204
rect 644 -3235 645 -3205
rect 645 -3235 675 -3205
rect 675 -3235 676 -3205
rect 644 -3236 676 -3235
rect 644 -3285 676 -3284
rect 644 -3315 645 -3285
rect 645 -3315 675 -3285
rect 675 -3315 676 -3285
rect 644 -3316 676 -3315
rect 644 -3396 676 -3364
rect 644 -3476 676 -3444
rect 644 -3525 676 -3524
rect 644 -3555 645 -3525
rect 645 -3555 675 -3525
rect 675 -3555 676 -3525
rect 644 -3556 676 -3555
rect 644 -3605 676 -3604
rect 644 -3635 645 -3605
rect 645 -3635 675 -3605
rect 675 -3635 676 -3605
rect 644 -3636 676 -3635
rect 644 -3685 676 -3684
rect 644 -3715 645 -3685
rect 645 -3715 675 -3685
rect 675 -3715 676 -3685
rect 644 -3716 676 -3715
rect 724 1035 756 1036
rect 724 1005 725 1035
rect 725 1005 755 1035
rect 755 1005 756 1035
rect 724 1004 756 1005
rect 724 955 756 956
rect 724 925 725 955
rect 725 925 755 955
rect 755 925 756 955
rect 724 924 756 925
rect 724 875 756 876
rect 724 845 725 875
rect 725 845 755 875
rect 755 845 756 875
rect 724 844 756 845
rect 724 764 756 796
rect 724 684 756 716
rect 724 635 756 636
rect 724 605 725 635
rect 725 605 755 635
rect 755 605 756 635
rect 724 604 756 605
rect 724 555 756 556
rect 724 525 725 555
rect 725 525 755 555
rect 755 525 756 555
rect 724 524 756 525
rect 724 444 756 476
rect 724 395 756 396
rect 724 365 725 395
rect 725 365 755 395
rect 755 365 756 395
rect 724 364 756 365
rect 724 284 756 316
rect 724 235 756 236
rect 724 205 725 235
rect 725 205 755 235
rect 755 205 756 235
rect 724 204 756 205
rect 724 124 756 156
rect 724 75 756 76
rect 724 45 725 75
rect 725 45 755 75
rect 755 45 756 75
rect 724 44 756 45
rect 724 -5 756 -4
rect 724 -35 725 -5
rect 725 -35 755 -5
rect 755 -35 756 -5
rect 724 -36 756 -35
rect 724 -85 756 -84
rect 724 -115 725 -85
rect 725 -115 755 -85
rect 755 -115 756 -85
rect 724 -116 756 -115
rect 724 -165 756 -164
rect 724 -195 725 -165
rect 725 -195 755 -165
rect 755 -195 756 -165
rect 724 -196 756 -195
rect 724 -245 756 -244
rect 724 -275 725 -245
rect 725 -275 755 -245
rect 755 -275 756 -245
rect 724 -276 756 -275
rect 724 -325 756 -324
rect 724 -355 725 -325
rect 725 -355 755 -325
rect 755 -355 756 -325
rect 724 -356 756 -355
rect 724 -436 756 -404
rect 724 -485 756 -484
rect 724 -515 725 -485
rect 725 -515 755 -485
rect 755 -515 756 -485
rect 724 -516 756 -515
rect 724 -596 756 -564
rect 724 -645 756 -644
rect 724 -675 725 -645
rect 725 -675 755 -645
rect 755 -675 756 -645
rect 724 -676 756 -675
rect 724 -756 756 -724
rect 724 -805 756 -804
rect 724 -835 725 -805
rect 725 -835 755 -805
rect 755 -835 756 -805
rect 724 -836 756 -835
rect 724 -885 756 -884
rect 724 -915 725 -885
rect 725 -915 755 -885
rect 755 -915 756 -885
rect 724 -916 756 -915
rect 724 -996 756 -964
rect 724 -1076 756 -1044
rect 724 -1125 756 -1124
rect 724 -1155 725 -1125
rect 725 -1155 755 -1125
rect 755 -1155 756 -1125
rect 724 -1156 756 -1155
rect 724 -1205 756 -1204
rect 724 -1235 725 -1205
rect 725 -1235 755 -1205
rect 755 -1235 756 -1205
rect 724 -1236 756 -1235
rect 724 -1285 756 -1284
rect 724 -1315 725 -1285
rect 725 -1315 755 -1285
rect 755 -1315 756 -1285
rect 724 -1316 756 -1315
rect 724 -1365 756 -1364
rect 724 -1395 725 -1365
rect 725 -1395 755 -1365
rect 755 -1395 756 -1365
rect 724 -1396 756 -1395
rect 724 -1445 756 -1444
rect 724 -1475 725 -1445
rect 725 -1475 755 -1445
rect 755 -1475 756 -1445
rect 724 -1476 756 -1475
rect 724 -1525 756 -1524
rect 724 -1555 725 -1525
rect 725 -1555 755 -1525
rect 755 -1555 756 -1525
rect 724 -1556 756 -1555
rect 724 -1636 756 -1604
rect 724 -1716 756 -1684
rect 724 -1765 756 -1764
rect 724 -1795 725 -1765
rect 725 -1795 755 -1765
rect 755 -1795 756 -1765
rect 724 -1796 756 -1795
rect 724 -1845 756 -1844
rect 724 -1875 725 -1845
rect 725 -1875 755 -1845
rect 755 -1875 756 -1845
rect 724 -1876 756 -1875
rect 724 -1956 756 -1924
rect 724 -2005 756 -2004
rect 724 -2035 725 -2005
rect 725 -2035 755 -2005
rect 755 -2035 756 -2005
rect 724 -2036 756 -2035
rect 724 -2116 756 -2084
rect 724 -2165 756 -2164
rect 724 -2195 725 -2165
rect 725 -2195 755 -2165
rect 755 -2195 756 -2165
rect 724 -2196 756 -2195
rect 724 -2276 756 -2244
rect 724 -2325 756 -2324
rect 724 -2355 725 -2325
rect 725 -2355 755 -2325
rect 755 -2355 756 -2325
rect 724 -2356 756 -2355
rect 724 -2405 756 -2404
rect 724 -2435 725 -2405
rect 725 -2435 755 -2405
rect 755 -2435 756 -2405
rect 724 -2436 756 -2435
rect 724 -2485 756 -2484
rect 724 -2515 725 -2485
rect 725 -2515 755 -2485
rect 755 -2515 756 -2485
rect 724 -2516 756 -2515
rect 724 -2565 756 -2564
rect 724 -2595 725 -2565
rect 725 -2595 755 -2565
rect 755 -2595 756 -2565
rect 724 -2596 756 -2595
rect 724 -2645 756 -2644
rect 724 -2675 725 -2645
rect 725 -2675 755 -2645
rect 755 -2675 756 -2645
rect 724 -2676 756 -2675
rect 724 -2725 756 -2724
rect 724 -2755 725 -2725
rect 725 -2755 755 -2725
rect 755 -2755 756 -2725
rect 724 -2756 756 -2755
rect 724 -2836 756 -2804
rect 724 -2885 756 -2884
rect 724 -2915 725 -2885
rect 725 -2915 755 -2885
rect 755 -2915 756 -2885
rect 724 -2916 756 -2915
rect 724 -2996 756 -2964
rect 724 -3045 756 -3044
rect 724 -3075 725 -3045
rect 725 -3075 755 -3045
rect 755 -3075 756 -3045
rect 724 -3076 756 -3075
rect 724 -3156 756 -3124
rect 724 -3205 756 -3204
rect 724 -3235 725 -3205
rect 725 -3235 755 -3205
rect 755 -3235 756 -3205
rect 724 -3236 756 -3235
rect 724 -3285 756 -3284
rect 724 -3315 725 -3285
rect 725 -3315 755 -3285
rect 755 -3315 756 -3285
rect 724 -3316 756 -3315
rect 724 -3396 756 -3364
rect 724 -3476 756 -3444
rect 724 -3525 756 -3524
rect 724 -3555 725 -3525
rect 725 -3555 755 -3525
rect 755 -3555 756 -3525
rect 724 -3556 756 -3555
rect 724 -3605 756 -3604
rect 724 -3635 725 -3605
rect 725 -3635 755 -3605
rect 755 -3635 756 -3605
rect 724 -3636 756 -3635
rect 724 -3685 756 -3684
rect 724 -3715 725 -3685
rect 725 -3715 755 -3685
rect 755 -3715 756 -3685
rect 724 -3716 756 -3715
rect 804 1035 836 1036
rect 804 1005 805 1035
rect 805 1005 835 1035
rect 835 1005 836 1035
rect 804 1004 836 1005
rect 804 955 836 956
rect 804 925 805 955
rect 805 925 835 955
rect 835 925 836 955
rect 804 924 836 925
rect 804 875 836 876
rect 804 845 805 875
rect 805 845 835 875
rect 835 845 836 875
rect 804 844 836 845
rect 804 764 836 796
rect 804 684 836 716
rect 804 635 836 636
rect 804 605 805 635
rect 805 605 835 635
rect 835 605 836 635
rect 804 604 836 605
rect 804 555 836 556
rect 804 525 805 555
rect 805 525 835 555
rect 835 525 836 555
rect 804 524 836 525
rect 804 444 836 476
rect 804 395 836 396
rect 804 365 805 395
rect 805 365 835 395
rect 835 365 836 395
rect 804 364 836 365
rect 804 284 836 316
rect 804 235 836 236
rect 804 205 805 235
rect 805 205 835 235
rect 835 205 836 235
rect 804 204 836 205
rect 804 124 836 156
rect 804 75 836 76
rect 804 45 805 75
rect 805 45 835 75
rect 835 45 836 75
rect 804 44 836 45
rect 804 -5 836 -4
rect 804 -35 805 -5
rect 805 -35 835 -5
rect 835 -35 836 -5
rect 804 -36 836 -35
rect 804 -85 836 -84
rect 804 -115 805 -85
rect 805 -115 835 -85
rect 835 -115 836 -85
rect 804 -116 836 -115
rect 804 -165 836 -164
rect 804 -195 805 -165
rect 805 -195 835 -165
rect 835 -195 836 -165
rect 804 -196 836 -195
rect 804 -245 836 -244
rect 804 -275 805 -245
rect 805 -275 835 -245
rect 835 -275 836 -245
rect 804 -276 836 -275
rect 804 -325 836 -324
rect 804 -355 805 -325
rect 805 -355 835 -325
rect 835 -355 836 -325
rect 804 -356 836 -355
rect 804 -436 836 -404
rect 804 -485 836 -484
rect 804 -515 805 -485
rect 805 -515 835 -485
rect 835 -515 836 -485
rect 804 -516 836 -515
rect 804 -596 836 -564
rect 804 -645 836 -644
rect 804 -675 805 -645
rect 805 -675 835 -645
rect 835 -675 836 -645
rect 804 -676 836 -675
rect 804 -756 836 -724
rect 804 -805 836 -804
rect 804 -835 805 -805
rect 805 -835 835 -805
rect 835 -835 836 -805
rect 804 -836 836 -835
rect 804 -885 836 -884
rect 804 -915 805 -885
rect 805 -915 835 -885
rect 835 -915 836 -885
rect 804 -916 836 -915
rect 804 -996 836 -964
rect 804 -1076 836 -1044
rect 804 -1125 836 -1124
rect 804 -1155 805 -1125
rect 805 -1155 835 -1125
rect 835 -1155 836 -1125
rect 804 -1156 836 -1155
rect 804 -1205 836 -1204
rect 804 -1235 805 -1205
rect 805 -1235 835 -1205
rect 835 -1235 836 -1205
rect 804 -1236 836 -1235
rect 804 -1285 836 -1284
rect 804 -1315 805 -1285
rect 805 -1315 835 -1285
rect 835 -1315 836 -1285
rect 804 -1316 836 -1315
rect 804 -1365 836 -1364
rect 804 -1395 805 -1365
rect 805 -1395 835 -1365
rect 835 -1395 836 -1365
rect 804 -1396 836 -1395
rect 804 -1445 836 -1444
rect 804 -1475 805 -1445
rect 805 -1475 835 -1445
rect 835 -1475 836 -1445
rect 804 -1476 836 -1475
rect 804 -1525 836 -1524
rect 804 -1555 805 -1525
rect 805 -1555 835 -1525
rect 835 -1555 836 -1525
rect 804 -1556 836 -1555
rect 804 -1636 836 -1604
rect 804 -1716 836 -1684
rect 804 -1765 836 -1764
rect 804 -1795 805 -1765
rect 805 -1795 835 -1765
rect 835 -1795 836 -1765
rect 804 -1796 836 -1795
rect 804 -1845 836 -1844
rect 804 -1875 805 -1845
rect 805 -1875 835 -1845
rect 835 -1875 836 -1845
rect 804 -1876 836 -1875
rect 804 -1956 836 -1924
rect 804 -2005 836 -2004
rect 804 -2035 805 -2005
rect 805 -2035 835 -2005
rect 835 -2035 836 -2005
rect 804 -2036 836 -2035
rect 804 -2116 836 -2084
rect 804 -2165 836 -2164
rect 804 -2195 805 -2165
rect 805 -2195 835 -2165
rect 835 -2195 836 -2165
rect 804 -2196 836 -2195
rect 804 -2276 836 -2244
rect 804 -2325 836 -2324
rect 804 -2355 805 -2325
rect 805 -2355 835 -2325
rect 835 -2355 836 -2325
rect 804 -2356 836 -2355
rect 804 -2405 836 -2404
rect 804 -2435 805 -2405
rect 805 -2435 835 -2405
rect 835 -2435 836 -2405
rect 804 -2436 836 -2435
rect 804 -2485 836 -2484
rect 804 -2515 805 -2485
rect 805 -2515 835 -2485
rect 835 -2515 836 -2485
rect 804 -2516 836 -2515
rect 804 -2565 836 -2564
rect 804 -2595 805 -2565
rect 805 -2595 835 -2565
rect 835 -2595 836 -2565
rect 804 -2596 836 -2595
rect 804 -2645 836 -2644
rect 804 -2675 805 -2645
rect 805 -2675 835 -2645
rect 835 -2675 836 -2645
rect 804 -2676 836 -2675
rect 804 -2725 836 -2724
rect 804 -2755 805 -2725
rect 805 -2755 835 -2725
rect 835 -2755 836 -2725
rect 804 -2756 836 -2755
rect 804 -2836 836 -2804
rect 804 -2885 836 -2884
rect 804 -2915 805 -2885
rect 805 -2915 835 -2885
rect 835 -2915 836 -2885
rect 804 -2916 836 -2915
rect 804 -2996 836 -2964
rect 804 -3045 836 -3044
rect 804 -3075 805 -3045
rect 805 -3075 835 -3045
rect 835 -3075 836 -3045
rect 804 -3076 836 -3075
rect 804 -3156 836 -3124
rect 804 -3205 836 -3204
rect 804 -3235 805 -3205
rect 805 -3235 835 -3205
rect 835 -3235 836 -3205
rect 804 -3236 836 -3235
rect 804 -3285 836 -3284
rect 804 -3315 805 -3285
rect 805 -3315 835 -3285
rect 835 -3315 836 -3285
rect 804 -3316 836 -3315
rect 804 -3396 836 -3364
rect 804 -3476 836 -3444
rect 804 -3525 836 -3524
rect 804 -3555 805 -3525
rect 805 -3555 835 -3525
rect 835 -3555 836 -3525
rect 804 -3556 836 -3555
rect 804 -3605 836 -3604
rect 804 -3635 805 -3605
rect 805 -3635 835 -3605
rect 835 -3635 836 -3605
rect 804 -3636 836 -3635
rect 804 -3685 836 -3684
rect 804 -3715 805 -3685
rect 805 -3715 835 -3685
rect 835 -3715 836 -3685
rect 804 -3716 836 -3715
rect 884 1035 916 1036
rect 884 1005 885 1035
rect 885 1005 915 1035
rect 915 1005 916 1035
rect 884 1004 916 1005
rect 884 955 916 956
rect 884 925 885 955
rect 885 925 915 955
rect 915 925 916 955
rect 884 924 916 925
rect 884 875 916 876
rect 884 845 885 875
rect 885 845 915 875
rect 915 845 916 875
rect 884 844 916 845
rect 884 764 916 796
rect 884 684 916 716
rect 884 635 916 636
rect 884 605 885 635
rect 885 605 915 635
rect 915 605 916 635
rect 884 604 916 605
rect 884 555 916 556
rect 884 525 885 555
rect 885 525 915 555
rect 915 525 916 555
rect 884 524 916 525
rect 884 444 916 476
rect 884 395 916 396
rect 884 365 885 395
rect 885 365 915 395
rect 915 365 916 395
rect 884 364 916 365
rect 884 284 916 316
rect 884 235 916 236
rect 884 205 885 235
rect 885 205 915 235
rect 915 205 916 235
rect 884 204 916 205
rect 884 124 916 156
rect 884 75 916 76
rect 884 45 885 75
rect 885 45 915 75
rect 915 45 916 75
rect 884 44 916 45
rect 884 -5 916 -4
rect 884 -35 885 -5
rect 885 -35 915 -5
rect 915 -35 916 -5
rect 884 -36 916 -35
rect 884 -85 916 -84
rect 884 -115 885 -85
rect 885 -115 915 -85
rect 915 -115 916 -85
rect 884 -116 916 -115
rect 884 -165 916 -164
rect 884 -195 885 -165
rect 885 -195 915 -165
rect 915 -195 916 -165
rect 884 -196 916 -195
rect 884 -245 916 -244
rect 884 -275 885 -245
rect 885 -275 915 -245
rect 915 -275 916 -245
rect 884 -276 916 -275
rect 884 -325 916 -324
rect 884 -355 885 -325
rect 885 -355 915 -325
rect 915 -355 916 -325
rect 884 -356 916 -355
rect 884 -436 916 -404
rect 884 -485 916 -484
rect 884 -515 885 -485
rect 885 -515 915 -485
rect 915 -515 916 -485
rect 884 -516 916 -515
rect 884 -596 916 -564
rect 884 -645 916 -644
rect 884 -675 885 -645
rect 885 -675 915 -645
rect 915 -675 916 -645
rect 884 -676 916 -675
rect 884 -756 916 -724
rect 884 -805 916 -804
rect 884 -835 885 -805
rect 885 -835 915 -805
rect 915 -835 916 -805
rect 884 -836 916 -835
rect 884 -885 916 -884
rect 884 -915 885 -885
rect 885 -915 915 -885
rect 915 -915 916 -885
rect 884 -916 916 -915
rect 884 -996 916 -964
rect 884 -1076 916 -1044
rect 884 -1125 916 -1124
rect 884 -1155 885 -1125
rect 885 -1155 915 -1125
rect 915 -1155 916 -1125
rect 884 -1156 916 -1155
rect 884 -1205 916 -1204
rect 884 -1235 885 -1205
rect 885 -1235 915 -1205
rect 915 -1235 916 -1205
rect 884 -1236 916 -1235
rect 884 -1285 916 -1284
rect 884 -1315 885 -1285
rect 885 -1315 915 -1285
rect 915 -1315 916 -1285
rect 884 -1316 916 -1315
rect 884 -1365 916 -1364
rect 884 -1395 885 -1365
rect 885 -1395 915 -1365
rect 915 -1395 916 -1365
rect 884 -1396 916 -1395
rect 884 -1445 916 -1444
rect 884 -1475 885 -1445
rect 885 -1475 915 -1445
rect 915 -1475 916 -1445
rect 884 -1476 916 -1475
rect 884 -1525 916 -1524
rect 884 -1555 885 -1525
rect 885 -1555 915 -1525
rect 915 -1555 916 -1525
rect 884 -1556 916 -1555
rect 884 -1636 916 -1604
rect 884 -1716 916 -1684
rect 884 -1765 916 -1764
rect 884 -1795 885 -1765
rect 885 -1795 915 -1765
rect 915 -1795 916 -1765
rect 884 -1796 916 -1795
rect 884 -1845 916 -1844
rect 884 -1875 885 -1845
rect 885 -1875 915 -1845
rect 915 -1875 916 -1845
rect 884 -1876 916 -1875
rect 884 -1956 916 -1924
rect 884 -2005 916 -2004
rect 884 -2035 885 -2005
rect 885 -2035 915 -2005
rect 915 -2035 916 -2005
rect 884 -2036 916 -2035
rect 884 -2116 916 -2084
rect 884 -2165 916 -2164
rect 884 -2195 885 -2165
rect 885 -2195 915 -2165
rect 915 -2195 916 -2165
rect 884 -2196 916 -2195
rect 884 -2276 916 -2244
rect 884 -2325 916 -2324
rect 884 -2355 885 -2325
rect 885 -2355 915 -2325
rect 915 -2355 916 -2325
rect 884 -2356 916 -2355
rect 884 -2405 916 -2404
rect 884 -2435 885 -2405
rect 885 -2435 915 -2405
rect 915 -2435 916 -2405
rect 884 -2436 916 -2435
rect 884 -2485 916 -2484
rect 884 -2515 885 -2485
rect 885 -2515 915 -2485
rect 915 -2515 916 -2485
rect 884 -2516 916 -2515
rect 884 -2565 916 -2564
rect 884 -2595 885 -2565
rect 885 -2595 915 -2565
rect 915 -2595 916 -2565
rect 884 -2596 916 -2595
rect 884 -2645 916 -2644
rect 884 -2675 885 -2645
rect 885 -2675 915 -2645
rect 915 -2675 916 -2645
rect 884 -2676 916 -2675
rect 884 -2725 916 -2724
rect 884 -2755 885 -2725
rect 885 -2755 915 -2725
rect 915 -2755 916 -2725
rect 884 -2756 916 -2755
rect 884 -2836 916 -2804
rect 884 -2885 916 -2884
rect 884 -2915 885 -2885
rect 885 -2915 915 -2885
rect 915 -2915 916 -2885
rect 884 -2916 916 -2915
rect 884 -2996 916 -2964
rect 884 -3045 916 -3044
rect 884 -3075 885 -3045
rect 885 -3075 915 -3045
rect 915 -3075 916 -3045
rect 884 -3076 916 -3075
rect 884 -3156 916 -3124
rect 884 -3205 916 -3204
rect 884 -3235 885 -3205
rect 885 -3235 915 -3205
rect 915 -3235 916 -3205
rect 884 -3236 916 -3235
rect 884 -3285 916 -3284
rect 884 -3315 885 -3285
rect 885 -3315 915 -3285
rect 915 -3315 916 -3285
rect 884 -3316 916 -3315
rect 884 -3396 916 -3364
rect 884 -3476 916 -3444
rect 884 -3525 916 -3524
rect 884 -3555 885 -3525
rect 885 -3555 915 -3525
rect 915 -3555 916 -3525
rect 884 -3556 916 -3555
rect 884 -3605 916 -3604
rect 884 -3635 885 -3605
rect 885 -3635 915 -3605
rect 915 -3635 916 -3605
rect 884 -3636 916 -3635
rect 884 -3685 916 -3684
rect 884 -3715 885 -3685
rect 885 -3715 915 -3685
rect 915 -3715 916 -3685
rect 884 -3716 916 -3715
rect 964 1035 996 1036
rect 964 1005 965 1035
rect 965 1005 995 1035
rect 995 1005 996 1035
rect 964 1004 996 1005
rect 964 955 996 956
rect 964 925 965 955
rect 965 925 995 955
rect 995 925 996 955
rect 964 924 996 925
rect 964 875 996 876
rect 964 845 965 875
rect 965 845 995 875
rect 995 845 996 875
rect 964 844 996 845
rect 964 764 996 796
rect 964 684 996 716
rect 964 635 996 636
rect 964 605 965 635
rect 965 605 995 635
rect 995 605 996 635
rect 964 604 996 605
rect 964 555 996 556
rect 964 525 965 555
rect 965 525 995 555
rect 995 525 996 555
rect 964 524 996 525
rect 964 444 996 476
rect 964 395 996 396
rect 964 365 965 395
rect 965 365 995 395
rect 995 365 996 395
rect 964 364 996 365
rect 964 284 996 316
rect 964 235 996 236
rect 964 205 965 235
rect 965 205 995 235
rect 995 205 996 235
rect 964 204 996 205
rect 964 124 996 156
rect 964 75 996 76
rect 964 45 965 75
rect 965 45 995 75
rect 995 45 996 75
rect 964 44 996 45
rect 964 -5 996 -4
rect 964 -35 965 -5
rect 965 -35 995 -5
rect 995 -35 996 -5
rect 964 -36 996 -35
rect 964 -85 996 -84
rect 964 -115 965 -85
rect 965 -115 995 -85
rect 995 -115 996 -85
rect 964 -116 996 -115
rect 964 -165 996 -164
rect 964 -195 965 -165
rect 965 -195 995 -165
rect 995 -195 996 -165
rect 964 -196 996 -195
rect 964 -245 996 -244
rect 964 -275 965 -245
rect 965 -275 995 -245
rect 995 -275 996 -245
rect 964 -276 996 -275
rect 964 -325 996 -324
rect 964 -355 965 -325
rect 965 -355 995 -325
rect 995 -355 996 -325
rect 964 -356 996 -355
rect 964 -436 996 -404
rect 964 -485 996 -484
rect 964 -515 965 -485
rect 965 -515 995 -485
rect 995 -515 996 -485
rect 964 -516 996 -515
rect 964 -596 996 -564
rect 964 -645 996 -644
rect 964 -675 965 -645
rect 965 -675 995 -645
rect 995 -675 996 -645
rect 964 -676 996 -675
rect 964 -756 996 -724
rect 964 -805 996 -804
rect 964 -835 965 -805
rect 965 -835 995 -805
rect 995 -835 996 -805
rect 964 -836 996 -835
rect 964 -885 996 -884
rect 964 -915 965 -885
rect 965 -915 995 -885
rect 995 -915 996 -885
rect 964 -916 996 -915
rect 964 -996 996 -964
rect 964 -1076 996 -1044
rect 964 -1125 996 -1124
rect 964 -1155 965 -1125
rect 965 -1155 995 -1125
rect 995 -1155 996 -1125
rect 964 -1156 996 -1155
rect 964 -1205 996 -1204
rect 964 -1235 965 -1205
rect 965 -1235 995 -1205
rect 995 -1235 996 -1205
rect 964 -1236 996 -1235
rect 964 -1285 996 -1284
rect 964 -1315 965 -1285
rect 965 -1315 995 -1285
rect 995 -1315 996 -1285
rect 964 -1316 996 -1315
rect 964 -1365 996 -1364
rect 964 -1395 965 -1365
rect 965 -1395 995 -1365
rect 995 -1395 996 -1365
rect 964 -1396 996 -1395
rect 964 -1445 996 -1444
rect 964 -1475 965 -1445
rect 965 -1475 995 -1445
rect 995 -1475 996 -1445
rect 964 -1476 996 -1475
rect 964 -1525 996 -1524
rect 964 -1555 965 -1525
rect 965 -1555 995 -1525
rect 995 -1555 996 -1525
rect 964 -1556 996 -1555
rect 964 -1636 996 -1604
rect 964 -1716 996 -1684
rect 964 -1765 996 -1764
rect 964 -1795 965 -1765
rect 965 -1795 995 -1765
rect 995 -1795 996 -1765
rect 964 -1796 996 -1795
rect 964 -1845 996 -1844
rect 964 -1875 965 -1845
rect 965 -1875 995 -1845
rect 995 -1875 996 -1845
rect 964 -1876 996 -1875
rect 964 -1956 996 -1924
rect 964 -2005 996 -2004
rect 964 -2035 965 -2005
rect 965 -2035 995 -2005
rect 995 -2035 996 -2005
rect 964 -2036 996 -2035
rect 964 -2116 996 -2084
rect 964 -2165 996 -2164
rect 964 -2195 965 -2165
rect 965 -2195 995 -2165
rect 995 -2195 996 -2165
rect 964 -2196 996 -2195
rect 964 -2276 996 -2244
rect 964 -2325 996 -2324
rect 964 -2355 965 -2325
rect 965 -2355 995 -2325
rect 995 -2355 996 -2325
rect 964 -2356 996 -2355
rect 964 -2405 996 -2404
rect 964 -2435 965 -2405
rect 965 -2435 995 -2405
rect 995 -2435 996 -2405
rect 964 -2436 996 -2435
rect 964 -2485 996 -2484
rect 964 -2515 965 -2485
rect 965 -2515 995 -2485
rect 995 -2515 996 -2485
rect 964 -2516 996 -2515
rect 964 -2565 996 -2564
rect 964 -2595 965 -2565
rect 965 -2595 995 -2565
rect 995 -2595 996 -2565
rect 964 -2596 996 -2595
rect 964 -2645 996 -2644
rect 964 -2675 965 -2645
rect 965 -2675 995 -2645
rect 995 -2675 996 -2645
rect 964 -2676 996 -2675
rect 964 -2725 996 -2724
rect 964 -2755 965 -2725
rect 965 -2755 995 -2725
rect 995 -2755 996 -2725
rect 964 -2756 996 -2755
rect 964 -2836 996 -2804
rect 964 -2885 996 -2884
rect 964 -2915 965 -2885
rect 965 -2915 995 -2885
rect 995 -2915 996 -2885
rect 964 -2916 996 -2915
rect 964 -2996 996 -2964
rect 964 -3045 996 -3044
rect 964 -3075 965 -3045
rect 965 -3075 995 -3045
rect 995 -3075 996 -3045
rect 964 -3076 996 -3075
rect 964 -3156 996 -3124
rect 964 -3205 996 -3204
rect 964 -3235 965 -3205
rect 965 -3235 995 -3205
rect 995 -3235 996 -3205
rect 964 -3236 996 -3235
rect 964 -3285 996 -3284
rect 964 -3315 965 -3285
rect 965 -3315 995 -3285
rect 995 -3315 996 -3285
rect 964 -3316 996 -3315
rect 964 -3396 996 -3364
rect 964 -3476 996 -3444
rect 964 -3525 996 -3524
rect 964 -3555 965 -3525
rect 965 -3555 995 -3525
rect 995 -3555 996 -3525
rect 964 -3556 996 -3555
rect 964 -3605 996 -3604
rect 964 -3635 965 -3605
rect 965 -3635 995 -3605
rect 995 -3635 996 -3605
rect 964 -3636 996 -3635
rect 964 -3685 996 -3684
rect 964 -3715 965 -3685
rect 965 -3715 995 -3685
rect 995 -3715 996 -3685
rect 964 -3716 996 -3715
rect 1044 1035 1076 1036
rect 1044 1005 1045 1035
rect 1045 1005 1075 1035
rect 1075 1005 1076 1035
rect 1044 1004 1076 1005
rect 1044 955 1076 956
rect 1044 925 1045 955
rect 1045 925 1075 955
rect 1075 925 1076 955
rect 1044 924 1076 925
rect 1044 875 1076 876
rect 1044 845 1045 875
rect 1045 845 1075 875
rect 1075 845 1076 875
rect 1044 844 1076 845
rect 1044 764 1076 796
rect 1044 684 1076 716
rect 1044 635 1076 636
rect 1044 605 1045 635
rect 1045 605 1075 635
rect 1075 605 1076 635
rect 1044 604 1076 605
rect 1044 555 1076 556
rect 1044 525 1045 555
rect 1045 525 1075 555
rect 1075 525 1076 555
rect 1044 524 1076 525
rect 1044 444 1076 476
rect 1044 395 1076 396
rect 1044 365 1045 395
rect 1045 365 1075 395
rect 1075 365 1076 395
rect 1044 364 1076 365
rect 1044 284 1076 316
rect 1044 235 1076 236
rect 1044 205 1045 235
rect 1045 205 1075 235
rect 1075 205 1076 235
rect 1044 204 1076 205
rect 1044 124 1076 156
rect 1044 75 1076 76
rect 1044 45 1045 75
rect 1045 45 1075 75
rect 1075 45 1076 75
rect 1044 44 1076 45
rect 1044 -5 1076 -4
rect 1044 -35 1045 -5
rect 1045 -35 1075 -5
rect 1075 -35 1076 -5
rect 1044 -36 1076 -35
rect 1044 -85 1076 -84
rect 1044 -115 1045 -85
rect 1045 -115 1075 -85
rect 1075 -115 1076 -85
rect 1044 -116 1076 -115
rect 1044 -165 1076 -164
rect 1044 -195 1045 -165
rect 1045 -195 1075 -165
rect 1075 -195 1076 -165
rect 1044 -196 1076 -195
rect 1044 -245 1076 -244
rect 1044 -275 1045 -245
rect 1045 -275 1075 -245
rect 1075 -275 1076 -245
rect 1044 -276 1076 -275
rect 1044 -325 1076 -324
rect 1044 -355 1045 -325
rect 1045 -355 1075 -325
rect 1075 -355 1076 -325
rect 1044 -356 1076 -355
rect 1044 -436 1076 -404
rect 1044 -485 1076 -484
rect 1044 -515 1045 -485
rect 1045 -515 1075 -485
rect 1075 -515 1076 -485
rect 1044 -516 1076 -515
rect 1044 -596 1076 -564
rect 1044 -645 1076 -644
rect 1044 -675 1045 -645
rect 1045 -675 1075 -645
rect 1075 -675 1076 -645
rect 1044 -676 1076 -675
rect 1044 -756 1076 -724
rect 1044 -805 1076 -804
rect 1044 -835 1045 -805
rect 1045 -835 1075 -805
rect 1075 -835 1076 -805
rect 1044 -836 1076 -835
rect 1044 -885 1076 -884
rect 1044 -915 1045 -885
rect 1045 -915 1075 -885
rect 1075 -915 1076 -885
rect 1044 -916 1076 -915
rect 1044 -996 1076 -964
rect 1044 -1076 1076 -1044
rect 1044 -1125 1076 -1124
rect 1044 -1155 1045 -1125
rect 1045 -1155 1075 -1125
rect 1075 -1155 1076 -1125
rect 1044 -1156 1076 -1155
rect 1044 -1205 1076 -1204
rect 1044 -1235 1045 -1205
rect 1045 -1235 1075 -1205
rect 1075 -1235 1076 -1205
rect 1044 -1236 1076 -1235
rect 1044 -1285 1076 -1284
rect 1044 -1315 1045 -1285
rect 1045 -1315 1075 -1285
rect 1075 -1315 1076 -1285
rect 1044 -1316 1076 -1315
rect 1044 -1365 1076 -1364
rect 1044 -1395 1045 -1365
rect 1045 -1395 1075 -1365
rect 1075 -1395 1076 -1365
rect 1044 -1396 1076 -1395
rect 1044 -1445 1076 -1444
rect 1044 -1475 1045 -1445
rect 1045 -1475 1075 -1445
rect 1075 -1475 1076 -1445
rect 1044 -1476 1076 -1475
rect 1044 -1525 1076 -1524
rect 1044 -1555 1045 -1525
rect 1045 -1555 1075 -1525
rect 1075 -1555 1076 -1525
rect 1044 -1556 1076 -1555
rect 1044 -1636 1076 -1604
rect 1044 -1716 1076 -1684
rect 1044 -1765 1076 -1764
rect 1044 -1795 1045 -1765
rect 1045 -1795 1075 -1765
rect 1075 -1795 1076 -1765
rect 1044 -1796 1076 -1795
rect 1044 -1845 1076 -1844
rect 1044 -1875 1045 -1845
rect 1045 -1875 1075 -1845
rect 1075 -1875 1076 -1845
rect 1044 -1876 1076 -1875
rect 1044 -1956 1076 -1924
rect 1044 -2005 1076 -2004
rect 1044 -2035 1045 -2005
rect 1045 -2035 1075 -2005
rect 1075 -2035 1076 -2005
rect 1044 -2036 1076 -2035
rect 1044 -2116 1076 -2084
rect 1044 -2165 1076 -2164
rect 1044 -2195 1045 -2165
rect 1045 -2195 1075 -2165
rect 1075 -2195 1076 -2165
rect 1044 -2196 1076 -2195
rect 1044 -2276 1076 -2244
rect 1044 -2325 1076 -2324
rect 1044 -2355 1045 -2325
rect 1045 -2355 1075 -2325
rect 1075 -2355 1076 -2325
rect 1044 -2356 1076 -2355
rect 1044 -2405 1076 -2404
rect 1044 -2435 1045 -2405
rect 1045 -2435 1075 -2405
rect 1075 -2435 1076 -2405
rect 1044 -2436 1076 -2435
rect 1044 -2485 1076 -2484
rect 1044 -2515 1045 -2485
rect 1045 -2515 1075 -2485
rect 1075 -2515 1076 -2485
rect 1044 -2516 1076 -2515
rect 1044 -2565 1076 -2564
rect 1044 -2595 1045 -2565
rect 1045 -2595 1075 -2565
rect 1075 -2595 1076 -2565
rect 1044 -2596 1076 -2595
rect 1044 -2645 1076 -2644
rect 1044 -2675 1045 -2645
rect 1045 -2675 1075 -2645
rect 1075 -2675 1076 -2645
rect 1044 -2676 1076 -2675
rect 1044 -2725 1076 -2724
rect 1044 -2755 1045 -2725
rect 1045 -2755 1075 -2725
rect 1075 -2755 1076 -2725
rect 1044 -2756 1076 -2755
rect 1044 -2836 1076 -2804
rect 1044 -2885 1076 -2884
rect 1044 -2915 1045 -2885
rect 1045 -2915 1075 -2885
rect 1075 -2915 1076 -2885
rect 1044 -2916 1076 -2915
rect 1044 -2996 1076 -2964
rect 1044 -3045 1076 -3044
rect 1044 -3075 1045 -3045
rect 1045 -3075 1075 -3045
rect 1075 -3075 1076 -3045
rect 1044 -3076 1076 -3075
rect 1044 -3156 1076 -3124
rect 1044 -3205 1076 -3204
rect 1044 -3235 1045 -3205
rect 1045 -3235 1075 -3205
rect 1075 -3235 1076 -3205
rect 1044 -3236 1076 -3235
rect 1044 -3285 1076 -3284
rect 1044 -3315 1045 -3285
rect 1045 -3315 1075 -3285
rect 1075 -3315 1076 -3285
rect 1044 -3316 1076 -3315
rect 1044 -3396 1076 -3364
rect 1044 -3476 1076 -3444
rect 1044 -3525 1076 -3524
rect 1044 -3555 1045 -3525
rect 1045 -3555 1075 -3525
rect 1075 -3555 1076 -3525
rect 1044 -3556 1076 -3555
rect 1044 -3605 1076 -3604
rect 1044 -3635 1045 -3605
rect 1045 -3635 1075 -3605
rect 1075 -3635 1076 -3605
rect 1044 -3636 1076 -3635
rect 1044 -3685 1076 -3684
rect 1044 -3715 1045 -3685
rect 1045 -3715 1075 -3685
rect 1075 -3715 1076 -3685
rect 1044 -3716 1076 -3715
rect 1124 1035 1156 1036
rect 1124 1005 1125 1035
rect 1125 1005 1155 1035
rect 1155 1005 1156 1035
rect 1124 1004 1156 1005
rect 1124 955 1156 956
rect 1124 925 1125 955
rect 1125 925 1155 955
rect 1155 925 1156 955
rect 1124 924 1156 925
rect 1124 875 1156 876
rect 1124 845 1125 875
rect 1125 845 1155 875
rect 1155 845 1156 875
rect 1124 844 1156 845
rect 1124 764 1156 796
rect 1124 684 1156 716
rect 1124 635 1156 636
rect 1124 605 1125 635
rect 1125 605 1155 635
rect 1155 605 1156 635
rect 1124 604 1156 605
rect 1124 555 1156 556
rect 1124 525 1125 555
rect 1125 525 1155 555
rect 1155 525 1156 555
rect 1124 524 1156 525
rect 1124 444 1156 476
rect 1124 395 1156 396
rect 1124 365 1125 395
rect 1125 365 1155 395
rect 1155 365 1156 395
rect 1124 364 1156 365
rect 1124 284 1156 316
rect 1124 235 1156 236
rect 1124 205 1125 235
rect 1125 205 1155 235
rect 1155 205 1156 235
rect 1124 204 1156 205
rect 1124 124 1156 156
rect 1124 75 1156 76
rect 1124 45 1125 75
rect 1125 45 1155 75
rect 1155 45 1156 75
rect 1124 44 1156 45
rect 1124 -5 1156 -4
rect 1124 -35 1125 -5
rect 1125 -35 1155 -5
rect 1155 -35 1156 -5
rect 1124 -36 1156 -35
rect 1124 -85 1156 -84
rect 1124 -115 1125 -85
rect 1125 -115 1155 -85
rect 1155 -115 1156 -85
rect 1124 -116 1156 -115
rect 1124 -165 1156 -164
rect 1124 -195 1125 -165
rect 1125 -195 1155 -165
rect 1155 -195 1156 -165
rect 1124 -196 1156 -195
rect 1124 -245 1156 -244
rect 1124 -275 1125 -245
rect 1125 -275 1155 -245
rect 1155 -275 1156 -245
rect 1124 -276 1156 -275
rect 1124 -325 1156 -324
rect 1124 -355 1125 -325
rect 1125 -355 1155 -325
rect 1155 -355 1156 -325
rect 1124 -356 1156 -355
rect 1124 -436 1156 -404
rect 1124 -485 1156 -484
rect 1124 -515 1125 -485
rect 1125 -515 1155 -485
rect 1155 -515 1156 -485
rect 1124 -516 1156 -515
rect 1124 -596 1156 -564
rect 1124 -645 1156 -644
rect 1124 -675 1125 -645
rect 1125 -675 1155 -645
rect 1155 -675 1156 -645
rect 1124 -676 1156 -675
rect 1124 -756 1156 -724
rect 1124 -805 1156 -804
rect 1124 -835 1125 -805
rect 1125 -835 1155 -805
rect 1155 -835 1156 -805
rect 1124 -836 1156 -835
rect 1124 -885 1156 -884
rect 1124 -915 1125 -885
rect 1125 -915 1155 -885
rect 1155 -915 1156 -885
rect 1124 -916 1156 -915
rect 1124 -996 1156 -964
rect 1124 -1076 1156 -1044
rect 1124 -1125 1156 -1124
rect 1124 -1155 1125 -1125
rect 1125 -1155 1155 -1125
rect 1155 -1155 1156 -1125
rect 1124 -1156 1156 -1155
rect 1124 -1205 1156 -1204
rect 1124 -1235 1125 -1205
rect 1125 -1235 1155 -1205
rect 1155 -1235 1156 -1205
rect 1124 -1236 1156 -1235
rect 1124 -1285 1156 -1284
rect 1124 -1315 1125 -1285
rect 1125 -1315 1155 -1285
rect 1155 -1315 1156 -1285
rect 1124 -1316 1156 -1315
rect 1124 -1365 1156 -1364
rect 1124 -1395 1125 -1365
rect 1125 -1395 1155 -1365
rect 1155 -1395 1156 -1365
rect 1124 -1396 1156 -1395
rect 1124 -1445 1156 -1444
rect 1124 -1475 1125 -1445
rect 1125 -1475 1155 -1445
rect 1155 -1475 1156 -1445
rect 1124 -1476 1156 -1475
rect 1124 -1525 1156 -1524
rect 1124 -1555 1125 -1525
rect 1125 -1555 1155 -1525
rect 1155 -1555 1156 -1525
rect 1124 -1556 1156 -1555
rect 1124 -1636 1156 -1604
rect 1124 -1716 1156 -1684
rect 1124 -1765 1156 -1764
rect 1124 -1795 1125 -1765
rect 1125 -1795 1155 -1765
rect 1155 -1795 1156 -1765
rect 1124 -1796 1156 -1795
rect 1124 -1845 1156 -1844
rect 1124 -1875 1125 -1845
rect 1125 -1875 1155 -1845
rect 1155 -1875 1156 -1845
rect 1124 -1876 1156 -1875
rect 1124 -1956 1156 -1924
rect 1124 -2005 1156 -2004
rect 1124 -2035 1125 -2005
rect 1125 -2035 1155 -2005
rect 1155 -2035 1156 -2005
rect 1124 -2036 1156 -2035
rect 1124 -2116 1156 -2084
rect 1124 -2165 1156 -2164
rect 1124 -2195 1125 -2165
rect 1125 -2195 1155 -2165
rect 1155 -2195 1156 -2165
rect 1124 -2196 1156 -2195
rect 1124 -2276 1156 -2244
rect 1124 -2325 1156 -2324
rect 1124 -2355 1125 -2325
rect 1125 -2355 1155 -2325
rect 1155 -2355 1156 -2325
rect 1124 -2356 1156 -2355
rect 1124 -2405 1156 -2404
rect 1124 -2435 1125 -2405
rect 1125 -2435 1155 -2405
rect 1155 -2435 1156 -2405
rect 1124 -2436 1156 -2435
rect 1124 -2485 1156 -2484
rect 1124 -2515 1125 -2485
rect 1125 -2515 1155 -2485
rect 1155 -2515 1156 -2485
rect 1124 -2516 1156 -2515
rect 1124 -2565 1156 -2564
rect 1124 -2595 1125 -2565
rect 1125 -2595 1155 -2565
rect 1155 -2595 1156 -2565
rect 1124 -2596 1156 -2595
rect 1124 -2645 1156 -2644
rect 1124 -2675 1125 -2645
rect 1125 -2675 1155 -2645
rect 1155 -2675 1156 -2645
rect 1124 -2676 1156 -2675
rect 1124 -2725 1156 -2724
rect 1124 -2755 1125 -2725
rect 1125 -2755 1155 -2725
rect 1155 -2755 1156 -2725
rect 1124 -2756 1156 -2755
rect 1124 -2836 1156 -2804
rect 1124 -2885 1156 -2884
rect 1124 -2915 1125 -2885
rect 1125 -2915 1155 -2885
rect 1155 -2915 1156 -2885
rect 1124 -2916 1156 -2915
rect 1124 -2996 1156 -2964
rect 1124 -3045 1156 -3044
rect 1124 -3075 1125 -3045
rect 1125 -3075 1155 -3045
rect 1155 -3075 1156 -3045
rect 1124 -3076 1156 -3075
rect 1124 -3156 1156 -3124
rect 1124 -3205 1156 -3204
rect 1124 -3235 1125 -3205
rect 1125 -3235 1155 -3205
rect 1155 -3235 1156 -3205
rect 1124 -3236 1156 -3235
rect 1124 -3285 1156 -3284
rect 1124 -3315 1125 -3285
rect 1125 -3315 1155 -3285
rect 1155 -3315 1156 -3285
rect 1124 -3316 1156 -3315
rect 1124 -3396 1156 -3364
rect 1124 -3476 1156 -3444
rect 1124 -3525 1156 -3524
rect 1124 -3555 1125 -3525
rect 1125 -3555 1155 -3525
rect 1155 -3555 1156 -3525
rect 1124 -3556 1156 -3555
rect 1124 -3605 1156 -3604
rect 1124 -3635 1125 -3605
rect 1125 -3635 1155 -3605
rect 1155 -3635 1156 -3605
rect 1124 -3636 1156 -3635
rect 1124 -3685 1156 -3684
rect 1124 -3715 1125 -3685
rect 1125 -3715 1155 -3685
rect 1155 -3715 1156 -3685
rect 1124 -3716 1156 -3715
rect 1204 1035 1236 1036
rect 1204 1005 1205 1035
rect 1205 1005 1235 1035
rect 1235 1005 1236 1035
rect 1204 1004 1236 1005
rect 1204 955 1236 956
rect 1204 925 1205 955
rect 1205 925 1235 955
rect 1235 925 1236 955
rect 1204 924 1236 925
rect 1204 875 1236 876
rect 1204 845 1205 875
rect 1205 845 1235 875
rect 1235 845 1236 875
rect 1204 844 1236 845
rect 1204 764 1236 796
rect 1204 684 1236 716
rect 1204 635 1236 636
rect 1204 605 1205 635
rect 1205 605 1235 635
rect 1235 605 1236 635
rect 1204 604 1236 605
rect 1204 555 1236 556
rect 1204 525 1205 555
rect 1205 525 1235 555
rect 1235 525 1236 555
rect 1204 524 1236 525
rect 1204 444 1236 476
rect 1204 395 1236 396
rect 1204 365 1205 395
rect 1205 365 1235 395
rect 1235 365 1236 395
rect 1204 364 1236 365
rect 1204 284 1236 316
rect 1204 235 1236 236
rect 1204 205 1205 235
rect 1205 205 1235 235
rect 1235 205 1236 235
rect 1204 204 1236 205
rect 1204 124 1236 156
rect 1204 75 1236 76
rect 1204 45 1205 75
rect 1205 45 1235 75
rect 1235 45 1236 75
rect 1204 44 1236 45
rect 1204 -5 1236 -4
rect 1204 -35 1205 -5
rect 1205 -35 1235 -5
rect 1235 -35 1236 -5
rect 1204 -36 1236 -35
rect 1204 -85 1236 -84
rect 1204 -115 1205 -85
rect 1205 -115 1235 -85
rect 1235 -115 1236 -85
rect 1204 -116 1236 -115
rect 1204 -165 1236 -164
rect 1204 -195 1205 -165
rect 1205 -195 1235 -165
rect 1235 -195 1236 -165
rect 1204 -196 1236 -195
rect 1204 -245 1236 -244
rect 1204 -275 1205 -245
rect 1205 -275 1235 -245
rect 1235 -275 1236 -245
rect 1204 -276 1236 -275
rect 1204 -325 1236 -324
rect 1204 -355 1205 -325
rect 1205 -355 1235 -325
rect 1235 -355 1236 -325
rect 1204 -356 1236 -355
rect 1204 -436 1236 -404
rect 1204 -485 1236 -484
rect 1204 -515 1205 -485
rect 1205 -515 1235 -485
rect 1235 -515 1236 -485
rect 1204 -516 1236 -515
rect 1204 -596 1236 -564
rect 1204 -645 1236 -644
rect 1204 -675 1205 -645
rect 1205 -675 1235 -645
rect 1235 -675 1236 -645
rect 1204 -676 1236 -675
rect 1204 -756 1236 -724
rect 1204 -805 1236 -804
rect 1204 -835 1205 -805
rect 1205 -835 1235 -805
rect 1235 -835 1236 -805
rect 1204 -836 1236 -835
rect 1204 -885 1236 -884
rect 1204 -915 1205 -885
rect 1205 -915 1235 -885
rect 1235 -915 1236 -885
rect 1204 -916 1236 -915
rect 1204 -996 1236 -964
rect 1204 -1076 1236 -1044
rect 1204 -1125 1236 -1124
rect 1204 -1155 1205 -1125
rect 1205 -1155 1235 -1125
rect 1235 -1155 1236 -1125
rect 1204 -1156 1236 -1155
rect 1204 -1205 1236 -1204
rect 1204 -1235 1205 -1205
rect 1205 -1235 1235 -1205
rect 1235 -1235 1236 -1205
rect 1204 -1236 1236 -1235
rect 1204 -1285 1236 -1284
rect 1204 -1315 1205 -1285
rect 1205 -1315 1235 -1285
rect 1235 -1315 1236 -1285
rect 1204 -1316 1236 -1315
rect 1204 -1365 1236 -1364
rect 1204 -1395 1205 -1365
rect 1205 -1395 1235 -1365
rect 1235 -1395 1236 -1365
rect 1204 -1396 1236 -1395
rect 1204 -1445 1236 -1444
rect 1204 -1475 1205 -1445
rect 1205 -1475 1235 -1445
rect 1235 -1475 1236 -1445
rect 1204 -1476 1236 -1475
rect 1204 -1525 1236 -1524
rect 1204 -1555 1205 -1525
rect 1205 -1555 1235 -1525
rect 1235 -1555 1236 -1525
rect 1204 -1556 1236 -1555
rect 1204 -1636 1236 -1604
rect 1204 -1716 1236 -1684
rect 1204 -1765 1236 -1764
rect 1204 -1795 1205 -1765
rect 1205 -1795 1235 -1765
rect 1235 -1795 1236 -1765
rect 1204 -1796 1236 -1795
rect 1204 -1845 1236 -1844
rect 1204 -1875 1205 -1845
rect 1205 -1875 1235 -1845
rect 1235 -1875 1236 -1845
rect 1204 -1876 1236 -1875
rect 1204 -1956 1236 -1924
rect 1204 -2005 1236 -2004
rect 1204 -2035 1205 -2005
rect 1205 -2035 1235 -2005
rect 1235 -2035 1236 -2005
rect 1204 -2036 1236 -2035
rect 1204 -2116 1236 -2084
rect 1204 -2165 1236 -2164
rect 1204 -2195 1205 -2165
rect 1205 -2195 1235 -2165
rect 1235 -2195 1236 -2165
rect 1204 -2196 1236 -2195
rect 1204 -2276 1236 -2244
rect 1204 -2325 1236 -2324
rect 1204 -2355 1205 -2325
rect 1205 -2355 1235 -2325
rect 1235 -2355 1236 -2325
rect 1204 -2356 1236 -2355
rect 1204 -2405 1236 -2404
rect 1204 -2435 1205 -2405
rect 1205 -2435 1235 -2405
rect 1235 -2435 1236 -2405
rect 1204 -2436 1236 -2435
rect 1204 -2485 1236 -2484
rect 1204 -2515 1205 -2485
rect 1205 -2515 1235 -2485
rect 1235 -2515 1236 -2485
rect 1204 -2516 1236 -2515
rect 1204 -2565 1236 -2564
rect 1204 -2595 1205 -2565
rect 1205 -2595 1235 -2565
rect 1235 -2595 1236 -2565
rect 1204 -2596 1236 -2595
rect 1204 -2645 1236 -2644
rect 1204 -2675 1205 -2645
rect 1205 -2675 1235 -2645
rect 1235 -2675 1236 -2645
rect 1204 -2676 1236 -2675
rect 1204 -2725 1236 -2724
rect 1204 -2755 1205 -2725
rect 1205 -2755 1235 -2725
rect 1235 -2755 1236 -2725
rect 1204 -2756 1236 -2755
rect 1204 -2836 1236 -2804
rect 1204 -2885 1236 -2884
rect 1204 -2915 1205 -2885
rect 1205 -2915 1235 -2885
rect 1235 -2915 1236 -2885
rect 1204 -2916 1236 -2915
rect 1204 -2996 1236 -2964
rect 1204 -3045 1236 -3044
rect 1204 -3075 1205 -3045
rect 1205 -3075 1235 -3045
rect 1235 -3075 1236 -3045
rect 1204 -3076 1236 -3075
rect 1204 -3156 1236 -3124
rect 1204 -3205 1236 -3204
rect 1204 -3235 1205 -3205
rect 1205 -3235 1235 -3205
rect 1235 -3235 1236 -3205
rect 1204 -3236 1236 -3235
rect 1204 -3285 1236 -3284
rect 1204 -3315 1205 -3285
rect 1205 -3315 1235 -3285
rect 1235 -3315 1236 -3285
rect 1204 -3316 1236 -3315
rect 1204 -3396 1236 -3364
rect 1204 -3476 1236 -3444
rect 1204 -3525 1236 -3524
rect 1204 -3555 1205 -3525
rect 1205 -3555 1235 -3525
rect 1235 -3555 1236 -3525
rect 1204 -3556 1236 -3555
rect 1204 -3605 1236 -3604
rect 1204 -3635 1205 -3605
rect 1205 -3635 1235 -3605
rect 1235 -3635 1236 -3605
rect 1204 -3636 1236 -3635
rect 1204 -3685 1236 -3684
rect 1204 -3715 1205 -3685
rect 1205 -3715 1235 -3685
rect 1235 -3715 1236 -3685
rect 1204 -3716 1236 -3715
rect 1284 1035 1316 1036
rect 1284 1005 1285 1035
rect 1285 1005 1315 1035
rect 1315 1005 1316 1035
rect 1284 1004 1316 1005
rect 1284 955 1316 956
rect 1284 925 1285 955
rect 1285 925 1315 955
rect 1315 925 1316 955
rect 1284 924 1316 925
rect 1284 875 1316 876
rect 1284 845 1285 875
rect 1285 845 1315 875
rect 1315 845 1316 875
rect 1284 844 1316 845
rect 1284 764 1316 796
rect 1284 684 1316 716
rect 1284 635 1316 636
rect 1284 605 1285 635
rect 1285 605 1315 635
rect 1315 605 1316 635
rect 1284 604 1316 605
rect 1284 555 1316 556
rect 1284 525 1285 555
rect 1285 525 1315 555
rect 1315 525 1316 555
rect 1284 524 1316 525
rect 1284 444 1316 476
rect 1284 395 1316 396
rect 1284 365 1285 395
rect 1285 365 1315 395
rect 1315 365 1316 395
rect 1284 364 1316 365
rect 1284 284 1316 316
rect 1284 235 1316 236
rect 1284 205 1285 235
rect 1285 205 1315 235
rect 1315 205 1316 235
rect 1284 204 1316 205
rect 1284 124 1316 156
rect 1284 75 1316 76
rect 1284 45 1285 75
rect 1285 45 1315 75
rect 1315 45 1316 75
rect 1284 44 1316 45
rect 1284 -5 1316 -4
rect 1284 -35 1285 -5
rect 1285 -35 1315 -5
rect 1315 -35 1316 -5
rect 1284 -36 1316 -35
rect 1284 -85 1316 -84
rect 1284 -115 1285 -85
rect 1285 -115 1315 -85
rect 1315 -115 1316 -85
rect 1284 -116 1316 -115
rect 1284 -165 1316 -164
rect 1284 -195 1285 -165
rect 1285 -195 1315 -165
rect 1315 -195 1316 -165
rect 1284 -196 1316 -195
rect 1284 -245 1316 -244
rect 1284 -275 1285 -245
rect 1285 -275 1315 -245
rect 1315 -275 1316 -245
rect 1284 -276 1316 -275
rect 1284 -325 1316 -324
rect 1284 -355 1285 -325
rect 1285 -355 1315 -325
rect 1315 -355 1316 -325
rect 1284 -356 1316 -355
rect 1284 -436 1316 -404
rect 1284 -485 1316 -484
rect 1284 -515 1285 -485
rect 1285 -515 1315 -485
rect 1315 -515 1316 -485
rect 1284 -516 1316 -515
rect 1284 -596 1316 -564
rect 1284 -645 1316 -644
rect 1284 -675 1285 -645
rect 1285 -675 1315 -645
rect 1315 -675 1316 -645
rect 1284 -676 1316 -675
rect 1284 -756 1316 -724
rect 1284 -805 1316 -804
rect 1284 -835 1285 -805
rect 1285 -835 1315 -805
rect 1315 -835 1316 -805
rect 1284 -836 1316 -835
rect 1284 -885 1316 -884
rect 1284 -915 1285 -885
rect 1285 -915 1315 -885
rect 1315 -915 1316 -885
rect 1284 -916 1316 -915
rect 1284 -996 1316 -964
rect 1284 -1076 1316 -1044
rect 1284 -1125 1316 -1124
rect 1284 -1155 1285 -1125
rect 1285 -1155 1315 -1125
rect 1315 -1155 1316 -1125
rect 1284 -1156 1316 -1155
rect 1284 -1205 1316 -1204
rect 1284 -1235 1285 -1205
rect 1285 -1235 1315 -1205
rect 1315 -1235 1316 -1205
rect 1284 -1236 1316 -1235
rect 1284 -1285 1316 -1284
rect 1284 -1315 1285 -1285
rect 1285 -1315 1315 -1285
rect 1315 -1315 1316 -1285
rect 1284 -1316 1316 -1315
rect 1284 -1365 1316 -1364
rect 1284 -1395 1285 -1365
rect 1285 -1395 1315 -1365
rect 1315 -1395 1316 -1365
rect 1284 -1396 1316 -1395
rect 1284 -1445 1316 -1444
rect 1284 -1475 1285 -1445
rect 1285 -1475 1315 -1445
rect 1315 -1475 1316 -1445
rect 1284 -1476 1316 -1475
rect 1284 -1525 1316 -1524
rect 1284 -1555 1285 -1525
rect 1285 -1555 1315 -1525
rect 1315 -1555 1316 -1525
rect 1284 -1556 1316 -1555
rect 1284 -1636 1316 -1604
rect 1284 -1716 1316 -1684
rect 1284 -1765 1316 -1764
rect 1284 -1795 1285 -1765
rect 1285 -1795 1315 -1765
rect 1315 -1795 1316 -1765
rect 1284 -1796 1316 -1795
rect 1284 -1845 1316 -1844
rect 1284 -1875 1285 -1845
rect 1285 -1875 1315 -1845
rect 1315 -1875 1316 -1845
rect 1284 -1876 1316 -1875
rect 1284 -1956 1316 -1924
rect 1284 -2005 1316 -2004
rect 1284 -2035 1285 -2005
rect 1285 -2035 1315 -2005
rect 1315 -2035 1316 -2005
rect 1284 -2036 1316 -2035
rect 1284 -2116 1316 -2084
rect 1284 -2165 1316 -2164
rect 1284 -2195 1285 -2165
rect 1285 -2195 1315 -2165
rect 1315 -2195 1316 -2165
rect 1284 -2196 1316 -2195
rect 1284 -2276 1316 -2244
rect 1284 -2325 1316 -2324
rect 1284 -2355 1285 -2325
rect 1285 -2355 1315 -2325
rect 1315 -2355 1316 -2325
rect 1284 -2356 1316 -2355
rect 1284 -2405 1316 -2404
rect 1284 -2435 1285 -2405
rect 1285 -2435 1315 -2405
rect 1315 -2435 1316 -2405
rect 1284 -2436 1316 -2435
rect 1284 -2485 1316 -2484
rect 1284 -2515 1285 -2485
rect 1285 -2515 1315 -2485
rect 1315 -2515 1316 -2485
rect 1284 -2516 1316 -2515
rect 1284 -2565 1316 -2564
rect 1284 -2595 1285 -2565
rect 1285 -2595 1315 -2565
rect 1315 -2595 1316 -2565
rect 1284 -2596 1316 -2595
rect 1284 -2645 1316 -2644
rect 1284 -2675 1285 -2645
rect 1285 -2675 1315 -2645
rect 1315 -2675 1316 -2645
rect 1284 -2676 1316 -2675
rect 1284 -2725 1316 -2724
rect 1284 -2755 1285 -2725
rect 1285 -2755 1315 -2725
rect 1315 -2755 1316 -2725
rect 1284 -2756 1316 -2755
rect 1284 -2836 1316 -2804
rect 1284 -2885 1316 -2884
rect 1284 -2915 1285 -2885
rect 1285 -2915 1315 -2885
rect 1315 -2915 1316 -2885
rect 1284 -2916 1316 -2915
rect 1284 -2996 1316 -2964
rect 1284 -3045 1316 -3044
rect 1284 -3075 1285 -3045
rect 1285 -3075 1315 -3045
rect 1315 -3075 1316 -3045
rect 1284 -3076 1316 -3075
rect 1284 -3156 1316 -3124
rect 1284 -3205 1316 -3204
rect 1284 -3235 1285 -3205
rect 1285 -3235 1315 -3205
rect 1315 -3235 1316 -3205
rect 1284 -3236 1316 -3235
rect 1284 -3285 1316 -3284
rect 1284 -3315 1285 -3285
rect 1285 -3315 1315 -3285
rect 1315 -3315 1316 -3285
rect 1284 -3316 1316 -3315
rect 1284 -3396 1316 -3364
rect 1284 -3476 1316 -3444
rect 1284 -3525 1316 -3524
rect 1284 -3555 1285 -3525
rect 1285 -3555 1315 -3525
rect 1315 -3555 1316 -3525
rect 1284 -3556 1316 -3555
rect 1284 -3605 1316 -3604
rect 1284 -3635 1285 -3605
rect 1285 -3635 1315 -3605
rect 1315 -3635 1316 -3605
rect 1284 -3636 1316 -3635
rect 1284 -3685 1316 -3684
rect 1284 -3715 1285 -3685
rect 1285 -3715 1315 -3685
rect 1315 -3715 1316 -3685
rect 1284 -3716 1316 -3715
rect 1364 1035 1396 1036
rect 1364 1005 1365 1035
rect 1365 1005 1395 1035
rect 1395 1005 1396 1035
rect 1364 1004 1396 1005
rect 1364 955 1396 956
rect 1364 925 1365 955
rect 1365 925 1395 955
rect 1395 925 1396 955
rect 1364 924 1396 925
rect 1364 875 1396 876
rect 1364 845 1365 875
rect 1365 845 1395 875
rect 1395 845 1396 875
rect 1364 844 1396 845
rect 1364 764 1396 796
rect 1364 684 1396 716
rect 1364 635 1396 636
rect 1364 605 1365 635
rect 1365 605 1395 635
rect 1395 605 1396 635
rect 1364 604 1396 605
rect 1364 555 1396 556
rect 1364 525 1365 555
rect 1365 525 1395 555
rect 1395 525 1396 555
rect 1364 524 1396 525
rect 1364 444 1396 476
rect 1364 395 1396 396
rect 1364 365 1365 395
rect 1365 365 1395 395
rect 1395 365 1396 395
rect 1364 364 1396 365
rect 1364 284 1396 316
rect 1364 235 1396 236
rect 1364 205 1365 235
rect 1365 205 1395 235
rect 1395 205 1396 235
rect 1364 204 1396 205
rect 1364 124 1396 156
rect 1364 75 1396 76
rect 1364 45 1365 75
rect 1365 45 1395 75
rect 1395 45 1396 75
rect 1364 44 1396 45
rect 1364 -5 1396 -4
rect 1364 -35 1365 -5
rect 1365 -35 1395 -5
rect 1395 -35 1396 -5
rect 1364 -36 1396 -35
rect 1364 -85 1396 -84
rect 1364 -115 1365 -85
rect 1365 -115 1395 -85
rect 1395 -115 1396 -85
rect 1364 -116 1396 -115
rect 1364 -165 1396 -164
rect 1364 -195 1365 -165
rect 1365 -195 1395 -165
rect 1395 -195 1396 -165
rect 1364 -196 1396 -195
rect 1364 -245 1396 -244
rect 1364 -275 1365 -245
rect 1365 -275 1395 -245
rect 1395 -275 1396 -245
rect 1364 -276 1396 -275
rect 1364 -325 1396 -324
rect 1364 -355 1365 -325
rect 1365 -355 1395 -325
rect 1395 -355 1396 -325
rect 1364 -356 1396 -355
rect 1364 -436 1396 -404
rect 1364 -485 1396 -484
rect 1364 -515 1365 -485
rect 1365 -515 1395 -485
rect 1395 -515 1396 -485
rect 1364 -516 1396 -515
rect 1364 -596 1396 -564
rect 1364 -645 1396 -644
rect 1364 -675 1365 -645
rect 1365 -675 1395 -645
rect 1395 -675 1396 -645
rect 1364 -676 1396 -675
rect 1364 -756 1396 -724
rect 1364 -805 1396 -804
rect 1364 -835 1365 -805
rect 1365 -835 1395 -805
rect 1395 -835 1396 -805
rect 1364 -836 1396 -835
rect 1364 -885 1396 -884
rect 1364 -915 1365 -885
rect 1365 -915 1395 -885
rect 1395 -915 1396 -885
rect 1364 -916 1396 -915
rect 1364 -996 1396 -964
rect 1364 -1076 1396 -1044
rect 1364 -1125 1396 -1124
rect 1364 -1155 1365 -1125
rect 1365 -1155 1395 -1125
rect 1395 -1155 1396 -1125
rect 1364 -1156 1396 -1155
rect 1364 -1205 1396 -1204
rect 1364 -1235 1365 -1205
rect 1365 -1235 1395 -1205
rect 1395 -1235 1396 -1205
rect 1364 -1236 1396 -1235
rect 1364 -1285 1396 -1284
rect 1364 -1315 1365 -1285
rect 1365 -1315 1395 -1285
rect 1395 -1315 1396 -1285
rect 1364 -1316 1396 -1315
rect 1364 -1365 1396 -1364
rect 1364 -1395 1365 -1365
rect 1365 -1395 1395 -1365
rect 1395 -1395 1396 -1365
rect 1364 -1396 1396 -1395
rect 1364 -1445 1396 -1444
rect 1364 -1475 1365 -1445
rect 1365 -1475 1395 -1445
rect 1395 -1475 1396 -1445
rect 1364 -1476 1396 -1475
rect 1364 -1525 1396 -1524
rect 1364 -1555 1365 -1525
rect 1365 -1555 1395 -1525
rect 1395 -1555 1396 -1525
rect 1364 -1556 1396 -1555
rect 1364 -1636 1396 -1604
rect 1364 -1716 1396 -1684
rect 1364 -1765 1396 -1764
rect 1364 -1795 1365 -1765
rect 1365 -1795 1395 -1765
rect 1395 -1795 1396 -1765
rect 1364 -1796 1396 -1795
rect 1364 -1845 1396 -1844
rect 1364 -1875 1365 -1845
rect 1365 -1875 1395 -1845
rect 1395 -1875 1396 -1845
rect 1364 -1876 1396 -1875
rect 1364 -1956 1396 -1924
rect 1364 -2005 1396 -2004
rect 1364 -2035 1365 -2005
rect 1365 -2035 1395 -2005
rect 1395 -2035 1396 -2005
rect 1364 -2036 1396 -2035
rect 1364 -2116 1396 -2084
rect 1364 -2165 1396 -2164
rect 1364 -2195 1365 -2165
rect 1365 -2195 1395 -2165
rect 1395 -2195 1396 -2165
rect 1364 -2196 1396 -2195
rect 1364 -2276 1396 -2244
rect 1364 -2325 1396 -2324
rect 1364 -2355 1365 -2325
rect 1365 -2355 1395 -2325
rect 1395 -2355 1396 -2325
rect 1364 -2356 1396 -2355
rect 1364 -2405 1396 -2404
rect 1364 -2435 1365 -2405
rect 1365 -2435 1395 -2405
rect 1395 -2435 1396 -2405
rect 1364 -2436 1396 -2435
rect 1364 -2485 1396 -2484
rect 1364 -2515 1365 -2485
rect 1365 -2515 1395 -2485
rect 1395 -2515 1396 -2485
rect 1364 -2516 1396 -2515
rect 1364 -2565 1396 -2564
rect 1364 -2595 1365 -2565
rect 1365 -2595 1395 -2565
rect 1395 -2595 1396 -2565
rect 1364 -2596 1396 -2595
rect 1364 -2645 1396 -2644
rect 1364 -2675 1365 -2645
rect 1365 -2675 1395 -2645
rect 1395 -2675 1396 -2645
rect 1364 -2676 1396 -2675
rect 1364 -2725 1396 -2724
rect 1364 -2755 1365 -2725
rect 1365 -2755 1395 -2725
rect 1395 -2755 1396 -2725
rect 1364 -2756 1396 -2755
rect 1364 -2836 1396 -2804
rect 1364 -2885 1396 -2884
rect 1364 -2915 1365 -2885
rect 1365 -2915 1395 -2885
rect 1395 -2915 1396 -2885
rect 1364 -2916 1396 -2915
rect 1364 -2996 1396 -2964
rect 1364 -3045 1396 -3044
rect 1364 -3075 1365 -3045
rect 1365 -3075 1395 -3045
rect 1395 -3075 1396 -3045
rect 1364 -3076 1396 -3075
rect 1364 -3156 1396 -3124
rect 1364 -3205 1396 -3204
rect 1364 -3235 1365 -3205
rect 1365 -3235 1395 -3205
rect 1395 -3235 1396 -3205
rect 1364 -3236 1396 -3235
rect 1364 -3285 1396 -3284
rect 1364 -3315 1365 -3285
rect 1365 -3315 1395 -3285
rect 1395 -3315 1396 -3285
rect 1364 -3316 1396 -3315
rect 1364 -3396 1396 -3364
rect 1364 -3476 1396 -3444
rect 1364 -3525 1396 -3524
rect 1364 -3555 1365 -3525
rect 1365 -3555 1395 -3525
rect 1395 -3555 1396 -3525
rect 1364 -3556 1396 -3555
rect 1364 -3605 1396 -3604
rect 1364 -3635 1365 -3605
rect 1365 -3635 1395 -3605
rect 1395 -3635 1396 -3605
rect 1364 -3636 1396 -3635
rect 1364 -3685 1396 -3684
rect 1364 -3715 1365 -3685
rect 1365 -3715 1395 -3685
rect 1395 -3715 1396 -3685
rect 1364 -3716 1396 -3715
rect 1444 1035 1476 1036
rect 1444 1005 1445 1035
rect 1445 1005 1475 1035
rect 1475 1005 1476 1035
rect 1444 1004 1476 1005
rect 1444 955 1476 956
rect 1444 925 1445 955
rect 1445 925 1475 955
rect 1475 925 1476 955
rect 1444 924 1476 925
rect 1444 875 1476 876
rect 1444 845 1445 875
rect 1445 845 1475 875
rect 1475 845 1476 875
rect 1444 844 1476 845
rect 1444 764 1476 796
rect 1444 684 1476 716
rect 1444 635 1476 636
rect 1444 605 1445 635
rect 1445 605 1475 635
rect 1475 605 1476 635
rect 1444 604 1476 605
rect 1444 555 1476 556
rect 1444 525 1445 555
rect 1445 525 1475 555
rect 1475 525 1476 555
rect 1444 524 1476 525
rect 1444 444 1476 476
rect 1444 395 1476 396
rect 1444 365 1445 395
rect 1445 365 1475 395
rect 1475 365 1476 395
rect 1444 364 1476 365
rect 1444 284 1476 316
rect 1444 235 1476 236
rect 1444 205 1445 235
rect 1445 205 1475 235
rect 1475 205 1476 235
rect 1444 204 1476 205
rect 1444 124 1476 156
rect 1444 75 1476 76
rect 1444 45 1445 75
rect 1445 45 1475 75
rect 1475 45 1476 75
rect 1444 44 1476 45
rect 1444 -5 1476 -4
rect 1444 -35 1445 -5
rect 1445 -35 1475 -5
rect 1475 -35 1476 -5
rect 1444 -36 1476 -35
rect 1444 -85 1476 -84
rect 1444 -115 1445 -85
rect 1445 -115 1475 -85
rect 1475 -115 1476 -85
rect 1444 -116 1476 -115
rect 1444 -165 1476 -164
rect 1444 -195 1445 -165
rect 1445 -195 1475 -165
rect 1475 -195 1476 -165
rect 1444 -196 1476 -195
rect 1444 -245 1476 -244
rect 1444 -275 1445 -245
rect 1445 -275 1475 -245
rect 1475 -275 1476 -245
rect 1444 -276 1476 -275
rect 1444 -325 1476 -324
rect 1444 -355 1445 -325
rect 1445 -355 1475 -325
rect 1475 -355 1476 -325
rect 1444 -356 1476 -355
rect 1444 -436 1476 -404
rect 1444 -485 1476 -484
rect 1444 -515 1445 -485
rect 1445 -515 1475 -485
rect 1475 -515 1476 -485
rect 1444 -516 1476 -515
rect 1444 -596 1476 -564
rect 1444 -645 1476 -644
rect 1444 -675 1445 -645
rect 1445 -675 1475 -645
rect 1475 -675 1476 -645
rect 1444 -676 1476 -675
rect 1444 -756 1476 -724
rect 1444 -805 1476 -804
rect 1444 -835 1445 -805
rect 1445 -835 1475 -805
rect 1475 -835 1476 -805
rect 1444 -836 1476 -835
rect 1444 -885 1476 -884
rect 1444 -915 1445 -885
rect 1445 -915 1475 -885
rect 1475 -915 1476 -885
rect 1444 -916 1476 -915
rect 1444 -996 1476 -964
rect 1444 -1076 1476 -1044
rect 1444 -1125 1476 -1124
rect 1444 -1155 1445 -1125
rect 1445 -1155 1475 -1125
rect 1475 -1155 1476 -1125
rect 1444 -1156 1476 -1155
rect 1444 -1205 1476 -1204
rect 1444 -1235 1445 -1205
rect 1445 -1235 1475 -1205
rect 1475 -1235 1476 -1205
rect 1444 -1236 1476 -1235
rect 1444 -1285 1476 -1284
rect 1444 -1315 1445 -1285
rect 1445 -1315 1475 -1285
rect 1475 -1315 1476 -1285
rect 1444 -1316 1476 -1315
rect 1444 -1365 1476 -1364
rect 1444 -1395 1445 -1365
rect 1445 -1395 1475 -1365
rect 1475 -1395 1476 -1365
rect 1444 -1396 1476 -1395
rect 1444 -1445 1476 -1444
rect 1444 -1475 1445 -1445
rect 1445 -1475 1475 -1445
rect 1475 -1475 1476 -1445
rect 1444 -1476 1476 -1475
rect 1444 -1525 1476 -1524
rect 1444 -1555 1445 -1525
rect 1445 -1555 1475 -1525
rect 1475 -1555 1476 -1525
rect 1444 -1556 1476 -1555
rect 1444 -1636 1476 -1604
rect 1444 -1716 1476 -1684
rect 1444 -1765 1476 -1764
rect 1444 -1795 1445 -1765
rect 1445 -1795 1475 -1765
rect 1475 -1795 1476 -1765
rect 1444 -1796 1476 -1795
rect 1444 -1845 1476 -1844
rect 1444 -1875 1445 -1845
rect 1445 -1875 1475 -1845
rect 1475 -1875 1476 -1845
rect 1444 -1876 1476 -1875
rect 1444 -1956 1476 -1924
rect 1444 -2005 1476 -2004
rect 1444 -2035 1445 -2005
rect 1445 -2035 1475 -2005
rect 1475 -2035 1476 -2005
rect 1444 -2036 1476 -2035
rect 1444 -2116 1476 -2084
rect 1444 -2165 1476 -2164
rect 1444 -2195 1445 -2165
rect 1445 -2195 1475 -2165
rect 1475 -2195 1476 -2165
rect 1444 -2196 1476 -2195
rect 1444 -2276 1476 -2244
rect 1444 -2325 1476 -2324
rect 1444 -2355 1445 -2325
rect 1445 -2355 1475 -2325
rect 1475 -2355 1476 -2325
rect 1444 -2356 1476 -2355
rect 1444 -2405 1476 -2404
rect 1444 -2435 1445 -2405
rect 1445 -2435 1475 -2405
rect 1475 -2435 1476 -2405
rect 1444 -2436 1476 -2435
rect 1444 -2485 1476 -2484
rect 1444 -2515 1445 -2485
rect 1445 -2515 1475 -2485
rect 1475 -2515 1476 -2485
rect 1444 -2516 1476 -2515
rect 1444 -2565 1476 -2564
rect 1444 -2595 1445 -2565
rect 1445 -2595 1475 -2565
rect 1475 -2595 1476 -2565
rect 1444 -2596 1476 -2595
rect 1444 -2645 1476 -2644
rect 1444 -2675 1445 -2645
rect 1445 -2675 1475 -2645
rect 1475 -2675 1476 -2645
rect 1444 -2676 1476 -2675
rect 1444 -2725 1476 -2724
rect 1444 -2755 1445 -2725
rect 1445 -2755 1475 -2725
rect 1475 -2755 1476 -2725
rect 1444 -2756 1476 -2755
rect 1444 -2836 1476 -2804
rect 1444 -2885 1476 -2884
rect 1444 -2915 1445 -2885
rect 1445 -2915 1475 -2885
rect 1475 -2915 1476 -2885
rect 1444 -2916 1476 -2915
rect 1444 -2996 1476 -2964
rect 1444 -3045 1476 -3044
rect 1444 -3075 1445 -3045
rect 1445 -3075 1475 -3045
rect 1475 -3075 1476 -3045
rect 1444 -3076 1476 -3075
rect 1444 -3156 1476 -3124
rect 1444 -3205 1476 -3204
rect 1444 -3235 1445 -3205
rect 1445 -3235 1475 -3205
rect 1475 -3235 1476 -3205
rect 1444 -3236 1476 -3235
rect 1444 -3285 1476 -3284
rect 1444 -3315 1445 -3285
rect 1445 -3315 1475 -3285
rect 1475 -3315 1476 -3285
rect 1444 -3316 1476 -3315
rect 1444 -3396 1476 -3364
rect 1444 -3476 1476 -3444
rect 1444 -3525 1476 -3524
rect 1444 -3555 1445 -3525
rect 1445 -3555 1475 -3525
rect 1475 -3555 1476 -3525
rect 1444 -3556 1476 -3555
rect 1444 -3605 1476 -3604
rect 1444 -3635 1445 -3605
rect 1445 -3635 1475 -3605
rect 1475 -3635 1476 -3605
rect 1444 -3636 1476 -3635
rect 1444 -3685 1476 -3684
rect 1444 -3715 1445 -3685
rect 1445 -3715 1475 -3685
rect 1475 -3715 1476 -3685
rect 1444 -3716 1476 -3715
rect 1524 1035 1556 1036
rect 1524 1005 1525 1035
rect 1525 1005 1555 1035
rect 1555 1005 1556 1035
rect 1524 1004 1556 1005
rect 1524 955 1556 956
rect 1524 925 1525 955
rect 1525 925 1555 955
rect 1555 925 1556 955
rect 1524 924 1556 925
rect 1524 875 1556 876
rect 1524 845 1525 875
rect 1525 845 1555 875
rect 1555 845 1556 875
rect 1524 844 1556 845
rect 1524 764 1556 796
rect 1524 684 1556 716
rect 1524 635 1556 636
rect 1524 605 1525 635
rect 1525 605 1555 635
rect 1555 605 1556 635
rect 1524 604 1556 605
rect 1524 555 1556 556
rect 1524 525 1525 555
rect 1525 525 1555 555
rect 1555 525 1556 555
rect 1524 524 1556 525
rect 1524 444 1556 476
rect 1524 395 1556 396
rect 1524 365 1525 395
rect 1525 365 1555 395
rect 1555 365 1556 395
rect 1524 364 1556 365
rect 1524 284 1556 316
rect 1524 235 1556 236
rect 1524 205 1525 235
rect 1525 205 1555 235
rect 1555 205 1556 235
rect 1524 204 1556 205
rect 1524 124 1556 156
rect 1524 75 1556 76
rect 1524 45 1525 75
rect 1525 45 1555 75
rect 1555 45 1556 75
rect 1524 44 1556 45
rect 1524 -5 1556 -4
rect 1524 -35 1525 -5
rect 1525 -35 1555 -5
rect 1555 -35 1556 -5
rect 1524 -36 1556 -35
rect 1524 -85 1556 -84
rect 1524 -115 1525 -85
rect 1525 -115 1555 -85
rect 1555 -115 1556 -85
rect 1524 -116 1556 -115
rect 1524 -165 1556 -164
rect 1524 -195 1525 -165
rect 1525 -195 1555 -165
rect 1555 -195 1556 -165
rect 1524 -196 1556 -195
rect 1524 -245 1556 -244
rect 1524 -275 1525 -245
rect 1525 -275 1555 -245
rect 1555 -275 1556 -245
rect 1524 -276 1556 -275
rect 1524 -325 1556 -324
rect 1524 -355 1525 -325
rect 1525 -355 1555 -325
rect 1555 -355 1556 -325
rect 1524 -356 1556 -355
rect 1524 -436 1556 -404
rect 1524 -485 1556 -484
rect 1524 -515 1525 -485
rect 1525 -515 1555 -485
rect 1555 -515 1556 -485
rect 1524 -516 1556 -515
rect 1524 -596 1556 -564
rect 1524 -645 1556 -644
rect 1524 -675 1525 -645
rect 1525 -675 1555 -645
rect 1555 -675 1556 -645
rect 1524 -676 1556 -675
rect 1524 -756 1556 -724
rect 1524 -805 1556 -804
rect 1524 -835 1525 -805
rect 1525 -835 1555 -805
rect 1555 -835 1556 -805
rect 1524 -836 1556 -835
rect 1524 -885 1556 -884
rect 1524 -915 1525 -885
rect 1525 -915 1555 -885
rect 1555 -915 1556 -885
rect 1524 -916 1556 -915
rect 1524 -996 1556 -964
rect 1524 -1076 1556 -1044
rect 1524 -1125 1556 -1124
rect 1524 -1155 1525 -1125
rect 1525 -1155 1555 -1125
rect 1555 -1155 1556 -1125
rect 1524 -1156 1556 -1155
rect 1524 -1205 1556 -1204
rect 1524 -1235 1525 -1205
rect 1525 -1235 1555 -1205
rect 1555 -1235 1556 -1205
rect 1524 -1236 1556 -1235
rect 1524 -1285 1556 -1284
rect 1524 -1315 1525 -1285
rect 1525 -1315 1555 -1285
rect 1555 -1315 1556 -1285
rect 1524 -1316 1556 -1315
rect 1524 -1365 1556 -1364
rect 1524 -1395 1525 -1365
rect 1525 -1395 1555 -1365
rect 1555 -1395 1556 -1365
rect 1524 -1396 1556 -1395
rect 1524 -1445 1556 -1444
rect 1524 -1475 1525 -1445
rect 1525 -1475 1555 -1445
rect 1555 -1475 1556 -1445
rect 1524 -1476 1556 -1475
rect 1524 -1525 1556 -1524
rect 1524 -1555 1525 -1525
rect 1525 -1555 1555 -1525
rect 1555 -1555 1556 -1525
rect 1524 -1556 1556 -1555
rect 1524 -1636 1556 -1604
rect 1524 -1716 1556 -1684
rect 1524 -1765 1556 -1764
rect 1524 -1795 1525 -1765
rect 1525 -1795 1555 -1765
rect 1555 -1795 1556 -1765
rect 1524 -1796 1556 -1795
rect 1524 -1845 1556 -1844
rect 1524 -1875 1525 -1845
rect 1525 -1875 1555 -1845
rect 1555 -1875 1556 -1845
rect 1524 -1876 1556 -1875
rect 1524 -1956 1556 -1924
rect 1524 -2005 1556 -2004
rect 1524 -2035 1525 -2005
rect 1525 -2035 1555 -2005
rect 1555 -2035 1556 -2005
rect 1524 -2036 1556 -2035
rect 1524 -2116 1556 -2084
rect 1524 -2165 1556 -2164
rect 1524 -2195 1525 -2165
rect 1525 -2195 1555 -2165
rect 1555 -2195 1556 -2165
rect 1524 -2196 1556 -2195
rect 1524 -2276 1556 -2244
rect 1524 -2325 1556 -2324
rect 1524 -2355 1525 -2325
rect 1525 -2355 1555 -2325
rect 1555 -2355 1556 -2325
rect 1524 -2356 1556 -2355
rect 1524 -2405 1556 -2404
rect 1524 -2435 1525 -2405
rect 1525 -2435 1555 -2405
rect 1555 -2435 1556 -2405
rect 1524 -2436 1556 -2435
rect 1524 -2485 1556 -2484
rect 1524 -2515 1525 -2485
rect 1525 -2515 1555 -2485
rect 1555 -2515 1556 -2485
rect 1524 -2516 1556 -2515
rect 1524 -2565 1556 -2564
rect 1524 -2595 1525 -2565
rect 1525 -2595 1555 -2565
rect 1555 -2595 1556 -2565
rect 1524 -2596 1556 -2595
rect 1524 -2645 1556 -2644
rect 1524 -2675 1525 -2645
rect 1525 -2675 1555 -2645
rect 1555 -2675 1556 -2645
rect 1524 -2676 1556 -2675
rect 1524 -2725 1556 -2724
rect 1524 -2755 1525 -2725
rect 1525 -2755 1555 -2725
rect 1555 -2755 1556 -2725
rect 1524 -2756 1556 -2755
rect 1524 -2836 1556 -2804
rect 1524 -2885 1556 -2884
rect 1524 -2915 1525 -2885
rect 1525 -2915 1555 -2885
rect 1555 -2915 1556 -2885
rect 1524 -2916 1556 -2915
rect 1524 -2996 1556 -2964
rect 1524 -3045 1556 -3044
rect 1524 -3075 1525 -3045
rect 1525 -3075 1555 -3045
rect 1555 -3075 1556 -3045
rect 1524 -3076 1556 -3075
rect 1524 -3156 1556 -3124
rect 1524 -3205 1556 -3204
rect 1524 -3235 1525 -3205
rect 1525 -3235 1555 -3205
rect 1555 -3235 1556 -3205
rect 1524 -3236 1556 -3235
rect 1524 -3285 1556 -3284
rect 1524 -3315 1525 -3285
rect 1525 -3315 1555 -3285
rect 1555 -3315 1556 -3285
rect 1524 -3316 1556 -3315
rect 1524 -3396 1556 -3364
rect 1524 -3476 1556 -3444
rect 1524 -3525 1556 -3524
rect 1524 -3555 1525 -3525
rect 1525 -3555 1555 -3525
rect 1555 -3555 1556 -3525
rect 1524 -3556 1556 -3555
rect 1524 -3605 1556 -3604
rect 1524 -3635 1525 -3605
rect 1525 -3635 1555 -3605
rect 1555 -3635 1556 -3605
rect 1524 -3636 1556 -3635
rect 1524 -3685 1556 -3684
rect 1524 -3715 1525 -3685
rect 1525 -3715 1555 -3685
rect 1555 -3715 1556 -3685
rect 1524 -3716 1556 -3715
rect 1604 1035 1636 1036
rect 1604 1005 1605 1035
rect 1605 1005 1635 1035
rect 1635 1005 1636 1035
rect 1604 1004 1636 1005
rect 1604 955 1636 956
rect 1604 925 1605 955
rect 1605 925 1635 955
rect 1635 925 1636 955
rect 1604 924 1636 925
rect 1604 875 1636 876
rect 1604 845 1605 875
rect 1605 845 1635 875
rect 1635 845 1636 875
rect 1604 844 1636 845
rect 1604 764 1636 796
rect 1604 684 1636 716
rect 1604 635 1636 636
rect 1604 605 1605 635
rect 1605 605 1635 635
rect 1635 605 1636 635
rect 1604 604 1636 605
rect 1604 555 1636 556
rect 1604 525 1605 555
rect 1605 525 1635 555
rect 1635 525 1636 555
rect 1604 524 1636 525
rect 1604 444 1636 476
rect 1604 395 1636 396
rect 1604 365 1605 395
rect 1605 365 1635 395
rect 1635 365 1636 395
rect 1604 364 1636 365
rect 1604 284 1636 316
rect 1604 235 1636 236
rect 1604 205 1605 235
rect 1605 205 1635 235
rect 1635 205 1636 235
rect 1604 204 1636 205
rect 1604 124 1636 156
rect 1604 75 1636 76
rect 1604 45 1605 75
rect 1605 45 1635 75
rect 1635 45 1636 75
rect 1604 44 1636 45
rect 1604 -5 1636 -4
rect 1604 -35 1605 -5
rect 1605 -35 1635 -5
rect 1635 -35 1636 -5
rect 1604 -36 1636 -35
rect 1604 -85 1636 -84
rect 1604 -115 1605 -85
rect 1605 -115 1635 -85
rect 1635 -115 1636 -85
rect 1604 -116 1636 -115
rect 1604 -165 1636 -164
rect 1604 -195 1605 -165
rect 1605 -195 1635 -165
rect 1635 -195 1636 -165
rect 1604 -196 1636 -195
rect 1604 -245 1636 -244
rect 1604 -275 1605 -245
rect 1605 -275 1635 -245
rect 1635 -275 1636 -245
rect 1604 -276 1636 -275
rect 1604 -325 1636 -324
rect 1604 -355 1605 -325
rect 1605 -355 1635 -325
rect 1635 -355 1636 -325
rect 1604 -356 1636 -355
rect 1604 -436 1636 -404
rect 1604 -485 1636 -484
rect 1604 -515 1605 -485
rect 1605 -515 1635 -485
rect 1635 -515 1636 -485
rect 1604 -516 1636 -515
rect 1604 -596 1636 -564
rect 1604 -645 1636 -644
rect 1604 -675 1605 -645
rect 1605 -675 1635 -645
rect 1635 -675 1636 -645
rect 1604 -676 1636 -675
rect 1604 -756 1636 -724
rect 1604 -805 1636 -804
rect 1604 -835 1605 -805
rect 1605 -835 1635 -805
rect 1635 -835 1636 -805
rect 1604 -836 1636 -835
rect 1604 -885 1636 -884
rect 1604 -915 1605 -885
rect 1605 -915 1635 -885
rect 1635 -915 1636 -885
rect 1604 -916 1636 -915
rect 1604 -996 1636 -964
rect 1604 -1076 1636 -1044
rect 1604 -1125 1636 -1124
rect 1604 -1155 1605 -1125
rect 1605 -1155 1635 -1125
rect 1635 -1155 1636 -1125
rect 1604 -1156 1636 -1155
rect 1604 -1205 1636 -1204
rect 1604 -1235 1605 -1205
rect 1605 -1235 1635 -1205
rect 1635 -1235 1636 -1205
rect 1604 -1236 1636 -1235
rect 1604 -1285 1636 -1284
rect 1604 -1315 1605 -1285
rect 1605 -1315 1635 -1285
rect 1635 -1315 1636 -1285
rect 1604 -1316 1636 -1315
rect 1604 -1365 1636 -1364
rect 1604 -1395 1605 -1365
rect 1605 -1395 1635 -1365
rect 1635 -1395 1636 -1365
rect 1604 -1396 1636 -1395
rect 1604 -1445 1636 -1444
rect 1604 -1475 1605 -1445
rect 1605 -1475 1635 -1445
rect 1635 -1475 1636 -1445
rect 1604 -1476 1636 -1475
rect 1604 -1525 1636 -1524
rect 1604 -1555 1605 -1525
rect 1605 -1555 1635 -1525
rect 1635 -1555 1636 -1525
rect 1604 -1556 1636 -1555
rect 1604 -1636 1636 -1604
rect 1604 -1716 1636 -1684
rect 1604 -1765 1636 -1764
rect 1604 -1795 1605 -1765
rect 1605 -1795 1635 -1765
rect 1635 -1795 1636 -1765
rect 1604 -1796 1636 -1795
rect 1604 -1845 1636 -1844
rect 1604 -1875 1605 -1845
rect 1605 -1875 1635 -1845
rect 1635 -1875 1636 -1845
rect 1604 -1876 1636 -1875
rect 1604 -1956 1636 -1924
rect 1604 -2005 1636 -2004
rect 1604 -2035 1605 -2005
rect 1605 -2035 1635 -2005
rect 1635 -2035 1636 -2005
rect 1604 -2036 1636 -2035
rect 1604 -2116 1636 -2084
rect 1604 -2165 1636 -2164
rect 1604 -2195 1605 -2165
rect 1605 -2195 1635 -2165
rect 1635 -2195 1636 -2165
rect 1604 -2196 1636 -2195
rect 1604 -2276 1636 -2244
rect 1604 -2325 1636 -2324
rect 1604 -2355 1605 -2325
rect 1605 -2355 1635 -2325
rect 1635 -2355 1636 -2325
rect 1604 -2356 1636 -2355
rect 1604 -2405 1636 -2404
rect 1604 -2435 1605 -2405
rect 1605 -2435 1635 -2405
rect 1635 -2435 1636 -2405
rect 1604 -2436 1636 -2435
rect 1604 -2485 1636 -2484
rect 1604 -2515 1605 -2485
rect 1605 -2515 1635 -2485
rect 1635 -2515 1636 -2485
rect 1604 -2516 1636 -2515
rect 1604 -2565 1636 -2564
rect 1604 -2595 1605 -2565
rect 1605 -2595 1635 -2565
rect 1635 -2595 1636 -2565
rect 1604 -2596 1636 -2595
rect 1604 -2645 1636 -2644
rect 1604 -2675 1605 -2645
rect 1605 -2675 1635 -2645
rect 1635 -2675 1636 -2645
rect 1604 -2676 1636 -2675
rect 1604 -2725 1636 -2724
rect 1604 -2755 1605 -2725
rect 1605 -2755 1635 -2725
rect 1635 -2755 1636 -2725
rect 1604 -2756 1636 -2755
rect 1604 -2836 1636 -2804
rect 1604 -2885 1636 -2884
rect 1604 -2915 1605 -2885
rect 1605 -2915 1635 -2885
rect 1635 -2915 1636 -2885
rect 1604 -2916 1636 -2915
rect 1604 -2996 1636 -2964
rect 1604 -3045 1636 -3044
rect 1604 -3075 1605 -3045
rect 1605 -3075 1635 -3045
rect 1635 -3075 1636 -3045
rect 1604 -3076 1636 -3075
rect 1604 -3156 1636 -3124
rect 1604 -3205 1636 -3204
rect 1604 -3235 1605 -3205
rect 1605 -3235 1635 -3205
rect 1635 -3235 1636 -3205
rect 1604 -3236 1636 -3235
rect 1604 -3285 1636 -3284
rect 1604 -3315 1605 -3285
rect 1605 -3315 1635 -3285
rect 1635 -3315 1636 -3285
rect 1604 -3316 1636 -3315
rect 1604 -3396 1636 -3364
rect 1604 -3476 1636 -3444
rect 1604 -3525 1636 -3524
rect 1604 -3555 1605 -3525
rect 1605 -3555 1635 -3525
rect 1635 -3555 1636 -3525
rect 1604 -3556 1636 -3555
rect 1604 -3605 1636 -3604
rect 1604 -3635 1605 -3605
rect 1605 -3635 1635 -3605
rect 1635 -3635 1636 -3605
rect 1604 -3636 1636 -3635
rect 1604 -3685 1636 -3684
rect 1604 -3715 1605 -3685
rect 1605 -3715 1635 -3685
rect 1635 -3715 1636 -3685
rect 1604 -3716 1636 -3715
rect 1684 1035 1716 1036
rect 1684 1005 1685 1035
rect 1685 1005 1715 1035
rect 1715 1005 1716 1035
rect 1684 1004 1716 1005
rect 1684 955 1716 956
rect 1684 925 1685 955
rect 1685 925 1715 955
rect 1715 925 1716 955
rect 1684 924 1716 925
rect 1684 875 1716 876
rect 1684 845 1685 875
rect 1685 845 1715 875
rect 1715 845 1716 875
rect 1684 844 1716 845
rect 1684 764 1716 796
rect 1684 684 1716 716
rect 1684 635 1716 636
rect 1684 605 1685 635
rect 1685 605 1715 635
rect 1715 605 1716 635
rect 1684 604 1716 605
rect 1684 555 1716 556
rect 1684 525 1685 555
rect 1685 525 1715 555
rect 1715 525 1716 555
rect 1684 524 1716 525
rect 1684 444 1716 476
rect 1684 395 1716 396
rect 1684 365 1685 395
rect 1685 365 1715 395
rect 1715 365 1716 395
rect 1684 364 1716 365
rect 1684 284 1716 316
rect 1684 235 1716 236
rect 1684 205 1685 235
rect 1685 205 1715 235
rect 1715 205 1716 235
rect 1684 204 1716 205
rect 1684 124 1716 156
rect 1684 75 1716 76
rect 1684 45 1685 75
rect 1685 45 1715 75
rect 1715 45 1716 75
rect 1684 44 1716 45
rect 1684 -5 1716 -4
rect 1684 -35 1685 -5
rect 1685 -35 1715 -5
rect 1715 -35 1716 -5
rect 1684 -36 1716 -35
rect 1684 -85 1716 -84
rect 1684 -115 1685 -85
rect 1685 -115 1715 -85
rect 1715 -115 1716 -85
rect 1684 -116 1716 -115
rect 1684 -165 1716 -164
rect 1684 -195 1685 -165
rect 1685 -195 1715 -165
rect 1715 -195 1716 -165
rect 1684 -196 1716 -195
rect 1684 -245 1716 -244
rect 1684 -275 1685 -245
rect 1685 -275 1715 -245
rect 1715 -275 1716 -245
rect 1684 -276 1716 -275
rect 1684 -325 1716 -324
rect 1684 -355 1685 -325
rect 1685 -355 1715 -325
rect 1715 -355 1716 -325
rect 1684 -356 1716 -355
rect 1684 -436 1716 -404
rect 1684 -485 1716 -484
rect 1684 -515 1685 -485
rect 1685 -515 1715 -485
rect 1715 -515 1716 -485
rect 1684 -516 1716 -515
rect 1684 -596 1716 -564
rect 1684 -645 1716 -644
rect 1684 -675 1685 -645
rect 1685 -675 1715 -645
rect 1715 -675 1716 -645
rect 1684 -676 1716 -675
rect 1684 -756 1716 -724
rect 1684 -805 1716 -804
rect 1684 -835 1685 -805
rect 1685 -835 1715 -805
rect 1715 -835 1716 -805
rect 1684 -836 1716 -835
rect 1684 -885 1716 -884
rect 1684 -915 1685 -885
rect 1685 -915 1715 -885
rect 1715 -915 1716 -885
rect 1684 -916 1716 -915
rect 1684 -996 1716 -964
rect 1684 -1076 1716 -1044
rect 1684 -1125 1716 -1124
rect 1684 -1155 1685 -1125
rect 1685 -1155 1715 -1125
rect 1715 -1155 1716 -1125
rect 1684 -1156 1716 -1155
rect 1684 -1205 1716 -1204
rect 1684 -1235 1685 -1205
rect 1685 -1235 1715 -1205
rect 1715 -1235 1716 -1205
rect 1684 -1236 1716 -1235
rect 1684 -1285 1716 -1284
rect 1684 -1315 1685 -1285
rect 1685 -1315 1715 -1285
rect 1715 -1315 1716 -1285
rect 1684 -1316 1716 -1315
rect 1684 -1365 1716 -1364
rect 1684 -1395 1685 -1365
rect 1685 -1395 1715 -1365
rect 1715 -1395 1716 -1365
rect 1684 -1396 1716 -1395
rect 1684 -1445 1716 -1444
rect 1684 -1475 1685 -1445
rect 1685 -1475 1715 -1445
rect 1715 -1475 1716 -1445
rect 1684 -1476 1716 -1475
rect 1684 -1525 1716 -1524
rect 1684 -1555 1685 -1525
rect 1685 -1555 1715 -1525
rect 1715 -1555 1716 -1525
rect 1684 -1556 1716 -1555
rect 1684 -1636 1716 -1604
rect 1684 -1716 1716 -1684
rect 1684 -1765 1716 -1764
rect 1684 -1795 1685 -1765
rect 1685 -1795 1715 -1765
rect 1715 -1795 1716 -1765
rect 1684 -1796 1716 -1795
rect 1684 -1845 1716 -1844
rect 1684 -1875 1685 -1845
rect 1685 -1875 1715 -1845
rect 1715 -1875 1716 -1845
rect 1684 -1876 1716 -1875
rect 1684 -1956 1716 -1924
rect 1684 -2005 1716 -2004
rect 1684 -2035 1685 -2005
rect 1685 -2035 1715 -2005
rect 1715 -2035 1716 -2005
rect 1684 -2036 1716 -2035
rect 1684 -2116 1716 -2084
rect 1684 -2165 1716 -2164
rect 1684 -2195 1685 -2165
rect 1685 -2195 1715 -2165
rect 1715 -2195 1716 -2165
rect 1684 -2196 1716 -2195
rect 1684 -2276 1716 -2244
rect 1684 -2325 1716 -2324
rect 1684 -2355 1685 -2325
rect 1685 -2355 1715 -2325
rect 1715 -2355 1716 -2325
rect 1684 -2356 1716 -2355
rect 1684 -2405 1716 -2404
rect 1684 -2435 1685 -2405
rect 1685 -2435 1715 -2405
rect 1715 -2435 1716 -2405
rect 1684 -2436 1716 -2435
rect 1684 -2485 1716 -2484
rect 1684 -2515 1685 -2485
rect 1685 -2515 1715 -2485
rect 1715 -2515 1716 -2485
rect 1684 -2516 1716 -2515
rect 1684 -2565 1716 -2564
rect 1684 -2595 1685 -2565
rect 1685 -2595 1715 -2565
rect 1715 -2595 1716 -2565
rect 1684 -2596 1716 -2595
rect 1684 -2645 1716 -2644
rect 1684 -2675 1685 -2645
rect 1685 -2675 1715 -2645
rect 1715 -2675 1716 -2645
rect 1684 -2676 1716 -2675
rect 1684 -2725 1716 -2724
rect 1684 -2755 1685 -2725
rect 1685 -2755 1715 -2725
rect 1715 -2755 1716 -2725
rect 1684 -2756 1716 -2755
rect 1684 -2836 1716 -2804
rect 1684 -2885 1716 -2884
rect 1684 -2915 1685 -2885
rect 1685 -2915 1715 -2885
rect 1715 -2915 1716 -2885
rect 1684 -2916 1716 -2915
rect 1684 -2996 1716 -2964
rect 1684 -3045 1716 -3044
rect 1684 -3075 1685 -3045
rect 1685 -3075 1715 -3045
rect 1715 -3075 1716 -3045
rect 1684 -3076 1716 -3075
rect 1684 -3156 1716 -3124
rect 1684 -3205 1716 -3204
rect 1684 -3235 1685 -3205
rect 1685 -3235 1715 -3205
rect 1715 -3235 1716 -3205
rect 1684 -3236 1716 -3235
rect 1684 -3285 1716 -3284
rect 1684 -3315 1685 -3285
rect 1685 -3315 1715 -3285
rect 1715 -3315 1716 -3285
rect 1684 -3316 1716 -3315
rect 1684 -3396 1716 -3364
rect 1684 -3476 1716 -3444
rect 1684 -3525 1716 -3524
rect 1684 -3555 1685 -3525
rect 1685 -3555 1715 -3525
rect 1715 -3555 1716 -3525
rect 1684 -3556 1716 -3555
rect 1684 -3605 1716 -3604
rect 1684 -3635 1685 -3605
rect 1685 -3635 1715 -3605
rect 1715 -3635 1716 -3605
rect 1684 -3636 1716 -3635
rect 1684 -3685 1716 -3684
rect 1684 -3715 1685 -3685
rect 1685 -3715 1715 -3685
rect 1715 -3715 1716 -3685
rect 1684 -3716 1716 -3715
rect 1764 1035 1796 1036
rect 1764 1005 1765 1035
rect 1765 1005 1795 1035
rect 1795 1005 1796 1035
rect 1764 1004 1796 1005
rect 1764 955 1796 956
rect 1764 925 1765 955
rect 1765 925 1795 955
rect 1795 925 1796 955
rect 1764 924 1796 925
rect 1764 875 1796 876
rect 1764 845 1765 875
rect 1765 845 1795 875
rect 1795 845 1796 875
rect 1764 844 1796 845
rect 1764 764 1796 796
rect 1764 684 1796 716
rect 1764 635 1796 636
rect 1764 605 1765 635
rect 1765 605 1795 635
rect 1795 605 1796 635
rect 1764 604 1796 605
rect 1764 555 1796 556
rect 1764 525 1765 555
rect 1765 525 1795 555
rect 1795 525 1796 555
rect 1764 524 1796 525
rect 1764 444 1796 476
rect 1764 395 1796 396
rect 1764 365 1765 395
rect 1765 365 1795 395
rect 1795 365 1796 395
rect 1764 364 1796 365
rect 1764 284 1796 316
rect 1764 235 1796 236
rect 1764 205 1765 235
rect 1765 205 1795 235
rect 1795 205 1796 235
rect 1764 204 1796 205
rect 1764 124 1796 156
rect 1764 75 1796 76
rect 1764 45 1765 75
rect 1765 45 1795 75
rect 1795 45 1796 75
rect 1764 44 1796 45
rect 1764 -5 1796 -4
rect 1764 -35 1765 -5
rect 1765 -35 1795 -5
rect 1795 -35 1796 -5
rect 1764 -36 1796 -35
rect 1764 -85 1796 -84
rect 1764 -115 1765 -85
rect 1765 -115 1795 -85
rect 1795 -115 1796 -85
rect 1764 -116 1796 -115
rect 1764 -165 1796 -164
rect 1764 -195 1765 -165
rect 1765 -195 1795 -165
rect 1795 -195 1796 -165
rect 1764 -196 1796 -195
rect 1764 -245 1796 -244
rect 1764 -275 1765 -245
rect 1765 -275 1795 -245
rect 1795 -275 1796 -245
rect 1764 -276 1796 -275
rect 1764 -325 1796 -324
rect 1764 -355 1765 -325
rect 1765 -355 1795 -325
rect 1795 -355 1796 -325
rect 1764 -356 1796 -355
rect 1764 -436 1796 -404
rect 1764 -485 1796 -484
rect 1764 -515 1765 -485
rect 1765 -515 1795 -485
rect 1795 -515 1796 -485
rect 1764 -516 1796 -515
rect 1764 -596 1796 -564
rect 1764 -645 1796 -644
rect 1764 -675 1765 -645
rect 1765 -675 1795 -645
rect 1795 -675 1796 -645
rect 1764 -676 1796 -675
rect 1764 -756 1796 -724
rect 1764 -805 1796 -804
rect 1764 -835 1765 -805
rect 1765 -835 1795 -805
rect 1795 -835 1796 -805
rect 1764 -836 1796 -835
rect 1764 -885 1796 -884
rect 1764 -915 1765 -885
rect 1765 -915 1795 -885
rect 1795 -915 1796 -885
rect 1764 -916 1796 -915
rect 1764 -996 1796 -964
rect 1764 -1076 1796 -1044
rect 1764 -1125 1796 -1124
rect 1764 -1155 1765 -1125
rect 1765 -1155 1795 -1125
rect 1795 -1155 1796 -1125
rect 1764 -1156 1796 -1155
rect 1764 -1205 1796 -1204
rect 1764 -1235 1765 -1205
rect 1765 -1235 1795 -1205
rect 1795 -1235 1796 -1205
rect 1764 -1236 1796 -1235
rect 1764 -1285 1796 -1284
rect 1764 -1315 1765 -1285
rect 1765 -1315 1795 -1285
rect 1795 -1315 1796 -1285
rect 1764 -1316 1796 -1315
rect 1764 -1365 1796 -1364
rect 1764 -1395 1765 -1365
rect 1765 -1395 1795 -1365
rect 1795 -1395 1796 -1365
rect 1764 -1396 1796 -1395
rect 1764 -1445 1796 -1444
rect 1764 -1475 1765 -1445
rect 1765 -1475 1795 -1445
rect 1795 -1475 1796 -1445
rect 1764 -1476 1796 -1475
rect 1764 -1525 1796 -1524
rect 1764 -1555 1765 -1525
rect 1765 -1555 1795 -1525
rect 1795 -1555 1796 -1525
rect 1764 -1556 1796 -1555
rect 1764 -1636 1796 -1604
rect 1764 -1716 1796 -1684
rect 1764 -1765 1796 -1764
rect 1764 -1795 1765 -1765
rect 1765 -1795 1795 -1765
rect 1795 -1795 1796 -1765
rect 1764 -1796 1796 -1795
rect 1764 -1845 1796 -1844
rect 1764 -1875 1765 -1845
rect 1765 -1875 1795 -1845
rect 1795 -1875 1796 -1845
rect 1764 -1876 1796 -1875
rect 1764 -1956 1796 -1924
rect 1764 -2005 1796 -2004
rect 1764 -2035 1765 -2005
rect 1765 -2035 1795 -2005
rect 1795 -2035 1796 -2005
rect 1764 -2036 1796 -2035
rect 1764 -2116 1796 -2084
rect 1764 -2165 1796 -2164
rect 1764 -2195 1765 -2165
rect 1765 -2195 1795 -2165
rect 1795 -2195 1796 -2165
rect 1764 -2196 1796 -2195
rect 1764 -2276 1796 -2244
rect 1764 -2325 1796 -2324
rect 1764 -2355 1765 -2325
rect 1765 -2355 1795 -2325
rect 1795 -2355 1796 -2325
rect 1764 -2356 1796 -2355
rect 1764 -2405 1796 -2404
rect 1764 -2435 1765 -2405
rect 1765 -2435 1795 -2405
rect 1795 -2435 1796 -2405
rect 1764 -2436 1796 -2435
rect 1764 -2485 1796 -2484
rect 1764 -2515 1765 -2485
rect 1765 -2515 1795 -2485
rect 1795 -2515 1796 -2485
rect 1764 -2516 1796 -2515
rect 1764 -2565 1796 -2564
rect 1764 -2595 1765 -2565
rect 1765 -2595 1795 -2565
rect 1795 -2595 1796 -2565
rect 1764 -2596 1796 -2595
rect 1764 -2645 1796 -2644
rect 1764 -2675 1765 -2645
rect 1765 -2675 1795 -2645
rect 1795 -2675 1796 -2645
rect 1764 -2676 1796 -2675
rect 1764 -2725 1796 -2724
rect 1764 -2755 1765 -2725
rect 1765 -2755 1795 -2725
rect 1795 -2755 1796 -2725
rect 1764 -2756 1796 -2755
rect 1764 -2836 1796 -2804
rect 1764 -2885 1796 -2884
rect 1764 -2915 1765 -2885
rect 1765 -2915 1795 -2885
rect 1795 -2915 1796 -2885
rect 1764 -2916 1796 -2915
rect 1764 -2996 1796 -2964
rect 1764 -3045 1796 -3044
rect 1764 -3075 1765 -3045
rect 1765 -3075 1795 -3045
rect 1795 -3075 1796 -3045
rect 1764 -3076 1796 -3075
rect 1764 -3156 1796 -3124
rect 1764 -3205 1796 -3204
rect 1764 -3235 1765 -3205
rect 1765 -3235 1795 -3205
rect 1795 -3235 1796 -3205
rect 1764 -3236 1796 -3235
rect 1764 -3285 1796 -3284
rect 1764 -3315 1765 -3285
rect 1765 -3315 1795 -3285
rect 1795 -3315 1796 -3285
rect 1764 -3316 1796 -3315
rect 1764 -3396 1796 -3364
rect 1764 -3476 1796 -3444
rect 1764 -3525 1796 -3524
rect 1764 -3555 1765 -3525
rect 1765 -3555 1795 -3525
rect 1795 -3555 1796 -3525
rect 1764 -3556 1796 -3555
rect 1764 -3605 1796 -3604
rect 1764 -3635 1765 -3605
rect 1765 -3635 1795 -3605
rect 1795 -3635 1796 -3605
rect 1764 -3636 1796 -3635
rect 1764 -3685 1796 -3684
rect 1764 -3715 1765 -3685
rect 1765 -3715 1795 -3685
rect 1795 -3715 1796 -3685
rect 1764 -3716 1796 -3715
rect 1844 1035 1876 1036
rect 1844 1005 1845 1035
rect 1845 1005 1875 1035
rect 1875 1005 1876 1035
rect 1844 1004 1876 1005
rect 1844 955 1876 956
rect 1844 925 1845 955
rect 1845 925 1875 955
rect 1875 925 1876 955
rect 1844 924 1876 925
rect 1844 875 1876 876
rect 1844 845 1845 875
rect 1845 845 1875 875
rect 1875 845 1876 875
rect 1844 844 1876 845
rect 1844 764 1876 796
rect 1844 684 1876 716
rect 1844 635 1876 636
rect 1844 605 1845 635
rect 1845 605 1875 635
rect 1875 605 1876 635
rect 1844 604 1876 605
rect 1844 555 1876 556
rect 1844 525 1845 555
rect 1845 525 1875 555
rect 1875 525 1876 555
rect 1844 524 1876 525
rect 1844 444 1876 476
rect 1844 395 1876 396
rect 1844 365 1845 395
rect 1845 365 1875 395
rect 1875 365 1876 395
rect 1844 364 1876 365
rect 1844 284 1876 316
rect 1844 235 1876 236
rect 1844 205 1845 235
rect 1845 205 1875 235
rect 1875 205 1876 235
rect 1844 204 1876 205
rect 1844 124 1876 156
rect 1844 75 1876 76
rect 1844 45 1845 75
rect 1845 45 1875 75
rect 1875 45 1876 75
rect 1844 44 1876 45
rect 1844 -5 1876 -4
rect 1844 -35 1845 -5
rect 1845 -35 1875 -5
rect 1875 -35 1876 -5
rect 1844 -36 1876 -35
rect 1844 -85 1876 -84
rect 1844 -115 1845 -85
rect 1845 -115 1875 -85
rect 1875 -115 1876 -85
rect 1844 -116 1876 -115
rect 1844 -165 1876 -164
rect 1844 -195 1845 -165
rect 1845 -195 1875 -165
rect 1875 -195 1876 -165
rect 1844 -196 1876 -195
rect 1844 -245 1876 -244
rect 1844 -275 1845 -245
rect 1845 -275 1875 -245
rect 1875 -275 1876 -245
rect 1844 -276 1876 -275
rect 1844 -325 1876 -324
rect 1844 -355 1845 -325
rect 1845 -355 1875 -325
rect 1875 -355 1876 -325
rect 1844 -356 1876 -355
rect 1844 -436 1876 -404
rect 1844 -485 1876 -484
rect 1844 -515 1845 -485
rect 1845 -515 1875 -485
rect 1875 -515 1876 -485
rect 1844 -516 1876 -515
rect 1844 -596 1876 -564
rect 1844 -645 1876 -644
rect 1844 -675 1845 -645
rect 1845 -675 1875 -645
rect 1875 -675 1876 -645
rect 1844 -676 1876 -675
rect 1844 -756 1876 -724
rect 1844 -805 1876 -804
rect 1844 -835 1845 -805
rect 1845 -835 1875 -805
rect 1875 -835 1876 -805
rect 1844 -836 1876 -835
rect 1844 -885 1876 -884
rect 1844 -915 1845 -885
rect 1845 -915 1875 -885
rect 1875 -915 1876 -885
rect 1844 -916 1876 -915
rect 1844 -996 1876 -964
rect 1844 -1076 1876 -1044
rect 1844 -1125 1876 -1124
rect 1844 -1155 1845 -1125
rect 1845 -1155 1875 -1125
rect 1875 -1155 1876 -1125
rect 1844 -1156 1876 -1155
rect 1844 -1205 1876 -1204
rect 1844 -1235 1845 -1205
rect 1845 -1235 1875 -1205
rect 1875 -1235 1876 -1205
rect 1844 -1236 1876 -1235
rect 1844 -1285 1876 -1284
rect 1844 -1315 1845 -1285
rect 1845 -1315 1875 -1285
rect 1875 -1315 1876 -1285
rect 1844 -1316 1876 -1315
rect 1844 -1365 1876 -1364
rect 1844 -1395 1845 -1365
rect 1845 -1395 1875 -1365
rect 1875 -1395 1876 -1365
rect 1844 -1396 1876 -1395
rect 1844 -1445 1876 -1444
rect 1844 -1475 1845 -1445
rect 1845 -1475 1875 -1445
rect 1875 -1475 1876 -1445
rect 1844 -1476 1876 -1475
rect 1844 -1525 1876 -1524
rect 1844 -1555 1845 -1525
rect 1845 -1555 1875 -1525
rect 1875 -1555 1876 -1525
rect 1844 -1556 1876 -1555
rect 1844 -1636 1876 -1604
rect 1844 -1716 1876 -1684
rect 1844 -1765 1876 -1764
rect 1844 -1795 1845 -1765
rect 1845 -1795 1875 -1765
rect 1875 -1795 1876 -1765
rect 1844 -1796 1876 -1795
rect 1844 -1845 1876 -1844
rect 1844 -1875 1845 -1845
rect 1845 -1875 1875 -1845
rect 1875 -1875 1876 -1845
rect 1844 -1876 1876 -1875
rect 1844 -1956 1876 -1924
rect 1844 -2005 1876 -2004
rect 1844 -2035 1845 -2005
rect 1845 -2035 1875 -2005
rect 1875 -2035 1876 -2005
rect 1844 -2036 1876 -2035
rect 1844 -2116 1876 -2084
rect 1844 -2165 1876 -2164
rect 1844 -2195 1845 -2165
rect 1845 -2195 1875 -2165
rect 1875 -2195 1876 -2165
rect 1844 -2196 1876 -2195
rect 1844 -2276 1876 -2244
rect 1844 -2325 1876 -2324
rect 1844 -2355 1845 -2325
rect 1845 -2355 1875 -2325
rect 1875 -2355 1876 -2325
rect 1844 -2356 1876 -2355
rect 1844 -2405 1876 -2404
rect 1844 -2435 1845 -2405
rect 1845 -2435 1875 -2405
rect 1875 -2435 1876 -2405
rect 1844 -2436 1876 -2435
rect 1844 -2485 1876 -2484
rect 1844 -2515 1845 -2485
rect 1845 -2515 1875 -2485
rect 1875 -2515 1876 -2485
rect 1844 -2516 1876 -2515
rect 1844 -2565 1876 -2564
rect 1844 -2595 1845 -2565
rect 1845 -2595 1875 -2565
rect 1875 -2595 1876 -2565
rect 1844 -2596 1876 -2595
rect 1844 -2645 1876 -2644
rect 1844 -2675 1845 -2645
rect 1845 -2675 1875 -2645
rect 1875 -2675 1876 -2645
rect 1844 -2676 1876 -2675
rect 1844 -2725 1876 -2724
rect 1844 -2755 1845 -2725
rect 1845 -2755 1875 -2725
rect 1875 -2755 1876 -2725
rect 1844 -2756 1876 -2755
rect 1844 -2836 1876 -2804
rect 1844 -2885 1876 -2884
rect 1844 -2915 1845 -2885
rect 1845 -2915 1875 -2885
rect 1875 -2915 1876 -2885
rect 1844 -2916 1876 -2915
rect 1844 -2996 1876 -2964
rect 1844 -3045 1876 -3044
rect 1844 -3075 1845 -3045
rect 1845 -3075 1875 -3045
rect 1875 -3075 1876 -3045
rect 1844 -3076 1876 -3075
rect 1844 -3156 1876 -3124
rect 1844 -3205 1876 -3204
rect 1844 -3235 1845 -3205
rect 1845 -3235 1875 -3205
rect 1875 -3235 1876 -3205
rect 1844 -3236 1876 -3235
rect 1844 -3285 1876 -3284
rect 1844 -3315 1845 -3285
rect 1845 -3315 1875 -3285
rect 1875 -3315 1876 -3285
rect 1844 -3316 1876 -3315
rect 1844 -3396 1876 -3364
rect 1844 -3476 1876 -3444
rect 1844 -3525 1876 -3524
rect 1844 -3555 1845 -3525
rect 1845 -3555 1875 -3525
rect 1875 -3555 1876 -3525
rect 1844 -3556 1876 -3555
rect 1844 -3605 1876 -3604
rect 1844 -3635 1845 -3605
rect 1845 -3635 1875 -3605
rect 1875 -3635 1876 -3605
rect 1844 -3636 1876 -3635
rect 1844 -3685 1876 -3684
rect 1844 -3715 1845 -3685
rect 1845 -3715 1875 -3685
rect 1875 -3715 1876 -3685
rect 1844 -3716 1876 -3715
rect 1924 1035 1956 1036
rect 1924 1005 1925 1035
rect 1925 1005 1955 1035
rect 1955 1005 1956 1035
rect 1924 1004 1956 1005
rect 1924 955 1956 956
rect 1924 925 1925 955
rect 1925 925 1955 955
rect 1955 925 1956 955
rect 1924 924 1956 925
rect 1924 875 1956 876
rect 1924 845 1925 875
rect 1925 845 1955 875
rect 1955 845 1956 875
rect 1924 844 1956 845
rect 1924 764 1956 796
rect 1924 684 1956 716
rect 1924 635 1956 636
rect 1924 605 1925 635
rect 1925 605 1955 635
rect 1955 605 1956 635
rect 1924 604 1956 605
rect 1924 555 1956 556
rect 1924 525 1925 555
rect 1925 525 1955 555
rect 1955 525 1956 555
rect 1924 524 1956 525
rect 1924 444 1956 476
rect 1924 395 1956 396
rect 1924 365 1925 395
rect 1925 365 1955 395
rect 1955 365 1956 395
rect 1924 364 1956 365
rect 1924 284 1956 316
rect 1924 235 1956 236
rect 1924 205 1925 235
rect 1925 205 1955 235
rect 1955 205 1956 235
rect 1924 204 1956 205
rect 1924 124 1956 156
rect 1924 75 1956 76
rect 1924 45 1925 75
rect 1925 45 1955 75
rect 1955 45 1956 75
rect 1924 44 1956 45
rect 1924 -5 1956 -4
rect 1924 -35 1925 -5
rect 1925 -35 1955 -5
rect 1955 -35 1956 -5
rect 1924 -36 1956 -35
rect 1924 -85 1956 -84
rect 1924 -115 1925 -85
rect 1925 -115 1955 -85
rect 1955 -115 1956 -85
rect 1924 -116 1956 -115
rect 1924 -165 1956 -164
rect 1924 -195 1925 -165
rect 1925 -195 1955 -165
rect 1955 -195 1956 -165
rect 1924 -196 1956 -195
rect 1924 -245 1956 -244
rect 1924 -275 1925 -245
rect 1925 -275 1955 -245
rect 1955 -275 1956 -245
rect 1924 -276 1956 -275
rect 1924 -325 1956 -324
rect 1924 -355 1925 -325
rect 1925 -355 1955 -325
rect 1955 -355 1956 -325
rect 1924 -356 1956 -355
rect 1924 -436 1956 -404
rect 1924 -485 1956 -484
rect 1924 -515 1925 -485
rect 1925 -515 1955 -485
rect 1955 -515 1956 -485
rect 1924 -516 1956 -515
rect 1924 -596 1956 -564
rect 1924 -645 1956 -644
rect 1924 -675 1925 -645
rect 1925 -675 1955 -645
rect 1955 -675 1956 -645
rect 1924 -676 1956 -675
rect 1924 -756 1956 -724
rect 1924 -805 1956 -804
rect 1924 -835 1925 -805
rect 1925 -835 1955 -805
rect 1955 -835 1956 -805
rect 1924 -836 1956 -835
rect 1924 -885 1956 -884
rect 1924 -915 1925 -885
rect 1925 -915 1955 -885
rect 1955 -915 1956 -885
rect 1924 -916 1956 -915
rect 1924 -996 1956 -964
rect 1924 -1076 1956 -1044
rect 1924 -1125 1956 -1124
rect 1924 -1155 1925 -1125
rect 1925 -1155 1955 -1125
rect 1955 -1155 1956 -1125
rect 1924 -1156 1956 -1155
rect 1924 -1205 1956 -1204
rect 1924 -1235 1925 -1205
rect 1925 -1235 1955 -1205
rect 1955 -1235 1956 -1205
rect 1924 -1236 1956 -1235
rect 1924 -1285 1956 -1284
rect 1924 -1315 1925 -1285
rect 1925 -1315 1955 -1285
rect 1955 -1315 1956 -1285
rect 1924 -1316 1956 -1315
rect 1924 -1365 1956 -1364
rect 1924 -1395 1925 -1365
rect 1925 -1395 1955 -1365
rect 1955 -1395 1956 -1365
rect 1924 -1396 1956 -1395
rect 1924 -1445 1956 -1444
rect 1924 -1475 1925 -1445
rect 1925 -1475 1955 -1445
rect 1955 -1475 1956 -1445
rect 1924 -1476 1956 -1475
rect 1924 -1525 1956 -1524
rect 1924 -1555 1925 -1525
rect 1925 -1555 1955 -1525
rect 1955 -1555 1956 -1525
rect 1924 -1556 1956 -1555
rect 1924 -1636 1956 -1604
rect 1924 -1716 1956 -1684
rect 1924 -1765 1956 -1764
rect 1924 -1795 1925 -1765
rect 1925 -1795 1955 -1765
rect 1955 -1795 1956 -1765
rect 1924 -1796 1956 -1795
rect 1924 -1845 1956 -1844
rect 1924 -1875 1925 -1845
rect 1925 -1875 1955 -1845
rect 1955 -1875 1956 -1845
rect 1924 -1876 1956 -1875
rect 1924 -1956 1956 -1924
rect 1924 -2005 1956 -2004
rect 1924 -2035 1925 -2005
rect 1925 -2035 1955 -2005
rect 1955 -2035 1956 -2005
rect 1924 -2036 1956 -2035
rect 1924 -2116 1956 -2084
rect 1924 -2165 1956 -2164
rect 1924 -2195 1925 -2165
rect 1925 -2195 1955 -2165
rect 1955 -2195 1956 -2165
rect 1924 -2196 1956 -2195
rect 1924 -2276 1956 -2244
rect 1924 -2325 1956 -2324
rect 1924 -2355 1925 -2325
rect 1925 -2355 1955 -2325
rect 1955 -2355 1956 -2325
rect 1924 -2356 1956 -2355
rect 1924 -2405 1956 -2404
rect 1924 -2435 1925 -2405
rect 1925 -2435 1955 -2405
rect 1955 -2435 1956 -2405
rect 1924 -2436 1956 -2435
rect 1924 -2485 1956 -2484
rect 1924 -2515 1925 -2485
rect 1925 -2515 1955 -2485
rect 1955 -2515 1956 -2485
rect 1924 -2516 1956 -2515
rect 1924 -2565 1956 -2564
rect 1924 -2595 1925 -2565
rect 1925 -2595 1955 -2565
rect 1955 -2595 1956 -2565
rect 1924 -2596 1956 -2595
rect 1924 -2645 1956 -2644
rect 1924 -2675 1925 -2645
rect 1925 -2675 1955 -2645
rect 1955 -2675 1956 -2645
rect 1924 -2676 1956 -2675
rect 1924 -2725 1956 -2724
rect 1924 -2755 1925 -2725
rect 1925 -2755 1955 -2725
rect 1955 -2755 1956 -2725
rect 1924 -2756 1956 -2755
rect 1924 -2836 1956 -2804
rect 1924 -2885 1956 -2884
rect 1924 -2915 1925 -2885
rect 1925 -2915 1955 -2885
rect 1955 -2915 1956 -2885
rect 1924 -2916 1956 -2915
rect 1924 -2996 1956 -2964
rect 1924 -3045 1956 -3044
rect 1924 -3075 1925 -3045
rect 1925 -3075 1955 -3045
rect 1955 -3075 1956 -3045
rect 1924 -3076 1956 -3075
rect 1924 -3156 1956 -3124
rect 1924 -3205 1956 -3204
rect 1924 -3235 1925 -3205
rect 1925 -3235 1955 -3205
rect 1955 -3235 1956 -3205
rect 1924 -3236 1956 -3235
rect 1924 -3285 1956 -3284
rect 1924 -3315 1925 -3285
rect 1925 -3315 1955 -3285
rect 1955 -3315 1956 -3285
rect 1924 -3316 1956 -3315
rect 1924 -3396 1956 -3364
rect 1924 -3476 1956 -3444
rect 1924 -3525 1956 -3524
rect 1924 -3555 1925 -3525
rect 1925 -3555 1955 -3525
rect 1955 -3555 1956 -3525
rect 1924 -3556 1956 -3555
rect 1924 -3605 1956 -3604
rect 1924 -3635 1925 -3605
rect 1925 -3635 1955 -3605
rect 1955 -3635 1956 -3605
rect 1924 -3636 1956 -3635
rect 1924 -3685 1956 -3684
rect 1924 -3715 1925 -3685
rect 1925 -3715 1955 -3685
rect 1955 -3715 1956 -3685
rect 1924 -3716 1956 -3715
rect 2004 1035 2036 1036
rect 2004 1005 2005 1035
rect 2005 1005 2035 1035
rect 2035 1005 2036 1035
rect 2004 1004 2036 1005
rect 2004 955 2036 956
rect 2004 925 2005 955
rect 2005 925 2035 955
rect 2035 925 2036 955
rect 2004 924 2036 925
rect 2004 875 2036 876
rect 2004 845 2005 875
rect 2005 845 2035 875
rect 2035 845 2036 875
rect 2004 844 2036 845
rect 2004 764 2036 796
rect 2004 684 2036 716
rect 2004 635 2036 636
rect 2004 605 2005 635
rect 2005 605 2035 635
rect 2035 605 2036 635
rect 2004 604 2036 605
rect 2004 555 2036 556
rect 2004 525 2005 555
rect 2005 525 2035 555
rect 2035 525 2036 555
rect 2004 524 2036 525
rect 2004 444 2036 476
rect 2004 395 2036 396
rect 2004 365 2005 395
rect 2005 365 2035 395
rect 2035 365 2036 395
rect 2004 364 2036 365
rect 2004 284 2036 316
rect 2004 235 2036 236
rect 2004 205 2005 235
rect 2005 205 2035 235
rect 2035 205 2036 235
rect 2004 204 2036 205
rect 2004 124 2036 156
rect 2004 75 2036 76
rect 2004 45 2005 75
rect 2005 45 2035 75
rect 2035 45 2036 75
rect 2004 44 2036 45
rect 2004 -5 2036 -4
rect 2004 -35 2005 -5
rect 2005 -35 2035 -5
rect 2035 -35 2036 -5
rect 2004 -36 2036 -35
rect 2004 -85 2036 -84
rect 2004 -115 2005 -85
rect 2005 -115 2035 -85
rect 2035 -115 2036 -85
rect 2004 -116 2036 -115
rect 2004 -165 2036 -164
rect 2004 -195 2005 -165
rect 2005 -195 2035 -165
rect 2035 -195 2036 -165
rect 2004 -196 2036 -195
rect 2004 -245 2036 -244
rect 2004 -275 2005 -245
rect 2005 -275 2035 -245
rect 2035 -275 2036 -245
rect 2004 -276 2036 -275
rect 2004 -325 2036 -324
rect 2004 -355 2005 -325
rect 2005 -355 2035 -325
rect 2035 -355 2036 -325
rect 2004 -356 2036 -355
rect 2004 -436 2036 -404
rect 2004 -485 2036 -484
rect 2004 -515 2005 -485
rect 2005 -515 2035 -485
rect 2035 -515 2036 -485
rect 2004 -516 2036 -515
rect 2004 -596 2036 -564
rect 2004 -645 2036 -644
rect 2004 -675 2005 -645
rect 2005 -675 2035 -645
rect 2035 -675 2036 -645
rect 2004 -676 2036 -675
rect 2004 -756 2036 -724
rect 2004 -805 2036 -804
rect 2004 -835 2005 -805
rect 2005 -835 2035 -805
rect 2035 -835 2036 -805
rect 2004 -836 2036 -835
rect 2004 -885 2036 -884
rect 2004 -915 2005 -885
rect 2005 -915 2035 -885
rect 2035 -915 2036 -885
rect 2004 -916 2036 -915
rect 2004 -996 2036 -964
rect 2004 -1076 2036 -1044
rect 2004 -1125 2036 -1124
rect 2004 -1155 2005 -1125
rect 2005 -1155 2035 -1125
rect 2035 -1155 2036 -1125
rect 2004 -1156 2036 -1155
rect 2004 -1205 2036 -1204
rect 2004 -1235 2005 -1205
rect 2005 -1235 2035 -1205
rect 2035 -1235 2036 -1205
rect 2004 -1236 2036 -1235
rect 2004 -1285 2036 -1284
rect 2004 -1315 2005 -1285
rect 2005 -1315 2035 -1285
rect 2035 -1315 2036 -1285
rect 2004 -1316 2036 -1315
rect 2004 -1365 2036 -1364
rect 2004 -1395 2005 -1365
rect 2005 -1395 2035 -1365
rect 2035 -1395 2036 -1365
rect 2004 -1396 2036 -1395
rect 2004 -1445 2036 -1444
rect 2004 -1475 2005 -1445
rect 2005 -1475 2035 -1445
rect 2035 -1475 2036 -1445
rect 2004 -1476 2036 -1475
rect 2004 -1525 2036 -1524
rect 2004 -1555 2005 -1525
rect 2005 -1555 2035 -1525
rect 2035 -1555 2036 -1525
rect 2004 -1556 2036 -1555
rect 2004 -1636 2036 -1604
rect 2004 -1716 2036 -1684
rect 2004 -1765 2036 -1764
rect 2004 -1795 2005 -1765
rect 2005 -1795 2035 -1765
rect 2035 -1795 2036 -1765
rect 2004 -1796 2036 -1795
rect 2004 -1845 2036 -1844
rect 2004 -1875 2005 -1845
rect 2005 -1875 2035 -1845
rect 2035 -1875 2036 -1845
rect 2004 -1876 2036 -1875
rect 2004 -1956 2036 -1924
rect 2004 -2005 2036 -2004
rect 2004 -2035 2005 -2005
rect 2005 -2035 2035 -2005
rect 2035 -2035 2036 -2005
rect 2004 -2036 2036 -2035
rect 2004 -2116 2036 -2084
rect 2004 -2165 2036 -2164
rect 2004 -2195 2005 -2165
rect 2005 -2195 2035 -2165
rect 2035 -2195 2036 -2165
rect 2004 -2196 2036 -2195
rect 2004 -2276 2036 -2244
rect 2004 -2325 2036 -2324
rect 2004 -2355 2005 -2325
rect 2005 -2355 2035 -2325
rect 2035 -2355 2036 -2325
rect 2004 -2356 2036 -2355
rect 2004 -2405 2036 -2404
rect 2004 -2435 2005 -2405
rect 2005 -2435 2035 -2405
rect 2035 -2435 2036 -2405
rect 2004 -2436 2036 -2435
rect 2004 -2485 2036 -2484
rect 2004 -2515 2005 -2485
rect 2005 -2515 2035 -2485
rect 2035 -2515 2036 -2485
rect 2004 -2516 2036 -2515
rect 2004 -2565 2036 -2564
rect 2004 -2595 2005 -2565
rect 2005 -2595 2035 -2565
rect 2035 -2595 2036 -2565
rect 2004 -2596 2036 -2595
rect 2004 -2645 2036 -2644
rect 2004 -2675 2005 -2645
rect 2005 -2675 2035 -2645
rect 2035 -2675 2036 -2645
rect 2004 -2676 2036 -2675
rect 2004 -2725 2036 -2724
rect 2004 -2755 2005 -2725
rect 2005 -2755 2035 -2725
rect 2035 -2755 2036 -2725
rect 2004 -2756 2036 -2755
rect 2004 -2836 2036 -2804
rect 2004 -2885 2036 -2884
rect 2004 -2915 2005 -2885
rect 2005 -2915 2035 -2885
rect 2035 -2915 2036 -2885
rect 2004 -2916 2036 -2915
rect 2004 -2996 2036 -2964
rect 2004 -3045 2036 -3044
rect 2004 -3075 2005 -3045
rect 2005 -3075 2035 -3045
rect 2035 -3075 2036 -3045
rect 2004 -3076 2036 -3075
rect 2004 -3156 2036 -3124
rect 2004 -3205 2036 -3204
rect 2004 -3235 2005 -3205
rect 2005 -3235 2035 -3205
rect 2035 -3235 2036 -3205
rect 2004 -3236 2036 -3235
rect 2004 -3285 2036 -3284
rect 2004 -3315 2005 -3285
rect 2005 -3315 2035 -3285
rect 2035 -3315 2036 -3285
rect 2004 -3316 2036 -3315
rect 2004 -3396 2036 -3364
rect 2004 -3476 2036 -3444
rect 2004 -3525 2036 -3524
rect 2004 -3555 2005 -3525
rect 2005 -3555 2035 -3525
rect 2035 -3555 2036 -3525
rect 2004 -3556 2036 -3555
rect 2004 -3605 2036 -3604
rect 2004 -3635 2005 -3605
rect 2005 -3635 2035 -3605
rect 2035 -3635 2036 -3605
rect 2004 -3636 2036 -3635
rect 2004 -3685 2036 -3684
rect 2004 -3715 2005 -3685
rect 2005 -3715 2035 -3685
rect 2035 -3715 2036 -3685
rect 2004 -3716 2036 -3715
rect 2084 1035 2116 1036
rect 2084 1005 2085 1035
rect 2085 1005 2115 1035
rect 2115 1005 2116 1035
rect 2084 1004 2116 1005
rect 2084 955 2116 956
rect 2084 925 2085 955
rect 2085 925 2115 955
rect 2115 925 2116 955
rect 2084 924 2116 925
rect 2084 875 2116 876
rect 2084 845 2085 875
rect 2085 845 2115 875
rect 2115 845 2116 875
rect 2084 844 2116 845
rect 2084 764 2116 796
rect 2084 684 2116 716
rect 2084 635 2116 636
rect 2084 605 2085 635
rect 2085 605 2115 635
rect 2115 605 2116 635
rect 2084 604 2116 605
rect 2084 555 2116 556
rect 2084 525 2085 555
rect 2085 525 2115 555
rect 2115 525 2116 555
rect 2084 524 2116 525
rect 2084 444 2116 476
rect 2084 395 2116 396
rect 2084 365 2085 395
rect 2085 365 2115 395
rect 2115 365 2116 395
rect 2084 364 2116 365
rect 2084 284 2116 316
rect 2084 235 2116 236
rect 2084 205 2085 235
rect 2085 205 2115 235
rect 2115 205 2116 235
rect 2084 204 2116 205
rect 2084 124 2116 156
rect 2084 75 2116 76
rect 2084 45 2085 75
rect 2085 45 2115 75
rect 2115 45 2116 75
rect 2084 44 2116 45
rect 2084 -5 2116 -4
rect 2084 -35 2085 -5
rect 2085 -35 2115 -5
rect 2115 -35 2116 -5
rect 2084 -36 2116 -35
rect 2084 -85 2116 -84
rect 2084 -115 2085 -85
rect 2085 -115 2115 -85
rect 2115 -115 2116 -85
rect 2084 -116 2116 -115
rect 2084 -165 2116 -164
rect 2084 -195 2085 -165
rect 2085 -195 2115 -165
rect 2115 -195 2116 -165
rect 2084 -196 2116 -195
rect 2084 -245 2116 -244
rect 2084 -275 2085 -245
rect 2085 -275 2115 -245
rect 2115 -275 2116 -245
rect 2084 -276 2116 -275
rect 2084 -325 2116 -324
rect 2084 -355 2085 -325
rect 2085 -355 2115 -325
rect 2115 -355 2116 -325
rect 2084 -356 2116 -355
rect 2084 -436 2116 -404
rect 2084 -485 2116 -484
rect 2084 -515 2085 -485
rect 2085 -515 2115 -485
rect 2115 -515 2116 -485
rect 2084 -516 2116 -515
rect 2084 -596 2116 -564
rect 2084 -645 2116 -644
rect 2084 -675 2085 -645
rect 2085 -675 2115 -645
rect 2115 -675 2116 -645
rect 2084 -676 2116 -675
rect 2084 -756 2116 -724
rect 2084 -805 2116 -804
rect 2084 -835 2085 -805
rect 2085 -835 2115 -805
rect 2115 -835 2116 -805
rect 2084 -836 2116 -835
rect 2084 -885 2116 -884
rect 2084 -915 2085 -885
rect 2085 -915 2115 -885
rect 2115 -915 2116 -885
rect 2084 -916 2116 -915
rect 2084 -996 2116 -964
rect 2084 -1076 2116 -1044
rect 2084 -1125 2116 -1124
rect 2084 -1155 2085 -1125
rect 2085 -1155 2115 -1125
rect 2115 -1155 2116 -1125
rect 2084 -1156 2116 -1155
rect 2084 -1205 2116 -1204
rect 2084 -1235 2085 -1205
rect 2085 -1235 2115 -1205
rect 2115 -1235 2116 -1205
rect 2084 -1236 2116 -1235
rect 2084 -1285 2116 -1284
rect 2084 -1315 2085 -1285
rect 2085 -1315 2115 -1285
rect 2115 -1315 2116 -1285
rect 2084 -1316 2116 -1315
rect 2084 -1365 2116 -1364
rect 2084 -1395 2085 -1365
rect 2085 -1395 2115 -1365
rect 2115 -1395 2116 -1365
rect 2084 -1396 2116 -1395
rect 2084 -1445 2116 -1444
rect 2084 -1475 2085 -1445
rect 2085 -1475 2115 -1445
rect 2115 -1475 2116 -1445
rect 2084 -1476 2116 -1475
rect 2084 -1525 2116 -1524
rect 2084 -1555 2085 -1525
rect 2085 -1555 2115 -1525
rect 2115 -1555 2116 -1525
rect 2084 -1556 2116 -1555
rect 2084 -1636 2116 -1604
rect 2084 -1716 2116 -1684
rect 2084 -1765 2116 -1764
rect 2084 -1795 2085 -1765
rect 2085 -1795 2115 -1765
rect 2115 -1795 2116 -1765
rect 2084 -1796 2116 -1795
rect 2084 -1845 2116 -1844
rect 2084 -1875 2085 -1845
rect 2085 -1875 2115 -1845
rect 2115 -1875 2116 -1845
rect 2084 -1876 2116 -1875
rect 2084 -1956 2116 -1924
rect 2084 -2005 2116 -2004
rect 2084 -2035 2085 -2005
rect 2085 -2035 2115 -2005
rect 2115 -2035 2116 -2005
rect 2084 -2036 2116 -2035
rect 2084 -2116 2116 -2084
rect 2084 -2165 2116 -2164
rect 2084 -2195 2085 -2165
rect 2085 -2195 2115 -2165
rect 2115 -2195 2116 -2165
rect 2084 -2196 2116 -2195
rect 2084 -2276 2116 -2244
rect 2084 -2325 2116 -2324
rect 2084 -2355 2085 -2325
rect 2085 -2355 2115 -2325
rect 2115 -2355 2116 -2325
rect 2084 -2356 2116 -2355
rect 2084 -2405 2116 -2404
rect 2084 -2435 2085 -2405
rect 2085 -2435 2115 -2405
rect 2115 -2435 2116 -2405
rect 2084 -2436 2116 -2435
rect 2084 -2485 2116 -2484
rect 2084 -2515 2085 -2485
rect 2085 -2515 2115 -2485
rect 2115 -2515 2116 -2485
rect 2084 -2516 2116 -2515
rect 2084 -2565 2116 -2564
rect 2084 -2595 2085 -2565
rect 2085 -2595 2115 -2565
rect 2115 -2595 2116 -2565
rect 2084 -2596 2116 -2595
rect 2084 -2645 2116 -2644
rect 2084 -2675 2085 -2645
rect 2085 -2675 2115 -2645
rect 2115 -2675 2116 -2645
rect 2084 -2676 2116 -2675
rect 2084 -2725 2116 -2724
rect 2084 -2755 2085 -2725
rect 2085 -2755 2115 -2725
rect 2115 -2755 2116 -2725
rect 2084 -2756 2116 -2755
rect 2084 -2836 2116 -2804
rect 2084 -2885 2116 -2884
rect 2084 -2915 2085 -2885
rect 2085 -2915 2115 -2885
rect 2115 -2915 2116 -2885
rect 2084 -2916 2116 -2915
rect 2084 -2996 2116 -2964
rect 2084 -3045 2116 -3044
rect 2084 -3075 2085 -3045
rect 2085 -3075 2115 -3045
rect 2115 -3075 2116 -3045
rect 2084 -3076 2116 -3075
rect 2084 -3156 2116 -3124
rect 2084 -3205 2116 -3204
rect 2084 -3235 2085 -3205
rect 2085 -3235 2115 -3205
rect 2115 -3235 2116 -3205
rect 2084 -3236 2116 -3235
rect 2084 -3285 2116 -3284
rect 2084 -3315 2085 -3285
rect 2085 -3315 2115 -3285
rect 2115 -3315 2116 -3285
rect 2084 -3316 2116 -3315
rect 2084 -3396 2116 -3364
rect 2084 -3476 2116 -3444
rect 2084 -3525 2116 -3524
rect 2084 -3555 2085 -3525
rect 2085 -3555 2115 -3525
rect 2115 -3555 2116 -3525
rect 2084 -3556 2116 -3555
rect 2084 -3605 2116 -3604
rect 2084 -3635 2085 -3605
rect 2085 -3635 2115 -3605
rect 2115 -3635 2116 -3605
rect 2084 -3636 2116 -3635
rect 2084 -3685 2116 -3684
rect 2084 -3715 2085 -3685
rect 2085 -3715 2115 -3685
rect 2115 -3715 2116 -3685
rect 2084 -3716 2116 -3715
rect 2164 1035 2196 1036
rect 2164 1005 2165 1035
rect 2165 1005 2195 1035
rect 2195 1005 2196 1035
rect 2164 1004 2196 1005
rect 2164 955 2196 956
rect 2164 925 2165 955
rect 2165 925 2195 955
rect 2195 925 2196 955
rect 2164 924 2196 925
rect 2164 875 2196 876
rect 2164 845 2165 875
rect 2165 845 2195 875
rect 2195 845 2196 875
rect 2164 844 2196 845
rect 2164 764 2196 796
rect 2164 684 2196 716
rect 2164 635 2196 636
rect 2164 605 2165 635
rect 2165 605 2195 635
rect 2195 605 2196 635
rect 2164 604 2196 605
rect 2164 555 2196 556
rect 2164 525 2165 555
rect 2165 525 2195 555
rect 2195 525 2196 555
rect 2164 524 2196 525
rect 2164 444 2196 476
rect 2164 395 2196 396
rect 2164 365 2165 395
rect 2165 365 2195 395
rect 2195 365 2196 395
rect 2164 364 2196 365
rect 2164 284 2196 316
rect 2164 235 2196 236
rect 2164 205 2165 235
rect 2165 205 2195 235
rect 2195 205 2196 235
rect 2164 204 2196 205
rect 2164 124 2196 156
rect 2164 75 2196 76
rect 2164 45 2165 75
rect 2165 45 2195 75
rect 2195 45 2196 75
rect 2164 44 2196 45
rect 2164 -5 2196 -4
rect 2164 -35 2165 -5
rect 2165 -35 2195 -5
rect 2195 -35 2196 -5
rect 2164 -36 2196 -35
rect 2164 -85 2196 -84
rect 2164 -115 2165 -85
rect 2165 -115 2195 -85
rect 2195 -115 2196 -85
rect 2164 -116 2196 -115
rect 2164 -165 2196 -164
rect 2164 -195 2165 -165
rect 2165 -195 2195 -165
rect 2195 -195 2196 -165
rect 2164 -196 2196 -195
rect 2164 -245 2196 -244
rect 2164 -275 2165 -245
rect 2165 -275 2195 -245
rect 2195 -275 2196 -245
rect 2164 -276 2196 -275
rect 2164 -325 2196 -324
rect 2164 -355 2165 -325
rect 2165 -355 2195 -325
rect 2195 -355 2196 -325
rect 2164 -356 2196 -355
rect 2164 -436 2196 -404
rect 2164 -485 2196 -484
rect 2164 -515 2165 -485
rect 2165 -515 2195 -485
rect 2195 -515 2196 -485
rect 2164 -516 2196 -515
rect 2164 -596 2196 -564
rect 2164 -645 2196 -644
rect 2164 -675 2165 -645
rect 2165 -675 2195 -645
rect 2195 -675 2196 -645
rect 2164 -676 2196 -675
rect 2164 -756 2196 -724
rect 2164 -805 2196 -804
rect 2164 -835 2165 -805
rect 2165 -835 2195 -805
rect 2195 -835 2196 -805
rect 2164 -836 2196 -835
rect 2164 -885 2196 -884
rect 2164 -915 2165 -885
rect 2165 -915 2195 -885
rect 2195 -915 2196 -885
rect 2164 -916 2196 -915
rect 2164 -996 2196 -964
rect 2164 -1076 2196 -1044
rect 2164 -1125 2196 -1124
rect 2164 -1155 2165 -1125
rect 2165 -1155 2195 -1125
rect 2195 -1155 2196 -1125
rect 2164 -1156 2196 -1155
rect 2164 -1205 2196 -1204
rect 2164 -1235 2165 -1205
rect 2165 -1235 2195 -1205
rect 2195 -1235 2196 -1205
rect 2164 -1236 2196 -1235
rect 2164 -1285 2196 -1284
rect 2164 -1315 2165 -1285
rect 2165 -1315 2195 -1285
rect 2195 -1315 2196 -1285
rect 2164 -1316 2196 -1315
rect 2164 -1365 2196 -1364
rect 2164 -1395 2165 -1365
rect 2165 -1395 2195 -1365
rect 2195 -1395 2196 -1365
rect 2164 -1396 2196 -1395
rect 2164 -1445 2196 -1444
rect 2164 -1475 2165 -1445
rect 2165 -1475 2195 -1445
rect 2195 -1475 2196 -1445
rect 2164 -1476 2196 -1475
rect 2164 -1525 2196 -1524
rect 2164 -1555 2165 -1525
rect 2165 -1555 2195 -1525
rect 2195 -1555 2196 -1525
rect 2164 -1556 2196 -1555
rect 2164 -1636 2196 -1604
rect 2164 -1716 2196 -1684
rect 2164 -1765 2196 -1764
rect 2164 -1795 2165 -1765
rect 2165 -1795 2195 -1765
rect 2195 -1795 2196 -1765
rect 2164 -1796 2196 -1795
rect 2164 -1845 2196 -1844
rect 2164 -1875 2165 -1845
rect 2165 -1875 2195 -1845
rect 2195 -1875 2196 -1845
rect 2164 -1876 2196 -1875
rect 2164 -1956 2196 -1924
rect 2164 -2005 2196 -2004
rect 2164 -2035 2165 -2005
rect 2165 -2035 2195 -2005
rect 2195 -2035 2196 -2005
rect 2164 -2036 2196 -2035
rect 2164 -2116 2196 -2084
rect 2164 -2165 2196 -2164
rect 2164 -2195 2165 -2165
rect 2165 -2195 2195 -2165
rect 2195 -2195 2196 -2165
rect 2164 -2196 2196 -2195
rect 2164 -2276 2196 -2244
rect 2164 -2325 2196 -2324
rect 2164 -2355 2165 -2325
rect 2165 -2355 2195 -2325
rect 2195 -2355 2196 -2325
rect 2164 -2356 2196 -2355
rect 2164 -2405 2196 -2404
rect 2164 -2435 2165 -2405
rect 2165 -2435 2195 -2405
rect 2195 -2435 2196 -2405
rect 2164 -2436 2196 -2435
rect 2164 -2485 2196 -2484
rect 2164 -2515 2165 -2485
rect 2165 -2515 2195 -2485
rect 2195 -2515 2196 -2485
rect 2164 -2516 2196 -2515
rect 2164 -2565 2196 -2564
rect 2164 -2595 2165 -2565
rect 2165 -2595 2195 -2565
rect 2195 -2595 2196 -2565
rect 2164 -2596 2196 -2595
rect 2164 -2645 2196 -2644
rect 2164 -2675 2165 -2645
rect 2165 -2675 2195 -2645
rect 2195 -2675 2196 -2645
rect 2164 -2676 2196 -2675
rect 2164 -2725 2196 -2724
rect 2164 -2755 2165 -2725
rect 2165 -2755 2195 -2725
rect 2195 -2755 2196 -2725
rect 2164 -2756 2196 -2755
rect 2164 -2836 2196 -2804
rect 2164 -2885 2196 -2884
rect 2164 -2915 2165 -2885
rect 2165 -2915 2195 -2885
rect 2195 -2915 2196 -2885
rect 2164 -2916 2196 -2915
rect 2164 -2996 2196 -2964
rect 2164 -3045 2196 -3044
rect 2164 -3075 2165 -3045
rect 2165 -3075 2195 -3045
rect 2195 -3075 2196 -3045
rect 2164 -3076 2196 -3075
rect 2164 -3156 2196 -3124
rect 2164 -3205 2196 -3204
rect 2164 -3235 2165 -3205
rect 2165 -3235 2195 -3205
rect 2195 -3235 2196 -3205
rect 2164 -3236 2196 -3235
rect 2164 -3285 2196 -3284
rect 2164 -3315 2165 -3285
rect 2165 -3315 2195 -3285
rect 2195 -3315 2196 -3285
rect 2164 -3316 2196 -3315
rect 2164 -3396 2196 -3364
rect 2164 -3476 2196 -3444
rect 2164 -3525 2196 -3524
rect 2164 -3555 2165 -3525
rect 2165 -3555 2195 -3525
rect 2195 -3555 2196 -3525
rect 2164 -3556 2196 -3555
rect 2164 -3605 2196 -3604
rect 2164 -3635 2165 -3605
rect 2165 -3635 2195 -3605
rect 2195 -3635 2196 -3605
rect 2164 -3636 2196 -3635
rect 2164 -3685 2196 -3684
rect 2164 -3715 2165 -3685
rect 2165 -3715 2195 -3685
rect 2195 -3715 2196 -3685
rect 2164 -3716 2196 -3715
rect 2244 1035 2276 1036
rect 2244 1005 2245 1035
rect 2245 1005 2275 1035
rect 2275 1005 2276 1035
rect 2244 1004 2276 1005
rect 2244 955 2276 956
rect 2244 925 2245 955
rect 2245 925 2275 955
rect 2275 925 2276 955
rect 2244 924 2276 925
rect 2244 875 2276 876
rect 2244 845 2245 875
rect 2245 845 2275 875
rect 2275 845 2276 875
rect 2244 844 2276 845
rect 2244 764 2276 796
rect 2244 684 2276 716
rect 2244 635 2276 636
rect 2244 605 2245 635
rect 2245 605 2275 635
rect 2275 605 2276 635
rect 2244 604 2276 605
rect 2244 555 2276 556
rect 2244 525 2245 555
rect 2245 525 2275 555
rect 2275 525 2276 555
rect 2244 524 2276 525
rect 2244 444 2276 476
rect 2244 395 2276 396
rect 2244 365 2245 395
rect 2245 365 2275 395
rect 2275 365 2276 395
rect 2244 364 2276 365
rect 2244 284 2276 316
rect 2244 235 2276 236
rect 2244 205 2245 235
rect 2245 205 2275 235
rect 2275 205 2276 235
rect 2244 204 2276 205
rect 2244 124 2276 156
rect 2244 75 2276 76
rect 2244 45 2245 75
rect 2245 45 2275 75
rect 2275 45 2276 75
rect 2244 44 2276 45
rect 2244 -5 2276 -4
rect 2244 -35 2245 -5
rect 2245 -35 2275 -5
rect 2275 -35 2276 -5
rect 2244 -36 2276 -35
rect 2244 -85 2276 -84
rect 2244 -115 2245 -85
rect 2245 -115 2275 -85
rect 2275 -115 2276 -85
rect 2244 -116 2276 -115
rect 2244 -165 2276 -164
rect 2244 -195 2245 -165
rect 2245 -195 2275 -165
rect 2275 -195 2276 -165
rect 2244 -196 2276 -195
rect 2244 -245 2276 -244
rect 2244 -275 2245 -245
rect 2245 -275 2275 -245
rect 2275 -275 2276 -245
rect 2244 -276 2276 -275
rect 2244 -325 2276 -324
rect 2244 -355 2245 -325
rect 2245 -355 2275 -325
rect 2275 -355 2276 -325
rect 2244 -356 2276 -355
rect 2244 -436 2276 -404
rect 2244 -485 2276 -484
rect 2244 -515 2245 -485
rect 2245 -515 2275 -485
rect 2275 -515 2276 -485
rect 2244 -516 2276 -515
rect 2244 -596 2276 -564
rect 2244 -645 2276 -644
rect 2244 -675 2245 -645
rect 2245 -675 2275 -645
rect 2275 -675 2276 -645
rect 2244 -676 2276 -675
rect 2244 -756 2276 -724
rect 2244 -805 2276 -804
rect 2244 -835 2245 -805
rect 2245 -835 2275 -805
rect 2275 -835 2276 -805
rect 2244 -836 2276 -835
rect 2244 -885 2276 -884
rect 2244 -915 2245 -885
rect 2245 -915 2275 -885
rect 2275 -915 2276 -885
rect 2244 -916 2276 -915
rect 2244 -996 2276 -964
rect 2244 -1076 2276 -1044
rect 2244 -1125 2276 -1124
rect 2244 -1155 2245 -1125
rect 2245 -1155 2275 -1125
rect 2275 -1155 2276 -1125
rect 2244 -1156 2276 -1155
rect 2244 -1205 2276 -1204
rect 2244 -1235 2245 -1205
rect 2245 -1235 2275 -1205
rect 2275 -1235 2276 -1205
rect 2244 -1236 2276 -1235
rect 2244 -1285 2276 -1284
rect 2244 -1315 2245 -1285
rect 2245 -1315 2275 -1285
rect 2275 -1315 2276 -1285
rect 2244 -1316 2276 -1315
rect 2244 -1365 2276 -1364
rect 2244 -1395 2245 -1365
rect 2245 -1395 2275 -1365
rect 2275 -1395 2276 -1365
rect 2244 -1396 2276 -1395
rect 2244 -1445 2276 -1444
rect 2244 -1475 2245 -1445
rect 2245 -1475 2275 -1445
rect 2275 -1475 2276 -1445
rect 2244 -1476 2276 -1475
rect 2244 -1525 2276 -1524
rect 2244 -1555 2245 -1525
rect 2245 -1555 2275 -1525
rect 2275 -1555 2276 -1525
rect 2244 -1556 2276 -1555
rect 2244 -1636 2276 -1604
rect 2244 -1716 2276 -1684
rect 2244 -1765 2276 -1764
rect 2244 -1795 2245 -1765
rect 2245 -1795 2275 -1765
rect 2275 -1795 2276 -1765
rect 2244 -1796 2276 -1795
rect 2244 -1845 2276 -1844
rect 2244 -1875 2245 -1845
rect 2245 -1875 2275 -1845
rect 2275 -1875 2276 -1845
rect 2244 -1876 2276 -1875
rect 2244 -1956 2276 -1924
rect 2244 -2005 2276 -2004
rect 2244 -2035 2245 -2005
rect 2245 -2035 2275 -2005
rect 2275 -2035 2276 -2005
rect 2244 -2036 2276 -2035
rect 2244 -2116 2276 -2084
rect 2244 -2165 2276 -2164
rect 2244 -2195 2245 -2165
rect 2245 -2195 2275 -2165
rect 2275 -2195 2276 -2165
rect 2244 -2196 2276 -2195
rect 2244 -2276 2276 -2244
rect 2244 -2325 2276 -2324
rect 2244 -2355 2245 -2325
rect 2245 -2355 2275 -2325
rect 2275 -2355 2276 -2325
rect 2244 -2356 2276 -2355
rect 2244 -2405 2276 -2404
rect 2244 -2435 2245 -2405
rect 2245 -2435 2275 -2405
rect 2275 -2435 2276 -2405
rect 2244 -2436 2276 -2435
rect 2244 -2485 2276 -2484
rect 2244 -2515 2245 -2485
rect 2245 -2515 2275 -2485
rect 2275 -2515 2276 -2485
rect 2244 -2516 2276 -2515
rect 2244 -2565 2276 -2564
rect 2244 -2595 2245 -2565
rect 2245 -2595 2275 -2565
rect 2275 -2595 2276 -2565
rect 2244 -2596 2276 -2595
rect 2244 -2645 2276 -2644
rect 2244 -2675 2245 -2645
rect 2245 -2675 2275 -2645
rect 2275 -2675 2276 -2645
rect 2244 -2676 2276 -2675
rect 2244 -2725 2276 -2724
rect 2244 -2755 2245 -2725
rect 2245 -2755 2275 -2725
rect 2275 -2755 2276 -2725
rect 2244 -2756 2276 -2755
rect 2244 -2836 2276 -2804
rect 2244 -2885 2276 -2884
rect 2244 -2915 2245 -2885
rect 2245 -2915 2275 -2885
rect 2275 -2915 2276 -2885
rect 2244 -2916 2276 -2915
rect 2244 -2996 2276 -2964
rect 2244 -3045 2276 -3044
rect 2244 -3075 2245 -3045
rect 2245 -3075 2275 -3045
rect 2275 -3075 2276 -3045
rect 2244 -3076 2276 -3075
rect 2244 -3156 2276 -3124
rect 2244 -3205 2276 -3204
rect 2244 -3235 2245 -3205
rect 2245 -3235 2275 -3205
rect 2275 -3235 2276 -3205
rect 2244 -3236 2276 -3235
rect 2244 -3285 2276 -3284
rect 2244 -3315 2245 -3285
rect 2245 -3315 2275 -3285
rect 2275 -3315 2276 -3285
rect 2244 -3316 2276 -3315
rect 2244 -3396 2276 -3364
rect 2244 -3476 2276 -3444
rect 2244 -3525 2276 -3524
rect 2244 -3555 2245 -3525
rect 2245 -3555 2275 -3525
rect 2275 -3555 2276 -3525
rect 2244 -3556 2276 -3555
rect 2244 -3605 2276 -3604
rect 2244 -3635 2245 -3605
rect 2245 -3635 2275 -3605
rect 2275 -3635 2276 -3605
rect 2244 -3636 2276 -3635
rect 2244 -3685 2276 -3684
rect 2244 -3715 2245 -3685
rect 2245 -3715 2275 -3685
rect 2275 -3715 2276 -3685
rect 2244 -3716 2276 -3715
rect 2324 1035 2356 1036
rect 2324 1005 2325 1035
rect 2325 1005 2355 1035
rect 2355 1005 2356 1035
rect 2324 1004 2356 1005
rect 2324 955 2356 956
rect 2324 925 2325 955
rect 2325 925 2355 955
rect 2355 925 2356 955
rect 2324 924 2356 925
rect 2324 875 2356 876
rect 2324 845 2325 875
rect 2325 845 2355 875
rect 2355 845 2356 875
rect 2324 844 2356 845
rect 2324 764 2356 796
rect 2324 684 2356 716
rect 2324 635 2356 636
rect 2324 605 2325 635
rect 2325 605 2355 635
rect 2355 605 2356 635
rect 2324 604 2356 605
rect 2324 555 2356 556
rect 2324 525 2325 555
rect 2325 525 2355 555
rect 2355 525 2356 555
rect 2324 524 2356 525
rect 2324 444 2356 476
rect 2324 395 2356 396
rect 2324 365 2325 395
rect 2325 365 2355 395
rect 2355 365 2356 395
rect 2324 364 2356 365
rect 2324 284 2356 316
rect 2324 235 2356 236
rect 2324 205 2325 235
rect 2325 205 2355 235
rect 2355 205 2356 235
rect 2324 204 2356 205
rect 2324 124 2356 156
rect 2324 75 2356 76
rect 2324 45 2325 75
rect 2325 45 2355 75
rect 2355 45 2356 75
rect 2324 44 2356 45
rect 2324 -5 2356 -4
rect 2324 -35 2325 -5
rect 2325 -35 2355 -5
rect 2355 -35 2356 -5
rect 2324 -36 2356 -35
rect 2324 -85 2356 -84
rect 2324 -115 2325 -85
rect 2325 -115 2355 -85
rect 2355 -115 2356 -85
rect 2324 -116 2356 -115
rect 2324 -165 2356 -164
rect 2324 -195 2325 -165
rect 2325 -195 2355 -165
rect 2355 -195 2356 -165
rect 2324 -196 2356 -195
rect 2324 -245 2356 -244
rect 2324 -275 2325 -245
rect 2325 -275 2355 -245
rect 2355 -275 2356 -245
rect 2324 -276 2356 -275
rect 2324 -325 2356 -324
rect 2324 -355 2325 -325
rect 2325 -355 2355 -325
rect 2355 -355 2356 -325
rect 2324 -356 2356 -355
rect 2324 -436 2356 -404
rect 2324 -485 2356 -484
rect 2324 -515 2325 -485
rect 2325 -515 2355 -485
rect 2355 -515 2356 -485
rect 2324 -516 2356 -515
rect 2324 -596 2356 -564
rect 2324 -645 2356 -644
rect 2324 -675 2325 -645
rect 2325 -675 2355 -645
rect 2355 -675 2356 -645
rect 2324 -676 2356 -675
rect 2324 -756 2356 -724
rect 2324 -805 2356 -804
rect 2324 -835 2325 -805
rect 2325 -835 2355 -805
rect 2355 -835 2356 -805
rect 2324 -836 2356 -835
rect 2324 -885 2356 -884
rect 2324 -915 2325 -885
rect 2325 -915 2355 -885
rect 2355 -915 2356 -885
rect 2324 -916 2356 -915
rect 2324 -996 2356 -964
rect 2324 -1076 2356 -1044
rect 2324 -1125 2356 -1124
rect 2324 -1155 2325 -1125
rect 2325 -1155 2355 -1125
rect 2355 -1155 2356 -1125
rect 2324 -1156 2356 -1155
rect 2324 -1205 2356 -1204
rect 2324 -1235 2325 -1205
rect 2325 -1235 2355 -1205
rect 2355 -1235 2356 -1205
rect 2324 -1236 2356 -1235
rect 2324 -1285 2356 -1284
rect 2324 -1315 2325 -1285
rect 2325 -1315 2355 -1285
rect 2355 -1315 2356 -1285
rect 2324 -1316 2356 -1315
rect 2324 -1365 2356 -1364
rect 2324 -1395 2325 -1365
rect 2325 -1395 2355 -1365
rect 2355 -1395 2356 -1365
rect 2324 -1396 2356 -1395
rect 2324 -1445 2356 -1444
rect 2324 -1475 2325 -1445
rect 2325 -1475 2355 -1445
rect 2355 -1475 2356 -1445
rect 2324 -1476 2356 -1475
rect 2324 -1525 2356 -1524
rect 2324 -1555 2325 -1525
rect 2325 -1555 2355 -1525
rect 2355 -1555 2356 -1525
rect 2324 -1556 2356 -1555
rect 2324 -1636 2356 -1604
rect 2324 -1716 2356 -1684
rect 2324 -1765 2356 -1764
rect 2324 -1795 2325 -1765
rect 2325 -1795 2355 -1765
rect 2355 -1795 2356 -1765
rect 2324 -1796 2356 -1795
rect 2324 -1845 2356 -1844
rect 2324 -1875 2325 -1845
rect 2325 -1875 2355 -1845
rect 2355 -1875 2356 -1845
rect 2324 -1876 2356 -1875
rect 2324 -1956 2356 -1924
rect 2324 -2005 2356 -2004
rect 2324 -2035 2325 -2005
rect 2325 -2035 2355 -2005
rect 2355 -2035 2356 -2005
rect 2324 -2036 2356 -2035
rect 2324 -2116 2356 -2084
rect 2324 -2165 2356 -2164
rect 2324 -2195 2325 -2165
rect 2325 -2195 2355 -2165
rect 2355 -2195 2356 -2165
rect 2324 -2196 2356 -2195
rect 2324 -2276 2356 -2244
rect 2324 -2325 2356 -2324
rect 2324 -2355 2325 -2325
rect 2325 -2355 2355 -2325
rect 2355 -2355 2356 -2325
rect 2324 -2356 2356 -2355
rect 2324 -2405 2356 -2404
rect 2324 -2435 2325 -2405
rect 2325 -2435 2355 -2405
rect 2355 -2435 2356 -2405
rect 2324 -2436 2356 -2435
rect 2324 -2485 2356 -2484
rect 2324 -2515 2325 -2485
rect 2325 -2515 2355 -2485
rect 2355 -2515 2356 -2485
rect 2324 -2516 2356 -2515
rect 2324 -2565 2356 -2564
rect 2324 -2595 2325 -2565
rect 2325 -2595 2355 -2565
rect 2355 -2595 2356 -2565
rect 2324 -2596 2356 -2595
rect 2324 -2645 2356 -2644
rect 2324 -2675 2325 -2645
rect 2325 -2675 2355 -2645
rect 2355 -2675 2356 -2645
rect 2324 -2676 2356 -2675
rect 2324 -2725 2356 -2724
rect 2324 -2755 2325 -2725
rect 2325 -2755 2355 -2725
rect 2355 -2755 2356 -2725
rect 2324 -2756 2356 -2755
rect 2324 -2836 2356 -2804
rect 2324 -2885 2356 -2884
rect 2324 -2915 2325 -2885
rect 2325 -2915 2355 -2885
rect 2355 -2915 2356 -2885
rect 2324 -2916 2356 -2915
rect 2324 -2996 2356 -2964
rect 2324 -3045 2356 -3044
rect 2324 -3075 2325 -3045
rect 2325 -3075 2355 -3045
rect 2355 -3075 2356 -3045
rect 2324 -3076 2356 -3075
rect 2324 -3156 2356 -3124
rect 2324 -3205 2356 -3204
rect 2324 -3235 2325 -3205
rect 2325 -3235 2355 -3205
rect 2355 -3235 2356 -3205
rect 2324 -3236 2356 -3235
rect 2324 -3285 2356 -3284
rect 2324 -3315 2325 -3285
rect 2325 -3315 2355 -3285
rect 2355 -3315 2356 -3285
rect 2324 -3316 2356 -3315
rect 2324 -3396 2356 -3364
rect 2324 -3476 2356 -3444
rect 2324 -3525 2356 -3524
rect 2324 -3555 2325 -3525
rect 2325 -3555 2355 -3525
rect 2355 -3555 2356 -3525
rect 2324 -3556 2356 -3555
rect 2324 -3605 2356 -3604
rect 2324 -3635 2325 -3605
rect 2325 -3635 2355 -3605
rect 2355 -3635 2356 -3605
rect 2324 -3636 2356 -3635
rect 2324 -3685 2356 -3684
rect 2324 -3715 2325 -3685
rect 2325 -3715 2355 -3685
rect 2355 -3715 2356 -3685
rect 2324 -3716 2356 -3715
rect 2404 1035 2436 1036
rect 2404 1005 2405 1035
rect 2405 1005 2435 1035
rect 2435 1005 2436 1035
rect 2404 1004 2436 1005
rect 2404 955 2436 956
rect 2404 925 2405 955
rect 2405 925 2435 955
rect 2435 925 2436 955
rect 2404 924 2436 925
rect 2404 875 2436 876
rect 2404 845 2405 875
rect 2405 845 2435 875
rect 2435 845 2436 875
rect 2404 844 2436 845
rect 2404 764 2436 796
rect 2404 684 2436 716
rect 2404 635 2436 636
rect 2404 605 2405 635
rect 2405 605 2435 635
rect 2435 605 2436 635
rect 2404 604 2436 605
rect 2404 555 2436 556
rect 2404 525 2405 555
rect 2405 525 2435 555
rect 2435 525 2436 555
rect 2404 524 2436 525
rect 2404 444 2436 476
rect 2404 395 2436 396
rect 2404 365 2405 395
rect 2405 365 2435 395
rect 2435 365 2436 395
rect 2404 364 2436 365
rect 2404 284 2436 316
rect 2404 235 2436 236
rect 2404 205 2405 235
rect 2405 205 2435 235
rect 2435 205 2436 235
rect 2404 204 2436 205
rect 2404 124 2436 156
rect 2404 75 2436 76
rect 2404 45 2405 75
rect 2405 45 2435 75
rect 2435 45 2436 75
rect 2404 44 2436 45
rect 2404 -5 2436 -4
rect 2404 -35 2405 -5
rect 2405 -35 2435 -5
rect 2435 -35 2436 -5
rect 2404 -36 2436 -35
rect 2404 -85 2436 -84
rect 2404 -115 2405 -85
rect 2405 -115 2435 -85
rect 2435 -115 2436 -85
rect 2404 -116 2436 -115
rect 2404 -165 2436 -164
rect 2404 -195 2405 -165
rect 2405 -195 2435 -165
rect 2435 -195 2436 -165
rect 2404 -196 2436 -195
rect 2404 -245 2436 -244
rect 2404 -275 2405 -245
rect 2405 -275 2435 -245
rect 2435 -275 2436 -245
rect 2404 -276 2436 -275
rect 2404 -325 2436 -324
rect 2404 -355 2405 -325
rect 2405 -355 2435 -325
rect 2435 -355 2436 -325
rect 2404 -356 2436 -355
rect 2404 -436 2436 -404
rect 2404 -485 2436 -484
rect 2404 -515 2405 -485
rect 2405 -515 2435 -485
rect 2435 -515 2436 -485
rect 2404 -516 2436 -515
rect 2404 -596 2436 -564
rect 2404 -645 2436 -644
rect 2404 -675 2405 -645
rect 2405 -675 2435 -645
rect 2435 -675 2436 -645
rect 2404 -676 2436 -675
rect 2404 -756 2436 -724
rect 2404 -805 2436 -804
rect 2404 -835 2405 -805
rect 2405 -835 2435 -805
rect 2435 -835 2436 -805
rect 2404 -836 2436 -835
rect 2404 -885 2436 -884
rect 2404 -915 2405 -885
rect 2405 -915 2435 -885
rect 2435 -915 2436 -885
rect 2404 -916 2436 -915
rect 2404 -996 2436 -964
rect 2404 -1076 2436 -1044
rect 2404 -1125 2436 -1124
rect 2404 -1155 2405 -1125
rect 2405 -1155 2435 -1125
rect 2435 -1155 2436 -1125
rect 2404 -1156 2436 -1155
rect 2404 -1205 2436 -1204
rect 2404 -1235 2405 -1205
rect 2405 -1235 2435 -1205
rect 2435 -1235 2436 -1205
rect 2404 -1236 2436 -1235
rect 2404 -1285 2436 -1284
rect 2404 -1315 2405 -1285
rect 2405 -1315 2435 -1285
rect 2435 -1315 2436 -1285
rect 2404 -1316 2436 -1315
rect 2404 -1365 2436 -1364
rect 2404 -1395 2405 -1365
rect 2405 -1395 2435 -1365
rect 2435 -1395 2436 -1365
rect 2404 -1396 2436 -1395
rect 2404 -1445 2436 -1444
rect 2404 -1475 2405 -1445
rect 2405 -1475 2435 -1445
rect 2435 -1475 2436 -1445
rect 2404 -1476 2436 -1475
rect 2404 -1525 2436 -1524
rect 2404 -1555 2405 -1525
rect 2405 -1555 2435 -1525
rect 2435 -1555 2436 -1525
rect 2404 -1556 2436 -1555
rect 2404 -1636 2436 -1604
rect 2404 -1716 2436 -1684
rect 2404 -1765 2436 -1764
rect 2404 -1795 2405 -1765
rect 2405 -1795 2435 -1765
rect 2435 -1795 2436 -1765
rect 2404 -1796 2436 -1795
rect 2404 -1845 2436 -1844
rect 2404 -1875 2405 -1845
rect 2405 -1875 2435 -1845
rect 2435 -1875 2436 -1845
rect 2404 -1876 2436 -1875
rect 2404 -1956 2436 -1924
rect 2404 -2005 2436 -2004
rect 2404 -2035 2405 -2005
rect 2405 -2035 2435 -2005
rect 2435 -2035 2436 -2005
rect 2404 -2036 2436 -2035
rect 2404 -2116 2436 -2084
rect 2404 -2165 2436 -2164
rect 2404 -2195 2405 -2165
rect 2405 -2195 2435 -2165
rect 2435 -2195 2436 -2165
rect 2404 -2196 2436 -2195
rect 2404 -2276 2436 -2244
rect 2404 -2325 2436 -2324
rect 2404 -2355 2405 -2325
rect 2405 -2355 2435 -2325
rect 2435 -2355 2436 -2325
rect 2404 -2356 2436 -2355
rect 2404 -2405 2436 -2404
rect 2404 -2435 2405 -2405
rect 2405 -2435 2435 -2405
rect 2435 -2435 2436 -2405
rect 2404 -2436 2436 -2435
rect 2404 -2485 2436 -2484
rect 2404 -2515 2405 -2485
rect 2405 -2515 2435 -2485
rect 2435 -2515 2436 -2485
rect 2404 -2516 2436 -2515
rect 2404 -2565 2436 -2564
rect 2404 -2595 2405 -2565
rect 2405 -2595 2435 -2565
rect 2435 -2595 2436 -2565
rect 2404 -2596 2436 -2595
rect 2404 -2645 2436 -2644
rect 2404 -2675 2405 -2645
rect 2405 -2675 2435 -2645
rect 2435 -2675 2436 -2645
rect 2404 -2676 2436 -2675
rect 2404 -2725 2436 -2724
rect 2404 -2755 2405 -2725
rect 2405 -2755 2435 -2725
rect 2435 -2755 2436 -2725
rect 2404 -2756 2436 -2755
rect 2404 -2836 2436 -2804
rect 2404 -2885 2436 -2884
rect 2404 -2915 2405 -2885
rect 2405 -2915 2435 -2885
rect 2435 -2915 2436 -2885
rect 2404 -2916 2436 -2915
rect 2404 -2996 2436 -2964
rect 2404 -3045 2436 -3044
rect 2404 -3075 2405 -3045
rect 2405 -3075 2435 -3045
rect 2435 -3075 2436 -3045
rect 2404 -3076 2436 -3075
rect 2404 -3156 2436 -3124
rect 2404 -3205 2436 -3204
rect 2404 -3235 2405 -3205
rect 2405 -3235 2435 -3205
rect 2435 -3235 2436 -3205
rect 2404 -3236 2436 -3235
rect 2404 -3285 2436 -3284
rect 2404 -3315 2405 -3285
rect 2405 -3315 2435 -3285
rect 2435 -3315 2436 -3285
rect 2404 -3316 2436 -3315
rect 2404 -3396 2436 -3364
rect 2404 -3476 2436 -3444
rect 2404 -3525 2436 -3524
rect 2404 -3555 2405 -3525
rect 2405 -3555 2435 -3525
rect 2435 -3555 2436 -3525
rect 2404 -3556 2436 -3555
rect 2404 -3605 2436 -3604
rect 2404 -3635 2405 -3605
rect 2405 -3635 2435 -3605
rect 2435 -3635 2436 -3605
rect 2404 -3636 2436 -3635
rect 2404 -3685 2436 -3684
rect 2404 -3715 2405 -3685
rect 2405 -3715 2435 -3685
rect 2435 -3715 2436 -3685
rect 2404 -3716 2436 -3715
rect 2484 1035 2516 1036
rect 2484 1005 2485 1035
rect 2485 1005 2515 1035
rect 2515 1005 2516 1035
rect 2484 1004 2516 1005
rect 2484 955 2516 956
rect 2484 925 2485 955
rect 2485 925 2515 955
rect 2515 925 2516 955
rect 2484 924 2516 925
rect 2484 875 2516 876
rect 2484 845 2485 875
rect 2485 845 2515 875
rect 2515 845 2516 875
rect 2484 844 2516 845
rect 2484 764 2516 796
rect 2484 684 2516 716
rect 2484 635 2516 636
rect 2484 605 2485 635
rect 2485 605 2515 635
rect 2515 605 2516 635
rect 2484 604 2516 605
rect 2484 555 2516 556
rect 2484 525 2485 555
rect 2485 525 2515 555
rect 2515 525 2516 555
rect 2484 524 2516 525
rect 2484 444 2516 476
rect 2484 395 2516 396
rect 2484 365 2485 395
rect 2485 365 2515 395
rect 2515 365 2516 395
rect 2484 364 2516 365
rect 2484 284 2516 316
rect 2484 235 2516 236
rect 2484 205 2485 235
rect 2485 205 2515 235
rect 2515 205 2516 235
rect 2484 204 2516 205
rect 2484 124 2516 156
rect 2484 75 2516 76
rect 2484 45 2485 75
rect 2485 45 2515 75
rect 2515 45 2516 75
rect 2484 44 2516 45
rect 2484 -5 2516 -4
rect 2484 -35 2485 -5
rect 2485 -35 2515 -5
rect 2515 -35 2516 -5
rect 2484 -36 2516 -35
rect 2484 -85 2516 -84
rect 2484 -115 2485 -85
rect 2485 -115 2515 -85
rect 2515 -115 2516 -85
rect 2484 -116 2516 -115
rect 2484 -165 2516 -164
rect 2484 -195 2485 -165
rect 2485 -195 2515 -165
rect 2515 -195 2516 -165
rect 2484 -196 2516 -195
rect 2484 -245 2516 -244
rect 2484 -275 2485 -245
rect 2485 -275 2515 -245
rect 2515 -275 2516 -245
rect 2484 -276 2516 -275
rect 2484 -325 2516 -324
rect 2484 -355 2485 -325
rect 2485 -355 2515 -325
rect 2515 -355 2516 -325
rect 2484 -356 2516 -355
rect 2484 -436 2516 -404
rect 2484 -485 2516 -484
rect 2484 -515 2485 -485
rect 2485 -515 2515 -485
rect 2515 -515 2516 -485
rect 2484 -516 2516 -515
rect 2484 -596 2516 -564
rect 2484 -645 2516 -644
rect 2484 -675 2485 -645
rect 2485 -675 2515 -645
rect 2515 -675 2516 -645
rect 2484 -676 2516 -675
rect 2484 -756 2516 -724
rect 2484 -805 2516 -804
rect 2484 -835 2485 -805
rect 2485 -835 2515 -805
rect 2515 -835 2516 -805
rect 2484 -836 2516 -835
rect 2484 -885 2516 -884
rect 2484 -915 2485 -885
rect 2485 -915 2515 -885
rect 2515 -915 2516 -885
rect 2484 -916 2516 -915
rect 2484 -996 2516 -964
rect 2484 -1076 2516 -1044
rect 2484 -1125 2516 -1124
rect 2484 -1155 2485 -1125
rect 2485 -1155 2515 -1125
rect 2515 -1155 2516 -1125
rect 2484 -1156 2516 -1155
rect 2484 -1205 2516 -1204
rect 2484 -1235 2485 -1205
rect 2485 -1235 2515 -1205
rect 2515 -1235 2516 -1205
rect 2484 -1236 2516 -1235
rect 2484 -1285 2516 -1284
rect 2484 -1315 2485 -1285
rect 2485 -1315 2515 -1285
rect 2515 -1315 2516 -1285
rect 2484 -1316 2516 -1315
rect 2484 -1365 2516 -1364
rect 2484 -1395 2485 -1365
rect 2485 -1395 2515 -1365
rect 2515 -1395 2516 -1365
rect 2484 -1396 2516 -1395
rect 2484 -1445 2516 -1444
rect 2484 -1475 2485 -1445
rect 2485 -1475 2515 -1445
rect 2515 -1475 2516 -1445
rect 2484 -1476 2516 -1475
rect 2484 -1525 2516 -1524
rect 2484 -1555 2485 -1525
rect 2485 -1555 2515 -1525
rect 2515 -1555 2516 -1525
rect 2484 -1556 2516 -1555
rect 2484 -1636 2516 -1604
rect 2484 -1716 2516 -1684
rect 2484 -1765 2516 -1764
rect 2484 -1795 2485 -1765
rect 2485 -1795 2515 -1765
rect 2515 -1795 2516 -1765
rect 2484 -1796 2516 -1795
rect 2484 -1845 2516 -1844
rect 2484 -1875 2485 -1845
rect 2485 -1875 2515 -1845
rect 2515 -1875 2516 -1845
rect 2484 -1876 2516 -1875
rect 2484 -1956 2516 -1924
rect 2484 -2005 2516 -2004
rect 2484 -2035 2485 -2005
rect 2485 -2035 2515 -2005
rect 2515 -2035 2516 -2005
rect 2484 -2036 2516 -2035
rect 2484 -2116 2516 -2084
rect 2484 -2165 2516 -2164
rect 2484 -2195 2485 -2165
rect 2485 -2195 2515 -2165
rect 2515 -2195 2516 -2165
rect 2484 -2196 2516 -2195
rect 2484 -2276 2516 -2244
rect 2484 -2325 2516 -2324
rect 2484 -2355 2485 -2325
rect 2485 -2355 2515 -2325
rect 2515 -2355 2516 -2325
rect 2484 -2356 2516 -2355
rect 2484 -2405 2516 -2404
rect 2484 -2435 2485 -2405
rect 2485 -2435 2515 -2405
rect 2515 -2435 2516 -2405
rect 2484 -2436 2516 -2435
rect 2484 -2485 2516 -2484
rect 2484 -2515 2485 -2485
rect 2485 -2515 2515 -2485
rect 2515 -2515 2516 -2485
rect 2484 -2516 2516 -2515
rect 2484 -2565 2516 -2564
rect 2484 -2595 2485 -2565
rect 2485 -2595 2515 -2565
rect 2515 -2595 2516 -2565
rect 2484 -2596 2516 -2595
rect 2484 -2645 2516 -2644
rect 2484 -2675 2485 -2645
rect 2485 -2675 2515 -2645
rect 2515 -2675 2516 -2645
rect 2484 -2676 2516 -2675
rect 2484 -2725 2516 -2724
rect 2484 -2755 2485 -2725
rect 2485 -2755 2515 -2725
rect 2515 -2755 2516 -2725
rect 2484 -2756 2516 -2755
rect 2484 -2836 2516 -2804
rect 2484 -2885 2516 -2884
rect 2484 -2915 2485 -2885
rect 2485 -2915 2515 -2885
rect 2515 -2915 2516 -2885
rect 2484 -2916 2516 -2915
rect 2484 -2996 2516 -2964
rect 2484 -3045 2516 -3044
rect 2484 -3075 2485 -3045
rect 2485 -3075 2515 -3045
rect 2515 -3075 2516 -3045
rect 2484 -3076 2516 -3075
rect 2484 -3156 2516 -3124
rect 2484 -3205 2516 -3204
rect 2484 -3235 2485 -3205
rect 2485 -3235 2515 -3205
rect 2515 -3235 2516 -3205
rect 2484 -3236 2516 -3235
rect 2484 -3285 2516 -3284
rect 2484 -3315 2485 -3285
rect 2485 -3315 2515 -3285
rect 2515 -3315 2516 -3285
rect 2484 -3316 2516 -3315
rect 2484 -3396 2516 -3364
rect 2484 -3476 2516 -3444
rect 2484 -3525 2516 -3524
rect 2484 -3555 2485 -3525
rect 2485 -3555 2515 -3525
rect 2515 -3555 2516 -3525
rect 2484 -3556 2516 -3555
rect 2484 -3605 2516 -3604
rect 2484 -3635 2485 -3605
rect 2485 -3635 2515 -3605
rect 2515 -3635 2516 -3605
rect 2484 -3636 2516 -3635
rect 2484 -3685 2516 -3684
rect 2484 -3715 2485 -3685
rect 2485 -3715 2515 -3685
rect 2515 -3715 2516 -3685
rect 2484 -3716 2516 -3715
rect 2564 1035 2596 1036
rect 2564 1005 2565 1035
rect 2565 1005 2595 1035
rect 2595 1005 2596 1035
rect 2564 1004 2596 1005
rect 2564 955 2596 956
rect 2564 925 2565 955
rect 2565 925 2595 955
rect 2595 925 2596 955
rect 2564 924 2596 925
rect 2564 875 2596 876
rect 2564 845 2565 875
rect 2565 845 2595 875
rect 2595 845 2596 875
rect 2564 844 2596 845
rect 2564 764 2596 796
rect 2564 684 2596 716
rect 2564 635 2596 636
rect 2564 605 2565 635
rect 2565 605 2595 635
rect 2595 605 2596 635
rect 2564 604 2596 605
rect 2564 555 2596 556
rect 2564 525 2565 555
rect 2565 525 2595 555
rect 2595 525 2596 555
rect 2564 524 2596 525
rect 2564 444 2596 476
rect 2564 395 2596 396
rect 2564 365 2565 395
rect 2565 365 2595 395
rect 2595 365 2596 395
rect 2564 364 2596 365
rect 2564 284 2596 316
rect 2564 235 2596 236
rect 2564 205 2565 235
rect 2565 205 2595 235
rect 2595 205 2596 235
rect 2564 204 2596 205
rect 2564 124 2596 156
rect 2564 75 2596 76
rect 2564 45 2565 75
rect 2565 45 2595 75
rect 2595 45 2596 75
rect 2564 44 2596 45
rect 2564 -5 2596 -4
rect 2564 -35 2565 -5
rect 2565 -35 2595 -5
rect 2595 -35 2596 -5
rect 2564 -36 2596 -35
rect 2564 -85 2596 -84
rect 2564 -115 2565 -85
rect 2565 -115 2595 -85
rect 2595 -115 2596 -85
rect 2564 -116 2596 -115
rect 2564 -165 2596 -164
rect 2564 -195 2565 -165
rect 2565 -195 2595 -165
rect 2595 -195 2596 -165
rect 2564 -196 2596 -195
rect 2564 -245 2596 -244
rect 2564 -275 2565 -245
rect 2565 -275 2595 -245
rect 2595 -275 2596 -245
rect 2564 -276 2596 -275
rect 2564 -325 2596 -324
rect 2564 -355 2565 -325
rect 2565 -355 2595 -325
rect 2595 -355 2596 -325
rect 2564 -356 2596 -355
rect 2564 -436 2596 -404
rect 2564 -485 2596 -484
rect 2564 -515 2565 -485
rect 2565 -515 2595 -485
rect 2595 -515 2596 -485
rect 2564 -516 2596 -515
rect 2564 -596 2596 -564
rect 2564 -645 2596 -644
rect 2564 -675 2565 -645
rect 2565 -675 2595 -645
rect 2595 -675 2596 -645
rect 2564 -676 2596 -675
rect 2564 -756 2596 -724
rect 2564 -805 2596 -804
rect 2564 -835 2565 -805
rect 2565 -835 2595 -805
rect 2595 -835 2596 -805
rect 2564 -836 2596 -835
rect 2564 -885 2596 -884
rect 2564 -915 2565 -885
rect 2565 -915 2595 -885
rect 2595 -915 2596 -885
rect 2564 -916 2596 -915
rect 2564 -996 2596 -964
rect 2564 -1076 2596 -1044
rect 2564 -1125 2596 -1124
rect 2564 -1155 2565 -1125
rect 2565 -1155 2595 -1125
rect 2595 -1155 2596 -1125
rect 2564 -1156 2596 -1155
rect 2564 -1205 2596 -1204
rect 2564 -1235 2565 -1205
rect 2565 -1235 2595 -1205
rect 2595 -1235 2596 -1205
rect 2564 -1236 2596 -1235
rect 2564 -1285 2596 -1284
rect 2564 -1315 2565 -1285
rect 2565 -1315 2595 -1285
rect 2595 -1315 2596 -1285
rect 2564 -1316 2596 -1315
rect 2564 -1365 2596 -1364
rect 2564 -1395 2565 -1365
rect 2565 -1395 2595 -1365
rect 2595 -1395 2596 -1365
rect 2564 -1396 2596 -1395
rect 2564 -1445 2596 -1444
rect 2564 -1475 2565 -1445
rect 2565 -1475 2595 -1445
rect 2595 -1475 2596 -1445
rect 2564 -1476 2596 -1475
rect 2564 -1525 2596 -1524
rect 2564 -1555 2565 -1525
rect 2565 -1555 2595 -1525
rect 2595 -1555 2596 -1525
rect 2564 -1556 2596 -1555
rect 2564 -1636 2596 -1604
rect 2564 -1716 2596 -1684
rect 2564 -1765 2596 -1764
rect 2564 -1795 2565 -1765
rect 2565 -1795 2595 -1765
rect 2595 -1795 2596 -1765
rect 2564 -1796 2596 -1795
rect 2564 -1845 2596 -1844
rect 2564 -1875 2565 -1845
rect 2565 -1875 2595 -1845
rect 2595 -1875 2596 -1845
rect 2564 -1876 2596 -1875
rect 2564 -1956 2596 -1924
rect 2564 -2005 2596 -2004
rect 2564 -2035 2565 -2005
rect 2565 -2035 2595 -2005
rect 2595 -2035 2596 -2005
rect 2564 -2036 2596 -2035
rect 2564 -2116 2596 -2084
rect 2564 -2165 2596 -2164
rect 2564 -2195 2565 -2165
rect 2565 -2195 2595 -2165
rect 2595 -2195 2596 -2165
rect 2564 -2196 2596 -2195
rect 2564 -2276 2596 -2244
rect 2564 -2325 2596 -2324
rect 2564 -2355 2565 -2325
rect 2565 -2355 2595 -2325
rect 2595 -2355 2596 -2325
rect 2564 -2356 2596 -2355
rect 2564 -2405 2596 -2404
rect 2564 -2435 2565 -2405
rect 2565 -2435 2595 -2405
rect 2595 -2435 2596 -2405
rect 2564 -2436 2596 -2435
rect 2564 -2485 2596 -2484
rect 2564 -2515 2565 -2485
rect 2565 -2515 2595 -2485
rect 2595 -2515 2596 -2485
rect 2564 -2516 2596 -2515
rect 2564 -2565 2596 -2564
rect 2564 -2595 2565 -2565
rect 2565 -2595 2595 -2565
rect 2595 -2595 2596 -2565
rect 2564 -2596 2596 -2595
rect 2564 -2645 2596 -2644
rect 2564 -2675 2565 -2645
rect 2565 -2675 2595 -2645
rect 2595 -2675 2596 -2645
rect 2564 -2676 2596 -2675
rect 2564 -2725 2596 -2724
rect 2564 -2755 2565 -2725
rect 2565 -2755 2595 -2725
rect 2595 -2755 2596 -2725
rect 2564 -2756 2596 -2755
rect 2564 -2836 2596 -2804
rect 2564 -2885 2596 -2884
rect 2564 -2915 2565 -2885
rect 2565 -2915 2595 -2885
rect 2595 -2915 2596 -2885
rect 2564 -2916 2596 -2915
rect 2564 -2996 2596 -2964
rect 2564 -3045 2596 -3044
rect 2564 -3075 2565 -3045
rect 2565 -3075 2595 -3045
rect 2595 -3075 2596 -3045
rect 2564 -3076 2596 -3075
rect 2564 -3156 2596 -3124
rect 2564 -3205 2596 -3204
rect 2564 -3235 2565 -3205
rect 2565 -3235 2595 -3205
rect 2595 -3235 2596 -3205
rect 2564 -3236 2596 -3235
rect 2564 -3285 2596 -3284
rect 2564 -3315 2565 -3285
rect 2565 -3315 2595 -3285
rect 2595 -3315 2596 -3285
rect 2564 -3316 2596 -3315
rect 2564 -3396 2596 -3364
rect 2564 -3476 2596 -3444
rect 2564 -3525 2596 -3524
rect 2564 -3555 2565 -3525
rect 2565 -3555 2595 -3525
rect 2595 -3555 2596 -3525
rect 2564 -3556 2596 -3555
rect 2564 -3605 2596 -3604
rect 2564 -3635 2565 -3605
rect 2565 -3635 2595 -3605
rect 2595 -3635 2596 -3605
rect 2564 -3636 2596 -3635
rect 2564 -3685 2596 -3684
rect 2564 -3715 2565 -3685
rect 2565 -3715 2595 -3685
rect 2595 -3715 2596 -3685
rect 2564 -3716 2596 -3715
rect 2644 1035 2676 1036
rect 2644 1005 2645 1035
rect 2645 1005 2675 1035
rect 2675 1005 2676 1035
rect 2644 1004 2676 1005
rect 2644 955 2676 956
rect 2644 925 2645 955
rect 2645 925 2675 955
rect 2675 925 2676 955
rect 2644 924 2676 925
rect 2644 875 2676 876
rect 2644 845 2645 875
rect 2645 845 2675 875
rect 2675 845 2676 875
rect 2644 844 2676 845
rect 2644 764 2676 796
rect 2644 684 2676 716
rect 2644 635 2676 636
rect 2644 605 2645 635
rect 2645 605 2675 635
rect 2675 605 2676 635
rect 2644 604 2676 605
rect 2644 555 2676 556
rect 2644 525 2645 555
rect 2645 525 2675 555
rect 2675 525 2676 555
rect 2644 524 2676 525
rect 2644 444 2676 476
rect 2644 395 2676 396
rect 2644 365 2645 395
rect 2645 365 2675 395
rect 2675 365 2676 395
rect 2644 364 2676 365
rect 2644 284 2676 316
rect 2644 235 2676 236
rect 2644 205 2645 235
rect 2645 205 2675 235
rect 2675 205 2676 235
rect 2644 204 2676 205
rect 2644 124 2676 156
rect 2644 75 2676 76
rect 2644 45 2645 75
rect 2645 45 2675 75
rect 2675 45 2676 75
rect 2644 44 2676 45
rect 2644 -5 2676 -4
rect 2644 -35 2645 -5
rect 2645 -35 2675 -5
rect 2675 -35 2676 -5
rect 2644 -36 2676 -35
rect 2644 -85 2676 -84
rect 2644 -115 2645 -85
rect 2645 -115 2675 -85
rect 2675 -115 2676 -85
rect 2644 -116 2676 -115
rect 2644 -165 2676 -164
rect 2644 -195 2645 -165
rect 2645 -195 2675 -165
rect 2675 -195 2676 -165
rect 2644 -196 2676 -195
rect 2644 -245 2676 -244
rect 2644 -275 2645 -245
rect 2645 -275 2675 -245
rect 2675 -275 2676 -245
rect 2644 -276 2676 -275
rect 2644 -325 2676 -324
rect 2644 -355 2645 -325
rect 2645 -355 2675 -325
rect 2675 -355 2676 -325
rect 2644 -356 2676 -355
rect 2644 -436 2676 -404
rect 2644 -485 2676 -484
rect 2644 -515 2645 -485
rect 2645 -515 2675 -485
rect 2675 -515 2676 -485
rect 2644 -516 2676 -515
rect 2644 -596 2676 -564
rect 2644 -645 2676 -644
rect 2644 -675 2645 -645
rect 2645 -675 2675 -645
rect 2675 -675 2676 -645
rect 2644 -676 2676 -675
rect 2644 -756 2676 -724
rect 2644 -805 2676 -804
rect 2644 -835 2645 -805
rect 2645 -835 2675 -805
rect 2675 -835 2676 -805
rect 2644 -836 2676 -835
rect 2644 -885 2676 -884
rect 2644 -915 2645 -885
rect 2645 -915 2675 -885
rect 2675 -915 2676 -885
rect 2644 -916 2676 -915
rect 2644 -996 2676 -964
rect 2644 -1076 2676 -1044
rect 2644 -1125 2676 -1124
rect 2644 -1155 2645 -1125
rect 2645 -1155 2675 -1125
rect 2675 -1155 2676 -1125
rect 2644 -1156 2676 -1155
rect 2644 -1205 2676 -1204
rect 2644 -1235 2645 -1205
rect 2645 -1235 2675 -1205
rect 2675 -1235 2676 -1205
rect 2644 -1236 2676 -1235
rect 2644 -1285 2676 -1284
rect 2644 -1315 2645 -1285
rect 2645 -1315 2675 -1285
rect 2675 -1315 2676 -1285
rect 2644 -1316 2676 -1315
rect 2644 -1365 2676 -1364
rect 2644 -1395 2645 -1365
rect 2645 -1395 2675 -1365
rect 2675 -1395 2676 -1365
rect 2644 -1396 2676 -1395
rect 2644 -1445 2676 -1444
rect 2644 -1475 2645 -1445
rect 2645 -1475 2675 -1445
rect 2675 -1475 2676 -1445
rect 2644 -1476 2676 -1475
rect 2644 -1525 2676 -1524
rect 2644 -1555 2645 -1525
rect 2645 -1555 2675 -1525
rect 2675 -1555 2676 -1525
rect 2644 -1556 2676 -1555
rect 2644 -1636 2676 -1604
rect 2644 -1716 2676 -1684
rect 2644 -1765 2676 -1764
rect 2644 -1795 2645 -1765
rect 2645 -1795 2675 -1765
rect 2675 -1795 2676 -1765
rect 2644 -1796 2676 -1795
rect 2644 -1845 2676 -1844
rect 2644 -1875 2645 -1845
rect 2645 -1875 2675 -1845
rect 2675 -1875 2676 -1845
rect 2644 -1876 2676 -1875
rect 2644 -1956 2676 -1924
rect 2644 -2005 2676 -2004
rect 2644 -2035 2645 -2005
rect 2645 -2035 2675 -2005
rect 2675 -2035 2676 -2005
rect 2644 -2036 2676 -2035
rect 2644 -2116 2676 -2084
rect 2644 -2165 2676 -2164
rect 2644 -2195 2645 -2165
rect 2645 -2195 2675 -2165
rect 2675 -2195 2676 -2165
rect 2644 -2196 2676 -2195
rect 2644 -2276 2676 -2244
rect 2644 -2325 2676 -2324
rect 2644 -2355 2645 -2325
rect 2645 -2355 2675 -2325
rect 2675 -2355 2676 -2325
rect 2644 -2356 2676 -2355
rect 2644 -2405 2676 -2404
rect 2644 -2435 2645 -2405
rect 2645 -2435 2675 -2405
rect 2675 -2435 2676 -2405
rect 2644 -2436 2676 -2435
rect 2644 -2485 2676 -2484
rect 2644 -2515 2645 -2485
rect 2645 -2515 2675 -2485
rect 2675 -2515 2676 -2485
rect 2644 -2516 2676 -2515
rect 2644 -2565 2676 -2564
rect 2644 -2595 2645 -2565
rect 2645 -2595 2675 -2565
rect 2675 -2595 2676 -2565
rect 2644 -2596 2676 -2595
rect 2644 -2645 2676 -2644
rect 2644 -2675 2645 -2645
rect 2645 -2675 2675 -2645
rect 2675 -2675 2676 -2645
rect 2644 -2676 2676 -2675
rect 2644 -2725 2676 -2724
rect 2644 -2755 2645 -2725
rect 2645 -2755 2675 -2725
rect 2675 -2755 2676 -2725
rect 2644 -2756 2676 -2755
rect 2644 -2836 2676 -2804
rect 2644 -2885 2676 -2884
rect 2644 -2915 2645 -2885
rect 2645 -2915 2675 -2885
rect 2675 -2915 2676 -2885
rect 2644 -2916 2676 -2915
rect 2644 -2996 2676 -2964
rect 2644 -3045 2676 -3044
rect 2644 -3075 2645 -3045
rect 2645 -3075 2675 -3045
rect 2675 -3075 2676 -3045
rect 2644 -3076 2676 -3075
rect 2644 -3156 2676 -3124
rect 2644 -3205 2676 -3204
rect 2644 -3235 2645 -3205
rect 2645 -3235 2675 -3205
rect 2675 -3235 2676 -3205
rect 2644 -3236 2676 -3235
rect 2644 -3285 2676 -3284
rect 2644 -3315 2645 -3285
rect 2645 -3315 2675 -3285
rect 2675 -3315 2676 -3285
rect 2644 -3316 2676 -3315
rect 2644 -3396 2676 -3364
rect 2644 -3476 2676 -3444
rect 2644 -3525 2676 -3524
rect 2644 -3555 2645 -3525
rect 2645 -3555 2675 -3525
rect 2675 -3555 2676 -3525
rect 2644 -3556 2676 -3555
rect 2644 -3605 2676 -3604
rect 2644 -3635 2645 -3605
rect 2645 -3635 2675 -3605
rect 2675 -3635 2676 -3605
rect 2644 -3636 2676 -3635
rect 2644 -3685 2676 -3684
rect 2644 -3715 2645 -3685
rect 2645 -3715 2675 -3685
rect 2675 -3715 2676 -3685
rect 2644 -3716 2676 -3715
rect 2724 1035 2756 1036
rect 2724 1005 2725 1035
rect 2725 1005 2755 1035
rect 2755 1005 2756 1035
rect 2724 1004 2756 1005
rect 2724 955 2756 956
rect 2724 925 2725 955
rect 2725 925 2755 955
rect 2755 925 2756 955
rect 2724 924 2756 925
rect 2724 875 2756 876
rect 2724 845 2725 875
rect 2725 845 2755 875
rect 2755 845 2756 875
rect 2724 844 2756 845
rect 2724 764 2756 796
rect 2724 684 2756 716
rect 2724 635 2756 636
rect 2724 605 2725 635
rect 2725 605 2755 635
rect 2755 605 2756 635
rect 2724 604 2756 605
rect 2724 555 2756 556
rect 2724 525 2725 555
rect 2725 525 2755 555
rect 2755 525 2756 555
rect 2724 524 2756 525
rect 2724 444 2756 476
rect 2724 395 2756 396
rect 2724 365 2725 395
rect 2725 365 2755 395
rect 2755 365 2756 395
rect 2724 364 2756 365
rect 2724 284 2756 316
rect 2724 235 2756 236
rect 2724 205 2725 235
rect 2725 205 2755 235
rect 2755 205 2756 235
rect 2724 204 2756 205
rect 2724 124 2756 156
rect 2724 75 2756 76
rect 2724 45 2725 75
rect 2725 45 2755 75
rect 2755 45 2756 75
rect 2724 44 2756 45
rect 2724 -5 2756 -4
rect 2724 -35 2725 -5
rect 2725 -35 2755 -5
rect 2755 -35 2756 -5
rect 2724 -36 2756 -35
rect 2724 -85 2756 -84
rect 2724 -115 2725 -85
rect 2725 -115 2755 -85
rect 2755 -115 2756 -85
rect 2724 -116 2756 -115
rect 2724 -165 2756 -164
rect 2724 -195 2725 -165
rect 2725 -195 2755 -165
rect 2755 -195 2756 -165
rect 2724 -196 2756 -195
rect 2724 -245 2756 -244
rect 2724 -275 2725 -245
rect 2725 -275 2755 -245
rect 2755 -275 2756 -245
rect 2724 -276 2756 -275
rect 2724 -325 2756 -324
rect 2724 -355 2725 -325
rect 2725 -355 2755 -325
rect 2755 -355 2756 -325
rect 2724 -356 2756 -355
rect 2724 -436 2756 -404
rect 2724 -485 2756 -484
rect 2724 -515 2725 -485
rect 2725 -515 2755 -485
rect 2755 -515 2756 -485
rect 2724 -516 2756 -515
rect 2724 -596 2756 -564
rect 2724 -645 2756 -644
rect 2724 -675 2725 -645
rect 2725 -675 2755 -645
rect 2755 -675 2756 -645
rect 2724 -676 2756 -675
rect 2724 -756 2756 -724
rect 2724 -805 2756 -804
rect 2724 -835 2725 -805
rect 2725 -835 2755 -805
rect 2755 -835 2756 -805
rect 2724 -836 2756 -835
rect 2724 -885 2756 -884
rect 2724 -915 2725 -885
rect 2725 -915 2755 -885
rect 2755 -915 2756 -885
rect 2724 -916 2756 -915
rect 2724 -996 2756 -964
rect 2724 -1076 2756 -1044
rect 2724 -1125 2756 -1124
rect 2724 -1155 2725 -1125
rect 2725 -1155 2755 -1125
rect 2755 -1155 2756 -1125
rect 2724 -1156 2756 -1155
rect 2724 -1205 2756 -1204
rect 2724 -1235 2725 -1205
rect 2725 -1235 2755 -1205
rect 2755 -1235 2756 -1205
rect 2724 -1236 2756 -1235
rect 2724 -1285 2756 -1284
rect 2724 -1315 2725 -1285
rect 2725 -1315 2755 -1285
rect 2755 -1315 2756 -1285
rect 2724 -1316 2756 -1315
rect 2724 -1365 2756 -1364
rect 2724 -1395 2725 -1365
rect 2725 -1395 2755 -1365
rect 2755 -1395 2756 -1365
rect 2724 -1396 2756 -1395
rect 2724 -1445 2756 -1444
rect 2724 -1475 2725 -1445
rect 2725 -1475 2755 -1445
rect 2755 -1475 2756 -1445
rect 2724 -1476 2756 -1475
rect 2724 -1525 2756 -1524
rect 2724 -1555 2725 -1525
rect 2725 -1555 2755 -1525
rect 2755 -1555 2756 -1525
rect 2724 -1556 2756 -1555
rect 2724 -1636 2756 -1604
rect 2724 -1716 2756 -1684
rect 2724 -1765 2756 -1764
rect 2724 -1795 2725 -1765
rect 2725 -1795 2755 -1765
rect 2755 -1795 2756 -1765
rect 2724 -1796 2756 -1795
rect 2724 -1845 2756 -1844
rect 2724 -1875 2725 -1845
rect 2725 -1875 2755 -1845
rect 2755 -1875 2756 -1845
rect 2724 -1876 2756 -1875
rect 2724 -1956 2756 -1924
rect 2724 -2005 2756 -2004
rect 2724 -2035 2725 -2005
rect 2725 -2035 2755 -2005
rect 2755 -2035 2756 -2005
rect 2724 -2036 2756 -2035
rect 2724 -2116 2756 -2084
rect 2724 -2165 2756 -2164
rect 2724 -2195 2725 -2165
rect 2725 -2195 2755 -2165
rect 2755 -2195 2756 -2165
rect 2724 -2196 2756 -2195
rect 2724 -2276 2756 -2244
rect 2724 -2325 2756 -2324
rect 2724 -2355 2725 -2325
rect 2725 -2355 2755 -2325
rect 2755 -2355 2756 -2325
rect 2724 -2356 2756 -2355
rect 2724 -2405 2756 -2404
rect 2724 -2435 2725 -2405
rect 2725 -2435 2755 -2405
rect 2755 -2435 2756 -2405
rect 2724 -2436 2756 -2435
rect 2724 -2485 2756 -2484
rect 2724 -2515 2725 -2485
rect 2725 -2515 2755 -2485
rect 2755 -2515 2756 -2485
rect 2724 -2516 2756 -2515
rect 2724 -2565 2756 -2564
rect 2724 -2595 2725 -2565
rect 2725 -2595 2755 -2565
rect 2755 -2595 2756 -2565
rect 2724 -2596 2756 -2595
rect 2724 -2645 2756 -2644
rect 2724 -2675 2725 -2645
rect 2725 -2675 2755 -2645
rect 2755 -2675 2756 -2645
rect 2724 -2676 2756 -2675
rect 2724 -2725 2756 -2724
rect 2724 -2755 2725 -2725
rect 2725 -2755 2755 -2725
rect 2755 -2755 2756 -2725
rect 2724 -2756 2756 -2755
rect 2724 -2836 2756 -2804
rect 2724 -2885 2756 -2884
rect 2724 -2915 2725 -2885
rect 2725 -2915 2755 -2885
rect 2755 -2915 2756 -2885
rect 2724 -2916 2756 -2915
rect 2724 -2996 2756 -2964
rect 2724 -3045 2756 -3044
rect 2724 -3075 2725 -3045
rect 2725 -3075 2755 -3045
rect 2755 -3075 2756 -3045
rect 2724 -3076 2756 -3075
rect 2724 -3156 2756 -3124
rect 2724 -3205 2756 -3204
rect 2724 -3235 2725 -3205
rect 2725 -3235 2755 -3205
rect 2755 -3235 2756 -3205
rect 2724 -3236 2756 -3235
rect 2724 -3285 2756 -3284
rect 2724 -3315 2725 -3285
rect 2725 -3315 2755 -3285
rect 2755 -3315 2756 -3285
rect 2724 -3316 2756 -3315
rect 2724 -3396 2756 -3364
rect 2724 -3476 2756 -3444
rect 2724 -3525 2756 -3524
rect 2724 -3555 2725 -3525
rect 2725 -3555 2755 -3525
rect 2755 -3555 2756 -3525
rect 2724 -3556 2756 -3555
rect 2724 -3605 2756 -3604
rect 2724 -3635 2725 -3605
rect 2725 -3635 2755 -3605
rect 2755 -3635 2756 -3605
rect 2724 -3636 2756 -3635
rect 2724 -3685 2756 -3684
rect 2724 -3715 2725 -3685
rect 2725 -3715 2755 -3685
rect 2755 -3715 2756 -3685
rect 2724 -3716 2756 -3715
rect 2804 1035 2836 1036
rect 2804 1005 2805 1035
rect 2805 1005 2835 1035
rect 2835 1005 2836 1035
rect 2804 1004 2836 1005
rect 2804 955 2836 956
rect 2804 925 2805 955
rect 2805 925 2835 955
rect 2835 925 2836 955
rect 2804 924 2836 925
rect 2804 875 2836 876
rect 2804 845 2805 875
rect 2805 845 2835 875
rect 2835 845 2836 875
rect 2804 844 2836 845
rect 2804 764 2836 796
rect 2804 684 2836 716
rect 2804 635 2836 636
rect 2804 605 2805 635
rect 2805 605 2835 635
rect 2835 605 2836 635
rect 2804 604 2836 605
rect 2804 555 2836 556
rect 2804 525 2805 555
rect 2805 525 2835 555
rect 2835 525 2836 555
rect 2804 524 2836 525
rect 2804 444 2836 476
rect 2804 395 2836 396
rect 2804 365 2805 395
rect 2805 365 2835 395
rect 2835 365 2836 395
rect 2804 364 2836 365
rect 2804 284 2836 316
rect 2804 235 2836 236
rect 2804 205 2805 235
rect 2805 205 2835 235
rect 2835 205 2836 235
rect 2804 204 2836 205
rect 2804 124 2836 156
rect 2804 75 2836 76
rect 2804 45 2805 75
rect 2805 45 2835 75
rect 2835 45 2836 75
rect 2804 44 2836 45
rect 2804 -5 2836 -4
rect 2804 -35 2805 -5
rect 2805 -35 2835 -5
rect 2835 -35 2836 -5
rect 2804 -36 2836 -35
rect 2804 -85 2836 -84
rect 2804 -115 2805 -85
rect 2805 -115 2835 -85
rect 2835 -115 2836 -85
rect 2804 -116 2836 -115
rect 2804 -165 2836 -164
rect 2804 -195 2805 -165
rect 2805 -195 2835 -165
rect 2835 -195 2836 -165
rect 2804 -196 2836 -195
rect 2804 -245 2836 -244
rect 2804 -275 2805 -245
rect 2805 -275 2835 -245
rect 2835 -275 2836 -245
rect 2804 -276 2836 -275
rect 2804 -325 2836 -324
rect 2804 -355 2805 -325
rect 2805 -355 2835 -325
rect 2835 -355 2836 -325
rect 2804 -356 2836 -355
rect 2804 -436 2836 -404
rect 2804 -485 2836 -484
rect 2804 -515 2805 -485
rect 2805 -515 2835 -485
rect 2835 -515 2836 -485
rect 2804 -516 2836 -515
rect 2804 -596 2836 -564
rect 2804 -645 2836 -644
rect 2804 -675 2805 -645
rect 2805 -675 2835 -645
rect 2835 -675 2836 -645
rect 2804 -676 2836 -675
rect 2804 -756 2836 -724
rect 2804 -805 2836 -804
rect 2804 -835 2805 -805
rect 2805 -835 2835 -805
rect 2835 -835 2836 -805
rect 2804 -836 2836 -835
rect 2804 -885 2836 -884
rect 2804 -915 2805 -885
rect 2805 -915 2835 -885
rect 2835 -915 2836 -885
rect 2804 -916 2836 -915
rect 2804 -996 2836 -964
rect 2804 -1076 2836 -1044
rect 2804 -1125 2836 -1124
rect 2804 -1155 2805 -1125
rect 2805 -1155 2835 -1125
rect 2835 -1155 2836 -1125
rect 2804 -1156 2836 -1155
rect 2804 -1205 2836 -1204
rect 2804 -1235 2805 -1205
rect 2805 -1235 2835 -1205
rect 2835 -1235 2836 -1205
rect 2804 -1236 2836 -1235
rect 2804 -1285 2836 -1284
rect 2804 -1315 2805 -1285
rect 2805 -1315 2835 -1285
rect 2835 -1315 2836 -1285
rect 2804 -1316 2836 -1315
rect 2804 -1365 2836 -1364
rect 2804 -1395 2805 -1365
rect 2805 -1395 2835 -1365
rect 2835 -1395 2836 -1365
rect 2804 -1396 2836 -1395
rect 2804 -1445 2836 -1444
rect 2804 -1475 2805 -1445
rect 2805 -1475 2835 -1445
rect 2835 -1475 2836 -1445
rect 2804 -1476 2836 -1475
rect 2804 -1525 2836 -1524
rect 2804 -1555 2805 -1525
rect 2805 -1555 2835 -1525
rect 2835 -1555 2836 -1525
rect 2804 -1556 2836 -1555
rect 2804 -1636 2836 -1604
rect 2804 -1716 2836 -1684
rect 2804 -1765 2836 -1764
rect 2804 -1795 2805 -1765
rect 2805 -1795 2835 -1765
rect 2835 -1795 2836 -1765
rect 2804 -1796 2836 -1795
rect 2804 -1845 2836 -1844
rect 2804 -1875 2805 -1845
rect 2805 -1875 2835 -1845
rect 2835 -1875 2836 -1845
rect 2804 -1876 2836 -1875
rect 2804 -1956 2836 -1924
rect 2804 -2005 2836 -2004
rect 2804 -2035 2805 -2005
rect 2805 -2035 2835 -2005
rect 2835 -2035 2836 -2005
rect 2804 -2036 2836 -2035
rect 2804 -2116 2836 -2084
rect 2804 -2165 2836 -2164
rect 2804 -2195 2805 -2165
rect 2805 -2195 2835 -2165
rect 2835 -2195 2836 -2165
rect 2804 -2196 2836 -2195
rect 2804 -2276 2836 -2244
rect 2804 -2325 2836 -2324
rect 2804 -2355 2805 -2325
rect 2805 -2355 2835 -2325
rect 2835 -2355 2836 -2325
rect 2804 -2356 2836 -2355
rect 2804 -2405 2836 -2404
rect 2804 -2435 2805 -2405
rect 2805 -2435 2835 -2405
rect 2835 -2435 2836 -2405
rect 2804 -2436 2836 -2435
rect 2804 -2485 2836 -2484
rect 2804 -2515 2805 -2485
rect 2805 -2515 2835 -2485
rect 2835 -2515 2836 -2485
rect 2804 -2516 2836 -2515
rect 2804 -2565 2836 -2564
rect 2804 -2595 2805 -2565
rect 2805 -2595 2835 -2565
rect 2835 -2595 2836 -2565
rect 2804 -2596 2836 -2595
rect 2804 -2645 2836 -2644
rect 2804 -2675 2805 -2645
rect 2805 -2675 2835 -2645
rect 2835 -2675 2836 -2645
rect 2804 -2676 2836 -2675
rect 2804 -2725 2836 -2724
rect 2804 -2755 2805 -2725
rect 2805 -2755 2835 -2725
rect 2835 -2755 2836 -2725
rect 2804 -2756 2836 -2755
rect 2804 -2836 2836 -2804
rect 2804 -2885 2836 -2884
rect 2804 -2915 2805 -2885
rect 2805 -2915 2835 -2885
rect 2835 -2915 2836 -2885
rect 2804 -2916 2836 -2915
rect 2804 -2996 2836 -2964
rect 2804 -3045 2836 -3044
rect 2804 -3075 2805 -3045
rect 2805 -3075 2835 -3045
rect 2835 -3075 2836 -3045
rect 2804 -3076 2836 -3075
rect 2804 -3156 2836 -3124
rect 2804 -3205 2836 -3204
rect 2804 -3235 2805 -3205
rect 2805 -3235 2835 -3205
rect 2835 -3235 2836 -3205
rect 2804 -3236 2836 -3235
rect 2804 -3285 2836 -3284
rect 2804 -3315 2805 -3285
rect 2805 -3315 2835 -3285
rect 2835 -3315 2836 -3285
rect 2804 -3316 2836 -3315
rect 2804 -3396 2836 -3364
rect 2804 -3476 2836 -3444
rect 2804 -3525 2836 -3524
rect 2804 -3555 2805 -3525
rect 2805 -3555 2835 -3525
rect 2835 -3555 2836 -3525
rect 2804 -3556 2836 -3555
rect 2804 -3605 2836 -3604
rect 2804 -3635 2805 -3605
rect 2805 -3635 2835 -3605
rect 2835 -3635 2836 -3605
rect 2804 -3636 2836 -3635
rect 2804 -3685 2836 -3684
rect 2804 -3715 2805 -3685
rect 2805 -3715 2835 -3685
rect 2835 -3715 2836 -3685
rect 2804 -3716 2836 -3715
rect 2884 1035 2916 1036
rect 2884 1005 2885 1035
rect 2885 1005 2915 1035
rect 2915 1005 2916 1035
rect 2884 1004 2916 1005
rect 2884 955 2916 956
rect 2884 925 2885 955
rect 2885 925 2915 955
rect 2915 925 2916 955
rect 2884 924 2916 925
rect 2884 875 2916 876
rect 2884 845 2885 875
rect 2885 845 2915 875
rect 2915 845 2916 875
rect 2884 844 2916 845
rect 2884 764 2916 796
rect 2884 684 2916 716
rect 2884 635 2916 636
rect 2884 605 2885 635
rect 2885 605 2915 635
rect 2915 605 2916 635
rect 2884 604 2916 605
rect 2884 555 2916 556
rect 2884 525 2885 555
rect 2885 525 2915 555
rect 2915 525 2916 555
rect 2884 524 2916 525
rect 2884 444 2916 476
rect 2884 395 2916 396
rect 2884 365 2885 395
rect 2885 365 2915 395
rect 2915 365 2916 395
rect 2884 364 2916 365
rect 2884 284 2916 316
rect 2884 235 2916 236
rect 2884 205 2885 235
rect 2885 205 2915 235
rect 2915 205 2916 235
rect 2884 204 2916 205
rect 2884 124 2916 156
rect 2884 75 2916 76
rect 2884 45 2885 75
rect 2885 45 2915 75
rect 2915 45 2916 75
rect 2884 44 2916 45
rect 2884 -5 2916 -4
rect 2884 -35 2885 -5
rect 2885 -35 2915 -5
rect 2915 -35 2916 -5
rect 2884 -36 2916 -35
rect 2884 -85 2916 -84
rect 2884 -115 2885 -85
rect 2885 -115 2915 -85
rect 2915 -115 2916 -85
rect 2884 -116 2916 -115
rect 2884 -165 2916 -164
rect 2884 -195 2885 -165
rect 2885 -195 2915 -165
rect 2915 -195 2916 -165
rect 2884 -196 2916 -195
rect 2884 -245 2916 -244
rect 2884 -275 2885 -245
rect 2885 -275 2915 -245
rect 2915 -275 2916 -245
rect 2884 -276 2916 -275
rect 2884 -325 2916 -324
rect 2884 -355 2885 -325
rect 2885 -355 2915 -325
rect 2915 -355 2916 -325
rect 2884 -356 2916 -355
rect 2884 -436 2916 -404
rect 2884 -485 2916 -484
rect 2884 -515 2885 -485
rect 2885 -515 2915 -485
rect 2915 -515 2916 -485
rect 2884 -516 2916 -515
rect 2884 -596 2916 -564
rect 2884 -645 2916 -644
rect 2884 -675 2885 -645
rect 2885 -675 2915 -645
rect 2915 -675 2916 -645
rect 2884 -676 2916 -675
rect 2884 -756 2916 -724
rect 2884 -805 2916 -804
rect 2884 -835 2885 -805
rect 2885 -835 2915 -805
rect 2915 -835 2916 -805
rect 2884 -836 2916 -835
rect 2884 -885 2916 -884
rect 2884 -915 2885 -885
rect 2885 -915 2915 -885
rect 2915 -915 2916 -885
rect 2884 -916 2916 -915
rect 2884 -996 2916 -964
rect 2884 -1076 2916 -1044
rect 2884 -1125 2916 -1124
rect 2884 -1155 2885 -1125
rect 2885 -1155 2915 -1125
rect 2915 -1155 2916 -1125
rect 2884 -1156 2916 -1155
rect 2884 -1205 2916 -1204
rect 2884 -1235 2885 -1205
rect 2885 -1235 2915 -1205
rect 2915 -1235 2916 -1205
rect 2884 -1236 2916 -1235
rect 2884 -1285 2916 -1284
rect 2884 -1315 2885 -1285
rect 2885 -1315 2915 -1285
rect 2915 -1315 2916 -1285
rect 2884 -1316 2916 -1315
rect 2884 -1365 2916 -1364
rect 2884 -1395 2885 -1365
rect 2885 -1395 2915 -1365
rect 2915 -1395 2916 -1365
rect 2884 -1396 2916 -1395
rect 2884 -1445 2916 -1444
rect 2884 -1475 2885 -1445
rect 2885 -1475 2915 -1445
rect 2915 -1475 2916 -1445
rect 2884 -1476 2916 -1475
rect 2884 -1525 2916 -1524
rect 2884 -1555 2885 -1525
rect 2885 -1555 2915 -1525
rect 2915 -1555 2916 -1525
rect 2884 -1556 2916 -1555
rect 2884 -1636 2916 -1604
rect 2884 -1716 2916 -1684
rect 2884 -1765 2916 -1764
rect 2884 -1795 2885 -1765
rect 2885 -1795 2915 -1765
rect 2915 -1795 2916 -1765
rect 2884 -1796 2916 -1795
rect 2884 -1845 2916 -1844
rect 2884 -1875 2885 -1845
rect 2885 -1875 2915 -1845
rect 2915 -1875 2916 -1845
rect 2884 -1876 2916 -1875
rect 2884 -1956 2916 -1924
rect 2884 -2005 2916 -2004
rect 2884 -2035 2885 -2005
rect 2885 -2035 2915 -2005
rect 2915 -2035 2916 -2005
rect 2884 -2036 2916 -2035
rect 2884 -2116 2916 -2084
rect 2884 -2165 2916 -2164
rect 2884 -2195 2885 -2165
rect 2885 -2195 2915 -2165
rect 2915 -2195 2916 -2165
rect 2884 -2196 2916 -2195
rect 2884 -2276 2916 -2244
rect 2884 -2325 2916 -2324
rect 2884 -2355 2885 -2325
rect 2885 -2355 2915 -2325
rect 2915 -2355 2916 -2325
rect 2884 -2356 2916 -2355
rect 2884 -2405 2916 -2404
rect 2884 -2435 2885 -2405
rect 2885 -2435 2915 -2405
rect 2915 -2435 2916 -2405
rect 2884 -2436 2916 -2435
rect 2884 -2485 2916 -2484
rect 2884 -2515 2885 -2485
rect 2885 -2515 2915 -2485
rect 2915 -2515 2916 -2485
rect 2884 -2516 2916 -2515
rect 2884 -2565 2916 -2564
rect 2884 -2595 2885 -2565
rect 2885 -2595 2915 -2565
rect 2915 -2595 2916 -2565
rect 2884 -2596 2916 -2595
rect 2884 -2645 2916 -2644
rect 2884 -2675 2885 -2645
rect 2885 -2675 2915 -2645
rect 2915 -2675 2916 -2645
rect 2884 -2676 2916 -2675
rect 2884 -2725 2916 -2724
rect 2884 -2755 2885 -2725
rect 2885 -2755 2915 -2725
rect 2915 -2755 2916 -2725
rect 2884 -2756 2916 -2755
rect 2884 -2836 2916 -2804
rect 2884 -2885 2916 -2884
rect 2884 -2915 2885 -2885
rect 2885 -2915 2915 -2885
rect 2915 -2915 2916 -2885
rect 2884 -2916 2916 -2915
rect 2884 -2996 2916 -2964
rect 2884 -3045 2916 -3044
rect 2884 -3075 2885 -3045
rect 2885 -3075 2915 -3045
rect 2915 -3075 2916 -3045
rect 2884 -3076 2916 -3075
rect 2884 -3156 2916 -3124
rect 2884 -3205 2916 -3204
rect 2884 -3235 2885 -3205
rect 2885 -3235 2915 -3205
rect 2915 -3235 2916 -3205
rect 2884 -3236 2916 -3235
rect 2884 -3285 2916 -3284
rect 2884 -3315 2885 -3285
rect 2885 -3315 2915 -3285
rect 2915 -3315 2916 -3285
rect 2884 -3316 2916 -3315
rect 2884 -3396 2916 -3364
rect 2884 -3476 2916 -3444
rect 2884 -3525 2916 -3524
rect 2884 -3555 2885 -3525
rect 2885 -3555 2915 -3525
rect 2915 -3555 2916 -3525
rect 2884 -3556 2916 -3555
rect 2884 -3605 2916 -3604
rect 2884 -3635 2885 -3605
rect 2885 -3635 2915 -3605
rect 2915 -3635 2916 -3605
rect 2884 -3636 2916 -3635
rect 2884 -3685 2916 -3684
rect 2884 -3715 2885 -3685
rect 2885 -3715 2915 -3685
rect 2915 -3715 2916 -3685
rect 2884 -3716 2916 -3715
rect 2964 1035 2996 1036
rect 2964 1005 2965 1035
rect 2965 1005 2995 1035
rect 2995 1005 2996 1035
rect 2964 1004 2996 1005
rect 2964 955 2996 956
rect 2964 925 2965 955
rect 2965 925 2995 955
rect 2995 925 2996 955
rect 2964 924 2996 925
rect 2964 875 2996 876
rect 2964 845 2965 875
rect 2965 845 2995 875
rect 2995 845 2996 875
rect 2964 844 2996 845
rect 2964 764 2996 796
rect 2964 684 2996 716
rect 2964 635 2996 636
rect 2964 605 2965 635
rect 2965 605 2995 635
rect 2995 605 2996 635
rect 2964 604 2996 605
rect 2964 555 2996 556
rect 2964 525 2965 555
rect 2965 525 2995 555
rect 2995 525 2996 555
rect 2964 524 2996 525
rect 2964 444 2996 476
rect 2964 395 2996 396
rect 2964 365 2965 395
rect 2965 365 2995 395
rect 2995 365 2996 395
rect 2964 364 2996 365
rect 2964 284 2996 316
rect 2964 235 2996 236
rect 2964 205 2965 235
rect 2965 205 2995 235
rect 2995 205 2996 235
rect 2964 204 2996 205
rect 2964 124 2996 156
rect 2964 75 2996 76
rect 2964 45 2965 75
rect 2965 45 2995 75
rect 2995 45 2996 75
rect 2964 44 2996 45
rect 2964 -5 2996 -4
rect 2964 -35 2965 -5
rect 2965 -35 2995 -5
rect 2995 -35 2996 -5
rect 2964 -36 2996 -35
rect 2964 -85 2996 -84
rect 2964 -115 2965 -85
rect 2965 -115 2995 -85
rect 2995 -115 2996 -85
rect 2964 -116 2996 -115
rect 2964 -165 2996 -164
rect 2964 -195 2965 -165
rect 2965 -195 2995 -165
rect 2995 -195 2996 -165
rect 2964 -196 2996 -195
rect 2964 -245 2996 -244
rect 2964 -275 2965 -245
rect 2965 -275 2995 -245
rect 2995 -275 2996 -245
rect 2964 -276 2996 -275
rect 2964 -325 2996 -324
rect 2964 -355 2965 -325
rect 2965 -355 2995 -325
rect 2995 -355 2996 -325
rect 2964 -356 2996 -355
rect 2964 -436 2996 -404
rect 2964 -485 2996 -484
rect 2964 -515 2965 -485
rect 2965 -515 2995 -485
rect 2995 -515 2996 -485
rect 2964 -516 2996 -515
rect 2964 -596 2996 -564
rect 2964 -645 2996 -644
rect 2964 -675 2965 -645
rect 2965 -675 2995 -645
rect 2995 -675 2996 -645
rect 2964 -676 2996 -675
rect 2964 -756 2996 -724
rect 2964 -805 2996 -804
rect 2964 -835 2965 -805
rect 2965 -835 2995 -805
rect 2995 -835 2996 -805
rect 2964 -836 2996 -835
rect 2964 -885 2996 -884
rect 2964 -915 2965 -885
rect 2965 -915 2995 -885
rect 2995 -915 2996 -885
rect 2964 -916 2996 -915
rect 2964 -996 2996 -964
rect 2964 -1076 2996 -1044
rect 2964 -1125 2996 -1124
rect 2964 -1155 2965 -1125
rect 2965 -1155 2995 -1125
rect 2995 -1155 2996 -1125
rect 2964 -1156 2996 -1155
rect 2964 -1205 2996 -1204
rect 2964 -1235 2965 -1205
rect 2965 -1235 2995 -1205
rect 2995 -1235 2996 -1205
rect 2964 -1236 2996 -1235
rect 2964 -1285 2996 -1284
rect 2964 -1315 2965 -1285
rect 2965 -1315 2995 -1285
rect 2995 -1315 2996 -1285
rect 2964 -1316 2996 -1315
rect 2964 -1365 2996 -1364
rect 2964 -1395 2965 -1365
rect 2965 -1395 2995 -1365
rect 2995 -1395 2996 -1365
rect 2964 -1396 2996 -1395
rect 2964 -1445 2996 -1444
rect 2964 -1475 2965 -1445
rect 2965 -1475 2995 -1445
rect 2995 -1475 2996 -1445
rect 2964 -1476 2996 -1475
rect 2964 -1525 2996 -1524
rect 2964 -1555 2965 -1525
rect 2965 -1555 2995 -1525
rect 2995 -1555 2996 -1525
rect 2964 -1556 2996 -1555
rect 2964 -1636 2996 -1604
rect 2964 -1716 2996 -1684
rect 2964 -1765 2996 -1764
rect 2964 -1795 2965 -1765
rect 2965 -1795 2995 -1765
rect 2995 -1795 2996 -1765
rect 2964 -1796 2996 -1795
rect 2964 -1845 2996 -1844
rect 2964 -1875 2965 -1845
rect 2965 -1875 2995 -1845
rect 2995 -1875 2996 -1845
rect 2964 -1876 2996 -1875
rect 2964 -1956 2996 -1924
rect 2964 -2005 2996 -2004
rect 2964 -2035 2965 -2005
rect 2965 -2035 2995 -2005
rect 2995 -2035 2996 -2005
rect 2964 -2036 2996 -2035
rect 2964 -2116 2996 -2084
rect 2964 -2165 2996 -2164
rect 2964 -2195 2965 -2165
rect 2965 -2195 2995 -2165
rect 2995 -2195 2996 -2165
rect 2964 -2196 2996 -2195
rect 2964 -2276 2996 -2244
rect 2964 -2325 2996 -2324
rect 2964 -2355 2965 -2325
rect 2965 -2355 2995 -2325
rect 2995 -2355 2996 -2325
rect 2964 -2356 2996 -2355
rect 2964 -2405 2996 -2404
rect 2964 -2435 2965 -2405
rect 2965 -2435 2995 -2405
rect 2995 -2435 2996 -2405
rect 2964 -2436 2996 -2435
rect 2964 -2485 2996 -2484
rect 2964 -2515 2965 -2485
rect 2965 -2515 2995 -2485
rect 2995 -2515 2996 -2485
rect 2964 -2516 2996 -2515
rect 2964 -2565 2996 -2564
rect 2964 -2595 2965 -2565
rect 2965 -2595 2995 -2565
rect 2995 -2595 2996 -2565
rect 2964 -2596 2996 -2595
rect 2964 -2645 2996 -2644
rect 2964 -2675 2965 -2645
rect 2965 -2675 2995 -2645
rect 2995 -2675 2996 -2645
rect 2964 -2676 2996 -2675
rect 2964 -2725 2996 -2724
rect 2964 -2755 2965 -2725
rect 2965 -2755 2995 -2725
rect 2995 -2755 2996 -2725
rect 2964 -2756 2996 -2755
rect 2964 -2836 2996 -2804
rect 2964 -2885 2996 -2884
rect 2964 -2915 2965 -2885
rect 2965 -2915 2995 -2885
rect 2995 -2915 2996 -2885
rect 2964 -2916 2996 -2915
rect 2964 -2996 2996 -2964
rect 2964 -3045 2996 -3044
rect 2964 -3075 2965 -3045
rect 2965 -3075 2995 -3045
rect 2995 -3075 2996 -3045
rect 2964 -3076 2996 -3075
rect 2964 -3156 2996 -3124
rect 2964 -3205 2996 -3204
rect 2964 -3235 2965 -3205
rect 2965 -3235 2995 -3205
rect 2995 -3235 2996 -3205
rect 2964 -3236 2996 -3235
rect 2964 -3285 2996 -3284
rect 2964 -3315 2965 -3285
rect 2965 -3315 2995 -3285
rect 2995 -3315 2996 -3285
rect 2964 -3316 2996 -3315
rect 2964 -3396 2996 -3364
rect 2964 -3476 2996 -3444
rect 2964 -3525 2996 -3524
rect 2964 -3555 2965 -3525
rect 2965 -3555 2995 -3525
rect 2995 -3555 2996 -3525
rect 2964 -3556 2996 -3555
rect 2964 -3605 2996 -3604
rect 2964 -3635 2965 -3605
rect 2965 -3635 2995 -3605
rect 2995 -3635 2996 -3605
rect 2964 -3636 2996 -3635
rect 2964 -3685 2996 -3684
rect 2964 -3715 2965 -3685
rect 2965 -3715 2995 -3685
rect 2995 -3715 2996 -3685
rect 2964 -3716 2996 -3715
rect 3044 1035 3076 1036
rect 3044 1005 3045 1035
rect 3045 1005 3075 1035
rect 3075 1005 3076 1035
rect 3044 1004 3076 1005
rect 3044 955 3076 956
rect 3044 925 3045 955
rect 3045 925 3075 955
rect 3075 925 3076 955
rect 3044 924 3076 925
rect 3044 875 3076 876
rect 3044 845 3045 875
rect 3045 845 3075 875
rect 3075 845 3076 875
rect 3044 844 3076 845
rect 3044 764 3076 796
rect 3044 684 3076 716
rect 3044 635 3076 636
rect 3044 605 3045 635
rect 3045 605 3075 635
rect 3075 605 3076 635
rect 3044 604 3076 605
rect 3044 555 3076 556
rect 3044 525 3045 555
rect 3045 525 3075 555
rect 3075 525 3076 555
rect 3044 524 3076 525
rect 3044 444 3076 476
rect 3044 395 3076 396
rect 3044 365 3045 395
rect 3045 365 3075 395
rect 3075 365 3076 395
rect 3044 364 3076 365
rect 3044 284 3076 316
rect 3044 235 3076 236
rect 3044 205 3045 235
rect 3045 205 3075 235
rect 3075 205 3076 235
rect 3044 204 3076 205
rect 3044 124 3076 156
rect 3044 75 3076 76
rect 3044 45 3045 75
rect 3045 45 3075 75
rect 3075 45 3076 75
rect 3044 44 3076 45
rect 3044 -5 3076 -4
rect 3044 -35 3045 -5
rect 3045 -35 3075 -5
rect 3075 -35 3076 -5
rect 3044 -36 3076 -35
rect 3044 -85 3076 -84
rect 3044 -115 3045 -85
rect 3045 -115 3075 -85
rect 3075 -115 3076 -85
rect 3044 -116 3076 -115
rect 3044 -165 3076 -164
rect 3044 -195 3045 -165
rect 3045 -195 3075 -165
rect 3075 -195 3076 -165
rect 3044 -196 3076 -195
rect 3044 -245 3076 -244
rect 3044 -275 3045 -245
rect 3045 -275 3075 -245
rect 3075 -275 3076 -245
rect 3044 -276 3076 -275
rect 3044 -325 3076 -324
rect 3044 -355 3045 -325
rect 3045 -355 3075 -325
rect 3075 -355 3076 -325
rect 3044 -356 3076 -355
rect 3044 -436 3076 -404
rect 3044 -485 3076 -484
rect 3044 -515 3045 -485
rect 3045 -515 3075 -485
rect 3075 -515 3076 -485
rect 3044 -516 3076 -515
rect 3044 -596 3076 -564
rect 3044 -645 3076 -644
rect 3044 -675 3045 -645
rect 3045 -675 3075 -645
rect 3075 -675 3076 -645
rect 3044 -676 3076 -675
rect 3044 -756 3076 -724
rect 3044 -805 3076 -804
rect 3044 -835 3045 -805
rect 3045 -835 3075 -805
rect 3075 -835 3076 -805
rect 3044 -836 3076 -835
rect 3044 -885 3076 -884
rect 3044 -915 3045 -885
rect 3045 -915 3075 -885
rect 3075 -915 3076 -885
rect 3044 -916 3076 -915
rect 3044 -996 3076 -964
rect 3044 -1076 3076 -1044
rect 3044 -1125 3076 -1124
rect 3044 -1155 3045 -1125
rect 3045 -1155 3075 -1125
rect 3075 -1155 3076 -1125
rect 3044 -1156 3076 -1155
rect 3044 -1205 3076 -1204
rect 3044 -1235 3045 -1205
rect 3045 -1235 3075 -1205
rect 3075 -1235 3076 -1205
rect 3044 -1236 3076 -1235
rect 3044 -1285 3076 -1284
rect 3044 -1315 3045 -1285
rect 3045 -1315 3075 -1285
rect 3075 -1315 3076 -1285
rect 3044 -1316 3076 -1315
rect 3044 -1365 3076 -1364
rect 3044 -1395 3045 -1365
rect 3045 -1395 3075 -1365
rect 3075 -1395 3076 -1365
rect 3044 -1396 3076 -1395
rect 3044 -1445 3076 -1444
rect 3044 -1475 3045 -1445
rect 3045 -1475 3075 -1445
rect 3075 -1475 3076 -1445
rect 3044 -1476 3076 -1475
rect 3044 -1525 3076 -1524
rect 3044 -1555 3045 -1525
rect 3045 -1555 3075 -1525
rect 3075 -1555 3076 -1525
rect 3044 -1556 3076 -1555
rect 3044 -1636 3076 -1604
rect 3044 -1716 3076 -1684
rect 3044 -1765 3076 -1764
rect 3044 -1795 3045 -1765
rect 3045 -1795 3075 -1765
rect 3075 -1795 3076 -1765
rect 3044 -1796 3076 -1795
rect 3044 -1845 3076 -1844
rect 3044 -1875 3045 -1845
rect 3045 -1875 3075 -1845
rect 3075 -1875 3076 -1845
rect 3044 -1876 3076 -1875
rect 3044 -1956 3076 -1924
rect 3044 -2005 3076 -2004
rect 3044 -2035 3045 -2005
rect 3045 -2035 3075 -2005
rect 3075 -2035 3076 -2005
rect 3044 -2036 3076 -2035
rect 3044 -2116 3076 -2084
rect 3044 -2165 3076 -2164
rect 3044 -2195 3045 -2165
rect 3045 -2195 3075 -2165
rect 3075 -2195 3076 -2165
rect 3044 -2196 3076 -2195
rect 3044 -2276 3076 -2244
rect 3044 -2325 3076 -2324
rect 3044 -2355 3045 -2325
rect 3045 -2355 3075 -2325
rect 3075 -2355 3076 -2325
rect 3044 -2356 3076 -2355
rect 3044 -2405 3076 -2404
rect 3044 -2435 3045 -2405
rect 3045 -2435 3075 -2405
rect 3075 -2435 3076 -2405
rect 3044 -2436 3076 -2435
rect 3044 -2485 3076 -2484
rect 3044 -2515 3045 -2485
rect 3045 -2515 3075 -2485
rect 3075 -2515 3076 -2485
rect 3044 -2516 3076 -2515
rect 3044 -2565 3076 -2564
rect 3044 -2595 3045 -2565
rect 3045 -2595 3075 -2565
rect 3075 -2595 3076 -2565
rect 3044 -2596 3076 -2595
rect 3044 -2645 3076 -2644
rect 3044 -2675 3045 -2645
rect 3045 -2675 3075 -2645
rect 3075 -2675 3076 -2645
rect 3044 -2676 3076 -2675
rect 3044 -2725 3076 -2724
rect 3044 -2755 3045 -2725
rect 3045 -2755 3075 -2725
rect 3075 -2755 3076 -2725
rect 3044 -2756 3076 -2755
rect 3044 -2836 3076 -2804
rect 3044 -2885 3076 -2884
rect 3044 -2915 3045 -2885
rect 3045 -2915 3075 -2885
rect 3075 -2915 3076 -2885
rect 3044 -2916 3076 -2915
rect 3044 -2996 3076 -2964
rect 3044 -3045 3076 -3044
rect 3044 -3075 3045 -3045
rect 3045 -3075 3075 -3045
rect 3075 -3075 3076 -3045
rect 3044 -3076 3076 -3075
rect 3044 -3156 3076 -3124
rect 3044 -3205 3076 -3204
rect 3044 -3235 3045 -3205
rect 3045 -3235 3075 -3205
rect 3075 -3235 3076 -3205
rect 3044 -3236 3076 -3235
rect 3044 -3285 3076 -3284
rect 3044 -3315 3045 -3285
rect 3045 -3315 3075 -3285
rect 3075 -3315 3076 -3285
rect 3044 -3316 3076 -3315
rect 3044 -3396 3076 -3364
rect 3044 -3476 3076 -3444
rect 3044 -3525 3076 -3524
rect 3044 -3555 3045 -3525
rect 3045 -3555 3075 -3525
rect 3075 -3555 3076 -3525
rect 3044 -3556 3076 -3555
rect 3044 -3605 3076 -3604
rect 3044 -3635 3045 -3605
rect 3045 -3635 3075 -3605
rect 3075 -3635 3076 -3605
rect 3044 -3636 3076 -3635
rect 3044 -3685 3076 -3684
rect 3044 -3715 3045 -3685
rect 3045 -3715 3075 -3685
rect 3075 -3715 3076 -3685
rect 3044 -3716 3076 -3715
rect 3124 1035 3156 1036
rect 3124 1005 3125 1035
rect 3125 1005 3155 1035
rect 3155 1005 3156 1035
rect 3124 1004 3156 1005
rect 3124 955 3156 956
rect 3124 925 3125 955
rect 3125 925 3155 955
rect 3155 925 3156 955
rect 3124 924 3156 925
rect 3124 875 3156 876
rect 3124 845 3125 875
rect 3125 845 3155 875
rect 3155 845 3156 875
rect 3124 844 3156 845
rect 3124 764 3156 796
rect 3124 684 3156 716
rect 3124 635 3156 636
rect 3124 605 3125 635
rect 3125 605 3155 635
rect 3155 605 3156 635
rect 3124 604 3156 605
rect 3124 555 3156 556
rect 3124 525 3125 555
rect 3125 525 3155 555
rect 3155 525 3156 555
rect 3124 524 3156 525
rect 3124 444 3156 476
rect 3124 395 3156 396
rect 3124 365 3125 395
rect 3125 365 3155 395
rect 3155 365 3156 395
rect 3124 364 3156 365
rect 3124 284 3156 316
rect 3124 235 3156 236
rect 3124 205 3125 235
rect 3125 205 3155 235
rect 3155 205 3156 235
rect 3124 204 3156 205
rect 3124 124 3156 156
rect 3124 75 3156 76
rect 3124 45 3125 75
rect 3125 45 3155 75
rect 3155 45 3156 75
rect 3124 44 3156 45
rect 3124 -5 3156 -4
rect 3124 -35 3125 -5
rect 3125 -35 3155 -5
rect 3155 -35 3156 -5
rect 3124 -36 3156 -35
rect 3124 -85 3156 -84
rect 3124 -115 3125 -85
rect 3125 -115 3155 -85
rect 3155 -115 3156 -85
rect 3124 -116 3156 -115
rect 3124 -165 3156 -164
rect 3124 -195 3125 -165
rect 3125 -195 3155 -165
rect 3155 -195 3156 -165
rect 3124 -196 3156 -195
rect 3124 -245 3156 -244
rect 3124 -275 3125 -245
rect 3125 -275 3155 -245
rect 3155 -275 3156 -245
rect 3124 -276 3156 -275
rect 3124 -325 3156 -324
rect 3124 -355 3125 -325
rect 3125 -355 3155 -325
rect 3155 -355 3156 -325
rect 3124 -356 3156 -355
rect 3124 -436 3156 -404
rect 3124 -485 3156 -484
rect 3124 -515 3125 -485
rect 3125 -515 3155 -485
rect 3155 -515 3156 -485
rect 3124 -516 3156 -515
rect 3124 -596 3156 -564
rect 3124 -645 3156 -644
rect 3124 -675 3125 -645
rect 3125 -675 3155 -645
rect 3155 -675 3156 -645
rect 3124 -676 3156 -675
rect 3124 -756 3156 -724
rect 3124 -805 3156 -804
rect 3124 -835 3125 -805
rect 3125 -835 3155 -805
rect 3155 -835 3156 -805
rect 3124 -836 3156 -835
rect 3124 -885 3156 -884
rect 3124 -915 3125 -885
rect 3125 -915 3155 -885
rect 3155 -915 3156 -885
rect 3124 -916 3156 -915
rect 3124 -996 3156 -964
rect 3124 -1076 3156 -1044
rect 3124 -1125 3156 -1124
rect 3124 -1155 3125 -1125
rect 3125 -1155 3155 -1125
rect 3155 -1155 3156 -1125
rect 3124 -1156 3156 -1155
rect 3124 -1205 3156 -1204
rect 3124 -1235 3125 -1205
rect 3125 -1235 3155 -1205
rect 3155 -1235 3156 -1205
rect 3124 -1236 3156 -1235
rect 3124 -1285 3156 -1284
rect 3124 -1315 3125 -1285
rect 3125 -1315 3155 -1285
rect 3155 -1315 3156 -1285
rect 3124 -1316 3156 -1315
rect 3124 -1365 3156 -1364
rect 3124 -1395 3125 -1365
rect 3125 -1395 3155 -1365
rect 3155 -1395 3156 -1365
rect 3124 -1396 3156 -1395
rect 3124 -1445 3156 -1444
rect 3124 -1475 3125 -1445
rect 3125 -1475 3155 -1445
rect 3155 -1475 3156 -1445
rect 3124 -1476 3156 -1475
rect 3124 -1525 3156 -1524
rect 3124 -1555 3125 -1525
rect 3125 -1555 3155 -1525
rect 3155 -1555 3156 -1525
rect 3124 -1556 3156 -1555
rect 3124 -1636 3156 -1604
rect 3124 -1716 3156 -1684
rect 3124 -1765 3156 -1764
rect 3124 -1795 3125 -1765
rect 3125 -1795 3155 -1765
rect 3155 -1795 3156 -1765
rect 3124 -1796 3156 -1795
rect 3124 -1845 3156 -1844
rect 3124 -1875 3125 -1845
rect 3125 -1875 3155 -1845
rect 3155 -1875 3156 -1845
rect 3124 -1876 3156 -1875
rect 3124 -1956 3156 -1924
rect 3124 -2005 3156 -2004
rect 3124 -2035 3125 -2005
rect 3125 -2035 3155 -2005
rect 3155 -2035 3156 -2005
rect 3124 -2036 3156 -2035
rect 3124 -2116 3156 -2084
rect 3124 -2165 3156 -2164
rect 3124 -2195 3125 -2165
rect 3125 -2195 3155 -2165
rect 3155 -2195 3156 -2165
rect 3124 -2196 3156 -2195
rect 3124 -2276 3156 -2244
rect 3124 -2325 3156 -2324
rect 3124 -2355 3125 -2325
rect 3125 -2355 3155 -2325
rect 3155 -2355 3156 -2325
rect 3124 -2356 3156 -2355
rect 3124 -2405 3156 -2404
rect 3124 -2435 3125 -2405
rect 3125 -2435 3155 -2405
rect 3155 -2435 3156 -2405
rect 3124 -2436 3156 -2435
rect 3124 -2485 3156 -2484
rect 3124 -2515 3125 -2485
rect 3125 -2515 3155 -2485
rect 3155 -2515 3156 -2485
rect 3124 -2516 3156 -2515
rect 3124 -2565 3156 -2564
rect 3124 -2595 3125 -2565
rect 3125 -2595 3155 -2565
rect 3155 -2595 3156 -2565
rect 3124 -2596 3156 -2595
rect 3124 -2645 3156 -2644
rect 3124 -2675 3125 -2645
rect 3125 -2675 3155 -2645
rect 3155 -2675 3156 -2645
rect 3124 -2676 3156 -2675
rect 3124 -2725 3156 -2724
rect 3124 -2755 3125 -2725
rect 3125 -2755 3155 -2725
rect 3155 -2755 3156 -2725
rect 3124 -2756 3156 -2755
rect 3124 -2836 3156 -2804
rect 3124 -2885 3156 -2884
rect 3124 -2915 3125 -2885
rect 3125 -2915 3155 -2885
rect 3155 -2915 3156 -2885
rect 3124 -2916 3156 -2915
rect 3124 -2996 3156 -2964
rect 3124 -3045 3156 -3044
rect 3124 -3075 3125 -3045
rect 3125 -3075 3155 -3045
rect 3155 -3075 3156 -3045
rect 3124 -3076 3156 -3075
rect 3124 -3156 3156 -3124
rect 3124 -3205 3156 -3204
rect 3124 -3235 3125 -3205
rect 3125 -3235 3155 -3205
rect 3155 -3235 3156 -3205
rect 3124 -3236 3156 -3235
rect 3124 -3285 3156 -3284
rect 3124 -3315 3125 -3285
rect 3125 -3315 3155 -3285
rect 3155 -3315 3156 -3285
rect 3124 -3316 3156 -3315
rect 3124 -3396 3156 -3364
rect 3124 -3476 3156 -3444
rect 3124 -3525 3156 -3524
rect 3124 -3555 3125 -3525
rect 3125 -3555 3155 -3525
rect 3155 -3555 3156 -3525
rect 3124 -3556 3156 -3555
rect 3124 -3605 3156 -3604
rect 3124 -3635 3125 -3605
rect 3125 -3635 3155 -3605
rect 3155 -3635 3156 -3605
rect 3124 -3636 3156 -3635
rect 3124 -3685 3156 -3684
rect 3124 -3715 3125 -3685
rect 3125 -3715 3155 -3685
rect 3155 -3715 3156 -3685
rect 3124 -3716 3156 -3715
rect 3204 1035 3236 1036
rect 3204 1005 3205 1035
rect 3205 1005 3235 1035
rect 3235 1005 3236 1035
rect 3204 1004 3236 1005
rect 3204 955 3236 956
rect 3204 925 3205 955
rect 3205 925 3235 955
rect 3235 925 3236 955
rect 3204 924 3236 925
rect 3204 875 3236 876
rect 3204 845 3205 875
rect 3205 845 3235 875
rect 3235 845 3236 875
rect 3204 844 3236 845
rect 3204 764 3236 796
rect 3204 684 3236 716
rect 3204 635 3236 636
rect 3204 605 3205 635
rect 3205 605 3235 635
rect 3235 605 3236 635
rect 3204 604 3236 605
rect 3204 555 3236 556
rect 3204 525 3205 555
rect 3205 525 3235 555
rect 3235 525 3236 555
rect 3204 524 3236 525
rect 3204 444 3236 476
rect 3204 395 3236 396
rect 3204 365 3205 395
rect 3205 365 3235 395
rect 3235 365 3236 395
rect 3204 364 3236 365
rect 3204 284 3236 316
rect 3204 235 3236 236
rect 3204 205 3205 235
rect 3205 205 3235 235
rect 3235 205 3236 235
rect 3204 204 3236 205
rect 3204 124 3236 156
rect 3204 75 3236 76
rect 3204 45 3205 75
rect 3205 45 3235 75
rect 3235 45 3236 75
rect 3204 44 3236 45
rect 3204 -5 3236 -4
rect 3204 -35 3205 -5
rect 3205 -35 3235 -5
rect 3235 -35 3236 -5
rect 3204 -36 3236 -35
rect 3204 -85 3236 -84
rect 3204 -115 3205 -85
rect 3205 -115 3235 -85
rect 3235 -115 3236 -85
rect 3204 -116 3236 -115
rect 3204 -165 3236 -164
rect 3204 -195 3205 -165
rect 3205 -195 3235 -165
rect 3235 -195 3236 -165
rect 3204 -196 3236 -195
rect 3204 -245 3236 -244
rect 3204 -275 3205 -245
rect 3205 -275 3235 -245
rect 3235 -275 3236 -245
rect 3204 -276 3236 -275
rect 3204 -325 3236 -324
rect 3204 -355 3205 -325
rect 3205 -355 3235 -325
rect 3235 -355 3236 -325
rect 3204 -356 3236 -355
rect 3204 -436 3236 -404
rect 3204 -485 3236 -484
rect 3204 -515 3205 -485
rect 3205 -515 3235 -485
rect 3235 -515 3236 -485
rect 3204 -516 3236 -515
rect 3204 -596 3236 -564
rect 3204 -645 3236 -644
rect 3204 -675 3205 -645
rect 3205 -675 3235 -645
rect 3235 -675 3236 -645
rect 3204 -676 3236 -675
rect 3204 -756 3236 -724
rect 3204 -805 3236 -804
rect 3204 -835 3205 -805
rect 3205 -835 3235 -805
rect 3235 -835 3236 -805
rect 3204 -836 3236 -835
rect 3204 -885 3236 -884
rect 3204 -915 3205 -885
rect 3205 -915 3235 -885
rect 3235 -915 3236 -885
rect 3204 -916 3236 -915
rect 3204 -996 3236 -964
rect 3204 -1076 3236 -1044
rect 3204 -1125 3236 -1124
rect 3204 -1155 3205 -1125
rect 3205 -1155 3235 -1125
rect 3235 -1155 3236 -1125
rect 3204 -1156 3236 -1155
rect 3204 -1205 3236 -1204
rect 3204 -1235 3205 -1205
rect 3205 -1235 3235 -1205
rect 3235 -1235 3236 -1205
rect 3204 -1236 3236 -1235
rect 3204 -1285 3236 -1284
rect 3204 -1315 3205 -1285
rect 3205 -1315 3235 -1285
rect 3235 -1315 3236 -1285
rect 3204 -1316 3236 -1315
rect 3204 -1365 3236 -1364
rect 3204 -1395 3205 -1365
rect 3205 -1395 3235 -1365
rect 3235 -1395 3236 -1365
rect 3204 -1396 3236 -1395
rect 3204 -1445 3236 -1444
rect 3204 -1475 3205 -1445
rect 3205 -1475 3235 -1445
rect 3235 -1475 3236 -1445
rect 3204 -1476 3236 -1475
rect 3204 -1525 3236 -1524
rect 3204 -1555 3205 -1525
rect 3205 -1555 3235 -1525
rect 3235 -1555 3236 -1525
rect 3204 -1556 3236 -1555
rect 3204 -1636 3236 -1604
rect 3204 -1716 3236 -1684
rect 3204 -1765 3236 -1764
rect 3204 -1795 3205 -1765
rect 3205 -1795 3235 -1765
rect 3235 -1795 3236 -1765
rect 3204 -1796 3236 -1795
rect 3204 -1845 3236 -1844
rect 3204 -1875 3205 -1845
rect 3205 -1875 3235 -1845
rect 3235 -1875 3236 -1845
rect 3204 -1876 3236 -1875
rect 3204 -1956 3236 -1924
rect 3204 -2005 3236 -2004
rect 3204 -2035 3205 -2005
rect 3205 -2035 3235 -2005
rect 3235 -2035 3236 -2005
rect 3204 -2036 3236 -2035
rect 3204 -2116 3236 -2084
rect 3204 -2165 3236 -2164
rect 3204 -2195 3205 -2165
rect 3205 -2195 3235 -2165
rect 3235 -2195 3236 -2165
rect 3204 -2196 3236 -2195
rect 3204 -2276 3236 -2244
rect 3204 -2325 3236 -2324
rect 3204 -2355 3205 -2325
rect 3205 -2355 3235 -2325
rect 3235 -2355 3236 -2325
rect 3204 -2356 3236 -2355
rect 3204 -2405 3236 -2404
rect 3204 -2435 3205 -2405
rect 3205 -2435 3235 -2405
rect 3235 -2435 3236 -2405
rect 3204 -2436 3236 -2435
rect 3204 -2485 3236 -2484
rect 3204 -2515 3205 -2485
rect 3205 -2515 3235 -2485
rect 3235 -2515 3236 -2485
rect 3204 -2516 3236 -2515
rect 3204 -2565 3236 -2564
rect 3204 -2595 3205 -2565
rect 3205 -2595 3235 -2565
rect 3235 -2595 3236 -2565
rect 3204 -2596 3236 -2595
rect 3204 -2645 3236 -2644
rect 3204 -2675 3205 -2645
rect 3205 -2675 3235 -2645
rect 3235 -2675 3236 -2645
rect 3204 -2676 3236 -2675
rect 3204 -2725 3236 -2724
rect 3204 -2755 3205 -2725
rect 3205 -2755 3235 -2725
rect 3235 -2755 3236 -2725
rect 3204 -2756 3236 -2755
rect 3204 -2836 3236 -2804
rect 3204 -2885 3236 -2884
rect 3204 -2915 3205 -2885
rect 3205 -2915 3235 -2885
rect 3235 -2915 3236 -2885
rect 3204 -2916 3236 -2915
rect 3204 -2996 3236 -2964
rect 3204 -3045 3236 -3044
rect 3204 -3075 3205 -3045
rect 3205 -3075 3235 -3045
rect 3235 -3075 3236 -3045
rect 3204 -3076 3236 -3075
rect 3204 -3156 3236 -3124
rect 3204 -3205 3236 -3204
rect 3204 -3235 3205 -3205
rect 3205 -3235 3235 -3205
rect 3235 -3235 3236 -3205
rect 3204 -3236 3236 -3235
rect 3204 -3285 3236 -3284
rect 3204 -3315 3205 -3285
rect 3205 -3315 3235 -3285
rect 3235 -3315 3236 -3285
rect 3204 -3316 3236 -3315
rect 3204 -3396 3236 -3364
rect 3204 -3476 3236 -3444
rect 3204 -3525 3236 -3524
rect 3204 -3555 3205 -3525
rect 3205 -3555 3235 -3525
rect 3235 -3555 3236 -3525
rect 3204 -3556 3236 -3555
rect 3204 -3605 3236 -3604
rect 3204 -3635 3205 -3605
rect 3205 -3635 3235 -3605
rect 3235 -3635 3236 -3605
rect 3204 -3636 3236 -3635
rect 3204 -3685 3236 -3684
rect 3204 -3715 3205 -3685
rect 3205 -3715 3235 -3685
rect 3235 -3715 3236 -3685
rect 3204 -3716 3236 -3715
rect 3284 1035 3316 1036
rect 3284 1005 3285 1035
rect 3285 1005 3315 1035
rect 3315 1005 3316 1035
rect 3284 1004 3316 1005
rect 3284 955 3316 956
rect 3284 925 3285 955
rect 3285 925 3315 955
rect 3315 925 3316 955
rect 3284 924 3316 925
rect 3284 875 3316 876
rect 3284 845 3285 875
rect 3285 845 3315 875
rect 3315 845 3316 875
rect 3284 844 3316 845
rect 3284 764 3316 796
rect 3284 684 3316 716
rect 3284 635 3316 636
rect 3284 605 3285 635
rect 3285 605 3315 635
rect 3315 605 3316 635
rect 3284 604 3316 605
rect 3284 555 3316 556
rect 3284 525 3285 555
rect 3285 525 3315 555
rect 3315 525 3316 555
rect 3284 524 3316 525
rect 3284 444 3316 476
rect 3284 395 3316 396
rect 3284 365 3285 395
rect 3285 365 3315 395
rect 3315 365 3316 395
rect 3284 364 3316 365
rect 3284 284 3316 316
rect 3284 235 3316 236
rect 3284 205 3285 235
rect 3285 205 3315 235
rect 3315 205 3316 235
rect 3284 204 3316 205
rect 3284 124 3316 156
rect 3284 75 3316 76
rect 3284 45 3285 75
rect 3285 45 3315 75
rect 3315 45 3316 75
rect 3284 44 3316 45
rect 3284 -5 3316 -4
rect 3284 -35 3285 -5
rect 3285 -35 3315 -5
rect 3315 -35 3316 -5
rect 3284 -36 3316 -35
rect 3284 -85 3316 -84
rect 3284 -115 3285 -85
rect 3285 -115 3315 -85
rect 3315 -115 3316 -85
rect 3284 -116 3316 -115
rect 3284 -165 3316 -164
rect 3284 -195 3285 -165
rect 3285 -195 3315 -165
rect 3315 -195 3316 -165
rect 3284 -196 3316 -195
rect 3284 -245 3316 -244
rect 3284 -275 3285 -245
rect 3285 -275 3315 -245
rect 3315 -275 3316 -245
rect 3284 -276 3316 -275
rect 3284 -325 3316 -324
rect 3284 -355 3285 -325
rect 3285 -355 3315 -325
rect 3315 -355 3316 -325
rect 3284 -356 3316 -355
rect 3284 -436 3316 -404
rect 3284 -485 3316 -484
rect 3284 -515 3285 -485
rect 3285 -515 3315 -485
rect 3315 -515 3316 -485
rect 3284 -516 3316 -515
rect 3284 -596 3316 -564
rect 3284 -645 3316 -644
rect 3284 -675 3285 -645
rect 3285 -675 3315 -645
rect 3315 -675 3316 -645
rect 3284 -676 3316 -675
rect 3284 -756 3316 -724
rect 3284 -805 3316 -804
rect 3284 -835 3285 -805
rect 3285 -835 3315 -805
rect 3315 -835 3316 -805
rect 3284 -836 3316 -835
rect 3284 -885 3316 -884
rect 3284 -915 3285 -885
rect 3285 -915 3315 -885
rect 3315 -915 3316 -885
rect 3284 -916 3316 -915
rect 3284 -996 3316 -964
rect 3284 -1076 3316 -1044
rect 3284 -1125 3316 -1124
rect 3284 -1155 3285 -1125
rect 3285 -1155 3315 -1125
rect 3315 -1155 3316 -1125
rect 3284 -1156 3316 -1155
rect 3284 -1205 3316 -1204
rect 3284 -1235 3285 -1205
rect 3285 -1235 3315 -1205
rect 3315 -1235 3316 -1205
rect 3284 -1236 3316 -1235
rect 3284 -1285 3316 -1284
rect 3284 -1315 3285 -1285
rect 3285 -1315 3315 -1285
rect 3315 -1315 3316 -1285
rect 3284 -1316 3316 -1315
rect 3284 -1365 3316 -1364
rect 3284 -1395 3285 -1365
rect 3285 -1395 3315 -1365
rect 3315 -1395 3316 -1365
rect 3284 -1396 3316 -1395
rect 3284 -1445 3316 -1444
rect 3284 -1475 3285 -1445
rect 3285 -1475 3315 -1445
rect 3315 -1475 3316 -1445
rect 3284 -1476 3316 -1475
rect 3284 -1525 3316 -1524
rect 3284 -1555 3285 -1525
rect 3285 -1555 3315 -1525
rect 3315 -1555 3316 -1525
rect 3284 -1556 3316 -1555
rect 3284 -1636 3316 -1604
rect 3284 -1716 3316 -1684
rect 3284 -1765 3316 -1764
rect 3284 -1795 3285 -1765
rect 3285 -1795 3315 -1765
rect 3315 -1795 3316 -1765
rect 3284 -1796 3316 -1795
rect 3284 -1845 3316 -1844
rect 3284 -1875 3285 -1845
rect 3285 -1875 3315 -1845
rect 3315 -1875 3316 -1845
rect 3284 -1876 3316 -1875
rect 3284 -1956 3316 -1924
rect 3284 -2005 3316 -2004
rect 3284 -2035 3285 -2005
rect 3285 -2035 3315 -2005
rect 3315 -2035 3316 -2005
rect 3284 -2036 3316 -2035
rect 3284 -2116 3316 -2084
rect 3284 -2165 3316 -2164
rect 3284 -2195 3285 -2165
rect 3285 -2195 3315 -2165
rect 3315 -2195 3316 -2165
rect 3284 -2196 3316 -2195
rect 3284 -2276 3316 -2244
rect 3284 -2325 3316 -2324
rect 3284 -2355 3285 -2325
rect 3285 -2355 3315 -2325
rect 3315 -2355 3316 -2325
rect 3284 -2356 3316 -2355
rect 3284 -2405 3316 -2404
rect 3284 -2435 3285 -2405
rect 3285 -2435 3315 -2405
rect 3315 -2435 3316 -2405
rect 3284 -2436 3316 -2435
rect 3284 -2485 3316 -2484
rect 3284 -2515 3285 -2485
rect 3285 -2515 3315 -2485
rect 3315 -2515 3316 -2485
rect 3284 -2516 3316 -2515
rect 3284 -2565 3316 -2564
rect 3284 -2595 3285 -2565
rect 3285 -2595 3315 -2565
rect 3315 -2595 3316 -2565
rect 3284 -2596 3316 -2595
rect 3284 -2645 3316 -2644
rect 3284 -2675 3285 -2645
rect 3285 -2675 3315 -2645
rect 3315 -2675 3316 -2645
rect 3284 -2676 3316 -2675
rect 3284 -2725 3316 -2724
rect 3284 -2755 3285 -2725
rect 3285 -2755 3315 -2725
rect 3315 -2755 3316 -2725
rect 3284 -2756 3316 -2755
rect 3284 -2836 3316 -2804
rect 3284 -2885 3316 -2884
rect 3284 -2915 3285 -2885
rect 3285 -2915 3315 -2885
rect 3315 -2915 3316 -2885
rect 3284 -2916 3316 -2915
rect 3284 -2996 3316 -2964
rect 3284 -3045 3316 -3044
rect 3284 -3075 3285 -3045
rect 3285 -3075 3315 -3045
rect 3315 -3075 3316 -3045
rect 3284 -3076 3316 -3075
rect 3284 -3156 3316 -3124
rect 3284 -3205 3316 -3204
rect 3284 -3235 3285 -3205
rect 3285 -3235 3315 -3205
rect 3315 -3235 3316 -3205
rect 3284 -3236 3316 -3235
rect 3284 -3285 3316 -3284
rect 3284 -3315 3285 -3285
rect 3285 -3315 3315 -3285
rect 3315 -3315 3316 -3285
rect 3284 -3316 3316 -3315
rect 3284 -3396 3316 -3364
rect 3284 -3476 3316 -3444
rect 3284 -3525 3316 -3524
rect 3284 -3555 3285 -3525
rect 3285 -3555 3315 -3525
rect 3315 -3555 3316 -3525
rect 3284 -3556 3316 -3555
rect 3284 -3605 3316 -3604
rect 3284 -3635 3285 -3605
rect 3285 -3635 3315 -3605
rect 3315 -3635 3316 -3605
rect 3284 -3636 3316 -3635
rect 3284 -3685 3316 -3684
rect 3284 -3715 3285 -3685
rect 3285 -3715 3315 -3685
rect 3315 -3715 3316 -3685
rect 3284 -3716 3316 -3715
rect 3364 1035 3396 1036
rect 3364 1005 3365 1035
rect 3365 1005 3395 1035
rect 3395 1005 3396 1035
rect 3364 1004 3396 1005
rect 3364 955 3396 956
rect 3364 925 3365 955
rect 3365 925 3395 955
rect 3395 925 3396 955
rect 3364 924 3396 925
rect 3364 875 3396 876
rect 3364 845 3365 875
rect 3365 845 3395 875
rect 3395 845 3396 875
rect 3364 844 3396 845
rect 3364 764 3396 796
rect 3364 684 3396 716
rect 3364 635 3396 636
rect 3364 605 3365 635
rect 3365 605 3395 635
rect 3395 605 3396 635
rect 3364 604 3396 605
rect 3364 555 3396 556
rect 3364 525 3365 555
rect 3365 525 3395 555
rect 3395 525 3396 555
rect 3364 524 3396 525
rect 3364 444 3396 476
rect 3364 395 3396 396
rect 3364 365 3365 395
rect 3365 365 3395 395
rect 3395 365 3396 395
rect 3364 364 3396 365
rect 3364 284 3396 316
rect 3364 235 3396 236
rect 3364 205 3365 235
rect 3365 205 3395 235
rect 3395 205 3396 235
rect 3364 204 3396 205
rect 3364 124 3396 156
rect 3364 75 3396 76
rect 3364 45 3365 75
rect 3365 45 3395 75
rect 3395 45 3396 75
rect 3364 44 3396 45
rect 3364 -5 3396 -4
rect 3364 -35 3365 -5
rect 3365 -35 3395 -5
rect 3395 -35 3396 -5
rect 3364 -36 3396 -35
rect 3364 -85 3396 -84
rect 3364 -115 3365 -85
rect 3365 -115 3395 -85
rect 3395 -115 3396 -85
rect 3364 -116 3396 -115
rect 3364 -165 3396 -164
rect 3364 -195 3365 -165
rect 3365 -195 3395 -165
rect 3395 -195 3396 -165
rect 3364 -196 3396 -195
rect 3364 -245 3396 -244
rect 3364 -275 3365 -245
rect 3365 -275 3395 -245
rect 3395 -275 3396 -245
rect 3364 -276 3396 -275
rect 3364 -325 3396 -324
rect 3364 -355 3365 -325
rect 3365 -355 3395 -325
rect 3395 -355 3396 -325
rect 3364 -356 3396 -355
rect 3364 -436 3396 -404
rect 3364 -485 3396 -484
rect 3364 -515 3365 -485
rect 3365 -515 3395 -485
rect 3395 -515 3396 -485
rect 3364 -516 3396 -515
rect 3364 -596 3396 -564
rect 3364 -645 3396 -644
rect 3364 -675 3365 -645
rect 3365 -675 3395 -645
rect 3395 -675 3396 -645
rect 3364 -676 3396 -675
rect 3364 -756 3396 -724
rect 3364 -805 3396 -804
rect 3364 -835 3365 -805
rect 3365 -835 3395 -805
rect 3395 -835 3396 -805
rect 3364 -836 3396 -835
rect 3364 -885 3396 -884
rect 3364 -915 3365 -885
rect 3365 -915 3395 -885
rect 3395 -915 3396 -885
rect 3364 -916 3396 -915
rect 3364 -996 3396 -964
rect 3364 -1076 3396 -1044
rect 3364 -1125 3396 -1124
rect 3364 -1155 3365 -1125
rect 3365 -1155 3395 -1125
rect 3395 -1155 3396 -1125
rect 3364 -1156 3396 -1155
rect 3364 -1205 3396 -1204
rect 3364 -1235 3365 -1205
rect 3365 -1235 3395 -1205
rect 3395 -1235 3396 -1205
rect 3364 -1236 3396 -1235
rect 3364 -1285 3396 -1284
rect 3364 -1315 3365 -1285
rect 3365 -1315 3395 -1285
rect 3395 -1315 3396 -1285
rect 3364 -1316 3396 -1315
rect 3364 -1365 3396 -1364
rect 3364 -1395 3365 -1365
rect 3365 -1395 3395 -1365
rect 3395 -1395 3396 -1365
rect 3364 -1396 3396 -1395
rect 3364 -1445 3396 -1444
rect 3364 -1475 3365 -1445
rect 3365 -1475 3395 -1445
rect 3395 -1475 3396 -1445
rect 3364 -1476 3396 -1475
rect 3364 -1525 3396 -1524
rect 3364 -1555 3365 -1525
rect 3365 -1555 3395 -1525
rect 3395 -1555 3396 -1525
rect 3364 -1556 3396 -1555
rect 3364 -1636 3396 -1604
rect 3364 -1716 3396 -1684
rect 3364 -1765 3396 -1764
rect 3364 -1795 3365 -1765
rect 3365 -1795 3395 -1765
rect 3395 -1795 3396 -1765
rect 3364 -1796 3396 -1795
rect 3364 -1845 3396 -1844
rect 3364 -1875 3365 -1845
rect 3365 -1875 3395 -1845
rect 3395 -1875 3396 -1845
rect 3364 -1876 3396 -1875
rect 3364 -1956 3396 -1924
rect 3364 -2005 3396 -2004
rect 3364 -2035 3365 -2005
rect 3365 -2035 3395 -2005
rect 3395 -2035 3396 -2005
rect 3364 -2036 3396 -2035
rect 3364 -2116 3396 -2084
rect 3364 -2165 3396 -2164
rect 3364 -2195 3365 -2165
rect 3365 -2195 3395 -2165
rect 3395 -2195 3396 -2165
rect 3364 -2196 3396 -2195
rect 3364 -2276 3396 -2244
rect 3364 -2325 3396 -2324
rect 3364 -2355 3365 -2325
rect 3365 -2355 3395 -2325
rect 3395 -2355 3396 -2325
rect 3364 -2356 3396 -2355
rect 3364 -2405 3396 -2404
rect 3364 -2435 3365 -2405
rect 3365 -2435 3395 -2405
rect 3395 -2435 3396 -2405
rect 3364 -2436 3396 -2435
rect 3364 -2485 3396 -2484
rect 3364 -2515 3365 -2485
rect 3365 -2515 3395 -2485
rect 3395 -2515 3396 -2485
rect 3364 -2516 3396 -2515
rect 3364 -2565 3396 -2564
rect 3364 -2595 3365 -2565
rect 3365 -2595 3395 -2565
rect 3395 -2595 3396 -2565
rect 3364 -2596 3396 -2595
rect 3364 -2645 3396 -2644
rect 3364 -2675 3365 -2645
rect 3365 -2675 3395 -2645
rect 3395 -2675 3396 -2645
rect 3364 -2676 3396 -2675
rect 3364 -2725 3396 -2724
rect 3364 -2755 3365 -2725
rect 3365 -2755 3395 -2725
rect 3395 -2755 3396 -2725
rect 3364 -2756 3396 -2755
rect 3364 -2836 3396 -2804
rect 3364 -2885 3396 -2884
rect 3364 -2915 3365 -2885
rect 3365 -2915 3395 -2885
rect 3395 -2915 3396 -2885
rect 3364 -2916 3396 -2915
rect 3364 -2996 3396 -2964
rect 3364 -3045 3396 -3044
rect 3364 -3075 3365 -3045
rect 3365 -3075 3395 -3045
rect 3395 -3075 3396 -3045
rect 3364 -3076 3396 -3075
rect 3364 -3156 3396 -3124
rect 3364 -3205 3396 -3204
rect 3364 -3235 3365 -3205
rect 3365 -3235 3395 -3205
rect 3395 -3235 3396 -3205
rect 3364 -3236 3396 -3235
rect 3364 -3285 3396 -3284
rect 3364 -3315 3365 -3285
rect 3365 -3315 3395 -3285
rect 3395 -3315 3396 -3285
rect 3364 -3316 3396 -3315
rect 3364 -3396 3396 -3364
rect 3364 -3476 3396 -3444
rect 3364 -3525 3396 -3524
rect 3364 -3555 3365 -3525
rect 3365 -3555 3395 -3525
rect 3395 -3555 3396 -3525
rect 3364 -3556 3396 -3555
rect 3364 -3605 3396 -3604
rect 3364 -3635 3365 -3605
rect 3365 -3635 3395 -3605
rect 3395 -3635 3396 -3605
rect 3364 -3636 3396 -3635
rect 3364 -3685 3396 -3684
rect 3364 -3715 3365 -3685
rect 3365 -3715 3395 -3685
rect 3395 -3715 3396 -3685
rect 3364 -3716 3396 -3715
rect 3444 1035 3476 1036
rect 3444 1005 3445 1035
rect 3445 1005 3475 1035
rect 3475 1005 3476 1035
rect 3444 1004 3476 1005
rect 3444 955 3476 956
rect 3444 925 3445 955
rect 3445 925 3475 955
rect 3475 925 3476 955
rect 3444 924 3476 925
rect 3444 875 3476 876
rect 3444 845 3445 875
rect 3445 845 3475 875
rect 3475 845 3476 875
rect 3444 844 3476 845
rect 3444 764 3476 796
rect 3444 684 3476 716
rect 3444 635 3476 636
rect 3444 605 3445 635
rect 3445 605 3475 635
rect 3475 605 3476 635
rect 3444 604 3476 605
rect 3444 555 3476 556
rect 3444 525 3445 555
rect 3445 525 3475 555
rect 3475 525 3476 555
rect 3444 524 3476 525
rect 3444 444 3476 476
rect 3444 395 3476 396
rect 3444 365 3445 395
rect 3445 365 3475 395
rect 3475 365 3476 395
rect 3444 364 3476 365
rect 3444 284 3476 316
rect 3444 235 3476 236
rect 3444 205 3445 235
rect 3445 205 3475 235
rect 3475 205 3476 235
rect 3444 204 3476 205
rect 3444 124 3476 156
rect 3444 75 3476 76
rect 3444 45 3445 75
rect 3445 45 3475 75
rect 3475 45 3476 75
rect 3444 44 3476 45
rect 3444 -5 3476 -4
rect 3444 -35 3445 -5
rect 3445 -35 3475 -5
rect 3475 -35 3476 -5
rect 3444 -36 3476 -35
rect 3444 -85 3476 -84
rect 3444 -115 3445 -85
rect 3445 -115 3475 -85
rect 3475 -115 3476 -85
rect 3444 -116 3476 -115
rect 3444 -165 3476 -164
rect 3444 -195 3445 -165
rect 3445 -195 3475 -165
rect 3475 -195 3476 -165
rect 3444 -196 3476 -195
rect 3444 -245 3476 -244
rect 3444 -275 3445 -245
rect 3445 -275 3475 -245
rect 3475 -275 3476 -245
rect 3444 -276 3476 -275
rect 3444 -325 3476 -324
rect 3444 -355 3445 -325
rect 3445 -355 3475 -325
rect 3475 -355 3476 -325
rect 3444 -356 3476 -355
rect 3444 -436 3476 -404
rect 3444 -485 3476 -484
rect 3444 -515 3445 -485
rect 3445 -515 3475 -485
rect 3475 -515 3476 -485
rect 3444 -516 3476 -515
rect 3444 -596 3476 -564
rect 3444 -645 3476 -644
rect 3444 -675 3445 -645
rect 3445 -675 3475 -645
rect 3475 -675 3476 -645
rect 3444 -676 3476 -675
rect 3444 -756 3476 -724
rect 3444 -805 3476 -804
rect 3444 -835 3445 -805
rect 3445 -835 3475 -805
rect 3475 -835 3476 -805
rect 3444 -836 3476 -835
rect 3444 -885 3476 -884
rect 3444 -915 3445 -885
rect 3445 -915 3475 -885
rect 3475 -915 3476 -885
rect 3444 -916 3476 -915
rect 3444 -996 3476 -964
rect 3444 -1076 3476 -1044
rect 3444 -1125 3476 -1124
rect 3444 -1155 3445 -1125
rect 3445 -1155 3475 -1125
rect 3475 -1155 3476 -1125
rect 3444 -1156 3476 -1155
rect 3444 -1205 3476 -1204
rect 3444 -1235 3445 -1205
rect 3445 -1235 3475 -1205
rect 3475 -1235 3476 -1205
rect 3444 -1236 3476 -1235
rect 3444 -1285 3476 -1284
rect 3444 -1315 3445 -1285
rect 3445 -1315 3475 -1285
rect 3475 -1315 3476 -1285
rect 3444 -1316 3476 -1315
rect 3444 -1365 3476 -1364
rect 3444 -1395 3445 -1365
rect 3445 -1395 3475 -1365
rect 3475 -1395 3476 -1365
rect 3444 -1396 3476 -1395
rect 3444 -1445 3476 -1444
rect 3444 -1475 3445 -1445
rect 3445 -1475 3475 -1445
rect 3475 -1475 3476 -1445
rect 3444 -1476 3476 -1475
rect 3444 -1525 3476 -1524
rect 3444 -1555 3445 -1525
rect 3445 -1555 3475 -1525
rect 3475 -1555 3476 -1525
rect 3444 -1556 3476 -1555
rect 3444 -1636 3476 -1604
rect 3444 -1716 3476 -1684
rect 3444 -1765 3476 -1764
rect 3444 -1795 3445 -1765
rect 3445 -1795 3475 -1765
rect 3475 -1795 3476 -1765
rect 3444 -1796 3476 -1795
rect 3444 -1845 3476 -1844
rect 3444 -1875 3445 -1845
rect 3445 -1875 3475 -1845
rect 3475 -1875 3476 -1845
rect 3444 -1876 3476 -1875
rect 3444 -1956 3476 -1924
rect 3444 -2005 3476 -2004
rect 3444 -2035 3445 -2005
rect 3445 -2035 3475 -2005
rect 3475 -2035 3476 -2005
rect 3444 -2036 3476 -2035
rect 3444 -2116 3476 -2084
rect 3444 -2165 3476 -2164
rect 3444 -2195 3445 -2165
rect 3445 -2195 3475 -2165
rect 3475 -2195 3476 -2165
rect 3444 -2196 3476 -2195
rect 3444 -2276 3476 -2244
rect 3444 -2325 3476 -2324
rect 3444 -2355 3445 -2325
rect 3445 -2355 3475 -2325
rect 3475 -2355 3476 -2325
rect 3444 -2356 3476 -2355
rect 3444 -2405 3476 -2404
rect 3444 -2435 3445 -2405
rect 3445 -2435 3475 -2405
rect 3475 -2435 3476 -2405
rect 3444 -2436 3476 -2435
rect 3444 -2485 3476 -2484
rect 3444 -2515 3445 -2485
rect 3445 -2515 3475 -2485
rect 3475 -2515 3476 -2485
rect 3444 -2516 3476 -2515
rect 3444 -2565 3476 -2564
rect 3444 -2595 3445 -2565
rect 3445 -2595 3475 -2565
rect 3475 -2595 3476 -2565
rect 3444 -2596 3476 -2595
rect 3444 -2645 3476 -2644
rect 3444 -2675 3445 -2645
rect 3445 -2675 3475 -2645
rect 3475 -2675 3476 -2645
rect 3444 -2676 3476 -2675
rect 3444 -2725 3476 -2724
rect 3444 -2755 3445 -2725
rect 3445 -2755 3475 -2725
rect 3475 -2755 3476 -2725
rect 3444 -2756 3476 -2755
rect 3444 -2836 3476 -2804
rect 3444 -2885 3476 -2884
rect 3444 -2915 3445 -2885
rect 3445 -2915 3475 -2885
rect 3475 -2915 3476 -2885
rect 3444 -2916 3476 -2915
rect 3444 -2996 3476 -2964
rect 3444 -3045 3476 -3044
rect 3444 -3075 3445 -3045
rect 3445 -3075 3475 -3045
rect 3475 -3075 3476 -3045
rect 3444 -3076 3476 -3075
rect 3444 -3156 3476 -3124
rect 3444 -3205 3476 -3204
rect 3444 -3235 3445 -3205
rect 3445 -3235 3475 -3205
rect 3475 -3235 3476 -3205
rect 3444 -3236 3476 -3235
rect 3444 -3285 3476 -3284
rect 3444 -3315 3445 -3285
rect 3445 -3315 3475 -3285
rect 3475 -3315 3476 -3285
rect 3444 -3316 3476 -3315
rect 3444 -3396 3476 -3364
rect 3444 -3476 3476 -3444
rect 3444 -3525 3476 -3524
rect 3444 -3555 3445 -3525
rect 3445 -3555 3475 -3525
rect 3475 -3555 3476 -3525
rect 3444 -3556 3476 -3555
rect 3444 -3605 3476 -3604
rect 3444 -3635 3445 -3605
rect 3445 -3635 3475 -3605
rect 3475 -3635 3476 -3605
rect 3444 -3636 3476 -3635
rect 3444 -3685 3476 -3684
rect 3444 -3715 3445 -3685
rect 3445 -3715 3475 -3685
rect 3475 -3715 3476 -3685
rect 3444 -3716 3476 -3715
rect 3524 1035 3556 1036
rect 3524 1005 3525 1035
rect 3525 1005 3555 1035
rect 3555 1005 3556 1035
rect 3524 1004 3556 1005
rect 3524 955 3556 956
rect 3524 925 3525 955
rect 3525 925 3555 955
rect 3555 925 3556 955
rect 3524 924 3556 925
rect 3524 875 3556 876
rect 3524 845 3525 875
rect 3525 845 3555 875
rect 3555 845 3556 875
rect 3524 844 3556 845
rect 3524 764 3556 796
rect 3524 684 3556 716
rect 3524 635 3556 636
rect 3524 605 3525 635
rect 3525 605 3555 635
rect 3555 605 3556 635
rect 3524 604 3556 605
rect 3524 555 3556 556
rect 3524 525 3525 555
rect 3525 525 3555 555
rect 3555 525 3556 555
rect 3524 524 3556 525
rect 3524 444 3556 476
rect 3524 395 3556 396
rect 3524 365 3525 395
rect 3525 365 3555 395
rect 3555 365 3556 395
rect 3524 364 3556 365
rect 3524 284 3556 316
rect 3524 235 3556 236
rect 3524 205 3525 235
rect 3525 205 3555 235
rect 3555 205 3556 235
rect 3524 204 3556 205
rect 3524 124 3556 156
rect 3524 75 3556 76
rect 3524 45 3525 75
rect 3525 45 3555 75
rect 3555 45 3556 75
rect 3524 44 3556 45
rect 3524 -5 3556 -4
rect 3524 -35 3525 -5
rect 3525 -35 3555 -5
rect 3555 -35 3556 -5
rect 3524 -36 3556 -35
rect 3524 -85 3556 -84
rect 3524 -115 3525 -85
rect 3525 -115 3555 -85
rect 3555 -115 3556 -85
rect 3524 -116 3556 -115
rect 3524 -165 3556 -164
rect 3524 -195 3525 -165
rect 3525 -195 3555 -165
rect 3555 -195 3556 -165
rect 3524 -196 3556 -195
rect 3524 -245 3556 -244
rect 3524 -275 3525 -245
rect 3525 -275 3555 -245
rect 3555 -275 3556 -245
rect 3524 -276 3556 -275
rect 3524 -325 3556 -324
rect 3524 -355 3525 -325
rect 3525 -355 3555 -325
rect 3555 -355 3556 -325
rect 3524 -356 3556 -355
rect 3524 -436 3556 -404
rect 3524 -485 3556 -484
rect 3524 -515 3525 -485
rect 3525 -515 3555 -485
rect 3555 -515 3556 -485
rect 3524 -516 3556 -515
rect 3524 -596 3556 -564
rect 3524 -645 3556 -644
rect 3524 -675 3525 -645
rect 3525 -675 3555 -645
rect 3555 -675 3556 -645
rect 3524 -676 3556 -675
rect 3524 -756 3556 -724
rect 3524 -805 3556 -804
rect 3524 -835 3525 -805
rect 3525 -835 3555 -805
rect 3555 -835 3556 -805
rect 3524 -836 3556 -835
rect 3524 -885 3556 -884
rect 3524 -915 3525 -885
rect 3525 -915 3555 -885
rect 3555 -915 3556 -885
rect 3524 -916 3556 -915
rect 3524 -996 3556 -964
rect 3524 -1076 3556 -1044
rect 3524 -1125 3556 -1124
rect 3524 -1155 3525 -1125
rect 3525 -1155 3555 -1125
rect 3555 -1155 3556 -1125
rect 3524 -1156 3556 -1155
rect 3524 -1205 3556 -1204
rect 3524 -1235 3525 -1205
rect 3525 -1235 3555 -1205
rect 3555 -1235 3556 -1205
rect 3524 -1236 3556 -1235
rect 3524 -1285 3556 -1284
rect 3524 -1315 3525 -1285
rect 3525 -1315 3555 -1285
rect 3555 -1315 3556 -1285
rect 3524 -1316 3556 -1315
rect 3524 -1365 3556 -1364
rect 3524 -1395 3525 -1365
rect 3525 -1395 3555 -1365
rect 3555 -1395 3556 -1365
rect 3524 -1396 3556 -1395
rect 3524 -1445 3556 -1444
rect 3524 -1475 3525 -1445
rect 3525 -1475 3555 -1445
rect 3555 -1475 3556 -1445
rect 3524 -1476 3556 -1475
rect 3524 -1525 3556 -1524
rect 3524 -1555 3525 -1525
rect 3525 -1555 3555 -1525
rect 3555 -1555 3556 -1525
rect 3524 -1556 3556 -1555
rect 3524 -1636 3556 -1604
rect 3524 -1716 3556 -1684
rect 3524 -1765 3556 -1764
rect 3524 -1795 3525 -1765
rect 3525 -1795 3555 -1765
rect 3555 -1795 3556 -1765
rect 3524 -1796 3556 -1795
rect 3524 -1845 3556 -1844
rect 3524 -1875 3525 -1845
rect 3525 -1875 3555 -1845
rect 3555 -1875 3556 -1845
rect 3524 -1876 3556 -1875
rect 3524 -1956 3556 -1924
rect 3524 -2005 3556 -2004
rect 3524 -2035 3525 -2005
rect 3525 -2035 3555 -2005
rect 3555 -2035 3556 -2005
rect 3524 -2036 3556 -2035
rect 3524 -2116 3556 -2084
rect 3524 -2165 3556 -2164
rect 3524 -2195 3525 -2165
rect 3525 -2195 3555 -2165
rect 3555 -2195 3556 -2165
rect 3524 -2196 3556 -2195
rect 3524 -2276 3556 -2244
rect 3524 -2325 3556 -2324
rect 3524 -2355 3525 -2325
rect 3525 -2355 3555 -2325
rect 3555 -2355 3556 -2325
rect 3524 -2356 3556 -2355
rect 3524 -2405 3556 -2404
rect 3524 -2435 3525 -2405
rect 3525 -2435 3555 -2405
rect 3555 -2435 3556 -2405
rect 3524 -2436 3556 -2435
rect 3524 -2485 3556 -2484
rect 3524 -2515 3525 -2485
rect 3525 -2515 3555 -2485
rect 3555 -2515 3556 -2485
rect 3524 -2516 3556 -2515
rect 3524 -2565 3556 -2564
rect 3524 -2595 3525 -2565
rect 3525 -2595 3555 -2565
rect 3555 -2595 3556 -2565
rect 3524 -2596 3556 -2595
rect 3524 -2645 3556 -2644
rect 3524 -2675 3525 -2645
rect 3525 -2675 3555 -2645
rect 3555 -2675 3556 -2645
rect 3524 -2676 3556 -2675
rect 3524 -2725 3556 -2724
rect 3524 -2755 3525 -2725
rect 3525 -2755 3555 -2725
rect 3555 -2755 3556 -2725
rect 3524 -2756 3556 -2755
rect 3524 -2836 3556 -2804
rect 3524 -2885 3556 -2884
rect 3524 -2915 3525 -2885
rect 3525 -2915 3555 -2885
rect 3555 -2915 3556 -2885
rect 3524 -2916 3556 -2915
rect 3524 -2996 3556 -2964
rect 3524 -3045 3556 -3044
rect 3524 -3075 3525 -3045
rect 3525 -3075 3555 -3045
rect 3555 -3075 3556 -3045
rect 3524 -3076 3556 -3075
rect 3524 -3156 3556 -3124
rect 3524 -3205 3556 -3204
rect 3524 -3235 3525 -3205
rect 3525 -3235 3555 -3205
rect 3555 -3235 3556 -3205
rect 3524 -3236 3556 -3235
rect 3524 -3285 3556 -3284
rect 3524 -3315 3525 -3285
rect 3525 -3315 3555 -3285
rect 3555 -3315 3556 -3285
rect 3524 -3316 3556 -3315
rect 3524 -3396 3556 -3364
rect 3524 -3476 3556 -3444
rect 3524 -3525 3556 -3524
rect 3524 -3555 3525 -3525
rect 3525 -3555 3555 -3525
rect 3555 -3555 3556 -3525
rect 3524 -3556 3556 -3555
rect 3524 -3605 3556 -3604
rect 3524 -3635 3525 -3605
rect 3525 -3635 3555 -3605
rect 3555 -3635 3556 -3605
rect 3524 -3636 3556 -3635
rect 3524 -3685 3556 -3684
rect 3524 -3715 3525 -3685
rect 3525 -3715 3555 -3685
rect 3555 -3715 3556 -3685
rect 3524 -3716 3556 -3715
rect 3604 1035 3636 1036
rect 3604 1005 3605 1035
rect 3605 1005 3635 1035
rect 3635 1005 3636 1035
rect 3604 1004 3636 1005
rect 3604 955 3636 956
rect 3604 925 3605 955
rect 3605 925 3635 955
rect 3635 925 3636 955
rect 3604 924 3636 925
rect 3604 875 3636 876
rect 3604 845 3605 875
rect 3605 845 3635 875
rect 3635 845 3636 875
rect 3604 844 3636 845
rect 3604 764 3636 796
rect 3604 684 3636 716
rect 3604 635 3636 636
rect 3604 605 3605 635
rect 3605 605 3635 635
rect 3635 605 3636 635
rect 3604 604 3636 605
rect 3604 555 3636 556
rect 3604 525 3605 555
rect 3605 525 3635 555
rect 3635 525 3636 555
rect 3604 524 3636 525
rect 3604 444 3636 476
rect 3604 395 3636 396
rect 3604 365 3605 395
rect 3605 365 3635 395
rect 3635 365 3636 395
rect 3604 364 3636 365
rect 3604 284 3636 316
rect 3604 235 3636 236
rect 3604 205 3605 235
rect 3605 205 3635 235
rect 3635 205 3636 235
rect 3604 204 3636 205
rect 3604 124 3636 156
rect 3604 75 3636 76
rect 3604 45 3605 75
rect 3605 45 3635 75
rect 3635 45 3636 75
rect 3604 44 3636 45
rect 3604 -5 3636 -4
rect 3604 -35 3605 -5
rect 3605 -35 3635 -5
rect 3635 -35 3636 -5
rect 3604 -36 3636 -35
rect 3604 -85 3636 -84
rect 3604 -115 3605 -85
rect 3605 -115 3635 -85
rect 3635 -115 3636 -85
rect 3604 -116 3636 -115
rect 3604 -165 3636 -164
rect 3604 -195 3605 -165
rect 3605 -195 3635 -165
rect 3635 -195 3636 -165
rect 3604 -196 3636 -195
rect 3604 -245 3636 -244
rect 3604 -275 3605 -245
rect 3605 -275 3635 -245
rect 3635 -275 3636 -245
rect 3604 -276 3636 -275
rect 3604 -325 3636 -324
rect 3604 -355 3605 -325
rect 3605 -355 3635 -325
rect 3635 -355 3636 -325
rect 3604 -356 3636 -355
rect 3604 -436 3636 -404
rect 3604 -485 3636 -484
rect 3604 -515 3605 -485
rect 3605 -515 3635 -485
rect 3635 -515 3636 -485
rect 3604 -516 3636 -515
rect 3604 -596 3636 -564
rect 3604 -645 3636 -644
rect 3604 -675 3605 -645
rect 3605 -675 3635 -645
rect 3635 -675 3636 -645
rect 3604 -676 3636 -675
rect 3604 -756 3636 -724
rect 3604 -805 3636 -804
rect 3604 -835 3605 -805
rect 3605 -835 3635 -805
rect 3635 -835 3636 -805
rect 3604 -836 3636 -835
rect 3604 -885 3636 -884
rect 3604 -915 3605 -885
rect 3605 -915 3635 -885
rect 3635 -915 3636 -885
rect 3604 -916 3636 -915
rect 3604 -996 3636 -964
rect 3604 -1076 3636 -1044
rect 3604 -1125 3636 -1124
rect 3604 -1155 3605 -1125
rect 3605 -1155 3635 -1125
rect 3635 -1155 3636 -1125
rect 3604 -1156 3636 -1155
rect 3604 -1205 3636 -1204
rect 3604 -1235 3605 -1205
rect 3605 -1235 3635 -1205
rect 3635 -1235 3636 -1205
rect 3604 -1236 3636 -1235
rect 3604 -1285 3636 -1284
rect 3604 -1315 3605 -1285
rect 3605 -1315 3635 -1285
rect 3635 -1315 3636 -1285
rect 3604 -1316 3636 -1315
rect 3604 -1365 3636 -1364
rect 3604 -1395 3605 -1365
rect 3605 -1395 3635 -1365
rect 3635 -1395 3636 -1365
rect 3604 -1396 3636 -1395
rect 3604 -1445 3636 -1444
rect 3604 -1475 3605 -1445
rect 3605 -1475 3635 -1445
rect 3635 -1475 3636 -1445
rect 3604 -1476 3636 -1475
rect 3604 -1525 3636 -1524
rect 3604 -1555 3605 -1525
rect 3605 -1555 3635 -1525
rect 3635 -1555 3636 -1525
rect 3604 -1556 3636 -1555
rect 3604 -1636 3636 -1604
rect 3604 -1716 3636 -1684
rect 3604 -1765 3636 -1764
rect 3604 -1795 3605 -1765
rect 3605 -1795 3635 -1765
rect 3635 -1795 3636 -1765
rect 3604 -1796 3636 -1795
rect 3604 -1845 3636 -1844
rect 3604 -1875 3605 -1845
rect 3605 -1875 3635 -1845
rect 3635 -1875 3636 -1845
rect 3604 -1876 3636 -1875
rect 3604 -1956 3636 -1924
rect 3604 -2005 3636 -2004
rect 3604 -2035 3605 -2005
rect 3605 -2035 3635 -2005
rect 3635 -2035 3636 -2005
rect 3604 -2036 3636 -2035
rect 3604 -2116 3636 -2084
rect 3604 -2165 3636 -2164
rect 3604 -2195 3605 -2165
rect 3605 -2195 3635 -2165
rect 3635 -2195 3636 -2165
rect 3604 -2196 3636 -2195
rect 3604 -2276 3636 -2244
rect 3604 -2325 3636 -2324
rect 3604 -2355 3605 -2325
rect 3605 -2355 3635 -2325
rect 3635 -2355 3636 -2325
rect 3604 -2356 3636 -2355
rect 3604 -2405 3636 -2404
rect 3604 -2435 3605 -2405
rect 3605 -2435 3635 -2405
rect 3635 -2435 3636 -2405
rect 3604 -2436 3636 -2435
rect 3604 -2485 3636 -2484
rect 3604 -2515 3605 -2485
rect 3605 -2515 3635 -2485
rect 3635 -2515 3636 -2485
rect 3604 -2516 3636 -2515
rect 3604 -2565 3636 -2564
rect 3604 -2595 3605 -2565
rect 3605 -2595 3635 -2565
rect 3635 -2595 3636 -2565
rect 3604 -2596 3636 -2595
rect 3604 -2645 3636 -2644
rect 3604 -2675 3605 -2645
rect 3605 -2675 3635 -2645
rect 3635 -2675 3636 -2645
rect 3604 -2676 3636 -2675
rect 3604 -2725 3636 -2724
rect 3604 -2755 3605 -2725
rect 3605 -2755 3635 -2725
rect 3635 -2755 3636 -2725
rect 3604 -2756 3636 -2755
rect 3604 -2836 3636 -2804
rect 3604 -2885 3636 -2884
rect 3604 -2915 3605 -2885
rect 3605 -2915 3635 -2885
rect 3635 -2915 3636 -2885
rect 3604 -2916 3636 -2915
rect 3604 -2996 3636 -2964
rect 3604 -3045 3636 -3044
rect 3604 -3075 3605 -3045
rect 3605 -3075 3635 -3045
rect 3635 -3075 3636 -3045
rect 3604 -3076 3636 -3075
rect 3604 -3156 3636 -3124
rect 3604 -3205 3636 -3204
rect 3604 -3235 3605 -3205
rect 3605 -3235 3635 -3205
rect 3635 -3235 3636 -3205
rect 3604 -3236 3636 -3235
rect 3604 -3285 3636 -3284
rect 3604 -3315 3605 -3285
rect 3605 -3315 3635 -3285
rect 3635 -3315 3636 -3285
rect 3604 -3316 3636 -3315
rect 3604 -3396 3636 -3364
rect 3604 -3476 3636 -3444
rect 3604 -3525 3636 -3524
rect 3604 -3555 3605 -3525
rect 3605 -3555 3635 -3525
rect 3635 -3555 3636 -3525
rect 3604 -3556 3636 -3555
rect 3604 -3605 3636 -3604
rect 3604 -3635 3605 -3605
rect 3605 -3635 3635 -3605
rect 3635 -3635 3636 -3605
rect 3604 -3636 3636 -3635
rect 3604 -3685 3636 -3684
rect 3604 -3715 3605 -3685
rect 3605 -3715 3635 -3685
rect 3635 -3715 3636 -3685
rect 3604 -3716 3636 -3715
rect 3684 1035 3716 1036
rect 3684 1005 3685 1035
rect 3685 1005 3715 1035
rect 3715 1005 3716 1035
rect 3684 1004 3716 1005
rect 3684 955 3716 956
rect 3684 925 3685 955
rect 3685 925 3715 955
rect 3715 925 3716 955
rect 3684 924 3716 925
rect 3684 875 3716 876
rect 3684 845 3685 875
rect 3685 845 3715 875
rect 3715 845 3716 875
rect 3684 844 3716 845
rect 3684 764 3716 796
rect 3684 684 3716 716
rect 3684 635 3716 636
rect 3684 605 3685 635
rect 3685 605 3715 635
rect 3715 605 3716 635
rect 3684 604 3716 605
rect 3684 555 3716 556
rect 3684 525 3685 555
rect 3685 525 3715 555
rect 3715 525 3716 555
rect 3684 524 3716 525
rect 3684 444 3716 476
rect 3684 395 3716 396
rect 3684 365 3685 395
rect 3685 365 3715 395
rect 3715 365 3716 395
rect 3684 364 3716 365
rect 3684 284 3716 316
rect 3684 235 3716 236
rect 3684 205 3685 235
rect 3685 205 3715 235
rect 3715 205 3716 235
rect 3684 204 3716 205
rect 3684 124 3716 156
rect 3684 75 3716 76
rect 3684 45 3685 75
rect 3685 45 3715 75
rect 3715 45 3716 75
rect 3684 44 3716 45
rect 3684 -5 3716 -4
rect 3684 -35 3685 -5
rect 3685 -35 3715 -5
rect 3715 -35 3716 -5
rect 3684 -36 3716 -35
rect 3684 -85 3716 -84
rect 3684 -115 3685 -85
rect 3685 -115 3715 -85
rect 3715 -115 3716 -85
rect 3684 -116 3716 -115
rect 3684 -165 3716 -164
rect 3684 -195 3685 -165
rect 3685 -195 3715 -165
rect 3715 -195 3716 -165
rect 3684 -196 3716 -195
rect 3684 -245 3716 -244
rect 3684 -275 3685 -245
rect 3685 -275 3715 -245
rect 3715 -275 3716 -245
rect 3684 -276 3716 -275
rect 3684 -325 3716 -324
rect 3684 -355 3685 -325
rect 3685 -355 3715 -325
rect 3715 -355 3716 -325
rect 3684 -356 3716 -355
rect 3684 -436 3716 -404
rect 3684 -485 3716 -484
rect 3684 -515 3685 -485
rect 3685 -515 3715 -485
rect 3715 -515 3716 -485
rect 3684 -516 3716 -515
rect 3684 -596 3716 -564
rect 3684 -645 3716 -644
rect 3684 -675 3685 -645
rect 3685 -675 3715 -645
rect 3715 -675 3716 -645
rect 3684 -676 3716 -675
rect 3684 -756 3716 -724
rect 3684 -805 3716 -804
rect 3684 -835 3685 -805
rect 3685 -835 3715 -805
rect 3715 -835 3716 -805
rect 3684 -836 3716 -835
rect 3684 -885 3716 -884
rect 3684 -915 3685 -885
rect 3685 -915 3715 -885
rect 3715 -915 3716 -885
rect 3684 -916 3716 -915
rect 3684 -996 3716 -964
rect 3684 -1076 3716 -1044
rect 3684 -1125 3716 -1124
rect 3684 -1155 3685 -1125
rect 3685 -1155 3715 -1125
rect 3715 -1155 3716 -1125
rect 3684 -1156 3716 -1155
rect 3684 -1205 3716 -1204
rect 3684 -1235 3685 -1205
rect 3685 -1235 3715 -1205
rect 3715 -1235 3716 -1205
rect 3684 -1236 3716 -1235
rect 3684 -1285 3716 -1284
rect 3684 -1315 3685 -1285
rect 3685 -1315 3715 -1285
rect 3715 -1315 3716 -1285
rect 3684 -1316 3716 -1315
rect 3684 -1365 3716 -1364
rect 3684 -1395 3685 -1365
rect 3685 -1395 3715 -1365
rect 3715 -1395 3716 -1365
rect 3684 -1396 3716 -1395
rect 3684 -1445 3716 -1444
rect 3684 -1475 3685 -1445
rect 3685 -1475 3715 -1445
rect 3715 -1475 3716 -1445
rect 3684 -1476 3716 -1475
rect 3684 -1525 3716 -1524
rect 3684 -1555 3685 -1525
rect 3685 -1555 3715 -1525
rect 3715 -1555 3716 -1525
rect 3684 -1556 3716 -1555
rect 3684 -1636 3716 -1604
rect 3684 -1716 3716 -1684
rect 3684 -1765 3716 -1764
rect 3684 -1795 3685 -1765
rect 3685 -1795 3715 -1765
rect 3715 -1795 3716 -1765
rect 3684 -1796 3716 -1795
rect 3684 -1845 3716 -1844
rect 3684 -1875 3685 -1845
rect 3685 -1875 3715 -1845
rect 3715 -1875 3716 -1845
rect 3684 -1876 3716 -1875
rect 3684 -1956 3716 -1924
rect 3684 -2005 3716 -2004
rect 3684 -2035 3685 -2005
rect 3685 -2035 3715 -2005
rect 3715 -2035 3716 -2005
rect 3684 -2036 3716 -2035
rect 3684 -2116 3716 -2084
rect 3684 -2165 3716 -2164
rect 3684 -2195 3685 -2165
rect 3685 -2195 3715 -2165
rect 3715 -2195 3716 -2165
rect 3684 -2196 3716 -2195
rect 3684 -2276 3716 -2244
rect 3684 -2325 3716 -2324
rect 3684 -2355 3685 -2325
rect 3685 -2355 3715 -2325
rect 3715 -2355 3716 -2325
rect 3684 -2356 3716 -2355
rect 3684 -2405 3716 -2404
rect 3684 -2435 3685 -2405
rect 3685 -2435 3715 -2405
rect 3715 -2435 3716 -2405
rect 3684 -2436 3716 -2435
rect 3684 -2485 3716 -2484
rect 3684 -2515 3685 -2485
rect 3685 -2515 3715 -2485
rect 3715 -2515 3716 -2485
rect 3684 -2516 3716 -2515
rect 3684 -2565 3716 -2564
rect 3684 -2595 3685 -2565
rect 3685 -2595 3715 -2565
rect 3715 -2595 3716 -2565
rect 3684 -2596 3716 -2595
rect 3684 -2645 3716 -2644
rect 3684 -2675 3685 -2645
rect 3685 -2675 3715 -2645
rect 3715 -2675 3716 -2645
rect 3684 -2676 3716 -2675
rect 3684 -2725 3716 -2724
rect 3684 -2755 3685 -2725
rect 3685 -2755 3715 -2725
rect 3715 -2755 3716 -2725
rect 3684 -2756 3716 -2755
rect 3684 -2836 3716 -2804
rect 3684 -2885 3716 -2884
rect 3684 -2915 3685 -2885
rect 3685 -2915 3715 -2885
rect 3715 -2915 3716 -2885
rect 3684 -2916 3716 -2915
rect 3684 -2996 3716 -2964
rect 3684 -3045 3716 -3044
rect 3684 -3075 3685 -3045
rect 3685 -3075 3715 -3045
rect 3715 -3075 3716 -3045
rect 3684 -3076 3716 -3075
rect 3684 -3156 3716 -3124
rect 3684 -3205 3716 -3204
rect 3684 -3235 3685 -3205
rect 3685 -3235 3715 -3205
rect 3715 -3235 3716 -3205
rect 3684 -3236 3716 -3235
rect 3684 -3285 3716 -3284
rect 3684 -3315 3685 -3285
rect 3685 -3315 3715 -3285
rect 3715 -3315 3716 -3285
rect 3684 -3316 3716 -3315
rect 3684 -3396 3716 -3364
rect 3684 -3476 3716 -3444
rect 3684 -3525 3716 -3524
rect 3684 -3555 3685 -3525
rect 3685 -3555 3715 -3525
rect 3715 -3555 3716 -3525
rect 3684 -3556 3716 -3555
rect 3684 -3605 3716 -3604
rect 3684 -3635 3685 -3605
rect 3685 -3635 3715 -3605
rect 3715 -3635 3716 -3605
rect 3684 -3636 3716 -3635
rect 3684 -3685 3716 -3684
rect 3684 -3715 3685 -3685
rect 3685 -3715 3715 -3685
rect 3715 -3715 3716 -3685
rect 3684 -3716 3716 -3715
rect 3764 1035 3796 1036
rect 3764 1005 3765 1035
rect 3765 1005 3795 1035
rect 3795 1005 3796 1035
rect 3764 1004 3796 1005
rect 3764 955 3796 956
rect 3764 925 3765 955
rect 3765 925 3795 955
rect 3795 925 3796 955
rect 3764 924 3796 925
rect 3764 875 3796 876
rect 3764 845 3765 875
rect 3765 845 3795 875
rect 3795 845 3796 875
rect 3764 844 3796 845
rect 3764 764 3796 796
rect 3764 684 3796 716
rect 3764 635 3796 636
rect 3764 605 3765 635
rect 3765 605 3795 635
rect 3795 605 3796 635
rect 3764 604 3796 605
rect 3764 555 3796 556
rect 3764 525 3765 555
rect 3765 525 3795 555
rect 3795 525 3796 555
rect 3764 524 3796 525
rect 3764 444 3796 476
rect 3764 395 3796 396
rect 3764 365 3765 395
rect 3765 365 3795 395
rect 3795 365 3796 395
rect 3764 364 3796 365
rect 3764 284 3796 316
rect 3764 235 3796 236
rect 3764 205 3765 235
rect 3765 205 3795 235
rect 3795 205 3796 235
rect 3764 204 3796 205
rect 3764 124 3796 156
rect 3764 75 3796 76
rect 3764 45 3765 75
rect 3765 45 3795 75
rect 3795 45 3796 75
rect 3764 44 3796 45
rect 3764 -5 3796 -4
rect 3764 -35 3765 -5
rect 3765 -35 3795 -5
rect 3795 -35 3796 -5
rect 3764 -36 3796 -35
rect 3764 -85 3796 -84
rect 3764 -115 3765 -85
rect 3765 -115 3795 -85
rect 3795 -115 3796 -85
rect 3764 -116 3796 -115
rect 3764 -165 3796 -164
rect 3764 -195 3765 -165
rect 3765 -195 3795 -165
rect 3795 -195 3796 -165
rect 3764 -196 3796 -195
rect 3764 -245 3796 -244
rect 3764 -275 3765 -245
rect 3765 -275 3795 -245
rect 3795 -275 3796 -245
rect 3764 -276 3796 -275
rect 3764 -325 3796 -324
rect 3764 -355 3765 -325
rect 3765 -355 3795 -325
rect 3795 -355 3796 -325
rect 3764 -356 3796 -355
rect 3764 -436 3796 -404
rect 3764 -485 3796 -484
rect 3764 -515 3765 -485
rect 3765 -515 3795 -485
rect 3795 -515 3796 -485
rect 3764 -516 3796 -515
rect 3764 -596 3796 -564
rect 3764 -645 3796 -644
rect 3764 -675 3765 -645
rect 3765 -675 3795 -645
rect 3795 -675 3796 -645
rect 3764 -676 3796 -675
rect 3764 -756 3796 -724
rect 3764 -805 3796 -804
rect 3764 -835 3765 -805
rect 3765 -835 3795 -805
rect 3795 -835 3796 -805
rect 3764 -836 3796 -835
rect 3764 -885 3796 -884
rect 3764 -915 3765 -885
rect 3765 -915 3795 -885
rect 3795 -915 3796 -885
rect 3764 -916 3796 -915
rect 3764 -996 3796 -964
rect 3764 -1076 3796 -1044
rect 3764 -1125 3796 -1124
rect 3764 -1155 3765 -1125
rect 3765 -1155 3795 -1125
rect 3795 -1155 3796 -1125
rect 3764 -1156 3796 -1155
rect 3764 -1205 3796 -1204
rect 3764 -1235 3765 -1205
rect 3765 -1235 3795 -1205
rect 3795 -1235 3796 -1205
rect 3764 -1236 3796 -1235
rect 3764 -1285 3796 -1284
rect 3764 -1315 3765 -1285
rect 3765 -1315 3795 -1285
rect 3795 -1315 3796 -1285
rect 3764 -1316 3796 -1315
rect 3764 -1365 3796 -1364
rect 3764 -1395 3765 -1365
rect 3765 -1395 3795 -1365
rect 3795 -1395 3796 -1365
rect 3764 -1396 3796 -1395
rect 3764 -1445 3796 -1444
rect 3764 -1475 3765 -1445
rect 3765 -1475 3795 -1445
rect 3795 -1475 3796 -1445
rect 3764 -1476 3796 -1475
rect 3764 -1525 3796 -1524
rect 3764 -1555 3765 -1525
rect 3765 -1555 3795 -1525
rect 3795 -1555 3796 -1525
rect 3764 -1556 3796 -1555
rect 3764 -1636 3796 -1604
rect 3764 -1716 3796 -1684
rect 3764 -1765 3796 -1764
rect 3764 -1795 3765 -1765
rect 3765 -1795 3795 -1765
rect 3795 -1795 3796 -1765
rect 3764 -1796 3796 -1795
rect 3764 -1845 3796 -1844
rect 3764 -1875 3765 -1845
rect 3765 -1875 3795 -1845
rect 3795 -1875 3796 -1845
rect 3764 -1876 3796 -1875
rect 3764 -1956 3796 -1924
rect 3764 -2005 3796 -2004
rect 3764 -2035 3765 -2005
rect 3765 -2035 3795 -2005
rect 3795 -2035 3796 -2005
rect 3764 -2036 3796 -2035
rect 3764 -2116 3796 -2084
rect 3764 -2165 3796 -2164
rect 3764 -2195 3765 -2165
rect 3765 -2195 3795 -2165
rect 3795 -2195 3796 -2165
rect 3764 -2196 3796 -2195
rect 3764 -2276 3796 -2244
rect 3764 -2325 3796 -2324
rect 3764 -2355 3765 -2325
rect 3765 -2355 3795 -2325
rect 3795 -2355 3796 -2325
rect 3764 -2356 3796 -2355
rect 3764 -2405 3796 -2404
rect 3764 -2435 3765 -2405
rect 3765 -2435 3795 -2405
rect 3795 -2435 3796 -2405
rect 3764 -2436 3796 -2435
rect 3764 -2485 3796 -2484
rect 3764 -2515 3765 -2485
rect 3765 -2515 3795 -2485
rect 3795 -2515 3796 -2485
rect 3764 -2516 3796 -2515
rect 3764 -2565 3796 -2564
rect 3764 -2595 3765 -2565
rect 3765 -2595 3795 -2565
rect 3795 -2595 3796 -2565
rect 3764 -2596 3796 -2595
rect 3764 -2645 3796 -2644
rect 3764 -2675 3765 -2645
rect 3765 -2675 3795 -2645
rect 3795 -2675 3796 -2645
rect 3764 -2676 3796 -2675
rect 3764 -2725 3796 -2724
rect 3764 -2755 3765 -2725
rect 3765 -2755 3795 -2725
rect 3795 -2755 3796 -2725
rect 3764 -2756 3796 -2755
rect 3764 -2836 3796 -2804
rect 3764 -2885 3796 -2884
rect 3764 -2915 3765 -2885
rect 3765 -2915 3795 -2885
rect 3795 -2915 3796 -2885
rect 3764 -2916 3796 -2915
rect 3764 -2996 3796 -2964
rect 3764 -3045 3796 -3044
rect 3764 -3075 3765 -3045
rect 3765 -3075 3795 -3045
rect 3795 -3075 3796 -3045
rect 3764 -3076 3796 -3075
rect 3764 -3156 3796 -3124
rect 3764 -3205 3796 -3204
rect 3764 -3235 3765 -3205
rect 3765 -3235 3795 -3205
rect 3795 -3235 3796 -3205
rect 3764 -3236 3796 -3235
rect 3764 -3285 3796 -3284
rect 3764 -3315 3765 -3285
rect 3765 -3315 3795 -3285
rect 3795 -3315 3796 -3285
rect 3764 -3316 3796 -3315
rect 3764 -3396 3796 -3364
rect 3764 -3476 3796 -3444
rect 3764 -3525 3796 -3524
rect 3764 -3555 3765 -3525
rect 3765 -3555 3795 -3525
rect 3795 -3555 3796 -3525
rect 3764 -3556 3796 -3555
rect 3764 -3605 3796 -3604
rect 3764 -3635 3765 -3605
rect 3765 -3635 3795 -3605
rect 3795 -3635 3796 -3605
rect 3764 -3636 3796 -3635
rect 3764 -3685 3796 -3684
rect 3764 -3715 3765 -3685
rect 3765 -3715 3795 -3685
rect 3795 -3715 3796 -3685
rect 3764 -3716 3796 -3715
rect 3844 1035 3876 1036
rect 3844 1005 3845 1035
rect 3845 1005 3875 1035
rect 3875 1005 3876 1035
rect 3844 1004 3876 1005
rect 3844 955 3876 956
rect 3844 925 3845 955
rect 3845 925 3875 955
rect 3875 925 3876 955
rect 3844 924 3876 925
rect 3844 875 3876 876
rect 3844 845 3845 875
rect 3845 845 3875 875
rect 3875 845 3876 875
rect 3844 844 3876 845
rect 3844 764 3876 796
rect 3844 684 3876 716
rect 3844 635 3876 636
rect 3844 605 3845 635
rect 3845 605 3875 635
rect 3875 605 3876 635
rect 3844 604 3876 605
rect 3844 555 3876 556
rect 3844 525 3845 555
rect 3845 525 3875 555
rect 3875 525 3876 555
rect 3844 524 3876 525
rect 3844 444 3876 476
rect 3844 395 3876 396
rect 3844 365 3845 395
rect 3845 365 3875 395
rect 3875 365 3876 395
rect 3844 364 3876 365
rect 3844 284 3876 316
rect 3844 235 3876 236
rect 3844 205 3845 235
rect 3845 205 3875 235
rect 3875 205 3876 235
rect 3844 204 3876 205
rect 3844 124 3876 156
rect 3844 75 3876 76
rect 3844 45 3845 75
rect 3845 45 3875 75
rect 3875 45 3876 75
rect 3844 44 3876 45
rect 3844 -5 3876 -4
rect 3844 -35 3845 -5
rect 3845 -35 3875 -5
rect 3875 -35 3876 -5
rect 3844 -36 3876 -35
rect 3844 -85 3876 -84
rect 3844 -115 3845 -85
rect 3845 -115 3875 -85
rect 3875 -115 3876 -85
rect 3844 -116 3876 -115
rect 3844 -165 3876 -164
rect 3844 -195 3845 -165
rect 3845 -195 3875 -165
rect 3875 -195 3876 -165
rect 3844 -196 3876 -195
rect 3844 -245 3876 -244
rect 3844 -275 3845 -245
rect 3845 -275 3875 -245
rect 3875 -275 3876 -245
rect 3844 -276 3876 -275
rect 3844 -325 3876 -324
rect 3844 -355 3845 -325
rect 3845 -355 3875 -325
rect 3875 -355 3876 -325
rect 3844 -356 3876 -355
rect 3844 -436 3876 -404
rect 3844 -485 3876 -484
rect 3844 -515 3845 -485
rect 3845 -515 3875 -485
rect 3875 -515 3876 -485
rect 3844 -516 3876 -515
rect 3844 -596 3876 -564
rect 3844 -645 3876 -644
rect 3844 -675 3845 -645
rect 3845 -675 3875 -645
rect 3875 -675 3876 -645
rect 3844 -676 3876 -675
rect 3844 -756 3876 -724
rect 3844 -805 3876 -804
rect 3844 -835 3845 -805
rect 3845 -835 3875 -805
rect 3875 -835 3876 -805
rect 3844 -836 3876 -835
rect 3844 -885 3876 -884
rect 3844 -915 3845 -885
rect 3845 -915 3875 -885
rect 3875 -915 3876 -885
rect 3844 -916 3876 -915
rect 3844 -996 3876 -964
rect 3844 -1076 3876 -1044
rect 3844 -1125 3876 -1124
rect 3844 -1155 3845 -1125
rect 3845 -1155 3875 -1125
rect 3875 -1155 3876 -1125
rect 3844 -1156 3876 -1155
rect 3844 -1205 3876 -1204
rect 3844 -1235 3845 -1205
rect 3845 -1235 3875 -1205
rect 3875 -1235 3876 -1205
rect 3844 -1236 3876 -1235
rect 3844 -1285 3876 -1284
rect 3844 -1315 3845 -1285
rect 3845 -1315 3875 -1285
rect 3875 -1315 3876 -1285
rect 3844 -1316 3876 -1315
rect 3844 -1365 3876 -1364
rect 3844 -1395 3845 -1365
rect 3845 -1395 3875 -1365
rect 3875 -1395 3876 -1365
rect 3844 -1396 3876 -1395
rect 3844 -1445 3876 -1444
rect 3844 -1475 3845 -1445
rect 3845 -1475 3875 -1445
rect 3875 -1475 3876 -1445
rect 3844 -1476 3876 -1475
rect 3844 -1525 3876 -1524
rect 3844 -1555 3845 -1525
rect 3845 -1555 3875 -1525
rect 3875 -1555 3876 -1525
rect 3844 -1556 3876 -1555
rect 3844 -1636 3876 -1604
rect 3844 -1716 3876 -1684
rect 3844 -1765 3876 -1764
rect 3844 -1795 3845 -1765
rect 3845 -1795 3875 -1765
rect 3875 -1795 3876 -1765
rect 3844 -1796 3876 -1795
rect 3844 -1845 3876 -1844
rect 3844 -1875 3845 -1845
rect 3845 -1875 3875 -1845
rect 3875 -1875 3876 -1845
rect 3844 -1876 3876 -1875
rect 3844 -1956 3876 -1924
rect 3844 -2005 3876 -2004
rect 3844 -2035 3845 -2005
rect 3845 -2035 3875 -2005
rect 3875 -2035 3876 -2005
rect 3844 -2036 3876 -2035
rect 3844 -2116 3876 -2084
rect 3844 -2165 3876 -2164
rect 3844 -2195 3845 -2165
rect 3845 -2195 3875 -2165
rect 3875 -2195 3876 -2165
rect 3844 -2196 3876 -2195
rect 3844 -2276 3876 -2244
rect 3844 -2325 3876 -2324
rect 3844 -2355 3845 -2325
rect 3845 -2355 3875 -2325
rect 3875 -2355 3876 -2325
rect 3844 -2356 3876 -2355
rect 3844 -2405 3876 -2404
rect 3844 -2435 3845 -2405
rect 3845 -2435 3875 -2405
rect 3875 -2435 3876 -2405
rect 3844 -2436 3876 -2435
rect 3844 -2485 3876 -2484
rect 3844 -2515 3845 -2485
rect 3845 -2515 3875 -2485
rect 3875 -2515 3876 -2485
rect 3844 -2516 3876 -2515
rect 3844 -2565 3876 -2564
rect 3844 -2595 3845 -2565
rect 3845 -2595 3875 -2565
rect 3875 -2595 3876 -2565
rect 3844 -2596 3876 -2595
rect 3844 -2645 3876 -2644
rect 3844 -2675 3845 -2645
rect 3845 -2675 3875 -2645
rect 3875 -2675 3876 -2645
rect 3844 -2676 3876 -2675
rect 3844 -2725 3876 -2724
rect 3844 -2755 3845 -2725
rect 3845 -2755 3875 -2725
rect 3875 -2755 3876 -2725
rect 3844 -2756 3876 -2755
rect 3844 -2836 3876 -2804
rect 3844 -2885 3876 -2884
rect 3844 -2915 3845 -2885
rect 3845 -2915 3875 -2885
rect 3875 -2915 3876 -2885
rect 3844 -2916 3876 -2915
rect 3844 -2996 3876 -2964
rect 3844 -3045 3876 -3044
rect 3844 -3075 3845 -3045
rect 3845 -3075 3875 -3045
rect 3875 -3075 3876 -3045
rect 3844 -3076 3876 -3075
rect 3844 -3156 3876 -3124
rect 3844 -3205 3876 -3204
rect 3844 -3235 3845 -3205
rect 3845 -3235 3875 -3205
rect 3875 -3235 3876 -3205
rect 3844 -3236 3876 -3235
rect 3844 -3285 3876 -3284
rect 3844 -3315 3845 -3285
rect 3845 -3315 3875 -3285
rect 3875 -3315 3876 -3285
rect 3844 -3316 3876 -3315
rect 3844 -3396 3876 -3364
rect 3844 -3476 3876 -3444
rect 3844 -3525 3876 -3524
rect 3844 -3555 3845 -3525
rect 3845 -3555 3875 -3525
rect 3875 -3555 3876 -3525
rect 3844 -3556 3876 -3555
rect 3844 -3605 3876 -3604
rect 3844 -3635 3845 -3605
rect 3845 -3635 3875 -3605
rect 3875 -3635 3876 -3605
rect 3844 -3636 3876 -3635
rect 3844 -3685 3876 -3684
rect 3844 -3715 3845 -3685
rect 3845 -3715 3875 -3685
rect 3875 -3715 3876 -3685
rect 3844 -3716 3876 -3715
rect 3924 1035 3956 1036
rect 3924 1005 3925 1035
rect 3925 1005 3955 1035
rect 3955 1005 3956 1035
rect 3924 1004 3956 1005
rect 3924 955 3956 956
rect 3924 925 3925 955
rect 3925 925 3955 955
rect 3955 925 3956 955
rect 3924 924 3956 925
rect 3924 875 3956 876
rect 3924 845 3925 875
rect 3925 845 3955 875
rect 3955 845 3956 875
rect 3924 844 3956 845
rect 3924 764 3956 796
rect 3924 684 3956 716
rect 3924 635 3956 636
rect 3924 605 3925 635
rect 3925 605 3955 635
rect 3955 605 3956 635
rect 3924 604 3956 605
rect 3924 555 3956 556
rect 3924 525 3925 555
rect 3925 525 3955 555
rect 3955 525 3956 555
rect 3924 524 3956 525
rect 3924 444 3956 476
rect 3924 395 3956 396
rect 3924 365 3925 395
rect 3925 365 3955 395
rect 3955 365 3956 395
rect 3924 364 3956 365
rect 3924 284 3956 316
rect 3924 235 3956 236
rect 3924 205 3925 235
rect 3925 205 3955 235
rect 3955 205 3956 235
rect 3924 204 3956 205
rect 3924 124 3956 156
rect 3924 75 3956 76
rect 3924 45 3925 75
rect 3925 45 3955 75
rect 3955 45 3956 75
rect 3924 44 3956 45
rect 3924 -5 3956 -4
rect 3924 -35 3925 -5
rect 3925 -35 3955 -5
rect 3955 -35 3956 -5
rect 3924 -36 3956 -35
rect 3924 -85 3956 -84
rect 3924 -115 3925 -85
rect 3925 -115 3955 -85
rect 3955 -115 3956 -85
rect 3924 -116 3956 -115
rect 3924 -165 3956 -164
rect 3924 -195 3925 -165
rect 3925 -195 3955 -165
rect 3955 -195 3956 -165
rect 3924 -196 3956 -195
rect 3924 -245 3956 -244
rect 3924 -275 3925 -245
rect 3925 -275 3955 -245
rect 3955 -275 3956 -245
rect 3924 -276 3956 -275
rect 3924 -325 3956 -324
rect 3924 -355 3925 -325
rect 3925 -355 3955 -325
rect 3955 -355 3956 -325
rect 3924 -356 3956 -355
rect 3924 -436 3956 -404
rect 3924 -485 3956 -484
rect 3924 -515 3925 -485
rect 3925 -515 3955 -485
rect 3955 -515 3956 -485
rect 3924 -516 3956 -515
rect 3924 -596 3956 -564
rect 3924 -645 3956 -644
rect 3924 -675 3925 -645
rect 3925 -675 3955 -645
rect 3955 -675 3956 -645
rect 3924 -676 3956 -675
rect 3924 -756 3956 -724
rect 3924 -805 3956 -804
rect 3924 -835 3925 -805
rect 3925 -835 3955 -805
rect 3955 -835 3956 -805
rect 3924 -836 3956 -835
rect 3924 -885 3956 -884
rect 3924 -915 3925 -885
rect 3925 -915 3955 -885
rect 3955 -915 3956 -885
rect 3924 -916 3956 -915
rect 3924 -996 3956 -964
rect 3924 -1076 3956 -1044
rect 3924 -1125 3956 -1124
rect 3924 -1155 3925 -1125
rect 3925 -1155 3955 -1125
rect 3955 -1155 3956 -1125
rect 3924 -1156 3956 -1155
rect 3924 -1205 3956 -1204
rect 3924 -1235 3925 -1205
rect 3925 -1235 3955 -1205
rect 3955 -1235 3956 -1205
rect 3924 -1236 3956 -1235
rect 3924 -1285 3956 -1284
rect 3924 -1315 3925 -1285
rect 3925 -1315 3955 -1285
rect 3955 -1315 3956 -1285
rect 3924 -1316 3956 -1315
rect 3924 -1365 3956 -1364
rect 3924 -1395 3925 -1365
rect 3925 -1395 3955 -1365
rect 3955 -1395 3956 -1365
rect 3924 -1396 3956 -1395
rect 3924 -1445 3956 -1444
rect 3924 -1475 3925 -1445
rect 3925 -1475 3955 -1445
rect 3955 -1475 3956 -1445
rect 3924 -1476 3956 -1475
rect 3924 -1525 3956 -1524
rect 3924 -1555 3925 -1525
rect 3925 -1555 3955 -1525
rect 3955 -1555 3956 -1525
rect 3924 -1556 3956 -1555
rect 3924 -1636 3956 -1604
rect 3924 -1716 3956 -1684
rect 3924 -1765 3956 -1764
rect 3924 -1795 3925 -1765
rect 3925 -1795 3955 -1765
rect 3955 -1795 3956 -1765
rect 3924 -1796 3956 -1795
rect 3924 -1845 3956 -1844
rect 3924 -1875 3925 -1845
rect 3925 -1875 3955 -1845
rect 3955 -1875 3956 -1845
rect 3924 -1876 3956 -1875
rect 3924 -1956 3956 -1924
rect 3924 -2005 3956 -2004
rect 3924 -2035 3925 -2005
rect 3925 -2035 3955 -2005
rect 3955 -2035 3956 -2005
rect 3924 -2036 3956 -2035
rect 3924 -2116 3956 -2084
rect 3924 -2165 3956 -2164
rect 3924 -2195 3925 -2165
rect 3925 -2195 3955 -2165
rect 3955 -2195 3956 -2165
rect 3924 -2196 3956 -2195
rect 3924 -2276 3956 -2244
rect 3924 -2325 3956 -2324
rect 3924 -2355 3925 -2325
rect 3925 -2355 3955 -2325
rect 3955 -2355 3956 -2325
rect 3924 -2356 3956 -2355
rect 3924 -2405 3956 -2404
rect 3924 -2435 3925 -2405
rect 3925 -2435 3955 -2405
rect 3955 -2435 3956 -2405
rect 3924 -2436 3956 -2435
rect 3924 -2485 3956 -2484
rect 3924 -2515 3925 -2485
rect 3925 -2515 3955 -2485
rect 3955 -2515 3956 -2485
rect 3924 -2516 3956 -2515
rect 3924 -2565 3956 -2564
rect 3924 -2595 3925 -2565
rect 3925 -2595 3955 -2565
rect 3955 -2595 3956 -2565
rect 3924 -2596 3956 -2595
rect 3924 -2645 3956 -2644
rect 3924 -2675 3925 -2645
rect 3925 -2675 3955 -2645
rect 3955 -2675 3956 -2645
rect 3924 -2676 3956 -2675
rect 3924 -2725 3956 -2724
rect 3924 -2755 3925 -2725
rect 3925 -2755 3955 -2725
rect 3955 -2755 3956 -2725
rect 3924 -2756 3956 -2755
rect 3924 -2836 3956 -2804
rect 3924 -2885 3956 -2884
rect 3924 -2915 3925 -2885
rect 3925 -2915 3955 -2885
rect 3955 -2915 3956 -2885
rect 3924 -2916 3956 -2915
rect 3924 -2996 3956 -2964
rect 3924 -3045 3956 -3044
rect 3924 -3075 3925 -3045
rect 3925 -3075 3955 -3045
rect 3955 -3075 3956 -3045
rect 3924 -3076 3956 -3075
rect 3924 -3156 3956 -3124
rect 3924 -3205 3956 -3204
rect 3924 -3235 3925 -3205
rect 3925 -3235 3955 -3205
rect 3955 -3235 3956 -3205
rect 3924 -3236 3956 -3235
rect 3924 -3285 3956 -3284
rect 3924 -3315 3925 -3285
rect 3925 -3315 3955 -3285
rect 3955 -3315 3956 -3285
rect 3924 -3316 3956 -3315
rect 3924 -3396 3956 -3364
rect 3924 -3476 3956 -3444
rect 3924 -3525 3956 -3524
rect 3924 -3555 3925 -3525
rect 3925 -3555 3955 -3525
rect 3955 -3555 3956 -3525
rect 3924 -3556 3956 -3555
rect 3924 -3605 3956 -3604
rect 3924 -3635 3925 -3605
rect 3925 -3635 3955 -3605
rect 3955 -3635 3956 -3605
rect 3924 -3636 3956 -3635
rect 3924 -3685 3956 -3684
rect 3924 -3715 3925 -3685
rect 3925 -3715 3955 -3685
rect 3955 -3715 3956 -3685
rect 3924 -3716 3956 -3715
rect 4004 1035 4036 1036
rect 4004 1005 4005 1035
rect 4005 1005 4035 1035
rect 4035 1005 4036 1035
rect 4004 1004 4036 1005
rect 4004 955 4036 956
rect 4004 925 4005 955
rect 4005 925 4035 955
rect 4035 925 4036 955
rect 4004 924 4036 925
rect 4004 875 4036 876
rect 4004 845 4005 875
rect 4005 845 4035 875
rect 4035 845 4036 875
rect 4004 844 4036 845
rect 4004 764 4036 796
rect 4004 684 4036 716
rect 4004 635 4036 636
rect 4004 605 4005 635
rect 4005 605 4035 635
rect 4035 605 4036 635
rect 4004 604 4036 605
rect 4004 555 4036 556
rect 4004 525 4005 555
rect 4005 525 4035 555
rect 4035 525 4036 555
rect 4004 524 4036 525
rect 4004 444 4036 476
rect 4004 395 4036 396
rect 4004 365 4005 395
rect 4005 365 4035 395
rect 4035 365 4036 395
rect 4004 364 4036 365
rect 4004 284 4036 316
rect 4004 235 4036 236
rect 4004 205 4005 235
rect 4005 205 4035 235
rect 4035 205 4036 235
rect 4004 204 4036 205
rect 4004 124 4036 156
rect 4004 75 4036 76
rect 4004 45 4005 75
rect 4005 45 4035 75
rect 4035 45 4036 75
rect 4004 44 4036 45
rect 4004 -5 4036 -4
rect 4004 -35 4005 -5
rect 4005 -35 4035 -5
rect 4035 -35 4036 -5
rect 4004 -36 4036 -35
rect 4004 -85 4036 -84
rect 4004 -115 4005 -85
rect 4005 -115 4035 -85
rect 4035 -115 4036 -85
rect 4004 -116 4036 -115
rect 4004 -165 4036 -164
rect 4004 -195 4005 -165
rect 4005 -195 4035 -165
rect 4035 -195 4036 -165
rect 4004 -196 4036 -195
rect 4004 -245 4036 -244
rect 4004 -275 4005 -245
rect 4005 -275 4035 -245
rect 4035 -275 4036 -245
rect 4004 -276 4036 -275
rect 4004 -325 4036 -324
rect 4004 -355 4005 -325
rect 4005 -355 4035 -325
rect 4035 -355 4036 -325
rect 4004 -356 4036 -355
rect 4004 -436 4036 -404
rect 4004 -485 4036 -484
rect 4004 -515 4005 -485
rect 4005 -515 4035 -485
rect 4035 -515 4036 -485
rect 4004 -516 4036 -515
rect 4004 -596 4036 -564
rect 4004 -645 4036 -644
rect 4004 -675 4005 -645
rect 4005 -675 4035 -645
rect 4035 -675 4036 -645
rect 4004 -676 4036 -675
rect 4004 -756 4036 -724
rect 4004 -805 4036 -804
rect 4004 -835 4005 -805
rect 4005 -835 4035 -805
rect 4035 -835 4036 -805
rect 4004 -836 4036 -835
rect 4004 -885 4036 -884
rect 4004 -915 4005 -885
rect 4005 -915 4035 -885
rect 4035 -915 4036 -885
rect 4004 -916 4036 -915
rect 4004 -996 4036 -964
rect 4004 -1076 4036 -1044
rect 4004 -1125 4036 -1124
rect 4004 -1155 4005 -1125
rect 4005 -1155 4035 -1125
rect 4035 -1155 4036 -1125
rect 4004 -1156 4036 -1155
rect 4004 -1205 4036 -1204
rect 4004 -1235 4005 -1205
rect 4005 -1235 4035 -1205
rect 4035 -1235 4036 -1205
rect 4004 -1236 4036 -1235
rect 4004 -1285 4036 -1284
rect 4004 -1315 4005 -1285
rect 4005 -1315 4035 -1285
rect 4035 -1315 4036 -1285
rect 4004 -1316 4036 -1315
rect 4004 -1365 4036 -1364
rect 4004 -1395 4005 -1365
rect 4005 -1395 4035 -1365
rect 4035 -1395 4036 -1365
rect 4004 -1396 4036 -1395
rect 4004 -1445 4036 -1444
rect 4004 -1475 4005 -1445
rect 4005 -1475 4035 -1445
rect 4035 -1475 4036 -1445
rect 4004 -1476 4036 -1475
rect 4004 -1525 4036 -1524
rect 4004 -1555 4005 -1525
rect 4005 -1555 4035 -1525
rect 4035 -1555 4036 -1525
rect 4004 -1556 4036 -1555
rect 4004 -1636 4036 -1604
rect 4004 -1716 4036 -1684
rect 4004 -1765 4036 -1764
rect 4004 -1795 4005 -1765
rect 4005 -1795 4035 -1765
rect 4035 -1795 4036 -1765
rect 4004 -1796 4036 -1795
rect 4004 -1845 4036 -1844
rect 4004 -1875 4005 -1845
rect 4005 -1875 4035 -1845
rect 4035 -1875 4036 -1845
rect 4004 -1876 4036 -1875
rect 4004 -1956 4036 -1924
rect 4004 -2005 4036 -2004
rect 4004 -2035 4005 -2005
rect 4005 -2035 4035 -2005
rect 4035 -2035 4036 -2005
rect 4004 -2036 4036 -2035
rect 4004 -2116 4036 -2084
rect 4004 -2165 4036 -2164
rect 4004 -2195 4005 -2165
rect 4005 -2195 4035 -2165
rect 4035 -2195 4036 -2165
rect 4004 -2196 4036 -2195
rect 4004 -2276 4036 -2244
rect 4004 -2325 4036 -2324
rect 4004 -2355 4005 -2325
rect 4005 -2355 4035 -2325
rect 4035 -2355 4036 -2325
rect 4004 -2356 4036 -2355
rect 4004 -2405 4036 -2404
rect 4004 -2435 4005 -2405
rect 4005 -2435 4035 -2405
rect 4035 -2435 4036 -2405
rect 4004 -2436 4036 -2435
rect 4004 -2485 4036 -2484
rect 4004 -2515 4005 -2485
rect 4005 -2515 4035 -2485
rect 4035 -2515 4036 -2485
rect 4004 -2516 4036 -2515
rect 4004 -2565 4036 -2564
rect 4004 -2595 4005 -2565
rect 4005 -2595 4035 -2565
rect 4035 -2595 4036 -2565
rect 4004 -2596 4036 -2595
rect 4004 -2645 4036 -2644
rect 4004 -2675 4005 -2645
rect 4005 -2675 4035 -2645
rect 4035 -2675 4036 -2645
rect 4004 -2676 4036 -2675
rect 4004 -2725 4036 -2724
rect 4004 -2755 4005 -2725
rect 4005 -2755 4035 -2725
rect 4035 -2755 4036 -2725
rect 4004 -2756 4036 -2755
rect 4004 -2836 4036 -2804
rect 4004 -2885 4036 -2884
rect 4004 -2915 4005 -2885
rect 4005 -2915 4035 -2885
rect 4035 -2915 4036 -2885
rect 4004 -2916 4036 -2915
rect 4004 -2996 4036 -2964
rect 4004 -3045 4036 -3044
rect 4004 -3075 4005 -3045
rect 4005 -3075 4035 -3045
rect 4035 -3075 4036 -3045
rect 4004 -3076 4036 -3075
rect 4004 -3156 4036 -3124
rect 4004 -3205 4036 -3204
rect 4004 -3235 4005 -3205
rect 4005 -3235 4035 -3205
rect 4035 -3235 4036 -3205
rect 4004 -3236 4036 -3235
rect 4004 -3285 4036 -3284
rect 4004 -3315 4005 -3285
rect 4005 -3315 4035 -3285
rect 4035 -3315 4036 -3285
rect 4004 -3316 4036 -3315
rect 4004 -3396 4036 -3364
rect 4004 -3476 4036 -3444
rect 4004 -3525 4036 -3524
rect 4004 -3555 4005 -3525
rect 4005 -3555 4035 -3525
rect 4035 -3555 4036 -3525
rect 4004 -3556 4036 -3555
rect 4004 -3605 4036 -3604
rect 4004 -3635 4005 -3605
rect 4005 -3635 4035 -3605
rect 4035 -3635 4036 -3605
rect 4004 -3636 4036 -3635
rect 4004 -3685 4036 -3684
rect 4004 -3715 4005 -3685
rect 4005 -3715 4035 -3685
rect 4035 -3715 4036 -3685
rect 4004 -3716 4036 -3715
rect 4084 1035 4116 1036
rect 4084 1005 4085 1035
rect 4085 1005 4115 1035
rect 4115 1005 4116 1035
rect 4084 1004 4116 1005
rect 4084 955 4116 956
rect 4084 925 4085 955
rect 4085 925 4115 955
rect 4115 925 4116 955
rect 4084 924 4116 925
rect 4084 875 4116 876
rect 4084 845 4085 875
rect 4085 845 4115 875
rect 4115 845 4116 875
rect 4084 844 4116 845
rect 4084 764 4116 796
rect 4084 684 4116 716
rect 4084 635 4116 636
rect 4084 605 4085 635
rect 4085 605 4115 635
rect 4115 605 4116 635
rect 4084 604 4116 605
rect 4084 555 4116 556
rect 4084 525 4085 555
rect 4085 525 4115 555
rect 4115 525 4116 555
rect 4084 524 4116 525
rect 4084 444 4116 476
rect 4084 395 4116 396
rect 4084 365 4085 395
rect 4085 365 4115 395
rect 4115 365 4116 395
rect 4084 364 4116 365
rect 4084 284 4116 316
rect 4084 235 4116 236
rect 4084 205 4085 235
rect 4085 205 4115 235
rect 4115 205 4116 235
rect 4084 204 4116 205
rect 4084 124 4116 156
rect 4084 75 4116 76
rect 4084 45 4085 75
rect 4085 45 4115 75
rect 4115 45 4116 75
rect 4084 44 4116 45
rect 4084 -5 4116 -4
rect 4084 -35 4085 -5
rect 4085 -35 4115 -5
rect 4115 -35 4116 -5
rect 4084 -36 4116 -35
rect 4084 -85 4116 -84
rect 4084 -115 4085 -85
rect 4085 -115 4115 -85
rect 4115 -115 4116 -85
rect 4084 -116 4116 -115
rect 4084 -165 4116 -164
rect 4084 -195 4085 -165
rect 4085 -195 4115 -165
rect 4115 -195 4116 -165
rect 4084 -196 4116 -195
rect 4084 -245 4116 -244
rect 4084 -275 4085 -245
rect 4085 -275 4115 -245
rect 4115 -275 4116 -245
rect 4084 -276 4116 -275
rect 4084 -325 4116 -324
rect 4084 -355 4085 -325
rect 4085 -355 4115 -325
rect 4115 -355 4116 -325
rect 4084 -356 4116 -355
rect 4084 -436 4116 -404
rect 4084 -485 4116 -484
rect 4084 -515 4085 -485
rect 4085 -515 4115 -485
rect 4115 -515 4116 -485
rect 4084 -516 4116 -515
rect 4084 -596 4116 -564
rect 4084 -645 4116 -644
rect 4084 -675 4085 -645
rect 4085 -675 4115 -645
rect 4115 -675 4116 -645
rect 4084 -676 4116 -675
rect 4084 -756 4116 -724
rect 4084 -805 4116 -804
rect 4084 -835 4085 -805
rect 4085 -835 4115 -805
rect 4115 -835 4116 -805
rect 4084 -836 4116 -835
rect 4084 -885 4116 -884
rect 4084 -915 4085 -885
rect 4085 -915 4115 -885
rect 4115 -915 4116 -885
rect 4084 -916 4116 -915
rect 4084 -996 4116 -964
rect 4084 -1076 4116 -1044
rect 4084 -1125 4116 -1124
rect 4084 -1155 4085 -1125
rect 4085 -1155 4115 -1125
rect 4115 -1155 4116 -1125
rect 4084 -1156 4116 -1155
rect 4084 -1205 4116 -1204
rect 4084 -1235 4085 -1205
rect 4085 -1235 4115 -1205
rect 4115 -1235 4116 -1205
rect 4084 -1236 4116 -1235
rect 4084 -1285 4116 -1284
rect 4084 -1315 4085 -1285
rect 4085 -1315 4115 -1285
rect 4115 -1315 4116 -1285
rect 4084 -1316 4116 -1315
rect 4084 -1365 4116 -1364
rect 4084 -1395 4085 -1365
rect 4085 -1395 4115 -1365
rect 4115 -1395 4116 -1365
rect 4084 -1396 4116 -1395
rect 4084 -1445 4116 -1444
rect 4084 -1475 4085 -1445
rect 4085 -1475 4115 -1445
rect 4115 -1475 4116 -1445
rect 4084 -1476 4116 -1475
rect 4084 -1525 4116 -1524
rect 4084 -1555 4085 -1525
rect 4085 -1555 4115 -1525
rect 4115 -1555 4116 -1525
rect 4084 -1556 4116 -1555
rect 4084 -1636 4116 -1604
rect 4084 -1716 4116 -1684
rect 4084 -1765 4116 -1764
rect 4084 -1795 4085 -1765
rect 4085 -1795 4115 -1765
rect 4115 -1795 4116 -1765
rect 4084 -1796 4116 -1795
rect 4084 -1845 4116 -1844
rect 4084 -1875 4085 -1845
rect 4085 -1875 4115 -1845
rect 4115 -1875 4116 -1845
rect 4084 -1876 4116 -1875
rect 4084 -1956 4116 -1924
rect 4084 -2005 4116 -2004
rect 4084 -2035 4085 -2005
rect 4085 -2035 4115 -2005
rect 4115 -2035 4116 -2005
rect 4084 -2036 4116 -2035
rect 4084 -2116 4116 -2084
rect 4084 -2165 4116 -2164
rect 4084 -2195 4085 -2165
rect 4085 -2195 4115 -2165
rect 4115 -2195 4116 -2165
rect 4084 -2196 4116 -2195
rect 4084 -2276 4116 -2244
rect 4084 -2325 4116 -2324
rect 4084 -2355 4085 -2325
rect 4085 -2355 4115 -2325
rect 4115 -2355 4116 -2325
rect 4084 -2356 4116 -2355
rect 4084 -2405 4116 -2404
rect 4084 -2435 4085 -2405
rect 4085 -2435 4115 -2405
rect 4115 -2435 4116 -2405
rect 4084 -2436 4116 -2435
rect 4084 -2485 4116 -2484
rect 4084 -2515 4085 -2485
rect 4085 -2515 4115 -2485
rect 4115 -2515 4116 -2485
rect 4084 -2516 4116 -2515
rect 4084 -2565 4116 -2564
rect 4084 -2595 4085 -2565
rect 4085 -2595 4115 -2565
rect 4115 -2595 4116 -2565
rect 4084 -2596 4116 -2595
rect 4084 -2645 4116 -2644
rect 4084 -2675 4085 -2645
rect 4085 -2675 4115 -2645
rect 4115 -2675 4116 -2645
rect 4084 -2676 4116 -2675
rect 4084 -2725 4116 -2724
rect 4084 -2755 4085 -2725
rect 4085 -2755 4115 -2725
rect 4115 -2755 4116 -2725
rect 4084 -2756 4116 -2755
rect 4084 -2836 4116 -2804
rect 4084 -2885 4116 -2884
rect 4084 -2915 4085 -2885
rect 4085 -2915 4115 -2885
rect 4115 -2915 4116 -2885
rect 4084 -2916 4116 -2915
rect 4084 -2996 4116 -2964
rect 4084 -3045 4116 -3044
rect 4084 -3075 4085 -3045
rect 4085 -3075 4115 -3045
rect 4115 -3075 4116 -3045
rect 4084 -3076 4116 -3075
rect 4084 -3156 4116 -3124
rect 4084 -3205 4116 -3204
rect 4084 -3235 4085 -3205
rect 4085 -3235 4115 -3205
rect 4115 -3235 4116 -3205
rect 4084 -3236 4116 -3235
rect 4084 -3285 4116 -3284
rect 4084 -3315 4085 -3285
rect 4085 -3315 4115 -3285
rect 4115 -3315 4116 -3285
rect 4084 -3316 4116 -3315
rect 4084 -3396 4116 -3364
rect 4084 -3476 4116 -3444
rect 4084 -3525 4116 -3524
rect 4084 -3555 4085 -3525
rect 4085 -3555 4115 -3525
rect 4115 -3555 4116 -3525
rect 4084 -3556 4116 -3555
rect 4084 -3605 4116 -3604
rect 4084 -3635 4085 -3605
rect 4085 -3635 4115 -3605
rect 4115 -3635 4116 -3605
rect 4084 -3636 4116 -3635
rect 4084 -3685 4116 -3684
rect 4084 -3715 4085 -3685
rect 4085 -3715 4115 -3685
rect 4115 -3715 4116 -3685
rect 4084 -3716 4116 -3715
rect 4164 1035 4196 1036
rect 4164 1005 4165 1035
rect 4165 1005 4195 1035
rect 4195 1005 4196 1035
rect 4164 1004 4196 1005
rect 4164 955 4196 956
rect 4164 925 4165 955
rect 4165 925 4195 955
rect 4195 925 4196 955
rect 4164 924 4196 925
rect 4164 875 4196 876
rect 4164 845 4165 875
rect 4165 845 4195 875
rect 4195 845 4196 875
rect 4164 844 4196 845
rect 4164 764 4196 796
rect 4164 684 4196 716
rect 4164 635 4196 636
rect 4164 605 4165 635
rect 4165 605 4195 635
rect 4195 605 4196 635
rect 4164 604 4196 605
rect 4164 555 4196 556
rect 4164 525 4165 555
rect 4165 525 4195 555
rect 4195 525 4196 555
rect 4164 524 4196 525
rect 4164 444 4196 476
rect 4164 395 4196 396
rect 4164 365 4165 395
rect 4165 365 4195 395
rect 4195 365 4196 395
rect 4164 364 4196 365
rect 4164 284 4196 316
rect 4164 235 4196 236
rect 4164 205 4165 235
rect 4165 205 4195 235
rect 4195 205 4196 235
rect 4164 204 4196 205
rect 4164 124 4196 156
rect 4164 75 4196 76
rect 4164 45 4165 75
rect 4165 45 4195 75
rect 4195 45 4196 75
rect 4164 44 4196 45
rect 4164 -5 4196 -4
rect 4164 -35 4165 -5
rect 4165 -35 4195 -5
rect 4195 -35 4196 -5
rect 4164 -36 4196 -35
rect 4164 -85 4196 -84
rect 4164 -115 4165 -85
rect 4165 -115 4195 -85
rect 4195 -115 4196 -85
rect 4164 -116 4196 -115
rect 4164 -165 4196 -164
rect 4164 -195 4165 -165
rect 4165 -195 4195 -165
rect 4195 -195 4196 -165
rect 4164 -196 4196 -195
rect 4164 -245 4196 -244
rect 4164 -275 4165 -245
rect 4165 -275 4195 -245
rect 4195 -275 4196 -245
rect 4164 -276 4196 -275
rect 4164 -325 4196 -324
rect 4164 -355 4165 -325
rect 4165 -355 4195 -325
rect 4195 -355 4196 -325
rect 4164 -356 4196 -355
rect 4164 -436 4196 -404
rect 4164 -485 4196 -484
rect 4164 -515 4165 -485
rect 4165 -515 4195 -485
rect 4195 -515 4196 -485
rect 4164 -516 4196 -515
rect 4164 -596 4196 -564
rect 4164 -645 4196 -644
rect 4164 -675 4165 -645
rect 4165 -675 4195 -645
rect 4195 -675 4196 -645
rect 4164 -676 4196 -675
rect 4164 -756 4196 -724
rect 4164 -805 4196 -804
rect 4164 -835 4165 -805
rect 4165 -835 4195 -805
rect 4195 -835 4196 -805
rect 4164 -836 4196 -835
rect 4164 -885 4196 -884
rect 4164 -915 4165 -885
rect 4165 -915 4195 -885
rect 4195 -915 4196 -885
rect 4164 -916 4196 -915
rect 4164 -996 4196 -964
rect 4164 -1076 4196 -1044
rect 4164 -1125 4196 -1124
rect 4164 -1155 4165 -1125
rect 4165 -1155 4195 -1125
rect 4195 -1155 4196 -1125
rect 4164 -1156 4196 -1155
rect 4164 -1205 4196 -1204
rect 4164 -1235 4165 -1205
rect 4165 -1235 4195 -1205
rect 4195 -1235 4196 -1205
rect 4164 -1236 4196 -1235
rect 4164 -1285 4196 -1284
rect 4164 -1315 4165 -1285
rect 4165 -1315 4195 -1285
rect 4195 -1315 4196 -1285
rect 4164 -1316 4196 -1315
rect 4164 -1365 4196 -1364
rect 4164 -1395 4165 -1365
rect 4165 -1395 4195 -1365
rect 4195 -1395 4196 -1365
rect 4164 -1396 4196 -1395
rect 4164 -1445 4196 -1444
rect 4164 -1475 4165 -1445
rect 4165 -1475 4195 -1445
rect 4195 -1475 4196 -1445
rect 4164 -1476 4196 -1475
rect 4164 -1525 4196 -1524
rect 4164 -1555 4165 -1525
rect 4165 -1555 4195 -1525
rect 4195 -1555 4196 -1525
rect 4164 -1556 4196 -1555
rect 4164 -1636 4196 -1604
rect 4164 -1716 4196 -1684
rect 4164 -1765 4196 -1764
rect 4164 -1795 4165 -1765
rect 4165 -1795 4195 -1765
rect 4195 -1795 4196 -1765
rect 4164 -1796 4196 -1795
rect 4164 -1845 4196 -1844
rect 4164 -1875 4165 -1845
rect 4165 -1875 4195 -1845
rect 4195 -1875 4196 -1845
rect 4164 -1876 4196 -1875
rect 4164 -1956 4196 -1924
rect 4164 -2005 4196 -2004
rect 4164 -2035 4165 -2005
rect 4165 -2035 4195 -2005
rect 4195 -2035 4196 -2005
rect 4164 -2036 4196 -2035
rect 4164 -2116 4196 -2084
rect 4164 -2165 4196 -2164
rect 4164 -2195 4165 -2165
rect 4165 -2195 4195 -2165
rect 4195 -2195 4196 -2165
rect 4164 -2196 4196 -2195
rect 4164 -2276 4196 -2244
rect 4164 -2325 4196 -2324
rect 4164 -2355 4165 -2325
rect 4165 -2355 4195 -2325
rect 4195 -2355 4196 -2325
rect 4164 -2356 4196 -2355
rect 4164 -2405 4196 -2404
rect 4164 -2435 4165 -2405
rect 4165 -2435 4195 -2405
rect 4195 -2435 4196 -2405
rect 4164 -2436 4196 -2435
rect 4164 -2485 4196 -2484
rect 4164 -2515 4165 -2485
rect 4165 -2515 4195 -2485
rect 4195 -2515 4196 -2485
rect 4164 -2516 4196 -2515
rect 4164 -2565 4196 -2564
rect 4164 -2595 4165 -2565
rect 4165 -2595 4195 -2565
rect 4195 -2595 4196 -2565
rect 4164 -2596 4196 -2595
rect 4164 -2645 4196 -2644
rect 4164 -2675 4165 -2645
rect 4165 -2675 4195 -2645
rect 4195 -2675 4196 -2645
rect 4164 -2676 4196 -2675
rect 4164 -2725 4196 -2724
rect 4164 -2755 4165 -2725
rect 4165 -2755 4195 -2725
rect 4195 -2755 4196 -2725
rect 4164 -2756 4196 -2755
rect 4164 -2836 4196 -2804
rect 4164 -2885 4196 -2884
rect 4164 -2915 4165 -2885
rect 4165 -2915 4195 -2885
rect 4195 -2915 4196 -2885
rect 4164 -2916 4196 -2915
rect 4164 -2996 4196 -2964
rect 4164 -3045 4196 -3044
rect 4164 -3075 4165 -3045
rect 4165 -3075 4195 -3045
rect 4195 -3075 4196 -3045
rect 4164 -3076 4196 -3075
rect 4164 -3156 4196 -3124
rect 4164 -3205 4196 -3204
rect 4164 -3235 4165 -3205
rect 4165 -3235 4195 -3205
rect 4195 -3235 4196 -3205
rect 4164 -3236 4196 -3235
rect 4164 -3285 4196 -3284
rect 4164 -3315 4165 -3285
rect 4165 -3315 4195 -3285
rect 4195 -3315 4196 -3285
rect 4164 -3316 4196 -3315
rect 4164 -3396 4196 -3364
rect 4164 -3476 4196 -3444
rect 4164 -3525 4196 -3524
rect 4164 -3555 4165 -3525
rect 4165 -3555 4195 -3525
rect 4195 -3555 4196 -3525
rect 4164 -3556 4196 -3555
rect 4164 -3605 4196 -3604
rect 4164 -3635 4165 -3605
rect 4165 -3635 4195 -3605
rect 4195 -3635 4196 -3605
rect 4164 -3636 4196 -3635
rect 4164 -3685 4196 -3684
rect 4164 -3715 4165 -3685
rect 4165 -3715 4195 -3685
rect 4195 -3715 4196 -3685
rect 4164 -3716 4196 -3715
rect 4244 1035 4276 1036
rect 4244 1005 4245 1035
rect 4245 1005 4275 1035
rect 4275 1005 4276 1035
rect 4244 1004 4276 1005
rect 4244 955 4276 956
rect 4244 925 4245 955
rect 4245 925 4275 955
rect 4275 925 4276 955
rect 4244 924 4276 925
rect 4244 875 4276 876
rect 4244 845 4245 875
rect 4245 845 4275 875
rect 4275 845 4276 875
rect 4244 844 4276 845
rect 4244 764 4276 796
rect 4244 684 4276 716
rect 4244 635 4276 636
rect 4244 605 4245 635
rect 4245 605 4275 635
rect 4275 605 4276 635
rect 4244 604 4276 605
rect 4244 555 4276 556
rect 4244 525 4245 555
rect 4245 525 4275 555
rect 4275 525 4276 555
rect 4244 524 4276 525
rect 4244 444 4276 476
rect 4244 395 4276 396
rect 4244 365 4245 395
rect 4245 365 4275 395
rect 4275 365 4276 395
rect 4244 364 4276 365
rect 4244 284 4276 316
rect 4244 235 4276 236
rect 4244 205 4245 235
rect 4245 205 4275 235
rect 4275 205 4276 235
rect 4244 204 4276 205
rect 4244 124 4276 156
rect 4244 75 4276 76
rect 4244 45 4245 75
rect 4245 45 4275 75
rect 4275 45 4276 75
rect 4244 44 4276 45
rect 4244 -5 4276 -4
rect 4244 -35 4245 -5
rect 4245 -35 4275 -5
rect 4275 -35 4276 -5
rect 4244 -36 4276 -35
rect 4244 -85 4276 -84
rect 4244 -115 4245 -85
rect 4245 -115 4275 -85
rect 4275 -115 4276 -85
rect 4244 -116 4276 -115
rect 4244 -165 4276 -164
rect 4244 -195 4245 -165
rect 4245 -195 4275 -165
rect 4275 -195 4276 -165
rect 4244 -196 4276 -195
rect 4244 -245 4276 -244
rect 4244 -275 4245 -245
rect 4245 -275 4275 -245
rect 4275 -275 4276 -245
rect 4244 -276 4276 -275
rect 4244 -325 4276 -324
rect 4244 -355 4245 -325
rect 4245 -355 4275 -325
rect 4275 -355 4276 -325
rect 4244 -356 4276 -355
rect 4244 -436 4276 -404
rect 4244 -485 4276 -484
rect 4244 -515 4245 -485
rect 4245 -515 4275 -485
rect 4275 -515 4276 -485
rect 4244 -516 4276 -515
rect 4244 -596 4276 -564
rect 4244 -645 4276 -644
rect 4244 -675 4245 -645
rect 4245 -675 4275 -645
rect 4275 -675 4276 -645
rect 4244 -676 4276 -675
rect 4244 -756 4276 -724
rect 4244 -805 4276 -804
rect 4244 -835 4245 -805
rect 4245 -835 4275 -805
rect 4275 -835 4276 -805
rect 4244 -836 4276 -835
rect 4244 -885 4276 -884
rect 4244 -915 4245 -885
rect 4245 -915 4275 -885
rect 4275 -915 4276 -885
rect 4244 -916 4276 -915
rect 4244 -996 4276 -964
rect 4244 -1076 4276 -1044
rect 4244 -1125 4276 -1124
rect 4244 -1155 4245 -1125
rect 4245 -1155 4275 -1125
rect 4275 -1155 4276 -1125
rect 4244 -1156 4276 -1155
rect 4244 -1205 4276 -1204
rect 4244 -1235 4245 -1205
rect 4245 -1235 4275 -1205
rect 4275 -1235 4276 -1205
rect 4244 -1236 4276 -1235
rect 4244 -1285 4276 -1284
rect 4244 -1315 4245 -1285
rect 4245 -1315 4275 -1285
rect 4275 -1315 4276 -1285
rect 4244 -1316 4276 -1315
rect 4244 -1365 4276 -1364
rect 4244 -1395 4245 -1365
rect 4245 -1395 4275 -1365
rect 4275 -1395 4276 -1365
rect 4244 -1396 4276 -1395
rect 4244 -1445 4276 -1444
rect 4244 -1475 4245 -1445
rect 4245 -1475 4275 -1445
rect 4275 -1475 4276 -1445
rect 4244 -1476 4276 -1475
rect 4244 -1525 4276 -1524
rect 4244 -1555 4245 -1525
rect 4245 -1555 4275 -1525
rect 4275 -1555 4276 -1525
rect 4244 -1556 4276 -1555
rect 4244 -1636 4276 -1604
rect 4244 -1716 4276 -1684
rect 4244 -1765 4276 -1764
rect 4244 -1795 4245 -1765
rect 4245 -1795 4275 -1765
rect 4275 -1795 4276 -1765
rect 4244 -1796 4276 -1795
rect 4244 -1845 4276 -1844
rect 4244 -1875 4245 -1845
rect 4245 -1875 4275 -1845
rect 4275 -1875 4276 -1845
rect 4244 -1876 4276 -1875
rect 4244 -1956 4276 -1924
rect 4244 -2005 4276 -2004
rect 4244 -2035 4245 -2005
rect 4245 -2035 4275 -2005
rect 4275 -2035 4276 -2005
rect 4244 -2036 4276 -2035
rect 4244 -2116 4276 -2084
rect 4244 -2165 4276 -2164
rect 4244 -2195 4245 -2165
rect 4245 -2195 4275 -2165
rect 4275 -2195 4276 -2165
rect 4244 -2196 4276 -2195
rect 4244 -2276 4276 -2244
rect 4244 -2325 4276 -2324
rect 4244 -2355 4245 -2325
rect 4245 -2355 4275 -2325
rect 4275 -2355 4276 -2325
rect 4244 -2356 4276 -2355
rect 4244 -2405 4276 -2404
rect 4244 -2435 4245 -2405
rect 4245 -2435 4275 -2405
rect 4275 -2435 4276 -2405
rect 4244 -2436 4276 -2435
rect 4244 -2485 4276 -2484
rect 4244 -2515 4245 -2485
rect 4245 -2515 4275 -2485
rect 4275 -2515 4276 -2485
rect 4244 -2516 4276 -2515
rect 4244 -2565 4276 -2564
rect 4244 -2595 4245 -2565
rect 4245 -2595 4275 -2565
rect 4275 -2595 4276 -2565
rect 4244 -2596 4276 -2595
rect 4244 -2645 4276 -2644
rect 4244 -2675 4245 -2645
rect 4245 -2675 4275 -2645
rect 4275 -2675 4276 -2645
rect 4244 -2676 4276 -2675
rect 4244 -2725 4276 -2724
rect 4244 -2755 4245 -2725
rect 4245 -2755 4275 -2725
rect 4275 -2755 4276 -2725
rect 4244 -2756 4276 -2755
rect 4244 -2836 4276 -2804
rect 4244 -2885 4276 -2884
rect 4244 -2915 4245 -2885
rect 4245 -2915 4275 -2885
rect 4275 -2915 4276 -2885
rect 4244 -2916 4276 -2915
rect 4244 -2996 4276 -2964
rect 4244 -3045 4276 -3044
rect 4244 -3075 4245 -3045
rect 4245 -3075 4275 -3045
rect 4275 -3075 4276 -3045
rect 4244 -3076 4276 -3075
rect 4244 -3156 4276 -3124
rect 4244 -3205 4276 -3204
rect 4244 -3235 4245 -3205
rect 4245 -3235 4275 -3205
rect 4275 -3235 4276 -3205
rect 4244 -3236 4276 -3235
rect 4244 -3285 4276 -3284
rect 4244 -3315 4245 -3285
rect 4245 -3315 4275 -3285
rect 4275 -3315 4276 -3285
rect 4244 -3316 4276 -3315
rect 4244 -3396 4276 -3364
rect 4244 -3476 4276 -3444
rect 4244 -3525 4276 -3524
rect 4244 -3555 4245 -3525
rect 4245 -3555 4275 -3525
rect 4275 -3555 4276 -3525
rect 4244 -3556 4276 -3555
rect 4244 -3605 4276 -3604
rect 4244 -3635 4245 -3605
rect 4245 -3635 4275 -3605
rect 4275 -3635 4276 -3605
rect 4244 -3636 4276 -3635
rect 4244 -3685 4276 -3684
rect 4244 -3715 4245 -3685
rect 4245 -3715 4275 -3685
rect 4275 -3715 4276 -3685
rect 4244 -3716 4276 -3715
rect 4324 1035 4356 1036
rect 4324 1005 4325 1035
rect 4325 1005 4355 1035
rect 4355 1005 4356 1035
rect 4324 1004 4356 1005
rect 4324 955 4356 956
rect 4324 925 4325 955
rect 4325 925 4355 955
rect 4355 925 4356 955
rect 4324 924 4356 925
rect 4324 875 4356 876
rect 4324 845 4325 875
rect 4325 845 4355 875
rect 4355 845 4356 875
rect 4324 844 4356 845
rect 4324 764 4356 796
rect 4324 684 4356 716
rect 4324 635 4356 636
rect 4324 605 4325 635
rect 4325 605 4355 635
rect 4355 605 4356 635
rect 4324 604 4356 605
rect 4324 555 4356 556
rect 4324 525 4325 555
rect 4325 525 4355 555
rect 4355 525 4356 555
rect 4324 524 4356 525
rect 4324 444 4356 476
rect 4324 395 4356 396
rect 4324 365 4325 395
rect 4325 365 4355 395
rect 4355 365 4356 395
rect 4324 364 4356 365
rect 4324 284 4356 316
rect 4324 235 4356 236
rect 4324 205 4325 235
rect 4325 205 4355 235
rect 4355 205 4356 235
rect 4324 204 4356 205
rect 4324 124 4356 156
rect 4324 75 4356 76
rect 4324 45 4325 75
rect 4325 45 4355 75
rect 4355 45 4356 75
rect 4324 44 4356 45
rect 4324 -5 4356 -4
rect 4324 -35 4325 -5
rect 4325 -35 4355 -5
rect 4355 -35 4356 -5
rect 4324 -36 4356 -35
rect 4324 -85 4356 -84
rect 4324 -115 4325 -85
rect 4325 -115 4355 -85
rect 4355 -115 4356 -85
rect 4324 -116 4356 -115
rect 4324 -165 4356 -164
rect 4324 -195 4325 -165
rect 4325 -195 4355 -165
rect 4355 -195 4356 -165
rect 4324 -196 4356 -195
rect 4324 -245 4356 -244
rect 4324 -275 4325 -245
rect 4325 -275 4355 -245
rect 4355 -275 4356 -245
rect 4324 -276 4356 -275
rect 4324 -325 4356 -324
rect 4324 -355 4325 -325
rect 4325 -355 4355 -325
rect 4355 -355 4356 -325
rect 4324 -356 4356 -355
rect 4324 -436 4356 -404
rect 4324 -485 4356 -484
rect 4324 -515 4325 -485
rect 4325 -515 4355 -485
rect 4355 -515 4356 -485
rect 4324 -516 4356 -515
rect 4324 -596 4356 -564
rect 4324 -645 4356 -644
rect 4324 -675 4325 -645
rect 4325 -675 4355 -645
rect 4355 -675 4356 -645
rect 4324 -676 4356 -675
rect 4324 -756 4356 -724
rect 4324 -805 4356 -804
rect 4324 -835 4325 -805
rect 4325 -835 4355 -805
rect 4355 -835 4356 -805
rect 4324 -836 4356 -835
rect 4324 -885 4356 -884
rect 4324 -915 4325 -885
rect 4325 -915 4355 -885
rect 4355 -915 4356 -885
rect 4324 -916 4356 -915
rect 4324 -996 4356 -964
rect 4324 -1076 4356 -1044
rect 4324 -1125 4356 -1124
rect 4324 -1155 4325 -1125
rect 4325 -1155 4355 -1125
rect 4355 -1155 4356 -1125
rect 4324 -1156 4356 -1155
rect 4324 -1205 4356 -1204
rect 4324 -1235 4325 -1205
rect 4325 -1235 4355 -1205
rect 4355 -1235 4356 -1205
rect 4324 -1236 4356 -1235
rect 4324 -1285 4356 -1284
rect 4324 -1315 4325 -1285
rect 4325 -1315 4355 -1285
rect 4355 -1315 4356 -1285
rect 4324 -1316 4356 -1315
rect 4324 -1365 4356 -1364
rect 4324 -1395 4325 -1365
rect 4325 -1395 4355 -1365
rect 4355 -1395 4356 -1365
rect 4324 -1396 4356 -1395
rect 4324 -1445 4356 -1444
rect 4324 -1475 4325 -1445
rect 4325 -1475 4355 -1445
rect 4355 -1475 4356 -1445
rect 4324 -1476 4356 -1475
rect 4324 -1525 4356 -1524
rect 4324 -1555 4325 -1525
rect 4325 -1555 4355 -1525
rect 4355 -1555 4356 -1525
rect 4324 -1556 4356 -1555
rect 4324 -1636 4356 -1604
rect 4324 -1716 4356 -1684
rect 4324 -1765 4356 -1764
rect 4324 -1795 4325 -1765
rect 4325 -1795 4355 -1765
rect 4355 -1795 4356 -1765
rect 4324 -1796 4356 -1795
rect 4324 -1845 4356 -1844
rect 4324 -1875 4325 -1845
rect 4325 -1875 4355 -1845
rect 4355 -1875 4356 -1845
rect 4324 -1876 4356 -1875
rect 4324 -1956 4356 -1924
rect 4324 -2005 4356 -2004
rect 4324 -2035 4325 -2005
rect 4325 -2035 4355 -2005
rect 4355 -2035 4356 -2005
rect 4324 -2036 4356 -2035
rect 4324 -2116 4356 -2084
rect 4324 -2165 4356 -2164
rect 4324 -2195 4325 -2165
rect 4325 -2195 4355 -2165
rect 4355 -2195 4356 -2165
rect 4324 -2196 4356 -2195
rect 4324 -2276 4356 -2244
rect 4324 -2325 4356 -2324
rect 4324 -2355 4325 -2325
rect 4325 -2355 4355 -2325
rect 4355 -2355 4356 -2325
rect 4324 -2356 4356 -2355
rect 4324 -2405 4356 -2404
rect 4324 -2435 4325 -2405
rect 4325 -2435 4355 -2405
rect 4355 -2435 4356 -2405
rect 4324 -2436 4356 -2435
rect 4324 -2485 4356 -2484
rect 4324 -2515 4325 -2485
rect 4325 -2515 4355 -2485
rect 4355 -2515 4356 -2485
rect 4324 -2516 4356 -2515
rect 4324 -2565 4356 -2564
rect 4324 -2595 4325 -2565
rect 4325 -2595 4355 -2565
rect 4355 -2595 4356 -2565
rect 4324 -2596 4356 -2595
rect 4324 -2645 4356 -2644
rect 4324 -2675 4325 -2645
rect 4325 -2675 4355 -2645
rect 4355 -2675 4356 -2645
rect 4324 -2676 4356 -2675
rect 4324 -2725 4356 -2724
rect 4324 -2755 4325 -2725
rect 4325 -2755 4355 -2725
rect 4355 -2755 4356 -2725
rect 4324 -2756 4356 -2755
rect 4324 -2836 4356 -2804
rect 4324 -2885 4356 -2884
rect 4324 -2915 4325 -2885
rect 4325 -2915 4355 -2885
rect 4355 -2915 4356 -2885
rect 4324 -2916 4356 -2915
rect 4324 -2996 4356 -2964
rect 4324 -3045 4356 -3044
rect 4324 -3075 4325 -3045
rect 4325 -3075 4355 -3045
rect 4355 -3075 4356 -3045
rect 4324 -3076 4356 -3075
rect 4324 -3156 4356 -3124
rect 4324 -3205 4356 -3204
rect 4324 -3235 4325 -3205
rect 4325 -3235 4355 -3205
rect 4355 -3235 4356 -3205
rect 4324 -3236 4356 -3235
rect 4324 -3285 4356 -3284
rect 4324 -3315 4325 -3285
rect 4325 -3315 4355 -3285
rect 4355 -3315 4356 -3285
rect 4324 -3316 4356 -3315
rect 4324 -3396 4356 -3364
rect 4324 -3476 4356 -3444
rect 4324 -3525 4356 -3524
rect 4324 -3555 4325 -3525
rect 4325 -3555 4355 -3525
rect 4355 -3555 4356 -3525
rect 4324 -3556 4356 -3555
rect 4324 -3605 4356 -3604
rect 4324 -3635 4325 -3605
rect 4325 -3635 4355 -3605
rect 4355 -3635 4356 -3605
rect 4324 -3636 4356 -3635
rect 4324 -3685 4356 -3684
rect 4324 -3715 4325 -3685
rect 4325 -3715 4355 -3685
rect 4355 -3715 4356 -3685
rect 4324 -3716 4356 -3715
rect 4404 1035 4436 1036
rect 4404 1005 4405 1035
rect 4405 1005 4435 1035
rect 4435 1005 4436 1035
rect 4404 1004 4436 1005
rect 4404 955 4436 956
rect 4404 925 4405 955
rect 4405 925 4435 955
rect 4435 925 4436 955
rect 4404 924 4436 925
rect 4404 875 4436 876
rect 4404 845 4405 875
rect 4405 845 4435 875
rect 4435 845 4436 875
rect 4404 844 4436 845
rect 4404 764 4436 796
rect 4404 684 4436 716
rect 4404 635 4436 636
rect 4404 605 4405 635
rect 4405 605 4435 635
rect 4435 605 4436 635
rect 4404 604 4436 605
rect 4404 555 4436 556
rect 4404 525 4405 555
rect 4405 525 4435 555
rect 4435 525 4436 555
rect 4404 524 4436 525
rect 4404 444 4436 476
rect 4404 395 4436 396
rect 4404 365 4405 395
rect 4405 365 4435 395
rect 4435 365 4436 395
rect 4404 364 4436 365
rect 4404 284 4436 316
rect 4404 235 4436 236
rect 4404 205 4405 235
rect 4405 205 4435 235
rect 4435 205 4436 235
rect 4404 204 4436 205
rect 4404 124 4436 156
rect 4404 75 4436 76
rect 4404 45 4405 75
rect 4405 45 4435 75
rect 4435 45 4436 75
rect 4404 44 4436 45
rect 4404 -5 4436 -4
rect 4404 -35 4405 -5
rect 4405 -35 4435 -5
rect 4435 -35 4436 -5
rect 4404 -36 4436 -35
rect 4404 -85 4436 -84
rect 4404 -115 4405 -85
rect 4405 -115 4435 -85
rect 4435 -115 4436 -85
rect 4404 -116 4436 -115
rect 4404 -165 4436 -164
rect 4404 -195 4405 -165
rect 4405 -195 4435 -165
rect 4435 -195 4436 -165
rect 4404 -196 4436 -195
rect 4404 -245 4436 -244
rect 4404 -275 4405 -245
rect 4405 -275 4435 -245
rect 4435 -275 4436 -245
rect 4404 -276 4436 -275
rect 4404 -325 4436 -324
rect 4404 -355 4405 -325
rect 4405 -355 4435 -325
rect 4435 -355 4436 -325
rect 4404 -356 4436 -355
rect 4404 -436 4436 -404
rect 4404 -485 4436 -484
rect 4404 -515 4405 -485
rect 4405 -515 4435 -485
rect 4435 -515 4436 -485
rect 4404 -516 4436 -515
rect 4404 -596 4436 -564
rect 4404 -645 4436 -644
rect 4404 -675 4405 -645
rect 4405 -675 4435 -645
rect 4435 -675 4436 -645
rect 4404 -676 4436 -675
rect 4404 -756 4436 -724
rect 4404 -805 4436 -804
rect 4404 -835 4405 -805
rect 4405 -835 4435 -805
rect 4435 -835 4436 -805
rect 4404 -836 4436 -835
rect 4404 -885 4436 -884
rect 4404 -915 4405 -885
rect 4405 -915 4435 -885
rect 4435 -915 4436 -885
rect 4404 -916 4436 -915
rect 4404 -996 4436 -964
rect 4404 -1076 4436 -1044
rect 4404 -1125 4436 -1124
rect 4404 -1155 4405 -1125
rect 4405 -1155 4435 -1125
rect 4435 -1155 4436 -1125
rect 4404 -1156 4436 -1155
rect 4404 -1205 4436 -1204
rect 4404 -1235 4405 -1205
rect 4405 -1235 4435 -1205
rect 4435 -1235 4436 -1205
rect 4404 -1236 4436 -1235
rect 4404 -1285 4436 -1284
rect 4404 -1315 4405 -1285
rect 4405 -1315 4435 -1285
rect 4435 -1315 4436 -1285
rect 4404 -1316 4436 -1315
rect 4404 -1365 4436 -1364
rect 4404 -1395 4405 -1365
rect 4405 -1395 4435 -1365
rect 4435 -1395 4436 -1365
rect 4404 -1396 4436 -1395
rect 4404 -1445 4436 -1444
rect 4404 -1475 4405 -1445
rect 4405 -1475 4435 -1445
rect 4435 -1475 4436 -1445
rect 4404 -1476 4436 -1475
rect 4404 -1525 4436 -1524
rect 4404 -1555 4405 -1525
rect 4405 -1555 4435 -1525
rect 4435 -1555 4436 -1525
rect 4404 -1556 4436 -1555
rect 4404 -1636 4436 -1604
rect 4404 -1716 4436 -1684
rect 4404 -1765 4436 -1764
rect 4404 -1795 4405 -1765
rect 4405 -1795 4435 -1765
rect 4435 -1795 4436 -1765
rect 4404 -1796 4436 -1795
rect 4404 -1845 4436 -1844
rect 4404 -1875 4405 -1845
rect 4405 -1875 4435 -1845
rect 4435 -1875 4436 -1845
rect 4404 -1876 4436 -1875
rect 4404 -1956 4436 -1924
rect 4404 -2005 4436 -2004
rect 4404 -2035 4405 -2005
rect 4405 -2035 4435 -2005
rect 4435 -2035 4436 -2005
rect 4404 -2036 4436 -2035
rect 4404 -2116 4436 -2084
rect 4404 -2165 4436 -2164
rect 4404 -2195 4405 -2165
rect 4405 -2195 4435 -2165
rect 4435 -2195 4436 -2165
rect 4404 -2196 4436 -2195
rect 4404 -2276 4436 -2244
rect 4404 -2325 4436 -2324
rect 4404 -2355 4405 -2325
rect 4405 -2355 4435 -2325
rect 4435 -2355 4436 -2325
rect 4404 -2356 4436 -2355
rect 4404 -2405 4436 -2404
rect 4404 -2435 4405 -2405
rect 4405 -2435 4435 -2405
rect 4435 -2435 4436 -2405
rect 4404 -2436 4436 -2435
rect 4404 -2485 4436 -2484
rect 4404 -2515 4405 -2485
rect 4405 -2515 4435 -2485
rect 4435 -2515 4436 -2485
rect 4404 -2516 4436 -2515
rect 4404 -2565 4436 -2564
rect 4404 -2595 4405 -2565
rect 4405 -2595 4435 -2565
rect 4435 -2595 4436 -2565
rect 4404 -2596 4436 -2595
rect 4404 -2645 4436 -2644
rect 4404 -2675 4405 -2645
rect 4405 -2675 4435 -2645
rect 4435 -2675 4436 -2645
rect 4404 -2676 4436 -2675
rect 4404 -2725 4436 -2724
rect 4404 -2755 4405 -2725
rect 4405 -2755 4435 -2725
rect 4435 -2755 4436 -2725
rect 4404 -2756 4436 -2755
rect 4404 -2836 4436 -2804
rect 4404 -2885 4436 -2884
rect 4404 -2915 4405 -2885
rect 4405 -2915 4435 -2885
rect 4435 -2915 4436 -2885
rect 4404 -2916 4436 -2915
rect 4404 -2996 4436 -2964
rect 4404 -3045 4436 -3044
rect 4404 -3075 4405 -3045
rect 4405 -3075 4435 -3045
rect 4435 -3075 4436 -3045
rect 4404 -3076 4436 -3075
rect 4404 -3156 4436 -3124
rect 4404 -3205 4436 -3204
rect 4404 -3235 4405 -3205
rect 4405 -3235 4435 -3205
rect 4435 -3235 4436 -3205
rect 4404 -3236 4436 -3235
rect 4404 -3285 4436 -3284
rect 4404 -3315 4405 -3285
rect 4405 -3315 4435 -3285
rect 4435 -3315 4436 -3285
rect 4404 -3316 4436 -3315
rect 4404 -3396 4436 -3364
rect 4404 -3476 4436 -3444
rect 4404 -3525 4436 -3524
rect 4404 -3555 4405 -3525
rect 4405 -3555 4435 -3525
rect 4435 -3555 4436 -3525
rect 4404 -3556 4436 -3555
rect 4404 -3605 4436 -3604
rect 4404 -3635 4405 -3605
rect 4405 -3635 4435 -3605
rect 4435 -3635 4436 -3605
rect 4404 -3636 4436 -3635
rect 4404 -3685 4436 -3684
rect 4404 -3715 4405 -3685
rect 4405 -3715 4435 -3685
rect 4435 -3715 4436 -3685
rect 4404 -3716 4436 -3715
rect 4484 1035 4516 1036
rect 4484 1005 4485 1035
rect 4485 1005 4515 1035
rect 4515 1005 4516 1035
rect 4484 1004 4516 1005
rect 4484 955 4516 956
rect 4484 925 4485 955
rect 4485 925 4515 955
rect 4515 925 4516 955
rect 4484 924 4516 925
rect 4484 875 4516 876
rect 4484 845 4485 875
rect 4485 845 4515 875
rect 4515 845 4516 875
rect 4484 844 4516 845
rect 4484 764 4516 796
rect 4484 684 4516 716
rect 4484 635 4516 636
rect 4484 605 4485 635
rect 4485 605 4515 635
rect 4515 605 4516 635
rect 4484 604 4516 605
rect 4484 555 4516 556
rect 4484 525 4485 555
rect 4485 525 4515 555
rect 4515 525 4516 555
rect 4484 524 4516 525
rect 4484 444 4516 476
rect 4484 395 4516 396
rect 4484 365 4485 395
rect 4485 365 4515 395
rect 4515 365 4516 395
rect 4484 364 4516 365
rect 4484 284 4516 316
rect 4484 235 4516 236
rect 4484 205 4485 235
rect 4485 205 4515 235
rect 4515 205 4516 235
rect 4484 204 4516 205
rect 4484 124 4516 156
rect 4484 75 4516 76
rect 4484 45 4485 75
rect 4485 45 4515 75
rect 4515 45 4516 75
rect 4484 44 4516 45
rect 4484 -5 4516 -4
rect 4484 -35 4485 -5
rect 4485 -35 4515 -5
rect 4515 -35 4516 -5
rect 4484 -36 4516 -35
rect 4484 -85 4516 -84
rect 4484 -115 4485 -85
rect 4485 -115 4515 -85
rect 4515 -115 4516 -85
rect 4484 -116 4516 -115
rect 4484 -165 4516 -164
rect 4484 -195 4485 -165
rect 4485 -195 4515 -165
rect 4515 -195 4516 -165
rect 4484 -196 4516 -195
rect 4484 -245 4516 -244
rect 4484 -275 4485 -245
rect 4485 -275 4515 -245
rect 4515 -275 4516 -245
rect 4484 -276 4516 -275
rect 4484 -325 4516 -324
rect 4484 -355 4485 -325
rect 4485 -355 4515 -325
rect 4515 -355 4516 -325
rect 4484 -356 4516 -355
rect 4484 -436 4516 -404
rect 4484 -485 4516 -484
rect 4484 -515 4485 -485
rect 4485 -515 4515 -485
rect 4515 -515 4516 -485
rect 4484 -516 4516 -515
rect 4484 -596 4516 -564
rect 4484 -645 4516 -644
rect 4484 -675 4485 -645
rect 4485 -675 4515 -645
rect 4515 -675 4516 -645
rect 4484 -676 4516 -675
rect 4484 -756 4516 -724
rect 4484 -805 4516 -804
rect 4484 -835 4485 -805
rect 4485 -835 4515 -805
rect 4515 -835 4516 -805
rect 4484 -836 4516 -835
rect 4484 -885 4516 -884
rect 4484 -915 4485 -885
rect 4485 -915 4515 -885
rect 4515 -915 4516 -885
rect 4484 -916 4516 -915
rect 4484 -996 4516 -964
rect 4484 -1076 4516 -1044
rect 4484 -1125 4516 -1124
rect 4484 -1155 4485 -1125
rect 4485 -1155 4515 -1125
rect 4515 -1155 4516 -1125
rect 4484 -1156 4516 -1155
rect 4484 -1205 4516 -1204
rect 4484 -1235 4485 -1205
rect 4485 -1235 4515 -1205
rect 4515 -1235 4516 -1205
rect 4484 -1236 4516 -1235
rect 4484 -1285 4516 -1284
rect 4484 -1315 4485 -1285
rect 4485 -1315 4515 -1285
rect 4515 -1315 4516 -1285
rect 4484 -1316 4516 -1315
rect 4484 -1365 4516 -1364
rect 4484 -1395 4485 -1365
rect 4485 -1395 4515 -1365
rect 4515 -1395 4516 -1365
rect 4484 -1396 4516 -1395
rect 4484 -1445 4516 -1444
rect 4484 -1475 4485 -1445
rect 4485 -1475 4515 -1445
rect 4515 -1475 4516 -1445
rect 4484 -1476 4516 -1475
rect 4484 -1525 4516 -1524
rect 4484 -1555 4485 -1525
rect 4485 -1555 4515 -1525
rect 4515 -1555 4516 -1525
rect 4484 -1556 4516 -1555
rect 4484 -1636 4516 -1604
rect 4484 -1716 4516 -1684
rect 4484 -1765 4516 -1764
rect 4484 -1795 4485 -1765
rect 4485 -1795 4515 -1765
rect 4515 -1795 4516 -1765
rect 4484 -1796 4516 -1795
rect 4484 -1845 4516 -1844
rect 4484 -1875 4485 -1845
rect 4485 -1875 4515 -1845
rect 4515 -1875 4516 -1845
rect 4484 -1876 4516 -1875
rect 4484 -1956 4516 -1924
rect 4484 -2005 4516 -2004
rect 4484 -2035 4485 -2005
rect 4485 -2035 4515 -2005
rect 4515 -2035 4516 -2005
rect 4484 -2036 4516 -2035
rect 4484 -2116 4516 -2084
rect 4484 -2165 4516 -2164
rect 4484 -2195 4485 -2165
rect 4485 -2195 4515 -2165
rect 4515 -2195 4516 -2165
rect 4484 -2196 4516 -2195
rect 4484 -2276 4516 -2244
rect 4484 -2325 4516 -2324
rect 4484 -2355 4485 -2325
rect 4485 -2355 4515 -2325
rect 4515 -2355 4516 -2325
rect 4484 -2356 4516 -2355
rect 4484 -2405 4516 -2404
rect 4484 -2435 4485 -2405
rect 4485 -2435 4515 -2405
rect 4515 -2435 4516 -2405
rect 4484 -2436 4516 -2435
rect 4484 -2485 4516 -2484
rect 4484 -2515 4485 -2485
rect 4485 -2515 4515 -2485
rect 4515 -2515 4516 -2485
rect 4484 -2516 4516 -2515
rect 4484 -2565 4516 -2564
rect 4484 -2595 4485 -2565
rect 4485 -2595 4515 -2565
rect 4515 -2595 4516 -2565
rect 4484 -2596 4516 -2595
rect 4484 -2645 4516 -2644
rect 4484 -2675 4485 -2645
rect 4485 -2675 4515 -2645
rect 4515 -2675 4516 -2645
rect 4484 -2676 4516 -2675
rect 4484 -2725 4516 -2724
rect 4484 -2755 4485 -2725
rect 4485 -2755 4515 -2725
rect 4515 -2755 4516 -2725
rect 4484 -2756 4516 -2755
rect 4484 -2836 4516 -2804
rect 4484 -2885 4516 -2884
rect 4484 -2915 4485 -2885
rect 4485 -2915 4515 -2885
rect 4515 -2915 4516 -2885
rect 4484 -2916 4516 -2915
rect 4484 -2996 4516 -2964
rect 4484 -3045 4516 -3044
rect 4484 -3075 4485 -3045
rect 4485 -3075 4515 -3045
rect 4515 -3075 4516 -3045
rect 4484 -3076 4516 -3075
rect 4484 -3156 4516 -3124
rect 4484 -3205 4516 -3204
rect 4484 -3235 4485 -3205
rect 4485 -3235 4515 -3205
rect 4515 -3235 4516 -3205
rect 4484 -3236 4516 -3235
rect 4484 -3285 4516 -3284
rect 4484 -3315 4485 -3285
rect 4485 -3315 4515 -3285
rect 4515 -3315 4516 -3285
rect 4484 -3316 4516 -3315
rect 4484 -3396 4516 -3364
rect 4484 -3476 4516 -3444
rect 4484 -3525 4516 -3524
rect 4484 -3555 4485 -3525
rect 4485 -3555 4515 -3525
rect 4515 -3555 4516 -3525
rect 4484 -3556 4516 -3555
rect 4484 -3605 4516 -3604
rect 4484 -3635 4485 -3605
rect 4485 -3635 4515 -3605
rect 4515 -3635 4516 -3605
rect 4484 -3636 4516 -3635
rect 4484 -3685 4516 -3684
rect 4484 -3715 4485 -3685
rect 4485 -3715 4515 -3685
rect 4515 -3715 4516 -3685
rect 4484 -3716 4516 -3715
rect 4564 1035 4596 1036
rect 4564 1005 4565 1035
rect 4565 1005 4595 1035
rect 4595 1005 4596 1035
rect 4564 1004 4596 1005
rect 4564 955 4596 956
rect 4564 925 4565 955
rect 4565 925 4595 955
rect 4595 925 4596 955
rect 4564 924 4596 925
rect 4564 875 4596 876
rect 4564 845 4565 875
rect 4565 845 4595 875
rect 4595 845 4596 875
rect 4564 844 4596 845
rect 4564 764 4596 796
rect 4564 684 4596 716
rect 4564 635 4596 636
rect 4564 605 4565 635
rect 4565 605 4595 635
rect 4595 605 4596 635
rect 4564 604 4596 605
rect 4564 555 4596 556
rect 4564 525 4565 555
rect 4565 525 4595 555
rect 4595 525 4596 555
rect 4564 524 4596 525
rect 4564 444 4596 476
rect 4564 395 4596 396
rect 4564 365 4565 395
rect 4565 365 4595 395
rect 4595 365 4596 395
rect 4564 364 4596 365
rect 4564 284 4596 316
rect 4564 235 4596 236
rect 4564 205 4565 235
rect 4565 205 4595 235
rect 4595 205 4596 235
rect 4564 204 4596 205
rect 4564 124 4596 156
rect 4564 75 4596 76
rect 4564 45 4565 75
rect 4565 45 4595 75
rect 4595 45 4596 75
rect 4564 44 4596 45
rect 4564 -5 4596 -4
rect 4564 -35 4565 -5
rect 4565 -35 4595 -5
rect 4595 -35 4596 -5
rect 4564 -36 4596 -35
rect 4564 -85 4596 -84
rect 4564 -115 4565 -85
rect 4565 -115 4595 -85
rect 4595 -115 4596 -85
rect 4564 -116 4596 -115
rect 4564 -165 4596 -164
rect 4564 -195 4565 -165
rect 4565 -195 4595 -165
rect 4595 -195 4596 -165
rect 4564 -196 4596 -195
rect 4564 -245 4596 -244
rect 4564 -275 4565 -245
rect 4565 -275 4595 -245
rect 4595 -275 4596 -245
rect 4564 -276 4596 -275
rect 4564 -325 4596 -324
rect 4564 -355 4565 -325
rect 4565 -355 4595 -325
rect 4595 -355 4596 -325
rect 4564 -356 4596 -355
rect 4564 -436 4596 -404
rect 4564 -485 4596 -484
rect 4564 -515 4565 -485
rect 4565 -515 4595 -485
rect 4595 -515 4596 -485
rect 4564 -516 4596 -515
rect 4564 -596 4596 -564
rect 4564 -645 4596 -644
rect 4564 -675 4565 -645
rect 4565 -675 4595 -645
rect 4595 -675 4596 -645
rect 4564 -676 4596 -675
rect 4564 -756 4596 -724
rect 4564 -805 4596 -804
rect 4564 -835 4565 -805
rect 4565 -835 4595 -805
rect 4595 -835 4596 -805
rect 4564 -836 4596 -835
rect 4564 -885 4596 -884
rect 4564 -915 4565 -885
rect 4565 -915 4595 -885
rect 4595 -915 4596 -885
rect 4564 -916 4596 -915
rect 4564 -996 4596 -964
rect 4564 -1076 4596 -1044
rect 4564 -1125 4596 -1124
rect 4564 -1155 4565 -1125
rect 4565 -1155 4595 -1125
rect 4595 -1155 4596 -1125
rect 4564 -1156 4596 -1155
rect 4564 -1205 4596 -1204
rect 4564 -1235 4565 -1205
rect 4565 -1235 4595 -1205
rect 4595 -1235 4596 -1205
rect 4564 -1236 4596 -1235
rect 4564 -1285 4596 -1284
rect 4564 -1315 4565 -1285
rect 4565 -1315 4595 -1285
rect 4595 -1315 4596 -1285
rect 4564 -1316 4596 -1315
rect 4564 -1365 4596 -1364
rect 4564 -1395 4565 -1365
rect 4565 -1395 4595 -1365
rect 4595 -1395 4596 -1365
rect 4564 -1396 4596 -1395
rect 4564 -1445 4596 -1444
rect 4564 -1475 4565 -1445
rect 4565 -1475 4595 -1445
rect 4595 -1475 4596 -1445
rect 4564 -1476 4596 -1475
rect 4564 -1525 4596 -1524
rect 4564 -1555 4565 -1525
rect 4565 -1555 4595 -1525
rect 4595 -1555 4596 -1525
rect 4564 -1556 4596 -1555
rect 4564 -1636 4596 -1604
rect 4564 -1716 4596 -1684
rect 4564 -1765 4596 -1764
rect 4564 -1795 4565 -1765
rect 4565 -1795 4595 -1765
rect 4595 -1795 4596 -1765
rect 4564 -1796 4596 -1795
rect 4564 -1845 4596 -1844
rect 4564 -1875 4565 -1845
rect 4565 -1875 4595 -1845
rect 4595 -1875 4596 -1845
rect 4564 -1876 4596 -1875
rect 4564 -1956 4596 -1924
rect 4564 -2005 4596 -2004
rect 4564 -2035 4565 -2005
rect 4565 -2035 4595 -2005
rect 4595 -2035 4596 -2005
rect 4564 -2036 4596 -2035
rect 4564 -2116 4596 -2084
rect 4564 -2165 4596 -2164
rect 4564 -2195 4565 -2165
rect 4565 -2195 4595 -2165
rect 4595 -2195 4596 -2165
rect 4564 -2196 4596 -2195
rect 4564 -2276 4596 -2244
rect 4564 -2325 4596 -2324
rect 4564 -2355 4565 -2325
rect 4565 -2355 4595 -2325
rect 4595 -2355 4596 -2325
rect 4564 -2356 4596 -2355
rect 4564 -2405 4596 -2404
rect 4564 -2435 4565 -2405
rect 4565 -2435 4595 -2405
rect 4595 -2435 4596 -2405
rect 4564 -2436 4596 -2435
rect 4564 -2485 4596 -2484
rect 4564 -2515 4565 -2485
rect 4565 -2515 4595 -2485
rect 4595 -2515 4596 -2485
rect 4564 -2516 4596 -2515
rect 4564 -2565 4596 -2564
rect 4564 -2595 4565 -2565
rect 4565 -2595 4595 -2565
rect 4595 -2595 4596 -2565
rect 4564 -2596 4596 -2595
rect 4564 -2645 4596 -2644
rect 4564 -2675 4565 -2645
rect 4565 -2675 4595 -2645
rect 4595 -2675 4596 -2645
rect 4564 -2676 4596 -2675
rect 4564 -2725 4596 -2724
rect 4564 -2755 4565 -2725
rect 4565 -2755 4595 -2725
rect 4595 -2755 4596 -2725
rect 4564 -2756 4596 -2755
rect 4564 -2836 4596 -2804
rect 4564 -2885 4596 -2884
rect 4564 -2915 4565 -2885
rect 4565 -2915 4595 -2885
rect 4595 -2915 4596 -2885
rect 4564 -2916 4596 -2915
rect 4564 -2996 4596 -2964
rect 4564 -3045 4596 -3044
rect 4564 -3075 4565 -3045
rect 4565 -3075 4595 -3045
rect 4595 -3075 4596 -3045
rect 4564 -3076 4596 -3075
rect 4564 -3156 4596 -3124
rect 4564 -3205 4596 -3204
rect 4564 -3235 4565 -3205
rect 4565 -3235 4595 -3205
rect 4595 -3235 4596 -3205
rect 4564 -3236 4596 -3235
rect 4564 -3285 4596 -3284
rect 4564 -3315 4565 -3285
rect 4565 -3315 4595 -3285
rect 4595 -3315 4596 -3285
rect 4564 -3316 4596 -3315
rect 4564 -3396 4596 -3364
rect 4564 -3476 4596 -3444
rect 4564 -3525 4596 -3524
rect 4564 -3555 4565 -3525
rect 4565 -3555 4595 -3525
rect 4595 -3555 4596 -3525
rect 4564 -3556 4596 -3555
rect 4564 -3605 4596 -3604
rect 4564 -3635 4565 -3605
rect 4565 -3635 4595 -3605
rect 4595 -3635 4596 -3605
rect 4564 -3636 4596 -3635
rect 4564 -3685 4596 -3684
rect 4564 -3715 4565 -3685
rect 4565 -3715 4595 -3685
rect 4595 -3715 4596 -3685
rect 4564 -3716 4596 -3715
rect 4644 1035 4676 1036
rect 4644 1005 4645 1035
rect 4645 1005 4675 1035
rect 4675 1005 4676 1035
rect 4644 1004 4676 1005
rect 4644 955 4676 956
rect 4644 925 4645 955
rect 4645 925 4675 955
rect 4675 925 4676 955
rect 4644 924 4676 925
rect 4644 875 4676 876
rect 4644 845 4645 875
rect 4645 845 4675 875
rect 4675 845 4676 875
rect 4644 844 4676 845
rect 4644 764 4676 796
rect 4644 684 4676 716
rect 4644 635 4676 636
rect 4644 605 4645 635
rect 4645 605 4675 635
rect 4675 605 4676 635
rect 4644 604 4676 605
rect 4644 555 4676 556
rect 4644 525 4645 555
rect 4645 525 4675 555
rect 4675 525 4676 555
rect 4644 524 4676 525
rect 4644 444 4676 476
rect 4644 395 4676 396
rect 4644 365 4645 395
rect 4645 365 4675 395
rect 4675 365 4676 395
rect 4644 364 4676 365
rect 4644 284 4676 316
rect 4644 235 4676 236
rect 4644 205 4645 235
rect 4645 205 4675 235
rect 4675 205 4676 235
rect 4644 204 4676 205
rect 4644 124 4676 156
rect 4644 75 4676 76
rect 4644 45 4645 75
rect 4645 45 4675 75
rect 4675 45 4676 75
rect 4644 44 4676 45
rect 4644 -5 4676 -4
rect 4644 -35 4645 -5
rect 4645 -35 4675 -5
rect 4675 -35 4676 -5
rect 4644 -36 4676 -35
rect 4644 -85 4676 -84
rect 4644 -115 4645 -85
rect 4645 -115 4675 -85
rect 4675 -115 4676 -85
rect 4644 -116 4676 -115
rect 4644 -165 4676 -164
rect 4644 -195 4645 -165
rect 4645 -195 4675 -165
rect 4675 -195 4676 -165
rect 4644 -196 4676 -195
rect 4644 -245 4676 -244
rect 4644 -275 4645 -245
rect 4645 -275 4675 -245
rect 4675 -275 4676 -245
rect 4644 -276 4676 -275
rect 4644 -325 4676 -324
rect 4644 -355 4645 -325
rect 4645 -355 4675 -325
rect 4675 -355 4676 -325
rect 4644 -356 4676 -355
rect 4644 -436 4676 -404
rect 4644 -485 4676 -484
rect 4644 -515 4645 -485
rect 4645 -515 4675 -485
rect 4675 -515 4676 -485
rect 4644 -516 4676 -515
rect 4644 -596 4676 -564
rect 4644 -645 4676 -644
rect 4644 -675 4645 -645
rect 4645 -675 4675 -645
rect 4675 -675 4676 -645
rect 4644 -676 4676 -675
rect 4644 -756 4676 -724
rect 4644 -805 4676 -804
rect 4644 -835 4645 -805
rect 4645 -835 4675 -805
rect 4675 -835 4676 -805
rect 4644 -836 4676 -835
rect 4644 -885 4676 -884
rect 4644 -915 4645 -885
rect 4645 -915 4675 -885
rect 4675 -915 4676 -885
rect 4644 -916 4676 -915
rect 4644 -996 4676 -964
rect 4644 -1076 4676 -1044
rect 4644 -1125 4676 -1124
rect 4644 -1155 4645 -1125
rect 4645 -1155 4675 -1125
rect 4675 -1155 4676 -1125
rect 4644 -1156 4676 -1155
rect 4644 -1205 4676 -1204
rect 4644 -1235 4645 -1205
rect 4645 -1235 4675 -1205
rect 4675 -1235 4676 -1205
rect 4644 -1236 4676 -1235
rect 4644 -1285 4676 -1284
rect 4644 -1315 4645 -1285
rect 4645 -1315 4675 -1285
rect 4675 -1315 4676 -1285
rect 4644 -1316 4676 -1315
rect 4644 -1365 4676 -1364
rect 4644 -1395 4645 -1365
rect 4645 -1395 4675 -1365
rect 4675 -1395 4676 -1365
rect 4644 -1396 4676 -1395
rect 4644 -1445 4676 -1444
rect 4644 -1475 4645 -1445
rect 4645 -1475 4675 -1445
rect 4675 -1475 4676 -1445
rect 4644 -1476 4676 -1475
rect 4644 -1525 4676 -1524
rect 4644 -1555 4645 -1525
rect 4645 -1555 4675 -1525
rect 4675 -1555 4676 -1525
rect 4644 -1556 4676 -1555
rect 4644 -1636 4676 -1604
rect 4644 -1716 4676 -1684
rect 4644 -1765 4676 -1764
rect 4644 -1795 4645 -1765
rect 4645 -1795 4675 -1765
rect 4675 -1795 4676 -1765
rect 4644 -1796 4676 -1795
rect 4644 -1845 4676 -1844
rect 4644 -1875 4645 -1845
rect 4645 -1875 4675 -1845
rect 4675 -1875 4676 -1845
rect 4644 -1876 4676 -1875
rect 4644 -1956 4676 -1924
rect 4644 -2005 4676 -2004
rect 4644 -2035 4645 -2005
rect 4645 -2035 4675 -2005
rect 4675 -2035 4676 -2005
rect 4644 -2036 4676 -2035
rect 4644 -2116 4676 -2084
rect 4644 -2165 4676 -2164
rect 4644 -2195 4645 -2165
rect 4645 -2195 4675 -2165
rect 4675 -2195 4676 -2165
rect 4644 -2196 4676 -2195
rect 4644 -2276 4676 -2244
rect 4644 -2325 4676 -2324
rect 4644 -2355 4645 -2325
rect 4645 -2355 4675 -2325
rect 4675 -2355 4676 -2325
rect 4644 -2356 4676 -2355
rect 4644 -2405 4676 -2404
rect 4644 -2435 4645 -2405
rect 4645 -2435 4675 -2405
rect 4675 -2435 4676 -2405
rect 4644 -2436 4676 -2435
rect 4644 -2485 4676 -2484
rect 4644 -2515 4645 -2485
rect 4645 -2515 4675 -2485
rect 4675 -2515 4676 -2485
rect 4644 -2516 4676 -2515
rect 4644 -2565 4676 -2564
rect 4644 -2595 4645 -2565
rect 4645 -2595 4675 -2565
rect 4675 -2595 4676 -2565
rect 4644 -2596 4676 -2595
rect 4644 -2645 4676 -2644
rect 4644 -2675 4645 -2645
rect 4645 -2675 4675 -2645
rect 4675 -2675 4676 -2645
rect 4644 -2676 4676 -2675
rect 4644 -2725 4676 -2724
rect 4644 -2755 4645 -2725
rect 4645 -2755 4675 -2725
rect 4675 -2755 4676 -2725
rect 4644 -2756 4676 -2755
rect 4644 -2836 4676 -2804
rect 4644 -2885 4676 -2884
rect 4644 -2915 4645 -2885
rect 4645 -2915 4675 -2885
rect 4675 -2915 4676 -2885
rect 4644 -2916 4676 -2915
rect 4644 -2996 4676 -2964
rect 4644 -3045 4676 -3044
rect 4644 -3075 4645 -3045
rect 4645 -3075 4675 -3045
rect 4675 -3075 4676 -3045
rect 4644 -3076 4676 -3075
rect 4644 -3156 4676 -3124
rect 4644 -3205 4676 -3204
rect 4644 -3235 4645 -3205
rect 4645 -3235 4675 -3205
rect 4675 -3235 4676 -3205
rect 4644 -3236 4676 -3235
rect 4644 -3285 4676 -3284
rect 4644 -3315 4645 -3285
rect 4645 -3315 4675 -3285
rect 4675 -3315 4676 -3285
rect 4644 -3316 4676 -3315
rect 4644 -3396 4676 -3364
rect 4644 -3476 4676 -3444
rect 4644 -3525 4676 -3524
rect 4644 -3555 4645 -3525
rect 4645 -3555 4675 -3525
rect 4675 -3555 4676 -3525
rect 4644 -3556 4676 -3555
rect 4644 -3605 4676 -3604
rect 4644 -3635 4645 -3605
rect 4645 -3635 4675 -3605
rect 4675 -3635 4676 -3605
rect 4644 -3636 4676 -3635
rect 4644 -3685 4676 -3684
rect 4644 -3715 4645 -3685
rect 4645 -3715 4675 -3685
rect 4675 -3715 4676 -3685
rect 4644 -3716 4676 -3715
rect 4724 1035 4756 1036
rect 4724 1005 4725 1035
rect 4725 1005 4755 1035
rect 4755 1005 4756 1035
rect 4724 1004 4756 1005
rect 4724 955 4756 956
rect 4724 925 4725 955
rect 4725 925 4755 955
rect 4755 925 4756 955
rect 4724 924 4756 925
rect 4724 875 4756 876
rect 4724 845 4725 875
rect 4725 845 4755 875
rect 4755 845 4756 875
rect 4724 844 4756 845
rect 4724 764 4756 796
rect 4724 684 4756 716
rect 4724 635 4756 636
rect 4724 605 4725 635
rect 4725 605 4755 635
rect 4755 605 4756 635
rect 4724 604 4756 605
rect 4724 555 4756 556
rect 4724 525 4725 555
rect 4725 525 4755 555
rect 4755 525 4756 555
rect 4724 524 4756 525
rect 4724 444 4756 476
rect 4724 395 4756 396
rect 4724 365 4725 395
rect 4725 365 4755 395
rect 4755 365 4756 395
rect 4724 364 4756 365
rect 4724 284 4756 316
rect 4724 235 4756 236
rect 4724 205 4725 235
rect 4725 205 4755 235
rect 4755 205 4756 235
rect 4724 204 4756 205
rect 4724 124 4756 156
rect 4724 75 4756 76
rect 4724 45 4725 75
rect 4725 45 4755 75
rect 4755 45 4756 75
rect 4724 44 4756 45
rect 4724 -5 4756 -4
rect 4724 -35 4725 -5
rect 4725 -35 4755 -5
rect 4755 -35 4756 -5
rect 4724 -36 4756 -35
rect 4724 -85 4756 -84
rect 4724 -115 4725 -85
rect 4725 -115 4755 -85
rect 4755 -115 4756 -85
rect 4724 -116 4756 -115
rect 4724 -165 4756 -164
rect 4724 -195 4725 -165
rect 4725 -195 4755 -165
rect 4755 -195 4756 -165
rect 4724 -196 4756 -195
rect 4724 -245 4756 -244
rect 4724 -275 4725 -245
rect 4725 -275 4755 -245
rect 4755 -275 4756 -245
rect 4724 -276 4756 -275
rect 4724 -325 4756 -324
rect 4724 -355 4725 -325
rect 4725 -355 4755 -325
rect 4755 -355 4756 -325
rect 4724 -356 4756 -355
rect 4724 -436 4756 -404
rect 4724 -485 4756 -484
rect 4724 -515 4725 -485
rect 4725 -515 4755 -485
rect 4755 -515 4756 -485
rect 4724 -516 4756 -515
rect 4724 -596 4756 -564
rect 4724 -645 4756 -644
rect 4724 -675 4725 -645
rect 4725 -675 4755 -645
rect 4755 -675 4756 -645
rect 4724 -676 4756 -675
rect 4724 -756 4756 -724
rect 4724 -805 4756 -804
rect 4724 -835 4725 -805
rect 4725 -835 4755 -805
rect 4755 -835 4756 -805
rect 4724 -836 4756 -835
rect 4724 -885 4756 -884
rect 4724 -915 4725 -885
rect 4725 -915 4755 -885
rect 4755 -915 4756 -885
rect 4724 -916 4756 -915
rect 4724 -996 4756 -964
rect 4724 -1076 4756 -1044
rect 4724 -1125 4756 -1124
rect 4724 -1155 4725 -1125
rect 4725 -1155 4755 -1125
rect 4755 -1155 4756 -1125
rect 4724 -1156 4756 -1155
rect 4724 -1205 4756 -1204
rect 4724 -1235 4725 -1205
rect 4725 -1235 4755 -1205
rect 4755 -1235 4756 -1205
rect 4724 -1236 4756 -1235
rect 4724 -1285 4756 -1284
rect 4724 -1315 4725 -1285
rect 4725 -1315 4755 -1285
rect 4755 -1315 4756 -1285
rect 4724 -1316 4756 -1315
rect 4724 -1365 4756 -1364
rect 4724 -1395 4725 -1365
rect 4725 -1395 4755 -1365
rect 4755 -1395 4756 -1365
rect 4724 -1396 4756 -1395
rect 4724 -1445 4756 -1444
rect 4724 -1475 4725 -1445
rect 4725 -1475 4755 -1445
rect 4755 -1475 4756 -1445
rect 4724 -1476 4756 -1475
rect 4724 -1525 4756 -1524
rect 4724 -1555 4725 -1525
rect 4725 -1555 4755 -1525
rect 4755 -1555 4756 -1525
rect 4724 -1556 4756 -1555
rect 4724 -1636 4756 -1604
rect 4724 -1716 4756 -1684
rect 4724 -1765 4756 -1764
rect 4724 -1795 4725 -1765
rect 4725 -1795 4755 -1765
rect 4755 -1795 4756 -1765
rect 4724 -1796 4756 -1795
rect 4724 -1845 4756 -1844
rect 4724 -1875 4725 -1845
rect 4725 -1875 4755 -1845
rect 4755 -1875 4756 -1845
rect 4724 -1876 4756 -1875
rect 4724 -1956 4756 -1924
rect 4724 -2005 4756 -2004
rect 4724 -2035 4725 -2005
rect 4725 -2035 4755 -2005
rect 4755 -2035 4756 -2005
rect 4724 -2036 4756 -2035
rect 4724 -2116 4756 -2084
rect 4724 -2165 4756 -2164
rect 4724 -2195 4725 -2165
rect 4725 -2195 4755 -2165
rect 4755 -2195 4756 -2165
rect 4724 -2196 4756 -2195
rect 4724 -2276 4756 -2244
rect 4724 -2325 4756 -2324
rect 4724 -2355 4725 -2325
rect 4725 -2355 4755 -2325
rect 4755 -2355 4756 -2325
rect 4724 -2356 4756 -2355
rect 4724 -2405 4756 -2404
rect 4724 -2435 4725 -2405
rect 4725 -2435 4755 -2405
rect 4755 -2435 4756 -2405
rect 4724 -2436 4756 -2435
rect 4724 -2485 4756 -2484
rect 4724 -2515 4725 -2485
rect 4725 -2515 4755 -2485
rect 4755 -2515 4756 -2485
rect 4724 -2516 4756 -2515
rect 4724 -2565 4756 -2564
rect 4724 -2595 4725 -2565
rect 4725 -2595 4755 -2565
rect 4755 -2595 4756 -2565
rect 4724 -2596 4756 -2595
rect 4724 -2645 4756 -2644
rect 4724 -2675 4725 -2645
rect 4725 -2675 4755 -2645
rect 4755 -2675 4756 -2645
rect 4724 -2676 4756 -2675
rect 4724 -2725 4756 -2724
rect 4724 -2755 4725 -2725
rect 4725 -2755 4755 -2725
rect 4755 -2755 4756 -2725
rect 4724 -2756 4756 -2755
rect 4724 -2836 4756 -2804
rect 4724 -2885 4756 -2884
rect 4724 -2915 4725 -2885
rect 4725 -2915 4755 -2885
rect 4755 -2915 4756 -2885
rect 4724 -2916 4756 -2915
rect 4724 -2996 4756 -2964
rect 4724 -3045 4756 -3044
rect 4724 -3075 4725 -3045
rect 4725 -3075 4755 -3045
rect 4755 -3075 4756 -3045
rect 4724 -3076 4756 -3075
rect 4724 -3156 4756 -3124
rect 4724 -3205 4756 -3204
rect 4724 -3235 4725 -3205
rect 4725 -3235 4755 -3205
rect 4755 -3235 4756 -3205
rect 4724 -3236 4756 -3235
rect 4724 -3285 4756 -3284
rect 4724 -3315 4725 -3285
rect 4725 -3315 4755 -3285
rect 4755 -3315 4756 -3285
rect 4724 -3316 4756 -3315
rect 4724 -3396 4756 -3364
rect 4724 -3476 4756 -3444
rect 4724 -3525 4756 -3524
rect 4724 -3555 4725 -3525
rect 4725 -3555 4755 -3525
rect 4755 -3555 4756 -3525
rect 4724 -3556 4756 -3555
rect 4724 -3605 4756 -3604
rect 4724 -3635 4725 -3605
rect 4725 -3635 4755 -3605
rect 4755 -3635 4756 -3605
rect 4724 -3636 4756 -3635
rect 4724 -3685 4756 -3684
rect 4724 -3715 4725 -3685
rect 4725 -3715 4755 -3685
rect 4755 -3715 4756 -3685
rect 4724 -3716 4756 -3715
rect 4804 1035 4836 1036
rect 4804 1005 4805 1035
rect 4805 1005 4835 1035
rect 4835 1005 4836 1035
rect 4804 1004 4836 1005
rect 4804 955 4836 956
rect 4804 925 4805 955
rect 4805 925 4835 955
rect 4835 925 4836 955
rect 4804 924 4836 925
rect 4804 875 4836 876
rect 4804 845 4805 875
rect 4805 845 4835 875
rect 4835 845 4836 875
rect 4804 844 4836 845
rect 4804 764 4836 796
rect 4804 684 4836 716
rect 4804 635 4836 636
rect 4804 605 4805 635
rect 4805 605 4835 635
rect 4835 605 4836 635
rect 4804 604 4836 605
rect 4804 555 4836 556
rect 4804 525 4805 555
rect 4805 525 4835 555
rect 4835 525 4836 555
rect 4804 524 4836 525
rect 4804 444 4836 476
rect 4804 395 4836 396
rect 4804 365 4805 395
rect 4805 365 4835 395
rect 4835 365 4836 395
rect 4804 364 4836 365
rect 4804 284 4836 316
rect 4804 235 4836 236
rect 4804 205 4805 235
rect 4805 205 4835 235
rect 4835 205 4836 235
rect 4804 204 4836 205
rect 4804 124 4836 156
rect 4804 75 4836 76
rect 4804 45 4805 75
rect 4805 45 4835 75
rect 4835 45 4836 75
rect 4804 44 4836 45
rect 4804 -5 4836 -4
rect 4804 -35 4805 -5
rect 4805 -35 4835 -5
rect 4835 -35 4836 -5
rect 4804 -36 4836 -35
rect 4804 -85 4836 -84
rect 4804 -115 4805 -85
rect 4805 -115 4835 -85
rect 4835 -115 4836 -85
rect 4804 -116 4836 -115
rect 4804 -165 4836 -164
rect 4804 -195 4805 -165
rect 4805 -195 4835 -165
rect 4835 -195 4836 -165
rect 4804 -196 4836 -195
rect 4804 -245 4836 -244
rect 4804 -275 4805 -245
rect 4805 -275 4835 -245
rect 4835 -275 4836 -245
rect 4804 -276 4836 -275
rect 4804 -325 4836 -324
rect 4804 -355 4805 -325
rect 4805 -355 4835 -325
rect 4835 -355 4836 -325
rect 4804 -356 4836 -355
rect 4804 -436 4836 -404
rect 4804 -485 4836 -484
rect 4804 -515 4805 -485
rect 4805 -515 4835 -485
rect 4835 -515 4836 -485
rect 4804 -516 4836 -515
rect 4804 -596 4836 -564
rect 4804 -645 4836 -644
rect 4804 -675 4805 -645
rect 4805 -675 4835 -645
rect 4835 -675 4836 -645
rect 4804 -676 4836 -675
rect 4804 -756 4836 -724
rect 4804 -805 4836 -804
rect 4804 -835 4805 -805
rect 4805 -835 4835 -805
rect 4835 -835 4836 -805
rect 4804 -836 4836 -835
rect 4804 -885 4836 -884
rect 4804 -915 4805 -885
rect 4805 -915 4835 -885
rect 4835 -915 4836 -885
rect 4804 -916 4836 -915
rect 4804 -996 4836 -964
rect 4804 -1076 4836 -1044
rect 4804 -1125 4836 -1124
rect 4804 -1155 4805 -1125
rect 4805 -1155 4835 -1125
rect 4835 -1155 4836 -1125
rect 4804 -1156 4836 -1155
rect 4804 -1205 4836 -1204
rect 4804 -1235 4805 -1205
rect 4805 -1235 4835 -1205
rect 4835 -1235 4836 -1205
rect 4804 -1236 4836 -1235
rect 4804 -1285 4836 -1284
rect 4804 -1315 4805 -1285
rect 4805 -1315 4835 -1285
rect 4835 -1315 4836 -1285
rect 4804 -1316 4836 -1315
rect 4804 -1365 4836 -1364
rect 4804 -1395 4805 -1365
rect 4805 -1395 4835 -1365
rect 4835 -1395 4836 -1365
rect 4804 -1396 4836 -1395
rect 4804 -1445 4836 -1444
rect 4804 -1475 4805 -1445
rect 4805 -1475 4835 -1445
rect 4835 -1475 4836 -1445
rect 4804 -1476 4836 -1475
rect 4804 -1525 4836 -1524
rect 4804 -1555 4805 -1525
rect 4805 -1555 4835 -1525
rect 4835 -1555 4836 -1525
rect 4804 -1556 4836 -1555
rect 4804 -1636 4836 -1604
rect 4804 -1716 4836 -1684
rect 4804 -1765 4836 -1764
rect 4804 -1795 4805 -1765
rect 4805 -1795 4835 -1765
rect 4835 -1795 4836 -1765
rect 4804 -1796 4836 -1795
rect 4804 -1845 4836 -1844
rect 4804 -1875 4805 -1845
rect 4805 -1875 4835 -1845
rect 4835 -1875 4836 -1845
rect 4804 -1876 4836 -1875
rect 4804 -1956 4836 -1924
rect 4804 -2005 4836 -2004
rect 4804 -2035 4805 -2005
rect 4805 -2035 4835 -2005
rect 4835 -2035 4836 -2005
rect 4804 -2036 4836 -2035
rect 4804 -2116 4836 -2084
rect 4804 -2165 4836 -2164
rect 4804 -2195 4805 -2165
rect 4805 -2195 4835 -2165
rect 4835 -2195 4836 -2165
rect 4804 -2196 4836 -2195
rect 4804 -2276 4836 -2244
rect 4804 -2325 4836 -2324
rect 4804 -2355 4805 -2325
rect 4805 -2355 4835 -2325
rect 4835 -2355 4836 -2325
rect 4804 -2356 4836 -2355
rect 4804 -2405 4836 -2404
rect 4804 -2435 4805 -2405
rect 4805 -2435 4835 -2405
rect 4835 -2435 4836 -2405
rect 4804 -2436 4836 -2435
rect 4804 -2485 4836 -2484
rect 4804 -2515 4805 -2485
rect 4805 -2515 4835 -2485
rect 4835 -2515 4836 -2485
rect 4804 -2516 4836 -2515
rect 4804 -2565 4836 -2564
rect 4804 -2595 4805 -2565
rect 4805 -2595 4835 -2565
rect 4835 -2595 4836 -2565
rect 4804 -2596 4836 -2595
rect 4804 -2645 4836 -2644
rect 4804 -2675 4805 -2645
rect 4805 -2675 4835 -2645
rect 4835 -2675 4836 -2645
rect 4804 -2676 4836 -2675
rect 4804 -2725 4836 -2724
rect 4804 -2755 4805 -2725
rect 4805 -2755 4835 -2725
rect 4835 -2755 4836 -2725
rect 4804 -2756 4836 -2755
rect 4804 -2836 4836 -2804
rect 4804 -2885 4836 -2884
rect 4804 -2915 4805 -2885
rect 4805 -2915 4835 -2885
rect 4835 -2915 4836 -2885
rect 4804 -2916 4836 -2915
rect 4804 -2996 4836 -2964
rect 4804 -3045 4836 -3044
rect 4804 -3075 4805 -3045
rect 4805 -3075 4835 -3045
rect 4835 -3075 4836 -3045
rect 4804 -3076 4836 -3075
rect 4804 -3156 4836 -3124
rect 4804 -3205 4836 -3204
rect 4804 -3235 4805 -3205
rect 4805 -3235 4835 -3205
rect 4835 -3235 4836 -3205
rect 4804 -3236 4836 -3235
rect 4804 -3285 4836 -3284
rect 4804 -3315 4805 -3285
rect 4805 -3315 4835 -3285
rect 4835 -3315 4836 -3285
rect 4804 -3316 4836 -3315
rect 4804 -3396 4836 -3364
rect 4804 -3476 4836 -3444
rect 4804 -3525 4836 -3524
rect 4804 -3555 4805 -3525
rect 4805 -3555 4835 -3525
rect 4835 -3555 4836 -3525
rect 4804 -3556 4836 -3555
rect 4804 -3605 4836 -3604
rect 4804 -3635 4805 -3605
rect 4805 -3635 4835 -3605
rect 4835 -3635 4836 -3605
rect 4804 -3636 4836 -3635
rect 4804 -3685 4836 -3684
rect 4804 -3715 4805 -3685
rect 4805 -3715 4835 -3685
rect 4835 -3715 4836 -3685
rect 4804 -3716 4836 -3715
rect 4884 1035 4916 1036
rect 4884 1005 4885 1035
rect 4885 1005 4915 1035
rect 4915 1005 4916 1035
rect 4884 1004 4916 1005
rect 4884 955 4916 956
rect 4884 925 4885 955
rect 4885 925 4915 955
rect 4915 925 4916 955
rect 4884 924 4916 925
rect 4884 875 4916 876
rect 4884 845 4885 875
rect 4885 845 4915 875
rect 4915 845 4916 875
rect 4884 844 4916 845
rect 4884 764 4916 796
rect 4884 684 4916 716
rect 4884 635 4916 636
rect 4884 605 4885 635
rect 4885 605 4915 635
rect 4915 605 4916 635
rect 4884 604 4916 605
rect 4884 555 4916 556
rect 4884 525 4885 555
rect 4885 525 4915 555
rect 4915 525 4916 555
rect 4884 524 4916 525
rect 4884 444 4916 476
rect 4884 395 4916 396
rect 4884 365 4885 395
rect 4885 365 4915 395
rect 4915 365 4916 395
rect 4884 364 4916 365
rect 4884 284 4916 316
rect 4884 235 4916 236
rect 4884 205 4885 235
rect 4885 205 4915 235
rect 4915 205 4916 235
rect 4884 204 4916 205
rect 4884 124 4916 156
rect 4884 75 4916 76
rect 4884 45 4885 75
rect 4885 45 4915 75
rect 4915 45 4916 75
rect 4884 44 4916 45
rect 4884 -5 4916 -4
rect 4884 -35 4885 -5
rect 4885 -35 4915 -5
rect 4915 -35 4916 -5
rect 4884 -36 4916 -35
rect 4884 -85 4916 -84
rect 4884 -115 4885 -85
rect 4885 -115 4915 -85
rect 4915 -115 4916 -85
rect 4884 -116 4916 -115
rect 4884 -165 4916 -164
rect 4884 -195 4885 -165
rect 4885 -195 4915 -165
rect 4915 -195 4916 -165
rect 4884 -196 4916 -195
rect 4884 -245 4916 -244
rect 4884 -275 4885 -245
rect 4885 -275 4915 -245
rect 4915 -275 4916 -245
rect 4884 -276 4916 -275
rect 4884 -325 4916 -324
rect 4884 -355 4885 -325
rect 4885 -355 4915 -325
rect 4915 -355 4916 -325
rect 4884 -356 4916 -355
rect 4884 -436 4916 -404
rect 4884 -485 4916 -484
rect 4884 -515 4885 -485
rect 4885 -515 4915 -485
rect 4915 -515 4916 -485
rect 4884 -516 4916 -515
rect 4884 -596 4916 -564
rect 4884 -645 4916 -644
rect 4884 -675 4885 -645
rect 4885 -675 4915 -645
rect 4915 -675 4916 -645
rect 4884 -676 4916 -675
rect 4884 -756 4916 -724
rect 4884 -805 4916 -804
rect 4884 -835 4885 -805
rect 4885 -835 4915 -805
rect 4915 -835 4916 -805
rect 4884 -836 4916 -835
rect 4884 -885 4916 -884
rect 4884 -915 4885 -885
rect 4885 -915 4915 -885
rect 4915 -915 4916 -885
rect 4884 -916 4916 -915
rect 4884 -996 4916 -964
rect 4884 -1076 4916 -1044
rect 4884 -1125 4916 -1124
rect 4884 -1155 4885 -1125
rect 4885 -1155 4915 -1125
rect 4915 -1155 4916 -1125
rect 4884 -1156 4916 -1155
rect 4884 -1205 4916 -1204
rect 4884 -1235 4885 -1205
rect 4885 -1235 4915 -1205
rect 4915 -1235 4916 -1205
rect 4884 -1236 4916 -1235
rect 4884 -1285 4916 -1284
rect 4884 -1315 4885 -1285
rect 4885 -1315 4915 -1285
rect 4915 -1315 4916 -1285
rect 4884 -1316 4916 -1315
rect 4884 -1365 4916 -1364
rect 4884 -1395 4885 -1365
rect 4885 -1395 4915 -1365
rect 4915 -1395 4916 -1365
rect 4884 -1396 4916 -1395
rect 4884 -1445 4916 -1444
rect 4884 -1475 4885 -1445
rect 4885 -1475 4915 -1445
rect 4915 -1475 4916 -1445
rect 4884 -1476 4916 -1475
rect 4884 -1525 4916 -1524
rect 4884 -1555 4885 -1525
rect 4885 -1555 4915 -1525
rect 4915 -1555 4916 -1525
rect 4884 -1556 4916 -1555
rect 4884 -1636 4916 -1604
rect 4884 -1716 4916 -1684
rect 4884 -1765 4916 -1764
rect 4884 -1795 4885 -1765
rect 4885 -1795 4915 -1765
rect 4915 -1795 4916 -1765
rect 4884 -1796 4916 -1795
rect 4884 -1845 4916 -1844
rect 4884 -1875 4885 -1845
rect 4885 -1875 4915 -1845
rect 4915 -1875 4916 -1845
rect 4884 -1876 4916 -1875
rect 4884 -1956 4916 -1924
rect 4884 -2005 4916 -2004
rect 4884 -2035 4885 -2005
rect 4885 -2035 4915 -2005
rect 4915 -2035 4916 -2005
rect 4884 -2036 4916 -2035
rect 4884 -2116 4916 -2084
rect 4884 -2165 4916 -2164
rect 4884 -2195 4885 -2165
rect 4885 -2195 4915 -2165
rect 4915 -2195 4916 -2165
rect 4884 -2196 4916 -2195
rect 4884 -2276 4916 -2244
rect 4884 -2325 4916 -2324
rect 4884 -2355 4885 -2325
rect 4885 -2355 4915 -2325
rect 4915 -2355 4916 -2325
rect 4884 -2356 4916 -2355
rect 4884 -2405 4916 -2404
rect 4884 -2435 4885 -2405
rect 4885 -2435 4915 -2405
rect 4915 -2435 4916 -2405
rect 4884 -2436 4916 -2435
rect 4884 -2485 4916 -2484
rect 4884 -2515 4885 -2485
rect 4885 -2515 4915 -2485
rect 4915 -2515 4916 -2485
rect 4884 -2516 4916 -2515
rect 4884 -2565 4916 -2564
rect 4884 -2595 4885 -2565
rect 4885 -2595 4915 -2565
rect 4915 -2595 4916 -2565
rect 4884 -2596 4916 -2595
rect 4884 -2645 4916 -2644
rect 4884 -2675 4885 -2645
rect 4885 -2675 4915 -2645
rect 4915 -2675 4916 -2645
rect 4884 -2676 4916 -2675
rect 4884 -2725 4916 -2724
rect 4884 -2755 4885 -2725
rect 4885 -2755 4915 -2725
rect 4915 -2755 4916 -2725
rect 4884 -2756 4916 -2755
rect 4884 -2836 4916 -2804
rect 4884 -2885 4916 -2884
rect 4884 -2915 4885 -2885
rect 4885 -2915 4915 -2885
rect 4915 -2915 4916 -2885
rect 4884 -2916 4916 -2915
rect 4884 -2996 4916 -2964
rect 4884 -3045 4916 -3044
rect 4884 -3075 4885 -3045
rect 4885 -3075 4915 -3045
rect 4915 -3075 4916 -3045
rect 4884 -3076 4916 -3075
rect 4884 -3156 4916 -3124
rect 4884 -3205 4916 -3204
rect 4884 -3235 4885 -3205
rect 4885 -3235 4915 -3205
rect 4915 -3235 4916 -3205
rect 4884 -3236 4916 -3235
rect 4884 -3285 4916 -3284
rect 4884 -3315 4885 -3285
rect 4885 -3315 4915 -3285
rect 4915 -3315 4916 -3285
rect 4884 -3316 4916 -3315
rect 4884 -3396 4916 -3364
rect 4884 -3476 4916 -3444
rect 4884 -3525 4916 -3524
rect 4884 -3555 4885 -3525
rect 4885 -3555 4915 -3525
rect 4915 -3555 4916 -3525
rect 4884 -3556 4916 -3555
rect 4884 -3605 4916 -3604
rect 4884 -3635 4885 -3605
rect 4885 -3635 4915 -3605
rect 4915 -3635 4916 -3605
rect 4884 -3636 4916 -3635
rect 4884 -3685 4916 -3684
rect 4884 -3715 4885 -3685
rect 4885 -3715 4915 -3685
rect 4915 -3715 4916 -3685
rect 4884 -3716 4916 -3715
rect 4964 1035 4996 1036
rect 4964 1005 4965 1035
rect 4965 1005 4995 1035
rect 4995 1005 4996 1035
rect 4964 1004 4996 1005
rect 4964 955 4996 956
rect 4964 925 4965 955
rect 4965 925 4995 955
rect 4995 925 4996 955
rect 4964 924 4996 925
rect 4964 875 4996 876
rect 4964 845 4965 875
rect 4965 845 4995 875
rect 4995 845 4996 875
rect 4964 844 4996 845
rect 4964 764 4996 796
rect 4964 684 4996 716
rect 4964 635 4996 636
rect 4964 605 4965 635
rect 4965 605 4995 635
rect 4995 605 4996 635
rect 4964 604 4996 605
rect 4964 555 4996 556
rect 4964 525 4965 555
rect 4965 525 4995 555
rect 4995 525 4996 555
rect 4964 524 4996 525
rect 4964 444 4996 476
rect 4964 395 4996 396
rect 4964 365 4965 395
rect 4965 365 4995 395
rect 4995 365 4996 395
rect 4964 364 4996 365
rect 4964 284 4996 316
rect 4964 235 4996 236
rect 4964 205 4965 235
rect 4965 205 4995 235
rect 4995 205 4996 235
rect 4964 204 4996 205
rect 4964 124 4996 156
rect 4964 75 4996 76
rect 4964 45 4965 75
rect 4965 45 4995 75
rect 4995 45 4996 75
rect 4964 44 4996 45
rect 4964 -5 4996 -4
rect 4964 -35 4965 -5
rect 4965 -35 4995 -5
rect 4995 -35 4996 -5
rect 4964 -36 4996 -35
rect 4964 -85 4996 -84
rect 4964 -115 4965 -85
rect 4965 -115 4995 -85
rect 4995 -115 4996 -85
rect 4964 -116 4996 -115
rect 4964 -165 4996 -164
rect 4964 -195 4965 -165
rect 4965 -195 4995 -165
rect 4995 -195 4996 -165
rect 4964 -196 4996 -195
rect 4964 -245 4996 -244
rect 4964 -275 4965 -245
rect 4965 -275 4995 -245
rect 4995 -275 4996 -245
rect 4964 -276 4996 -275
rect 4964 -325 4996 -324
rect 4964 -355 4965 -325
rect 4965 -355 4995 -325
rect 4995 -355 4996 -325
rect 4964 -356 4996 -355
rect 4964 -436 4996 -404
rect 4964 -485 4996 -484
rect 4964 -515 4965 -485
rect 4965 -515 4995 -485
rect 4995 -515 4996 -485
rect 4964 -516 4996 -515
rect 4964 -596 4996 -564
rect 4964 -645 4996 -644
rect 4964 -675 4965 -645
rect 4965 -675 4995 -645
rect 4995 -675 4996 -645
rect 4964 -676 4996 -675
rect 4964 -756 4996 -724
rect 4964 -805 4996 -804
rect 4964 -835 4965 -805
rect 4965 -835 4995 -805
rect 4995 -835 4996 -805
rect 4964 -836 4996 -835
rect 4964 -885 4996 -884
rect 4964 -915 4965 -885
rect 4965 -915 4995 -885
rect 4995 -915 4996 -885
rect 4964 -916 4996 -915
rect 4964 -996 4996 -964
rect 4964 -1076 4996 -1044
rect 4964 -1125 4996 -1124
rect 4964 -1155 4965 -1125
rect 4965 -1155 4995 -1125
rect 4995 -1155 4996 -1125
rect 4964 -1156 4996 -1155
rect 4964 -1205 4996 -1204
rect 4964 -1235 4965 -1205
rect 4965 -1235 4995 -1205
rect 4995 -1235 4996 -1205
rect 4964 -1236 4996 -1235
rect 4964 -1285 4996 -1284
rect 4964 -1315 4965 -1285
rect 4965 -1315 4995 -1285
rect 4995 -1315 4996 -1285
rect 4964 -1316 4996 -1315
rect 4964 -1365 4996 -1364
rect 4964 -1395 4965 -1365
rect 4965 -1395 4995 -1365
rect 4995 -1395 4996 -1365
rect 4964 -1396 4996 -1395
rect 4964 -1445 4996 -1444
rect 4964 -1475 4965 -1445
rect 4965 -1475 4995 -1445
rect 4995 -1475 4996 -1445
rect 4964 -1476 4996 -1475
rect 4964 -1525 4996 -1524
rect 4964 -1555 4965 -1525
rect 4965 -1555 4995 -1525
rect 4995 -1555 4996 -1525
rect 4964 -1556 4996 -1555
rect 4964 -1636 4996 -1604
rect 4964 -1716 4996 -1684
rect 4964 -1765 4996 -1764
rect 4964 -1795 4965 -1765
rect 4965 -1795 4995 -1765
rect 4995 -1795 4996 -1765
rect 4964 -1796 4996 -1795
rect 4964 -1845 4996 -1844
rect 4964 -1875 4965 -1845
rect 4965 -1875 4995 -1845
rect 4995 -1875 4996 -1845
rect 4964 -1876 4996 -1875
rect 4964 -1956 4996 -1924
rect 4964 -2005 4996 -2004
rect 4964 -2035 4965 -2005
rect 4965 -2035 4995 -2005
rect 4995 -2035 4996 -2005
rect 4964 -2036 4996 -2035
rect 4964 -2116 4996 -2084
rect 4964 -2165 4996 -2164
rect 4964 -2195 4965 -2165
rect 4965 -2195 4995 -2165
rect 4995 -2195 4996 -2165
rect 4964 -2196 4996 -2195
rect 4964 -2276 4996 -2244
rect 4964 -2325 4996 -2324
rect 4964 -2355 4965 -2325
rect 4965 -2355 4995 -2325
rect 4995 -2355 4996 -2325
rect 4964 -2356 4996 -2355
rect 4964 -2405 4996 -2404
rect 4964 -2435 4965 -2405
rect 4965 -2435 4995 -2405
rect 4995 -2435 4996 -2405
rect 4964 -2436 4996 -2435
rect 4964 -2485 4996 -2484
rect 4964 -2515 4965 -2485
rect 4965 -2515 4995 -2485
rect 4995 -2515 4996 -2485
rect 4964 -2516 4996 -2515
rect 4964 -2565 4996 -2564
rect 4964 -2595 4965 -2565
rect 4965 -2595 4995 -2565
rect 4995 -2595 4996 -2565
rect 4964 -2596 4996 -2595
rect 4964 -2645 4996 -2644
rect 4964 -2675 4965 -2645
rect 4965 -2675 4995 -2645
rect 4995 -2675 4996 -2645
rect 4964 -2676 4996 -2675
rect 4964 -2725 4996 -2724
rect 4964 -2755 4965 -2725
rect 4965 -2755 4995 -2725
rect 4995 -2755 4996 -2725
rect 4964 -2756 4996 -2755
rect 4964 -2836 4996 -2804
rect 4964 -2885 4996 -2884
rect 4964 -2915 4965 -2885
rect 4965 -2915 4995 -2885
rect 4995 -2915 4996 -2885
rect 4964 -2916 4996 -2915
rect 4964 -2996 4996 -2964
rect 4964 -3045 4996 -3044
rect 4964 -3075 4965 -3045
rect 4965 -3075 4995 -3045
rect 4995 -3075 4996 -3045
rect 4964 -3076 4996 -3075
rect 4964 -3156 4996 -3124
rect 4964 -3205 4996 -3204
rect 4964 -3235 4965 -3205
rect 4965 -3235 4995 -3205
rect 4995 -3235 4996 -3205
rect 4964 -3236 4996 -3235
rect 4964 -3285 4996 -3284
rect 4964 -3315 4965 -3285
rect 4965 -3315 4995 -3285
rect 4995 -3315 4996 -3285
rect 4964 -3316 4996 -3315
rect 4964 -3396 4996 -3364
rect 4964 -3476 4996 -3444
rect 4964 -3525 4996 -3524
rect 4964 -3555 4965 -3525
rect 4965 -3555 4995 -3525
rect 4995 -3555 4996 -3525
rect 4964 -3556 4996 -3555
rect 4964 -3605 4996 -3604
rect 4964 -3635 4965 -3605
rect 4965 -3635 4995 -3605
rect 4995 -3635 4996 -3605
rect 4964 -3636 4996 -3635
rect 4964 -3685 4996 -3684
rect 4964 -3715 4965 -3685
rect 4965 -3715 4995 -3685
rect 4995 -3715 4996 -3685
rect 4964 -3716 4996 -3715
rect 5044 1035 5076 1036
rect 5044 1005 5045 1035
rect 5045 1005 5075 1035
rect 5075 1005 5076 1035
rect 5044 1004 5076 1005
rect 5044 955 5076 956
rect 5044 925 5045 955
rect 5045 925 5075 955
rect 5075 925 5076 955
rect 5044 924 5076 925
rect 5044 875 5076 876
rect 5044 845 5045 875
rect 5045 845 5075 875
rect 5075 845 5076 875
rect 5044 844 5076 845
rect 5044 764 5076 796
rect 5044 684 5076 716
rect 5044 635 5076 636
rect 5044 605 5045 635
rect 5045 605 5075 635
rect 5075 605 5076 635
rect 5044 604 5076 605
rect 5044 555 5076 556
rect 5044 525 5045 555
rect 5045 525 5075 555
rect 5075 525 5076 555
rect 5044 524 5076 525
rect 5044 444 5076 476
rect 5044 395 5076 396
rect 5044 365 5045 395
rect 5045 365 5075 395
rect 5075 365 5076 395
rect 5044 364 5076 365
rect 5044 284 5076 316
rect 5044 235 5076 236
rect 5044 205 5045 235
rect 5045 205 5075 235
rect 5075 205 5076 235
rect 5044 204 5076 205
rect 5044 124 5076 156
rect 5044 75 5076 76
rect 5044 45 5045 75
rect 5045 45 5075 75
rect 5075 45 5076 75
rect 5044 44 5076 45
rect 5044 -5 5076 -4
rect 5044 -35 5045 -5
rect 5045 -35 5075 -5
rect 5075 -35 5076 -5
rect 5044 -36 5076 -35
rect 5044 -85 5076 -84
rect 5044 -115 5045 -85
rect 5045 -115 5075 -85
rect 5075 -115 5076 -85
rect 5044 -116 5076 -115
rect 5044 -165 5076 -164
rect 5044 -195 5045 -165
rect 5045 -195 5075 -165
rect 5075 -195 5076 -165
rect 5044 -196 5076 -195
rect 5044 -245 5076 -244
rect 5044 -275 5045 -245
rect 5045 -275 5075 -245
rect 5075 -275 5076 -245
rect 5044 -276 5076 -275
rect 5044 -325 5076 -324
rect 5044 -355 5045 -325
rect 5045 -355 5075 -325
rect 5075 -355 5076 -325
rect 5044 -356 5076 -355
rect 5044 -436 5076 -404
rect 5044 -485 5076 -484
rect 5044 -515 5045 -485
rect 5045 -515 5075 -485
rect 5075 -515 5076 -485
rect 5044 -516 5076 -515
rect 5044 -596 5076 -564
rect 5044 -645 5076 -644
rect 5044 -675 5045 -645
rect 5045 -675 5075 -645
rect 5075 -675 5076 -645
rect 5044 -676 5076 -675
rect 5044 -756 5076 -724
rect 5044 -805 5076 -804
rect 5044 -835 5045 -805
rect 5045 -835 5075 -805
rect 5075 -835 5076 -805
rect 5044 -836 5076 -835
rect 5044 -885 5076 -884
rect 5044 -915 5045 -885
rect 5045 -915 5075 -885
rect 5075 -915 5076 -885
rect 5044 -916 5076 -915
rect 5044 -996 5076 -964
rect 5044 -1076 5076 -1044
rect 5044 -1125 5076 -1124
rect 5044 -1155 5045 -1125
rect 5045 -1155 5075 -1125
rect 5075 -1155 5076 -1125
rect 5044 -1156 5076 -1155
rect 5044 -1205 5076 -1204
rect 5044 -1235 5045 -1205
rect 5045 -1235 5075 -1205
rect 5075 -1235 5076 -1205
rect 5044 -1236 5076 -1235
rect 5044 -1285 5076 -1284
rect 5044 -1315 5045 -1285
rect 5045 -1315 5075 -1285
rect 5075 -1315 5076 -1285
rect 5044 -1316 5076 -1315
rect 5044 -1365 5076 -1364
rect 5044 -1395 5045 -1365
rect 5045 -1395 5075 -1365
rect 5075 -1395 5076 -1365
rect 5044 -1396 5076 -1395
rect 5044 -1445 5076 -1444
rect 5044 -1475 5045 -1445
rect 5045 -1475 5075 -1445
rect 5075 -1475 5076 -1445
rect 5044 -1476 5076 -1475
rect 5044 -1525 5076 -1524
rect 5044 -1555 5045 -1525
rect 5045 -1555 5075 -1525
rect 5075 -1555 5076 -1525
rect 5044 -1556 5076 -1555
rect 5044 -1636 5076 -1604
rect 5044 -1716 5076 -1684
rect 5044 -1765 5076 -1764
rect 5044 -1795 5045 -1765
rect 5045 -1795 5075 -1765
rect 5075 -1795 5076 -1765
rect 5044 -1796 5076 -1795
rect 5044 -1845 5076 -1844
rect 5044 -1875 5045 -1845
rect 5045 -1875 5075 -1845
rect 5075 -1875 5076 -1845
rect 5044 -1876 5076 -1875
rect 5044 -1956 5076 -1924
rect 5044 -2005 5076 -2004
rect 5044 -2035 5045 -2005
rect 5045 -2035 5075 -2005
rect 5075 -2035 5076 -2005
rect 5044 -2036 5076 -2035
rect 5044 -2116 5076 -2084
rect 5044 -2165 5076 -2164
rect 5044 -2195 5045 -2165
rect 5045 -2195 5075 -2165
rect 5075 -2195 5076 -2165
rect 5044 -2196 5076 -2195
rect 5044 -2276 5076 -2244
rect 5044 -2325 5076 -2324
rect 5044 -2355 5045 -2325
rect 5045 -2355 5075 -2325
rect 5075 -2355 5076 -2325
rect 5044 -2356 5076 -2355
rect 5044 -2405 5076 -2404
rect 5044 -2435 5045 -2405
rect 5045 -2435 5075 -2405
rect 5075 -2435 5076 -2405
rect 5044 -2436 5076 -2435
rect 5044 -2485 5076 -2484
rect 5044 -2515 5045 -2485
rect 5045 -2515 5075 -2485
rect 5075 -2515 5076 -2485
rect 5044 -2516 5076 -2515
rect 5044 -2565 5076 -2564
rect 5044 -2595 5045 -2565
rect 5045 -2595 5075 -2565
rect 5075 -2595 5076 -2565
rect 5044 -2596 5076 -2595
rect 5044 -2645 5076 -2644
rect 5044 -2675 5045 -2645
rect 5045 -2675 5075 -2645
rect 5075 -2675 5076 -2645
rect 5044 -2676 5076 -2675
rect 5044 -2725 5076 -2724
rect 5044 -2755 5045 -2725
rect 5045 -2755 5075 -2725
rect 5075 -2755 5076 -2725
rect 5044 -2756 5076 -2755
rect 5044 -2836 5076 -2804
rect 5044 -2885 5076 -2884
rect 5044 -2915 5045 -2885
rect 5045 -2915 5075 -2885
rect 5075 -2915 5076 -2885
rect 5044 -2916 5076 -2915
rect 5044 -2996 5076 -2964
rect 5044 -3045 5076 -3044
rect 5044 -3075 5045 -3045
rect 5045 -3075 5075 -3045
rect 5075 -3075 5076 -3045
rect 5044 -3076 5076 -3075
rect 5044 -3156 5076 -3124
rect 5044 -3205 5076 -3204
rect 5044 -3235 5045 -3205
rect 5045 -3235 5075 -3205
rect 5075 -3235 5076 -3205
rect 5044 -3236 5076 -3235
rect 5044 -3285 5076 -3284
rect 5044 -3315 5045 -3285
rect 5045 -3315 5075 -3285
rect 5075 -3315 5076 -3285
rect 5044 -3316 5076 -3315
rect 5044 -3396 5076 -3364
rect 5044 -3476 5076 -3444
rect 5044 -3525 5076 -3524
rect 5044 -3555 5045 -3525
rect 5045 -3555 5075 -3525
rect 5075 -3555 5076 -3525
rect 5044 -3556 5076 -3555
rect 5044 -3605 5076 -3604
rect 5044 -3635 5045 -3605
rect 5045 -3635 5075 -3605
rect 5075 -3635 5076 -3605
rect 5044 -3636 5076 -3635
rect 5044 -3685 5076 -3684
rect 5044 -3715 5045 -3685
rect 5045 -3715 5075 -3685
rect 5075 -3715 5076 -3685
rect 5044 -3716 5076 -3715
rect 5124 1035 5156 1036
rect 5124 1005 5125 1035
rect 5125 1005 5155 1035
rect 5155 1005 5156 1035
rect 5124 1004 5156 1005
rect 5124 955 5156 956
rect 5124 925 5125 955
rect 5125 925 5155 955
rect 5155 925 5156 955
rect 5124 924 5156 925
rect 5124 875 5156 876
rect 5124 845 5125 875
rect 5125 845 5155 875
rect 5155 845 5156 875
rect 5124 844 5156 845
rect 5124 764 5156 796
rect 5124 684 5156 716
rect 5124 635 5156 636
rect 5124 605 5125 635
rect 5125 605 5155 635
rect 5155 605 5156 635
rect 5124 604 5156 605
rect 5124 555 5156 556
rect 5124 525 5125 555
rect 5125 525 5155 555
rect 5155 525 5156 555
rect 5124 524 5156 525
rect 5124 444 5156 476
rect 5124 395 5156 396
rect 5124 365 5125 395
rect 5125 365 5155 395
rect 5155 365 5156 395
rect 5124 364 5156 365
rect 5124 284 5156 316
rect 5124 235 5156 236
rect 5124 205 5125 235
rect 5125 205 5155 235
rect 5155 205 5156 235
rect 5124 204 5156 205
rect 5124 124 5156 156
rect 5124 75 5156 76
rect 5124 45 5125 75
rect 5125 45 5155 75
rect 5155 45 5156 75
rect 5124 44 5156 45
rect 5124 -5 5156 -4
rect 5124 -35 5125 -5
rect 5125 -35 5155 -5
rect 5155 -35 5156 -5
rect 5124 -36 5156 -35
rect 5124 -85 5156 -84
rect 5124 -115 5125 -85
rect 5125 -115 5155 -85
rect 5155 -115 5156 -85
rect 5124 -116 5156 -115
rect 5124 -165 5156 -164
rect 5124 -195 5125 -165
rect 5125 -195 5155 -165
rect 5155 -195 5156 -165
rect 5124 -196 5156 -195
rect 5124 -245 5156 -244
rect 5124 -275 5125 -245
rect 5125 -275 5155 -245
rect 5155 -275 5156 -245
rect 5124 -276 5156 -275
rect 5124 -325 5156 -324
rect 5124 -355 5125 -325
rect 5125 -355 5155 -325
rect 5155 -355 5156 -325
rect 5124 -356 5156 -355
rect 5124 -436 5156 -404
rect 5124 -485 5156 -484
rect 5124 -515 5125 -485
rect 5125 -515 5155 -485
rect 5155 -515 5156 -485
rect 5124 -516 5156 -515
rect 5124 -596 5156 -564
rect 5124 -645 5156 -644
rect 5124 -675 5125 -645
rect 5125 -675 5155 -645
rect 5155 -675 5156 -645
rect 5124 -676 5156 -675
rect 5124 -756 5156 -724
rect 5124 -805 5156 -804
rect 5124 -835 5125 -805
rect 5125 -835 5155 -805
rect 5155 -835 5156 -805
rect 5124 -836 5156 -835
rect 5124 -885 5156 -884
rect 5124 -915 5125 -885
rect 5125 -915 5155 -885
rect 5155 -915 5156 -885
rect 5124 -916 5156 -915
rect 5124 -996 5156 -964
rect 5124 -1076 5156 -1044
rect 5124 -1125 5156 -1124
rect 5124 -1155 5125 -1125
rect 5125 -1155 5155 -1125
rect 5155 -1155 5156 -1125
rect 5124 -1156 5156 -1155
rect 5124 -1205 5156 -1204
rect 5124 -1235 5125 -1205
rect 5125 -1235 5155 -1205
rect 5155 -1235 5156 -1205
rect 5124 -1236 5156 -1235
rect 5124 -1285 5156 -1284
rect 5124 -1315 5125 -1285
rect 5125 -1315 5155 -1285
rect 5155 -1315 5156 -1285
rect 5124 -1316 5156 -1315
rect 5124 -1365 5156 -1364
rect 5124 -1395 5125 -1365
rect 5125 -1395 5155 -1365
rect 5155 -1395 5156 -1365
rect 5124 -1396 5156 -1395
rect 5124 -1445 5156 -1444
rect 5124 -1475 5125 -1445
rect 5125 -1475 5155 -1445
rect 5155 -1475 5156 -1445
rect 5124 -1476 5156 -1475
rect 5124 -1525 5156 -1524
rect 5124 -1555 5125 -1525
rect 5125 -1555 5155 -1525
rect 5155 -1555 5156 -1525
rect 5124 -1556 5156 -1555
rect 5124 -1636 5156 -1604
rect 5124 -1716 5156 -1684
rect 5124 -1765 5156 -1764
rect 5124 -1795 5125 -1765
rect 5125 -1795 5155 -1765
rect 5155 -1795 5156 -1765
rect 5124 -1796 5156 -1795
rect 5124 -1845 5156 -1844
rect 5124 -1875 5125 -1845
rect 5125 -1875 5155 -1845
rect 5155 -1875 5156 -1845
rect 5124 -1876 5156 -1875
rect 5124 -1956 5156 -1924
rect 5124 -2005 5156 -2004
rect 5124 -2035 5125 -2005
rect 5125 -2035 5155 -2005
rect 5155 -2035 5156 -2005
rect 5124 -2036 5156 -2035
rect 5124 -2116 5156 -2084
rect 5124 -2165 5156 -2164
rect 5124 -2195 5125 -2165
rect 5125 -2195 5155 -2165
rect 5155 -2195 5156 -2165
rect 5124 -2196 5156 -2195
rect 5124 -2276 5156 -2244
rect 5124 -2325 5156 -2324
rect 5124 -2355 5125 -2325
rect 5125 -2355 5155 -2325
rect 5155 -2355 5156 -2325
rect 5124 -2356 5156 -2355
rect 5124 -2405 5156 -2404
rect 5124 -2435 5125 -2405
rect 5125 -2435 5155 -2405
rect 5155 -2435 5156 -2405
rect 5124 -2436 5156 -2435
rect 5124 -2485 5156 -2484
rect 5124 -2515 5125 -2485
rect 5125 -2515 5155 -2485
rect 5155 -2515 5156 -2485
rect 5124 -2516 5156 -2515
rect 5124 -2565 5156 -2564
rect 5124 -2595 5125 -2565
rect 5125 -2595 5155 -2565
rect 5155 -2595 5156 -2565
rect 5124 -2596 5156 -2595
rect 5124 -2645 5156 -2644
rect 5124 -2675 5125 -2645
rect 5125 -2675 5155 -2645
rect 5155 -2675 5156 -2645
rect 5124 -2676 5156 -2675
rect 5124 -2725 5156 -2724
rect 5124 -2755 5125 -2725
rect 5125 -2755 5155 -2725
rect 5155 -2755 5156 -2725
rect 5124 -2756 5156 -2755
rect 5124 -2836 5156 -2804
rect 5124 -2885 5156 -2884
rect 5124 -2915 5125 -2885
rect 5125 -2915 5155 -2885
rect 5155 -2915 5156 -2885
rect 5124 -2916 5156 -2915
rect 5124 -2996 5156 -2964
rect 5124 -3045 5156 -3044
rect 5124 -3075 5125 -3045
rect 5125 -3075 5155 -3045
rect 5155 -3075 5156 -3045
rect 5124 -3076 5156 -3075
rect 5124 -3156 5156 -3124
rect 5124 -3205 5156 -3204
rect 5124 -3235 5125 -3205
rect 5125 -3235 5155 -3205
rect 5155 -3235 5156 -3205
rect 5124 -3236 5156 -3235
rect 5124 -3285 5156 -3284
rect 5124 -3315 5125 -3285
rect 5125 -3315 5155 -3285
rect 5155 -3315 5156 -3285
rect 5124 -3316 5156 -3315
rect 5124 -3396 5156 -3364
rect 5124 -3476 5156 -3444
rect 5124 -3525 5156 -3524
rect 5124 -3555 5125 -3525
rect 5125 -3555 5155 -3525
rect 5155 -3555 5156 -3525
rect 5124 -3556 5156 -3555
rect 5124 -3605 5156 -3604
rect 5124 -3635 5125 -3605
rect 5125 -3635 5155 -3605
rect 5155 -3635 5156 -3605
rect 5124 -3636 5156 -3635
rect 5124 -3685 5156 -3684
rect 5124 -3715 5125 -3685
rect 5125 -3715 5155 -3685
rect 5155 -3715 5156 -3685
rect 5124 -3716 5156 -3715
rect 5204 1035 5236 1036
rect 5204 1005 5205 1035
rect 5205 1005 5235 1035
rect 5235 1005 5236 1035
rect 5204 1004 5236 1005
rect 5204 955 5236 956
rect 5204 925 5205 955
rect 5205 925 5235 955
rect 5235 925 5236 955
rect 5204 924 5236 925
rect 5204 875 5236 876
rect 5204 845 5205 875
rect 5205 845 5235 875
rect 5235 845 5236 875
rect 5204 844 5236 845
rect 5204 764 5236 796
rect 5204 684 5236 716
rect 5204 635 5236 636
rect 5204 605 5205 635
rect 5205 605 5235 635
rect 5235 605 5236 635
rect 5204 604 5236 605
rect 5204 555 5236 556
rect 5204 525 5205 555
rect 5205 525 5235 555
rect 5235 525 5236 555
rect 5204 524 5236 525
rect 5204 444 5236 476
rect 5204 395 5236 396
rect 5204 365 5205 395
rect 5205 365 5235 395
rect 5235 365 5236 395
rect 5204 364 5236 365
rect 5204 284 5236 316
rect 5204 235 5236 236
rect 5204 205 5205 235
rect 5205 205 5235 235
rect 5235 205 5236 235
rect 5204 204 5236 205
rect 5204 124 5236 156
rect 5204 75 5236 76
rect 5204 45 5205 75
rect 5205 45 5235 75
rect 5235 45 5236 75
rect 5204 44 5236 45
rect 5204 -5 5236 -4
rect 5204 -35 5205 -5
rect 5205 -35 5235 -5
rect 5235 -35 5236 -5
rect 5204 -36 5236 -35
rect 5204 -85 5236 -84
rect 5204 -115 5205 -85
rect 5205 -115 5235 -85
rect 5235 -115 5236 -85
rect 5204 -116 5236 -115
rect 5204 -165 5236 -164
rect 5204 -195 5205 -165
rect 5205 -195 5235 -165
rect 5235 -195 5236 -165
rect 5204 -196 5236 -195
rect 5204 -245 5236 -244
rect 5204 -275 5205 -245
rect 5205 -275 5235 -245
rect 5235 -275 5236 -245
rect 5204 -276 5236 -275
rect 5204 -325 5236 -324
rect 5204 -355 5205 -325
rect 5205 -355 5235 -325
rect 5235 -355 5236 -325
rect 5204 -356 5236 -355
rect 5204 -436 5236 -404
rect 5204 -485 5236 -484
rect 5204 -515 5205 -485
rect 5205 -515 5235 -485
rect 5235 -515 5236 -485
rect 5204 -516 5236 -515
rect 5204 -596 5236 -564
rect 5204 -645 5236 -644
rect 5204 -675 5205 -645
rect 5205 -675 5235 -645
rect 5235 -675 5236 -645
rect 5204 -676 5236 -675
rect 5204 -756 5236 -724
rect 5204 -805 5236 -804
rect 5204 -835 5205 -805
rect 5205 -835 5235 -805
rect 5235 -835 5236 -805
rect 5204 -836 5236 -835
rect 5204 -885 5236 -884
rect 5204 -915 5205 -885
rect 5205 -915 5235 -885
rect 5235 -915 5236 -885
rect 5204 -916 5236 -915
rect 5204 -996 5236 -964
rect 5204 -1076 5236 -1044
rect 5204 -1125 5236 -1124
rect 5204 -1155 5205 -1125
rect 5205 -1155 5235 -1125
rect 5235 -1155 5236 -1125
rect 5204 -1156 5236 -1155
rect 5204 -1205 5236 -1204
rect 5204 -1235 5205 -1205
rect 5205 -1235 5235 -1205
rect 5235 -1235 5236 -1205
rect 5204 -1236 5236 -1235
rect 5204 -1285 5236 -1284
rect 5204 -1315 5205 -1285
rect 5205 -1315 5235 -1285
rect 5235 -1315 5236 -1285
rect 5204 -1316 5236 -1315
rect 5204 -1365 5236 -1364
rect 5204 -1395 5205 -1365
rect 5205 -1395 5235 -1365
rect 5235 -1395 5236 -1365
rect 5204 -1396 5236 -1395
rect 5204 -1445 5236 -1444
rect 5204 -1475 5205 -1445
rect 5205 -1475 5235 -1445
rect 5235 -1475 5236 -1445
rect 5204 -1476 5236 -1475
rect 5204 -1525 5236 -1524
rect 5204 -1555 5205 -1525
rect 5205 -1555 5235 -1525
rect 5235 -1555 5236 -1525
rect 5204 -1556 5236 -1555
rect 5204 -1636 5236 -1604
rect 5204 -1716 5236 -1684
rect 5204 -1765 5236 -1764
rect 5204 -1795 5205 -1765
rect 5205 -1795 5235 -1765
rect 5235 -1795 5236 -1765
rect 5204 -1796 5236 -1795
rect 5204 -1845 5236 -1844
rect 5204 -1875 5205 -1845
rect 5205 -1875 5235 -1845
rect 5235 -1875 5236 -1845
rect 5204 -1876 5236 -1875
rect 5204 -1956 5236 -1924
rect 5204 -2005 5236 -2004
rect 5204 -2035 5205 -2005
rect 5205 -2035 5235 -2005
rect 5235 -2035 5236 -2005
rect 5204 -2036 5236 -2035
rect 5204 -2116 5236 -2084
rect 5204 -2165 5236 -2164
rect 5204 -2195 5205 -2165
rect 5205 -2195 5235 -2165
rect 5235 -2195 5236 -2165
rect 5204 -2196 5236 -2195
rect 5204 -2276 5236 -2244
rect 5204 -2325 5236 -2324
rect 5204 -2355 5205 -2325
rect 5205 -2355 5235 -2325
rect 5235 -2355 5236 -2325
rect 5204 -2356 5236 -2355
rect 5204 -2405 5236 -2404
rect 5204 -2435 5205 -2405
rect 5205 -2435 5235 -2405
rect 5235 -2435 5236 -2405
rect 5204 -2436 5236 -2435
rect 5204 -2485 5236 -2484
rect 5204 -2515 5205 -2485
rect 5205 -2515 5235 -2485
rect 5235 -2515 5236 -2485
rect 5204 -2516 5236 -2515
rect 5204 -2565 5236 -2564
rect 5204 -2595 5205 -2565
rect 5205 -2595 5235 -2565
rect 5235 -2595 5236 -2565
rect 5204 -2596 5236 -2595
rect 5204 -2645 5236 -2644
rect 5204 -2675 5205 -2645
rect 5205 -2675 5235 -2645
rect 5235 -2675 5236 -2645
rect 5204 -2676 5236 -2675
rect 5204 -2725 5236 -2724
rect 5204 -2755 5205 -2725
rect 5205 -2755 5235 -2725
rect 5235 -2755 5236 -2725
rect 5204 -2756 5236 -2755
rect 5204 -2836 5236 -2804
rect 5204 -2885 5236 -2884
rect 5204 -2915 5205 -2885
rect 5205 -2915 5235 -2885
rect 5235 -2915 5236 -2885
rect 5204 -2916 5236 -2915
rect 5204 -2996 5236 -2964
rect 5204 -3045 5236 -3044
rect 5204 -3075 5205 -3045
rect 5205 -3075 5235 -3045
rect 5235 -3075 5236 -3045
rect 5204 -3076 5236 -3075
rect 5204 -3156 5236 -3124
rect 5204 -3205 5236 -3204
rect 5204 -3235 5205 -3205
rect 5205 -3235 5235 -3205
rect 5235 -3235 5236 -3205
rect 5204 -3236 5236 -3235
rect 5204 -3285 5236 -3284
rect 5204 -3315 5205 -3285
rect 5205 -3315 5235 -3285
rect 5235 -3315 5236 -3285
rect 5204 -3316 5236 -3315
rect 5204 -3396 5236 -3364
rect 5204 -3476 5236 -3444
rect 5204 -3525 5236 -3524
rect 5204 -3555 5205 -3525
rect 5205 -3555 5235 -3525
rect 5235 -3555 5236 -3525
rect 5204 -3556 5236 -3555
rect 5204 -3605 5236 -3604
rect 5204 -3635 5205 -3605
rect 5205 -3635 5235 -3605
rect 5235 -3635 5236 -3605
rect 5204 -3636 5236 -3635
rect 5204 -3685 5236 -3684
rect 5204 -3715 5205 -3685
rect 5205 -3715 5235 -3685
rect 5235 -3715 5236 -3685
rect 5204 -3716 5236 -3715
rect 5284 1035 5316 1036
rect 5284 1005 5285 1035
rect 5285 1005 5315 1035
rect 5315 1005 5316 1035
rect 5284 1004 5316 1005
rect 5284 955 5316 956
rect 5284 925 5285 955
rect 5285 925 5315 955
rect 5315 925 5316 955
rect 5284 924 5316 925
rect 5284 875 5316 876
rect 5284 845 5285 875
rect 5285 845 5315 875
rect 5315 845 5316 875
rect 5284 844 5316 845
rect 5284 764 5316 796
rect 5284 684 5316 716
rect 5284 635 5316 636
rect 5284 605 5285 635
rect 5285 605 5315 635
rect 5315 605 5316 635
rect 5284 604 5316 605
rect 5284 555 5316 556
rect 5284 525 5285 555
rect 5285 525 5315 555
rect 5315 525 5316 555
rect 5284 524 5316 525
rect 5284 444 5316 476
rect 5284 395 5316 396
rect 5284 365 5285 395
rect 5285 365 5315 395
rect 5315 365 5316 395
rect 5284 364 5316 365
rect 5284 284 5316 316
rect 5284 235 5316 236
rect 5284 205 5285 235
rect 5285 205 5315 235
rect 5315 205 5316 235
rect 5284 204 5316 205
rect 5284 124 5316 156
rect 5284 75 5316 76
rect 5284 45 5285 75
rect 5285 45 5315 75
rect 5315 45 5316 75
rect 5284 44 5316 45
rect 5284 -5 5316 -4
rect 5284 -35 5285 -5
rect 5285 -35 5315 -5
rect 5315 -35 5316 -5
rect 5284 -36 5316 -35
rect 5284 -85 5316 -84
rect 5284 -115 5285 -85
rect 5285 -115 5315 -85
rect 5315 -115 5316 -85
rect 5284 -116 5316 -115
rect 5284 -165 5316 -164
rect 5284 -195 5285 -165
rect 5285 -195 5315 -165
rect 5315 -195 5316 -165
rect 5284 -196 5316 -195
rect 5284 -245 5316 -244
rect 5284 -275 5285 -245
rect 5285 -275 5315 -245
rect 5315 -275 5316 -245
rect 5284 -276 5316 -275
rect 5284 -325 5316 -324
rect 5284 -355 5285 -325
rect 5285 -355 5315 -325
rect 5315 -355 5316 -325
rect 5284 -356 5316 -355
rect 5284 -436 5316 -404
rect 5284 -485 5316 -484
rect 5284 -515 5285 -485
rect 5285 -515 5315 -485
rect 5315 -515 5316 -485
rect 5284 -516 5316 -515
rect 5284 -596 5316 -564
rect 5284 -645 5316 -644
rect 5284 -675 5285 -645
rect 5285 -675 5315 -645
rect 5315 -675 5316 -645
rect 5284 -676 5316 -675
rect 5284 -756 5316 -724
rect 5284 -805 5316 -804
rect 5284 -835 5285 -805
rect 5285 -835 5315 -805
rect 5315 -835 5316 -805
rect 5284 -836 5316 -835
rect 5284 -885 5316 -884
rect 5284 -915 5285 -885
rect 5285 -915 5315 -885
rect 5315 -915 5316 -885
rect 5284 -916 5316 -915
rect 5284 -996 5316 -964
rect 5284 -1076 5316 -1044
rect 5284 -1125 5316 -1124
rect 5284 -1155 5285 -1125
rect 5285 -1155 5315 -1125
rect 5315 -1155 5316 -1125
rect 5284 -1156 5316 -1155
rect 5284 -1205 5316 -1204
rect 5284 -1235 5285 -1205
rect 5285 -1235 5315 -1205
rect 5315 -1235 5316 -1205
rect 5284 -1236 5316 -1235
rect 5284 -1285 5316 -1284
rect 5284 -1315 5285 -1285
rect 5285 -1315 5315 -1285
rect 5315 -1315 5316 -1285
rect 5284 -1316 5316 -1315
rect 5284 -1365 5316 -1364
rect 5284 -1395 5285 -1365
rect 5285 -1395 5315 -1365
rect 5315 -1395 5316 -1365
rect 5284 -1396 5316 -1395
rect 5284 -1445 5316 -1444
rect 5284 -1475 5285 -1445
rect 5285 -1475 5315 -1445
rect 5315 -1475 5316 -1445
rect 5284 -1476 5316 -1475
rect 5284 -1525 5316 -1524
rect 5284 -1555 5285 -1525
rect 5285 -1555 5315 -1525
rect 5315 -1555 5316 -1525
rect 5284 -1556 5316 -1555
rect 5284 -1636 5316 -1604
rect 5284 -1716 5316 -1684
rect 5284 -1765 5316 -1764
rect 5284 -1795 5285 -1765
rect 5285 -1795 5315 -1765
rect 5315 -1795 5316 -1765
rect 5284 -1796 5316 -1795
rect 5284 -1845 5316 -1844
rect 5284 -1875 5285 -1845
rect 5285 -1875 5315 -1845
rect 5315 -1875 5316 -1845
rect 5284 -1876 5316 -1875
rect 5284 -1956 5316 -1924
rect 5284 -2005 5316 -2004
rect 5284 -2035 5285 -2005
rect 5285 -2035 5315 -2005
rect 5315 -2035 5316 -2005
rect 5284 -2036 5316 -2035
rect 5284 -2116 5316 -2084
rect 5284 -2165 5316 -2164
rect 5284 -2195 5285 -2165
rect 5285 -2195 5315 -2165
rect 5315 -2195 5316 -2165
rect 5284 -2196 5316 -2195
rect 5284 -2276 5316 -2244
rect 5284 -2325 5316 -2324
rect 5284 -2355 5285 -2325
rect 5285 -2355 5315 -2325
rect 5315 -2355 5316 -2325
rect 5284 -2356 5316 -2355
rect 5284 -2405 5316 -2404
rect 5284 -2435 5285 -2405
rect 5285 -2435 5315 -2405
rect 5315 -2435 5316 -2405
rect 5284 -2436 5316 -2435
rect 5284 -2485 5316 -2484
rect 5284 -2515 5285 -2485
rect 5285 -2515 5315 -2485
rect 5315 -2515 5316 -2485
rect 5284 -2516 5316 -2515
rect 5284 -2565 5316 -2564
rect 5284 -2595 5285 -2565
rect 5285 -2595 5315 -2565
rect 5315 -2595 5316 -2565
rect 5284 -2596 5316 -2595
rect 5284 -2645 5316 -2644
rect 5284 -2675 5285 -2645
rect 5285 -2675 5315 -2645
rect 5315 -2675 5316 -2645
rect 5284 -2676 5316 -2675
rect 5284 -2725 5316 -2724
rect 5284 -2755 5285 -2725
rect 5285 -2755 5315 -2725
rect 5315 -2755 5316 -2725
rect 5284 -2756 5316 -2755
rect 5284 -2836 5316 -2804
rect 5284 -2885 5316 -2884
rect 5284 -2915 5285 -2885
rect 5285 -2915 5315 -2885
rect 5315 -2915 5316 -2885
rect 5284 -2916 5316 -2915
rect 5284 -2996 5316 -2964
rect 5284 -3045 5316 -3044
rect 5284 -3075 5285 -3045
rect 5285 -3075 5315 -3045
rect 5315 -3075 5316 -3045
rect 5284 -3076 5316 -3075
rect 5284 -3156 5316 -3124
rect 5284 -3205 5316 -3204
rect 5284 -3235 5285 -3205
rect 5285 -3235 5315 -3205
rect 5315 -3235 5316 -3205
rect 5284 -3236 5316 -3235
rect 5284 -3285 5316 -3284
rect 5284 -3315 5285 -3285
rect 5285 -3315 5315 -3285
rect 5315 -3315 5316 -3285
rect 5284 -3316 5316 -3315
rect 5284 -3396 5316 -3364
rect 5284 -3476 5316 -3444
rect 5284 -3525 5316 -3524
rect 5284 -3555 5285 -3525
rect 5285 -3555 5315 -3525
rect 5315 -3555 5316 -3525
rect 5284 -3556 5316 -3555
rect 5284 -3605 5316 -3604
rect 5284 -3635 5285 -3605
rect 5285 -3635 5315 -3605
rect 5315 -3635 5316 -3605
rect 5284 -3636 5316 -3635
rect 5284 -3685 5316 -3684
rect 5284 -3715 5285 -3685
rect 5285 -3715 5315 -3685
rect 5315 -3715 5316 -3685
rect 5284 -3716 5316 -3715
rect 5364 1035 5396 1036
rect 5364 1005 5365 1035
rect 5365 1005 5395 1035
rect 5395 1005 5396 1035
rect 5364 1004 5396 1005
rect 5364 955 5396 956
rect 5364 925 5365 955
rect 5365 925 5395 955
rect 5395 925 5396 955
rect 5364 924 5396 925
rect 5364 875 5396 876
rect 5364 845 5365 875
rect 5365 845 5395 875
rect 5395 845 5396 875
rect 5364 844 5396 845
rect 5364 764 5396 796
rect 5364 684 5396 716
rect 5364 635 5396 636
rect 5364 605 5365 635
rect 5365 605 5395 635
rect 5395 605 5396 635
rect 5364 604 5396 605
rect 5364 555 5396 556
rect 5364 525 5365 555
rect 5365 525 5395 555
rect 5395 525 5396 555
rect 5364 524 5396 525
rect 5364 444 5396 476
rect 5364 395 5396 396
rect 5364 365 5365 395
rect 5365 365 5395 395
rect 5395 365 5396 395
rect 5364 364 5396 365
rect 5364 284 5396 316
rect 5364 235 5396 236
rect 5364 205 5365 235
rect 5365 205 5395 235
rect 5395 205 5396 235
rect 5364 204 5396 205
rect 5364 124 5396 156
rect 5364 75 5396 76
rect 5364 45 5365 75
rect 5365 45 5395 75
rect 5395 45 5396 75
rect 5364 44 5396 45
rect 5364 -5 5396 -4
rect 5364 -35 5365 -5
rect 5365 -35 5395 -5
rect 5395 -35 5396 -5
rect 5364 -36 5396 -35
rect 5364 -85 5396 -84
rect 5364 -115 5365 -85
rect 5365 -115 5395 -85
rect 5395 -115 5396 -85
rect 5364 -116 5396 -115
rect 5364 -165 5396 -164
rect 5364 -195 5365 -165
rect 5365 -195 5395 -165
rect 5395 -195 5396 -165
rect 5364 -196 5396 -195
rect 5364 -245 5396 -244
rect 5364 -275 5365 -245
rect 5365 -275 5395 -245
rect 5395 -275 5396 -245
rect 5364 -276 5396 -275
rect 5364 -325 5396 -324
rect 5364 -355 5365 -325
rect 5365 -355 5395 -325
rect 5395 -355 5396 -325
rect 5364 -356 5396 -355
rect 5364 -436 5396 -404
rect 5364 -485 5396 -484
rect 5364 -515 5365 -485
rect 5365 -515 5395 -485
rect 5395 -515 5396 -485
rect 5364 -516 5396 -515
rect 5364 -596 5396 -564
rect 5364 -645 5396 -644
rect 5364 -675 5365 -645
rect 5365 -675 5395 -645
rect 5395 -675 5396 -645
rect 5364 -676 5396 -675
rect 5364 -756 5396 -724
rect 5364 -805 5396 -804
rect 5364 -835 5365 -805
rect 5365 -835 5395 -805
rect 5395 -835 5396 -805
rect 5364 -836 5396 -835
rect 5364 -885 5396 -884
rect 5364 -915 5365 -885
rect 5365 -915 5395 -885
rect 5395 -915 5396 -885
rect 5364 -916 5396 -915
rect 5364 -996 5396 -964
rect 5364 -1076 5396 -1044
rect 5364 -1125 5396 -1124
rect 5364 -1155 5365 -1125
rect 5365 -1155 5395 -1125
rect 5395 -1155 5396 -1125
rect 5364 -1156 5396 -1155
rect 5364 -1205 5396 -1204
rect 5364 -1235 5365 -1205
rect 5365 -1235 5395 -1205
rect 5395 -1235 5396 -1205
rect 5364 -1236 5396 -1235
rect 5364 -1285 5396 -1284
rect 5364 -1315 5365 -1285
rect 5365 -1315 5395 -1285
rect 5395 -1315 5396 -1285
rect 5364 -1316 5396 -1315
rect 5364 -1365 5396 -1364
rect 5364 -1395 5365 -1365
rect 5365 -1395 5395 -1365
rect 5395 -1395 5396 -1365
rect 5364 -1396 5396 -1395
rect 5364 -1445 5396 -1444
rect 5364 -1475 5365 -1445
rect 5365 -1475 5395 -1445
rect 5395 -1475 5396 -1445
rect 5364 -1476 5396 -1475
rect 5364 -1525 5396 -1524
rect 5364 -1555 5365 -1525
rect 5365 -1555 5395 -1525
rect 5395 -1555 5396 -1525
rect 5364 -1556 5396 -1555
rect 5364 -1636 5396 -1604
rect 5364 -1716 5396 -1684
rect 5364 -1765 5396 -1764
rect 5364 -1795 5365 -1765
rect 5365 -1795 5395 -1765
rect 5395 -1795 5396 -1765
rect 5364 -1796 5396 -1795
rect 5364 -1845 5396 -1844
rect 5364 -1875 5365 -1845
rect 5365 -1875 5395 -1845
rect 5395 -1875 5396 -1845
rect 5364 -1876 5396 -1875
rect 5364 -1956 5396 -1924
rect 5364 -2005 5396 -2004
rect 5364 -2035 5365 -2005
rect 5365 -2035 5395 -2005
rect 5395 -2035 5396 -2005
rect 5364 -2036 5396 -2035
rect 5364 -2116 5396 -2084
rect 5364 -2165 5396 -2164
rect 5364 -2195 5365 -2165
rect 5365 -2195 5395 -2165
rect 5395 -2195 5396 -2165
rect 5364 -2196 5396 -2195
rect 5364 -2276 5396 -2244
rect 5364 -2325 5396 -2324
rect 5364 -2355 5365 -2325
rect 5365 -2355 5395 -2325
rect 5395 -2355 5396 -2325
rect 5364 -2356 5396 -2355
rect 5364 -2405 5396 -2404
rect 5364 -2435 5365 -2405
rect 5365 -2435 5395 -2405
rect 5395 -2435 5396 -2405
rect 5364 -2436 5396 -2435
rect 5364 -2485 5396 -2484
rect 5364 -2515 5365 -2485
rect 5365 -2515 5395 -2485
rect 5395 -2515 5396 -2485
rect 5364 -2516 5396 -2515
rect 5364 -2565 5396 -2564
rect 5364 -2595 5365 -2565
rect 5365 -2595 5395 -2565
rect 5395 -2595 5396 -2565
rect 5364 -2596 5396 -2595
rect 5364 -2645 5396 -2644
rect 5364 -2675 5365 -2645
rect 5365 -2675 5395 -2645
rect 5395 -2675 5396 -2645
rect 5364 -2676 5396 -2675
rect 5364 -2725 5396 -2724
rect 5364 -2755 5365 -2725
rect 5365 -2755 5395 -2725
rect 5395 -2755 5396 -2725
rect 5364 -2756 5396 -2755
rect 5364 -2836 5396 -2804
rect 5364 -2885 5396 -2884
rect 5364 -2915 5365 -2885
rect 5365 -2915 5395 -2885
rect 5395 -2915 5396 -2885
rect 5364 -2916 5396 -2915
rect 5364 -2996 5396 -2964
rect 5364 -3045 5396 -3044
rect 5364 -3075 5365 -3045
rect 5365 -3075 5395 -3045
rect 5395 -3075 5396 -3045
rect 5364 -3076 5396 -3075
rect 5364 -3156 5396 -3124
rect 5364 -3205 5396 -3204
rect 5364 -3235 5365 -3205
rect 5365 -3235 5395 -3205
rect 5395 -3235 5396 -3205
rect 5364 -3236 5396 -3235
rect 5364 -3285 5396 -3284
rect 5364 -3315 5365 -3285
rect 5365 -3315 5395 -3285
rect 5395 -3315 5396 -3285
rect 5364 -3316 5396 -3315
rect 5364 -3396 5396 -3364
rect 5364 -3476 5396 -3444
rect 5364 -3525 5396 -3524
rect 5364 -3555 5365 -3525
rect 5365 -3555 5395 -3525
rect 5395 -3555 5396 -3525
rect 5364 -3556 5396 -3555
rect 5364 -3605 5396 -3604
rect 5364 -3635 5365 -3605
rect 5365 -3635 5395 -3605
rect 5395 -3635 5396 -3605
rect 5364 -3636 5396 -3635
rect 5364 -3685 5396 -3684
rect 5364 -3715 5365 -3685
rect 5365 -3715 5395 -3685
rect 5395 -3715 5396 -3685
rect 5364 -3716 5396 -3715
rect 5444 1035 5476 1036
rect 5444 1005 5445 1035
rect 5445 1005 5475 1035
rect 5475 1005 5476 1035
rect 5444 1004 5476 1005
rect 5444 955 5476 956
rect 5444 925 5445 955
rect 5445 925 5475 955
rect 5475 925 5476 955
rect 5444 924 5476 925
rect 5444 875 5476 876
rect 5444 845 5445 875
rect 5445 845 5475 875
rect 5475 845 5476 875
rect 5444 844 5476 845
rect 5444 764 5476 796
rect 5444 684 5476 716
rect 5444 635 5476 636
rect 5444 605 5445 635
rect 5445 605 5475 635
rect 5475 605 5476 635
rect 5444 604 5476 605
rect 5444 555 5476 556
rect 5444 525 5445 555
rect 5445 525 5475 555
rect 5475 525 5476 555
rect 5444 524 5476 525
rect 5444 444 5476 476
rect 5444 395 5476 396
rect 5444 365 5445 395
rect 5445 365 5475 395
rect 5475 365 5476 395
rect 5444 364 5476 365
rect 5444 284 5476 316
rect 5444 235 5476 236
rect 5444 205 5445 235
rect 5445 205 5475 235
rect 5475 205 5476 235
rect 5444 204 5476 205
rect 5444 124 5476 156
rect 5444 75 5476 76
rect 5444 45 5445 75
rect 5445 45 5475 75
rect 5475 45 5476 75
rect 5444 44 5476 45
rect 5444 -5 5476 -4
rect 5444 -35 5445 -5
rect 5445 -35 5475 -5
rect 5475 -35 5476 -5
rect 5444 -36 5476 -35
rect 5444 -85 5476 -84
rect 5444 -115 5445 -85
rect 5445 -115 5475 -85
rect 5475 -115 5476 -85
rect 5444 -116 5476 -115
rect 5444 -165 5476 -164
rect 5444 -195 5445 -165
rect 5445 -195 5475 -165
rect 5475 -195 5476 -165
rect 5444 -196 5476 -195
rect 5444 -245 5476 -244
rect 5444 -275 5445 -245
rect 5445 -275 5475 -245
rect 5475 -275 5476 -245
rect 5444 -276 5476 -275
rect 5444 -325 5476 -324
rect 5444 -355 5445 -325
rect 5445 -355 5475 -325
rect 5475 -355 5476 -325
rect 5444 -356 5476 -355
rect 5444 -436 5476 -404
rect 5444 -485 5476 -484
rect 5444 -515 5445 -485
rect 5445 -515 5475 -485
rect 5475 -515 5476 -485
rect 5444 -516 5476 -515
rect 5444 -596 5476 -564
rect 5444 -645 5476 -644
rect 5444 -675 5445 -645
rect 5445 -675 5475 -645
rect 5475 -675 5476 -645
rect 5444 -676 5476 -675
rect 5444 -756 5476 -724
rect 5444 -805 5476 -804
rect 5444 -835 5445 -805
rect 5445 -835 5475 -805
rect 5475 -835 5476 -805
rect 5444 -836 5476 -835
rect 5444 -885 5476 -884
rect 5444 -915 5445 -885
rect 5445 -915 5475 -885
rect 5475 -915 5476 -885
rect 5444 -916 5476 -915
rect 5444 -996 5476 -964
rect 5444 -1076 5476 -1044
rect 5444 -1125 5476 -1124
rect 5444 -1155 5445 -1125
rect 5445 -1155 5475 -1125
rect 5475 -1155 5476 -1125
rect 5444 -1156 5476 -1155
rect 5444 -1205 5476 -1204
rect 5444 -1235 5445 -1205
rect 5445 -1235 5475 -1205
rect 5475 -1235 5476 -1205
rect 5444 -1236 5476 -1235
rect 5444 -1285 5476 -1284
rect 5444 -1315 5445 -1285
rect 5445 -1315 5475 -1285
rect 5475 -1315 5476 -1285
rect 5444 -1316 5476 -1315
rect 5444 -1365 5476 -1364
rect 5444 -1395 5445 -1365
rect 5445 -1395 5475 -1365
rect 5475 -1395 5476 -1365
rect 5444 -1396 5476 -1395
rect 5444 -1445 5476 -1444
rect 5444 -1475 5445 -1445
rect 5445 -1475 5475 -1445
rect 5475 -1475 5476 -1445
rect 5444 -1476 5476 -1475
rect 5444 -1525 5476 -1524
rect 5444 -1555 5445 -1525
rect 5445 -1555 5475 -1525
rect 5475 -1555 5476 -1525
rect 5444 -1556 5476 -1555
rect 5444 -1636 5476 -1604
rect 5444 -1716 5476 -1684
rect 5444 -1765 5476 -1764
rect 5444 -1795 5445 -1765
rect 5445 -1795 5475 -1765
rect 5475 -1795 5476 -1765
rect 5444 -1796 5476 -1795
rect 5444 -1845 5476 -1844
rect 5444 -1875 5445 -1845
rect 5445 -1875 5475 -1845
rect 5475 -1875 5476 -1845
rect 5444 -1876 5476 -1875
rect 5444 -1956 5476 -1924
rect 5444 -2005 5476 -2004
rect 5444 -2035 5445 -2005
rect 5445 -2035 5475 -2005
rect 5475 -2035 5476 -2005
rect 5444 -2036 5476 -2035
rect 5444 -2116 5476 -2084
rect 5444 -2165 5476 -2164
rect 5444 -2195 5445 -2165
rect 5445 -2195 5475 -2165
rect 5475 -2195 5476 -2165
rect 5444 -2196 5476 -2195
rect 5444 -2276 5476 -2244
rect 5444 -2325 5476 -2324
rect 5444 -2355 5445 -2325
rect 5445 -2355 5475 -2325
rect 5475 -2355 5476 -2325
rect 5444 -2356 5476 -2355
rect 5444 -2405 5476 -2404
rect 5444 -2435 5445 -2405
rect 5445 -2435 5475 -2405
rect 5475 -2435 5476 -2405
rect 5444 -2436 5476 -2435
rect 5444 -2485 5476 -2484
rect 5444 -2515 5445 -2485
rect 5445 -2515 5475 -2485
rect 5475 -2515 5476 -2485
rect 5444 -2516 5476 -2515
rect 5444 -2565 5476 -2564
rect 5444 -2595 5445 -2565
rect 5445 -2595 5475 -2565
rect 5475 -2595 5476 -2565
rect 5444 -2596 5476 -2595
rect 5444 -2645 5476 -2644
rect 5444 -2675 5445 -2645
rect 5445 -2675 5475 -2645
rect 5475 -2675 5476 -2645
rect 5444 -2676 5476 -2675
rect 5444 -2725 5476 -2724
rect 5444 -2755 5445 -2725
rect 5445 -2755 5475 -2725
rect 5475 -2755 5476 -2725
rect 5444 -2756 5476 -2755
rect 5444 -2836 5476 -2804
rect 5444 -2885 5476 -2884
rect 5444 -2915 5445 -2885
rect 5445 -2915 5475 -2885
rect 5475 -2915 5476 -2885
rect 5444 -2916 5476 -2915
rect 5444 -2996 5476 -2964
rect 5444 -3045 5476 -3044
rect 5444 -3075 5445 -3045
rect 5445 -3075 5475 -3045
rect 5475 -3075 5476 -3045
rect 5444 -3076 5476 -3075
rect 5444 -3156 5476 -3124
rect 5444 -3205 5476 -3204
rect 5444 -3235 5445 -3205
rect 5445 -3235 5475 -3205
rect 5475 -3235 5476 -3205
rect 5444 -3236 5476 -3235
rect 5444 -3285 5476 -3284
rect 5444 -3315 5445 -3285
rect 5445 -3315 5475 -3285
rect 5475 -3315 5476 -3285
rect 5444 -3316 5476 -3315
rect 5444 -3396 5476 -3364
rect 5444 -3476 5476 -3444
rect 5444 -3525 5476 -3524
rect 5444 -3555 5445 -3525
rect 5445 -3555 5475 -3525
rect 5475 -3555 5476 -3525
rect 5444 -3556 5476 -3555
rect 5444 -3605 5476 -3604
rect 5444 -3635 5445 -3605
rect 5445 -3635 5475 -3605
rect 5475 -3635 5476 -3605
rect 5444 -3636 5476 -3635
rect 5444 -3685 5476 -3684
rect 5444 -3715 5445 -3685
rect 5445 -3715 5475 -3685
rect 5475 -3715 5476 -3685
rect 5444 -3716 5476 -3715
rect 5524 1035 5556 1036
rect 5524 1005 5525 1035
rect 5525 1005 5555 1035
rect 5555 1005 5556 1035
rect 5524 1004 5556 1005
rect 5524 955 5556 956
rect 5524 925 5525 955
rect 5525 925 5555 955
rect 5555 925 5556 955
rect 5524 924 5556 925
rect 5524 875 5556 876
rect 5524 845 5525 875
rect 5525 845 5555 875
rect 5555 845 5556 875
rect 5524 844 5556 845
rect 5524 764 5556 796
rect 5524 684 5556 716
rect 5524 635 5556 636
rect 5524 605 5525 635
rect 5525 605 5555 635
rect 5555 605 5556 635
rect 5524 604 5556 605
rect 5524 555 5556 556
rect 5524 525 5525 555
rect 5525 525 5555 555
rect 5555 525 5556 555
rect 5524 524 5556 525
rect 5524 444 5556 476
rect 5524 395 5556 396
rect 5524 365 5525 395
rect 5525 365 5555 395
rect 5555 365 5556 395
rect 5524 364 5556 365
rect 5524 284 5556 316
rect 5524 235 5556 236
rect 5524 205 5525 235
rect 5525 205 5555 235
rect 5555 205 5556 235
rect 5524 204 5556 205
rect 5524 124 5556 156
rect 5524 75 5556 76
rect 5524 45 5525 75
rect 5525 45 5555 75
rect 5555 45 5556 75
rect 5524 44 5556 45
rect 5524 -5 5556 -4
rect 5524 -35 5525 -5
rect 5525 -35 5555 -5
rect 5555 -35 5556 -5
rect 5524 -36 5556 -35
rect 5524 -85 5556 -84
rect 5524 -115 5525 -85
rect 5525 -115 5555 -85
rect 5555 -115 5556 -85
rect 5524 -116 5556 -115
rect 5524 -165 5556 -164
rect 5524 -195 5525 -165
rect 5525 -195 5555 -165
rect 5555 -195 5556 -165
rect 5524 -196 5556 -195
rect 5524 -245 5556 -244
rect 5524 -275 5525 -245
rect 5525 -275 5555 -245
rect 5555 -275 5556 -245
rect 5524 -276 5556 -275
rect 5524 -325 5556 -324
rect 5524 -355 5525 -325
rect 5525 -355 5555 -325
rect 5555 -355 5556 -325
rect 5524 -356 5556 -355
rect 5524 -436 5556 -404
rect 5524 -485 5556 -484
rect 5524 -515 5525 -485
rect 5525 -515 5555 -485
rect 5555 -515 5556 -485
rect 5524 -516 5556 -515
rect 5524 -596 5556 -564
rect 5524 -645 5556 -644
rect 5524 -675 5525 -645
rect 5525 -675 5555 -645
rect 5555 -675 5556 -645
rect 5524 -676 5556 -675
rect 5524 -756 5556 -724
rect 5524 -805 5556 -804
rect 5524 -835 5525 -805
rect 5525 -835 5555 -805
rect 5555 -835 5556 -805
rect 5524 -836 5556 -835
rect 5524 -885 5556 -884
rect 5524 -915 5525 -885
rect 5525 -915 5555 -885
rect 5555 -915 5556 -885
rect 5524 -916 5556 -915
rect 5524 -996 5556 -964
rect 5524 -1076 5556 -1044
rect 5524 -1125 5556 -1124
rect 5524 -1155 5525 -1125
rect 5525 -1155 5555 -1125
rect 5555 -1155 5556 -1125
rect 5524 -1156 5556 -1155
rect 5524 -1205 5556 -1204
rect 5524 -1235 5525 -1205
rect 5525 -1235 5555 -1205
rect 5555 -1235 5556 -1205
rect 5524 -1236 5556 -1235
rect 5524 -1285 5556 -1284
rect 5524 -1315 5525 -1285
rect 5525 -1315 5555 -1285
rect 5555 -1315 5556 -1285
rect 5524 -1316 5556 -1315
rect 5524 -1365 5556 -1364
rect 5524 -1395 5525 -1365
rect 5525 -1395 5555 -1365
rect 5555 -1395 5556 -1365
rect 5524 -1396 5556 -1395
rect 5524 -1445 5556 -1444
rect 5524 -1475 5525 -1445
rect 5525 -1475 5555 -1445
rect 5555 -1475 5556 -1445
rect 5524 -1476 5556 -1475
rect 5524 -1525 5556 -1524
rect 5524 -1555 5525 -1525
rect 5525 -1555 5555 -1525
rect 5555 -1555 5556 -1525
rect 5524 -1556 5556 -1555
rect 5524 -1636 5556 -1604
rect 5524 -1716 5556 -1684
rect 5524 -1765 5556 -1764
rect 5524 -1795 5525 -1765
rect 5525 -1795 5555 -1765
rect 5555 -1795 5556 -1765
rect 5524 -1796 5556 -1795
rect 5524 -1845 5556 -1844
rect 5524 -1875 5525 -1845
rect 5525 -1875 5555 -1845
rect 5555 -1875 5556 -1845
rect 5524 -1876 5556 -1875
rect 5524 -1956 5556 -1924
rect 5524 -2005 5556 -2004
rect 5524 -2035 5525 -2005
rect 5525 -2035 5555 -2005
rect 5555 -2035 5556 -2005
rect 5524 -2036 5556 -2035
rect 5524 -2116 5556 -2084
rect 5524 -2165 5556 -2164
rect 5524 -2195 5525 -2165
rect 5525 -2195 5555 -2165
rect 5555 -2195 5556 -2165
rect 5524 -2196 5556 -2195
rect 5524 -2276 5556 -2244
rect 5524 -2325 5556 -2324
rect 5524 -2355 5525 -2325
rect 5525 -2355 5555 -2325
rect 5555 -2355 5556 -2325
rect 5524 -2356 5556 -2355
rect 5524 -2405 5556 -2404
rect 5524 -2435 5525 -2405
rect 5525 -2435 5555 -2405
rect 5555 -2435 5556 -2405
rect 5524 -2436 5556 -2435
rect 5524 -2485 5556 -2484
rect 5524 -2515 5525 -2485
rect 5525 -2515 5555 -2485
rect 5555 -2515 5556 -2485
rect 5524 -2516 5556 -2515
rect 5524 -2565 5556 -2564
rect 5524 -2595 5525 -2565
rect 5525 -2595 5555 -2565
rect 5555 -2595 5556 -2565
rect 5524 -2596 5556 -2595
rect 5524 -2645 5556 -2644
rect 5524 -2675 5525 -2645
rect 5525 -2675 5555 -2645
rect 5555 -2675 5556 -2645
rect 5524 -2676 5556 -2675
rect 5524 -2725 5556 -2724
rect 5524 -2755 5525 -2725
rect 5525 -2755 5555 -2725
rect 5555 -2755 5556 -2725
rect 5524 -2756 5556 -2755
rect 5524 -2836 5556 -2804
rect 5524 -2885 5556 -2884
rect 5524 -2915 5525 -2885
rect 5525 -2915 5555 -2885
rect 5555 -2915 5556 -2885
rect 5524 -2916 5556 -2915
rect 5524 -2996 5556 -2964
rect 5524 -3045 5556 -3044
rect 5524 -3075 5525 -3045
rect 5525 -3075 5555 -3045
rect 5555 -3075 5556 -3045
rect 5524 -3076 5556 -3075
rect 5524 -3156 5556 -3124
rect 5524 -3205 5556 -3204
rect 5524 -3235 5525 -3205
rect 5525 -3235 5555 -3205
rect 5555 -3235 5556 -3205
rect 5524 -3236 5556 -3235
rect 5524 -3285 5556 -3284
rect 5524 -3315 5525 -3285
rect 5525 -3315 5555 -3285
rect 5555 -3315 5556 -3285
rect 5524 -3316 5556 -3315
rect 5524 -3396 5556 -3364
rect 5524 -3476 5556 -3444
rect 5524 -3525 5556 -3524
rect 5524 -3555 5525 -3525
rect 5525 -3555 5555 -3525
rect 5555 -3555 5556 -3525
rect 5524 -3556 5556 -3555
rect 5524 -3605 5556 -3604
rect 5524 -3635 5525 -3605
rect 5525 -3635 5555 -3605
rect 5555 -3635 5556 -3605
rect 5524 -3636 5556 -3635
rect 5524 -3685 5556 -3684
rect 5524 -3715 5525 -3685
rect 5525 -3715 5555 -3685
rect 5555 -3715 5556 -3685
rect 5524 -3716 5556 -3715
rect 5604 1035 5636 1036
rect 5604 1005 5605 1035
rect 5605 1005 5635 1035
rect 5635 1005 5636 1035
rect 5604 1004 5636 1005
rect 5604 955 5636 956
rect 5604 925 5605 955
rect 5605 925 5635 955
rect 5635 925 5636 955
rect 5604 924 5636 925
rect 5604 875 5636 876
rect 5604 845 5605 875
rect 5605 845 5635 875
rect 5635 845 5636 875
rect 5604 844 5636 845
rect 5604 764 5636 796
rect 5604 684 5636 716
rect 5604 635 5636 636
rect 5604 605 5605 635
rect 5605 605 5635 635
rect 5635 605 5636 635
rect 5604 604 5636 605
rect 5604 555 5636 556
rect 5604 525 5605 555
rect 5605 525 5635 555
rect 5635 525 5636 555
rect 5604 524 5636 525
rect 5604 444 5636 476
rect 5604 395 5636 396
rect 5604 365 5605 395
rect 5605 365 5635 395
rect 5635 365 5636 395
rect 5604 364 5636 365
rect 5604 284 5636 316
rect 5604 235 5636 236
rect 5604 205 5605 235
rect 5605 205 5635 235
rect 5635 205 5636 235
rect 5604 204 5636 205
rect 5604 124 5636 156
rect 5604 75 5636 76
rect 5604 45 5605 75
rect 5605 45 5635 75
rect 5635 45 5636 75
rect 5604 44 5636 45
rect 5604 -5 5636 -4
rect 5604 -35 5605 -5
rect 5605 -35 5635 -5
rect 5635 -35 5636 -5
rect 5604 -36 5636 -35
rect 5604 -85 5636 -84
rect 5604 -115 5605 -85
rect 5605 -115 5635 -85
rect 5635 -115 5636 -85
rect 5604 -116 5636 -115
rect 5604 -165 5636 -164
rect 5604 -195 5605 -165
rect 5605 -195 5635 -165
rect 5635 -195 5636 -165
rect 5604 -196 5636 -195
rect 5604 -245 5636 -244
rect 5604 -275 5605 -245
rect 5605 -275 5635 -245
rect 5635 -275 5636 -245
rect 5604 -276 5636 -275
rect 5604 -325 5636 -324
rect 5604 -355 5605 -325
rect 5605 -355 5635 -325
rect 5635 -355 5636 -325
rect 5604 -356 5636 -355
rect 5604 -436 5636 -404
rect 5604 -485 5636 -484
rect 5604 -515 5605 -485
rect 5605 -515 5635 -485
rect 5635 -515 5636 -485
rect 5604 -516 5636 -515
rect 5604 -596 5636 -564
rect 5604 -645 5636 -644
rect 5604 -675 5605 -645
rect 5605 -675 5635 -645
rect 5635 -675 5636 -645
rect 5604 -676 5636 -675
rect 5604 -756 5636 -724
rect 5604 -805 5636 -804
rect 5604 -835 5605 -805
rect 5605 -835 5635 -805
rect 5635 -835 5636 -805
rect 5604 -836 5636 -835
rect 5604 -885 5636 -884
rect 5604 -915 5605 -885
rect 5605 -915 5635 -885
rect 5635 -915 5636 -885
rect 5604 -916 5636 -915
rect 5604 -996 5636 -964
rect 5604 -1076 5636 -1044
rect 5604 -1125 5636 -1124
rect 5604 -1155 5605 -1125
rect 5605 -1155 5635 -1125
rect 5635 -1155 5636 -1125
rect 5604 -1156 5636 -1155
rect 5604 -1205 5636 -1204
rect 5604 -1235 5605 -1205
rect 5605 -1235 5635 -1205
rect 5635 -1235 5636 -1205
rect 5604 -1236 5636 -1235
rect 5604 -1285 5636 -1284
rect 5604 -1315 5605 -1285
rect 5605 -1315 5635 -1285
rect 5635 -1315 5636 -1285
rect 5604 -1316 5636 -1315
rect 5604 -1365 5636 -1364
rect 5604 -1395 5605 -1365
rect 5605 -1395 5635 -1365
rect 5635 -1395 5636 -1365
rect 5604 -1396 5636 -1395
rect 5604 -1445 5636 -1444
rect 5604 -1475 5605 -1445
rect 5605 -1475 5635 -1445
rect 5635 -1475 5636 -1445
rect 5604 -1476 5636 -1475
rect 5604 -1525 5636 -1524
rect 5604 -1555 5605 -1525
rect 5605 -1555 5635 -1525
rect 5635 -1555 5636 -1525
rect 5604 -1556 5636 -1555
rect 5604 -1636 5636 -1604
rect 5604 -1716 5636 -1684
rect 5604 -1765 5636 -1764
rect 5604 -1795 5605 -1765
rect 5605 -1795 5635 -1765
rect 5635 -1795 5636 -1765
rect 5604 -1796 5636 -1795
rect 5604 -1845 5636 -1844
rect 5604 -1875 5605 -1845
rect 5605 -1875 5635 -1845
rect 5635 -1875 5636 -1845
rect 5604 -1876 5636 -1875
rect 5604 -1956 5636 -1924
rect 5604 -2005 5636 -2004
rect 5604 -2035 5605 -2005
rect 5605 -2035 5635 -2005
rect 5635 -2035 5636 -2005
rect 5604 -2036 5636 -2035
rect 5604 -2116 5636 -2084
rect 5604 -2165 5636 -2164
rect 5604 -2195 5605 -2165
rect 5605 -2195 5635 -2165
rect 5635 -2195 5636 -2165
rect 5604 -2196 5636 -2195
rect 5604 -2276 5636 -2244
rect 5604 -2325 5636 -2324
rect 5604 -2355 5605 -2325
rect 5605 -2355 5635 -2325
rect 5635 -2355 5636 -2325
rect 5604 -2356 5636 -2355
rect 5604 -2405 5636 -2404
rect 5604 -2435 5605 -2405
rect 5605 -2435 5635 -2405
rect 5635 -2435 5636 -2405
rect 5604 -2436 5636 -2435
rect 5604 -2485 5636 -2484
rect 5604 -2515 5605 -2485
rect 5605 -2515 5635 -2485
rect 5635 -2515 5636 -2485
rect 5604 -2516 5636 -2515
rect 5604 -2565 5636 -2564
rect 5604 -2595 5605 -2565
rect 5605 -2595 5635 -2565
rect 5635 -2595 5636 -2565
rect 5604 -2596 5636 -2595
rect 5604 -2645 5636 -2644
rect 5604 -2675 5605 -2645
rect 5605 -2675 5635 -2645
rect 5635 -2675 5636 -2645
rect 5604 -2676 5636 -2675
rect 5604 -2725 5636 -2724
rect 5604 -2755 5605 -2725
rect 5605 -2755 5635 -2725
rect 5635 -2755 5636 -2725
rect 5604 -2756 5636 -2755
rect 5604 -2836 5636 -2804
rect 5604 -2885 5636 -2884
rect 5604 -2915 5605 -2885
rect 5605 -2915 5635 -2885
rect 5635 -2915 5636 -2885
rect 5604 -2916 5636 -2915
rect 5604 -2996 5636 -2964
rect 5604 -3045 5636 -3044
rect 5604 -3075 5605 -3045
rect 5605 -3075 5635 -3045
rect 5635 -3075 5636 -3045
rect 5604 -3076 5636 -3075
rect 5604 -3156 5636 -3124
rect 5604 -3205 5636 -3204
rect 5604 -3235 5605 -3205
rect 5605 -3235 5635 -3205
rect 5635 -3235 5636 -3205
rect 5604 -3236 5636 -3235
rect 5604 -3285 5636 -3284
rect 5604 -3315 5605 -3285
rect 5605 -3315 5635 -3285
rect 5635 -3315 5636 -3285
rect 5604 -3316 5636 -3315
rect 5604 -3396 5636 -3364
rect 5604 -3476 5636 -3444
rect 5604 -3525 5636 -3524
rect 5604 -3555 5605 -3525
rect 5605 -3555 5635 -3525
rect 5635 -3555 5636 -3525
rect 5604 -3556 5636 -3555
rect 5604 -3605 5636 -3604
rect 5604 -3635 5605 -3605
rect 5605 -3635 5635 -3605
rect 5635 -3635 5636 -3605
rect 5604 -3636 5636 -3635
rect 5604 -3685 5636 -3684
rect 5604 -3715 5605 -3685
rect 5605 -3715 5635 -3685
rect 5635 -3715 5636 -3685
rect 5604 -3716 5636 -3715
rect 5684 1035 5716 1036
rect 5684 1005 5685 1035
rect 5685 1005 5715 1035
rect 5715 1005 5716 1035
rect 5684 1004 5716 1005
rect 5684 955 5716 956
rect 5684 925 5685 955
rect 5685 925 5715 955
rect 5715 925 5716 955
rect 5684 924 5716 925
rect 5684 875 5716 876
rect 5684 845 5685 875
rect 5685 845 5715 875
rect 5715 845 5716 875
rect 5684 844 5716 845
rect 5684 764 5716 796
rect 5684 684 5716 716
rect 5684 635 5716 636
rect 5684 605 5685 635
rect 5685 605 5715 635
rect 5715 605 5716 635
rect 5684 604 5716 605
rect 5684 555 5716 556
rect 5684 525 5685 555
rect 5685 525 5715 555
rect 5715 525 5716 555
rect 5684 524 5716 525
rect 5684 444 5716 476
rect 5684 395 5716 396
rect 5684 365 5685 395
rect 5685 365 5715 395
rect 5715 365 5716 395
rect 5684 364 5716 365
rect 5684 284 5716 316
rect 5684 235 5716 236
rect 5684 205 5685 235
rect 5685 205 5715 235
rect 5715 205 5716 235
rect 5684 204 5716 205
rect 5684 124 5716 156
rect 5684 75 5716 76
rect 5684 45 5685 75
rect 5685 45 5715 75
rect 5715 45 5716 75
rect 5684 44 5716 45
rect 5684 -5 5716 -4
rect 5684 -35 5685 -5
rect 5685 -35 5715 -5
rect 5715 -35 5716 -5
rect 5684 -36 5716 -35
rect 5684 -85 5716 -84
rect 5684 -115 5685 -85
rect 5685 -115 5715 -85
rect 5715 -115 5716 -85
rect 5684 -116 5716 -115
rect 5684 -165 5716 -164
rect 5684 -195 5685 -165
rect 5685 -195 5715 -165
rect 5715 -195 5716 -165
rect 5684 -196 5716 -195
rect 5684 -245 5716 -244
rect 5684 -275 5685 -245
rect 5685 -275 5715 -245
rect 5715 -275 5716 -245
rect 5684 -276 5716 -275
rect 5684 -325 5716 -324
rect 5684 -355 5685 -325
rect 5685 -355 5715 -325
rect 5715 -355 5716 -325
rect 5684 -356 5716 -355
rect 5684 -436 5716 -404
rect 5684 -485 5716 -484
rect 5684 -515 5685 -485
rect 5685 -515 5715 -485
rect 5715 -515 5716 -485
rect 5684 -516 5716 -515
rect 5684 -596 5716 -564
rect 5684 -645 5716 -644
rect 5684 -675 5685 -645
rect 5685 -675 5715 -645
rect 5715 -675 5716 -645
rect 5684 -676 5716 -675
rect 5684 -756 5716 -724
rect 5684 -805 5716 -804
rect 5684 -835 5685 -805
rect 5685 -835 5715 -805
rect 5715 -835 5716 -805
rect 5684 -836 5716 -835
rect 5684 -885 5716 -884
rect 5684 -915 5685 -885
rect 5685 -915 5715 -885
rect 5715 -915 5716 -885
rect 5684 -916 5716 -915
rect 5684 -996 5716 -964
rect 5684 -1076 5716 -1044
rect 5684 -1125 5716 -1124
rect 5684 -1155 5685 -1125
rect 5685 -1155 5715 -1125
rect 5715 -1155 5716 -1125
rect 5684 -1156 5716 -1155
rect 5684 -1205 5716 -1204
rect 5684 -1235 5685 -1205
rect 5685 -1235 5715 -1205
rect 5715 -1235 5716 -1205
rect 5684 -1236 5716 -1235
rect 5684 -1285 5716 -1284
rect 5684 -1315 5685 -1285
rect 5685 -1315 5715 -1285
rect 5715 -1315 5716 -1285
rect 5684 -1316 5716 -1315
rect 5684 -1365 5716 -1364
rect 5684 -1395 5685 -1365
rect 5685 -1395 5715 -1365
rect 5715 -1395 5716 -1365
rect 5684 -1396 5716 -1395
rect 5684 -1445 5716 -1444
rect 5684 -1475 5685 -1445
rect 5685 -1475 5715 -1445
rect 5715 -1475 5716 -1445
rect 5684 -1476 5716 -1475
rect 5684 -1525 5716 -1524
rect 5684 -1555 5685 -1525
rect 5685 -1555 5715 -1525
rect 5715 -1555 5716 -1525
rect 5684 -1556 5716 -1555
rect 5684 -1636 5716 -1604
rect 5684 -1716 5716 -1684
rect 5684 -1765 5716 -1764
rect 5684 -1795 5685 -1765
rect 5685 -1795 5715 -1765
rect 5715 -1795 5716 -1765
rect 5684 -1796 5716 -1795
rect 5684 -1845 5716 -1844
rect 5684 -1875 5685 -1845
rect 5685 -1875 5715 -1845
rect 5715 -1875 5716 -1845
rect 5684 -1876 5716 -1875
rect 5684 -1956 5716 -1924
rect 5684 -2005 5716 -2004
rect 5684 -2035 5685 -2005
rect 5685 -2035 5715 -2005
rect 5715 -2035 5716 -2005
rect 5684 -2036 5716 -2035
rect 5684 -2116 5716 -2084
rect 5684 -2165 5716 -2164
rect 5684 -2195 5685 -2165
rect 5685 -2195 5715 -2165
rect 5715 -2195 5716 -2165
rect 5684 -2196 5716 -2195
rect 5684 -2276 5716 -2244
rect 5684 -2325 5716 -2324
rect 5684 -2355 5685 -2325
rect 5685 -2355 5715 -2325
rect 5715 -2355 5716 -2325
rect 5684 -2356 5716 -2355
rect 5684 -2405 5716 -2404
rect 5684 -2435 5685 -2405
rect 5685 -2435 5715 -2405
rect 5715 -2435 5716 -2405
rect 5684 -2436 5716 -2435
rect 5684 -2485 5716 -2484
rect 5684 -2515 5685 -2485
rect 5685 -2515 5715 -2485
rect 5715 -2515 5716 -2485
rect 5684 -2516 5716 -2515
rect 5684 -2565 5716 -2564
rect 5684 -2595 5685 -2565
rect 5685 -2595 5715 -2565
rect 5715 -2595 5716 -2565
rect 5684 -2596 5716 -2595
rect 5684 -2645 5716 -2644
rect 5684 -2675 5685 -2645
rect 5685 -2675 5715 -2645
rect 5715 -2675 5716 -2645
rect 5684 -2676 5716 -2675
rect 5684 -2725 5716 -2724
rect 5684 -2755 5685 -2725
rect 5685 -2755 5715 -2725
rect 5715 -2755 5716 -2725
rect 5684 -2756 5716 -2755
rect 5684 -2836 5716 -2804
rect 5684 -2885 5716 -2884
rect 5684 -2915 5685 -2885
rect 5685 -2915 5715 -2885
rect 5715 -2915 5716 -2885
rect 5684 -2916 5716 -2915
rect 5684 -2996 5716 -2964
rect 5684 -3045 5716 -3044
rect 5684 -3075 5685 -3045
rect 5685 -3075 5715 -3045
rect 5715 -3075 5716 -3045
rect 5684 -3076 5716 -3075
rect 5684 -3156 5716 -3124
rect 5684 -3205 5716 -3204
rect 5684 -3235 5685 -3205
rect 5685 -3235 5715 -3205
rect 5715 -3235 5716 -3205
rect 5684 -3236 5716 -3235
rect 5684 -3285 5716 -3284
rect 5684 -3315 5685 -3285
rect 5685 -3315 5715 -3285
rect 5715 -3315 5716 -3285
rect 5684 -3316 5716 -3315
rect 5684 -3396 5716 -3364
rect 5684 -3476 5716 -3444
rect 5684 -3525 5716 -3524
rect 5684 -3555 5685 -3525
rect 5685 -3555 5715 -3525
rect 5715 -3555 5716 -3525
rect 5684 -3556 5716 -3555
rect 5684 -3605 5716 -3604
rect 5684 -3635 5685 -3605
rect 5685 -3635 5715 -3605
rect 5715 -3635 5716 -3605
rect 5684 -3636 5716 -3635
rect 5684 -3685 5716 -3684
rect 5684 -3715 5685 -3685
rect 5685 -3715 5715 -3685
rect 5715 -3715 5716 -3685
rect 5684 -3716 5716 -3715
rect 5764 1035 5796 1036
rect 5764 1005 5765 1035
rect 5765 1005 5795 1035
rect 5795 1005 5796 1035
rect 5764 1004 5796 1005
rect 5764 955 5796 956
rect 5764 925 5765 955
rect 5765 925 5795 955
rect 5795 925 5796 955
rect 5764 924 5796 925
rect 5764 875 5796 876
rect 5764 845 5765 875
rect 5765 845 5795 875
rect 5795 845 5796 875
rect 5764 844 5796 845
rect 5764 764 5796 796
rect 5764 684 5796 716
rect 5764 635 5796 636
rect 5764 605 5765 635
rect 5765 605 5795 635
rect 5795 605 5796 635
rect 5764 604 5796 605
rect 5764 555 5796 556
rect 5764 525 5765 555
rect 5765 525 5795 555
rect 5795 525 5796 555
rect 5764 524 5796 525
rect 5764 444 5796 476
rect 5764 395 5796 396
rect 5764 365 5765 395
rect 5765 365 5795 395
rect 5795 365 5796 395
rect 5764 364 5796 365
rect 5764 284 5796 316
rect 5764 235 5796 236
rect 5764 205 5765 235
rect 5765 205 5795 235
rect 5795 205 5796 235
rect 5764 204 5796 205
rect 5764 124 5796 156
rect 5764 75 5796 76
rect 5764 45 5765 75
rect 5765 45 5795 75
rect 5795 45 5796 75
rect 5764 44 5796 45
rect 5764 -5 5796 -4
rect 5764 -35 5765 -5
rect 5765 -35 5795 -5
rect 5795 -35 5796 -5
rect 5764 -36 5796 -35
rect 5764 -85 5796 -84
rect 5764 -115 5765 -85
rect 5765 -115 5795 -85
rect 5795 -115 5796 -85
rect 5764 -116 5796 -115
rect 5764 -165 5796 -164
rect 5764 -195 5765 -165
rect 5765 -195 5795 -165
rect 5795 -195 5796 -165
rect 5764 -196 5796 -195
rect 5764 -245 5796 -244
rect 5764 -275 5765 -245
rect 5765 -275 5795 -245
rect 5795 -275 5796 -245
rect 5764 -276 5796 -275
rect 5764 -325 5796 -324
rect 5764 -355 5765 -325
rect 5765 -355 5795 -325
rect 5795 -355 5796 -325
rect 5764 -356 5796 -355
rect 5764 -436 5796 -404
rect 5764 -485 5796 -484
rect 5764 -515 5765 -485
rect 5765 -515 5795 -485
rect 5795 -515 5796 -485
rect 5764 -516 5796 -515
rect 5764 -596 5796 -564
rect 5764 -645 5796 -644
rect 5764 -675 5765 -645
rect 5765 -675 5795 -645
rect 5795 -675 5796 -645
rect 5764 -676 5796 -675
rect 5764 -756 5796 -724
rect 5764 -805 5796 -804
rect 5764 -835 5765 -805
rect 5765 -835 5795 -805
rect 5795 -835 5796 -805
rect 5764 -836 5796 -835
rect 5764 -885 5796 -884
rect 5764 -915 5765 -885
rect 5765 -915 5795 -885
rect 5795 -915 5796 -885
rect 5764 -916 5796 -915
rect 5764 -996 5796 -964
rect 5764 -1076 5796 -1044
rect 5764 -1125 5796 -1124
rect 5764 -1155 5765 -1125
rect 5765 -1155 5795 -1125
rect 5795 -1155 5796 -1125
rect 5764 -1156 5796 -1155
rect 5764 -1205 5796 -1204
rect 5764 -1235 5765 -1205
rect 5765 -1235 5795 -1205
rect 5795 -1235 5796 -1205
rect 5764 -1236 5796 -1235
rect 5764 -1285 5796 -1284
rect 5764 -1315 5765 -1285
rect 5765 -1315 5795 -1285
rect 5795 -1315 5796 -1285
rect 5764 -1316 5796 -1315
rect 5764 -1365 5796 -1364
rect 5764 -1395 5765 -1365
rect 5765 -1395 5795 -1365
rect 5795 -1395 5796 -1365
rect 5764 -1396 5796 -1395
rect 5764 -1445 5796 -1444
rect 5764 -1475 5765 -1445
rect 5765 -1475 5795 -1445
rect 5795 -1475 5796 -1445
rect 5764 -1476 5796 -1475
rect 5764 -1525 5796 -1524
rect 5764 -1555 5765 -1525
rect 5765 -1555 5795 -1525
rect 5795 -1555 5796 -1525
rect 5764 -1556 5796 -1555
rect 5764 -1636 5796 -1604
rect 5764 -1716 5796 -1684
rect 5764 -1765 5796 -1764
rect 5764 -1795 5765 -1765
rect 5765 -1795 5795 -1765
rect 5795 -1795 5796 -1765
rect 5764 -1796 5796 -1795
rect 5764 -1845 5796 -1844
rect 5764 -1875 5765 -1845
rect 5765 -1875 5795 -1845
rect 5795 -1875 5796 -1845
rect 5764 -1876 5796 -1875
rect 5764 -1956 5796 -1924
rect 5764 -2005 5796 -2004
rect 5764 -2035 5765 -2005
rect 5765 -2035 5795 -2005
rect 5795 -2035 5796 -2005
rect 5764 -2036 5796 -2035
rect 5764 -2116 5796 -2084
rect 5764 -2165 5796 -2164
rect 5764 -2195 5765 -2165
rect 5765 -2195 5795 -2165
rect 5795 -2195 5796 -2165
rect 5764 -2196 5796 -2195
rect 5764 -2276 5796 -2244
rect 5764 -2325 5796 -2324
rect 5764 -2355 5765 -2325
rect 5765 -2355 5795 -2325
rect 5795 -2355 5796 -2325
rect 5764 -2356 5796 -2355
rect 5764 -2405 5796 -2404
rect 5764 -2435 5765 -2405
rect 5765 -2435 5795 -2405
rect 5795 -2435 5796 -2405
rect 5764 -2436 5796 -2435
rect 5764 -2485 5796 -2484
rect 5764 -2515 5765 -2485
rect 5765 -2515 5795 -2485
rect 5795 -2515 5796 -2485
rect 5764 -2516 5796 -2515
rect 5764 -2565 5796 -2564
rect 5764 -2595 5765 -2565
rect 5765 -2595 5795 -2565
rect 5795 -2595 5796 -2565
rect 5764 -2596 5796 -2595
rect 5764 -2645 5796 -2644
rect 5764 -2675 5765 -2645
rect 5765 -2675 5795 -2645
rect 5795 -2675 5796 -2645
rect 5764 -2676 5796 -2675
rect 5764 -2725 5796 -2724
rect 5764 -2755 5765 -2725
rect 5765 -2755 5795 -2725
rect 5795 -2755 5796 -2725
rect 5764 -2756 5796 -2755
rect 5764 -2836 5796 -2804
rect 5764 -2885 5796 -2884
rect 5764 -2915 5765 -2885
rect 5765 -2915 5795 -2885
rect 5795 -2915 5796 -2885
rect 5764 -2916 5796 -2915
rect 5764 -2996 5796 -2964
rect 5764 -3045 5796 -3044
rect 5764 -3075 5765 -3045
rect 5765 -3075 5795 -3045
rect 5795 -3075 5796 -3045
rect 5764 -3076 5796 -3075
rect 5764 -3156 5796 -3124
rect 5764 -3205 5796 -3204
rect 5764 -3235 5765 -3205
rect 5765 -3235 5795 -3205
rect 5795 -3235 5796 -3205
rect 5764 -3236 5796 -3235
rect 5764 -3285 5796 -3284
rect 5764 -3315 5765 -3285
rect 5765 -3315 5795 -3285
rect 5795 -3315 5796 -3285
rect 5764 -3316 5796 -3315
rect 5764 -3396 5796 -3364
rect 5764 -3476 5796 -3444
rect 5764 -3525 5796 -3524
rect 5764 -3555 5765 -3525
rect 5765 -3555 5795 -3525
rect 5795 -3555 5796 -3525
rect 5764 -3556 5796 -3555
rect 5764 -3605 5796 -3604
rect 5764 -3635 5765 -3605
rect 5765 -3635 5795 -3605
rect 5795 -3635 5796 -3605
rect 5764 -3636 5796 -3635
rect 5764 -3685 5796 -3684
rect 5764 -3715 5765 -3685
rect 5765 -3715 5795 -3685
rect 5795 -3715 5796 -3685
rect 5764 -3716 5796 -3715
rect 5844 1035 5876 1036
rect 5844 1005 5845 1035
rect 5845 1005 5875 1035
rect 5875 1005 5876 1035
rect 5844 1004 5876 1005
rect 5844 955 5876 956
rect 5844 925 5845 955
rect 5845 925 5875 955
rect 5875 925 5876 955
rect 5844 924 5876 925
rect 5844 875 5876 876
rect 5844 845 5845 875
rect 5845 845 5875 875
rect 5875 845 5876 875
rect 5844 844 5876 845
rect 5844 764 5876 796
rect 5844 684 5876 716
rect 5844 635 5876 636
rect 5844 605 5845 635
rect 5845 605 5875 635
rect 5875 605 5876 635
rect 5844 604 5876 605
rect 5844 555 5876 556
rect 5844 525 5845 555
rect 5845 525 5875 555
rect 5875 525 5876 555
rect 5844 524 5876 525
rect 5844 444 5876 476
rect 5844 395 5876 396
rect 5844 365 5845 395
rect 5845 365 5875 395
rect 5875 365 5876 395
rect 5844 364 5876 365
rect 5844 284 5876 316
rect 5844 235 5876 236
rect 5844 205 5845 235
rect 5845 205 5875 235
rect 5875 205 5876 235
rect 5844 204 5876 205
rect 5844 124 5876 156
rect 5844 75 5876 76
rect 5844 45 5845 75
rect 5845 45 5875 75
rect 5875 45 5876 75
rect 5844 44 5876 45
rect 5844 -5 5876 -4
rect 5844 -35 5845 -5
rect 5845 -35 5875 -5
rect 5875 -35 5876 -5
rect 5844 -36 5876 -35
rect 5844 -85 5876 -84
rect 5844 -115 5845 -85
rect 5845 -115 5875 -85
rect 5875 -115 5876 -85
rect 5844 -116 5876 -115
rect 5844 -165 5876 -164
rect 5844 -195 5845 -165
rect 5845 -195 5875 -165
rect 5875 -195 5876 -165
rect 5844 -196 5876 -195
rect 5844 -245 5876 -244
rect 5844 -275 5845 -245
rect 5845 -275 5875 -245
rect 5875 -275 5876 -245
rect 5844 -276 5876 -275
rect 5844 -325 5876 -324
rect 5844 -355 5845 -325
rect 5845 -355 5875 -325
rect 5875 -355 5876 -325
rect 5844 -356 5876 -355
rect 5844 -436 5876 -404
rect 5844 -485 5876 -484
rect 5844 -515 5845 -485
rect 5845 -515 5875 -485
rect 5875 -515 5876 -485
rect 5844 -516 5876 -515
rect 5844 -596 5876 -564
rect 5844 -645 5876 -644
rect 5844 -675 5845 -645
rect 5845 -675 5875 -645
rect 5875 -675 5876 -645
rect 5844 -676 5876 -675
rect 5844 -756 5876 -724
rect 5844 -805 5876 -804
rect 5844 -835 5845 -805
rect 5845 -835 5875 -805
rect 5875 -835 5876 -805
rect 5844 -836 5876 -835
rect 5844 -885 5876 -884
rect 5844 -915 5845 -885
rect 5845 -915 5875 -885
rect 5875 -915 5876 -885
rect 5844 -916 5876 -915
rect 5844 -996 5876 -964
rect 5844 -1076 5876 -1044
rect 5844 -1125 5876 -1124
rect 5844 -1155 5845 -1125
rect 5845 -1155 5875 -1125
rect 5875 -1155 5876 -1125
rect 5844 -1156 5876 -1155
rect 5844 -1205 5876 -1204
rect 5844 -1235 5845 -1205
rect 5845 -1235 5875 -1205
rect 5875 -1235 5876 -1205
rect 5844 -1236 5876 -1235
rect 5844 -1285 5876 -1284
rect 5844 -1315 5845 -1285
rect 5845 -1315 5875 -1285
rect 5875 -1315 5876 -1285
rect 5844 -1316 5876 -1315
rect 5844 -1365 5876 -1364
rect 5844 -1395 5845 -1365
rect 5845 -1395 5875 -1365
rect 5875 -1395 5876 -1365
rect 5844 -1396 5876 -1395
rect 5844 -1445 5876 -1444
rect 5844 -1475 5845 -1445
rect 5845 -1475 5875 -1445
rect 5875 -1475 5876 -1445
rect 5844 -1476 5876 -1475
rect 5844 -1525 5876 -1524
rect 5844 -1555 5845 -1525
rect 5845 -1555 5875 -1525
rect 5875 -1555 5876 -1525
rect 5844 -1556 5876 -1555
rect 5844 -1636 5876 -1604
rect 5844 -1716 5876 -1684
rect 5844 -1765 5876 -1764
rect 5844 -1795 5845 -1765
rect 5845 -1795 5875 -1765
rect 5875 -1795 5876 -1765
rect 5844 -1796 5876 -1795
rect 5844 -1845 5876 -1844
rect 5844 -1875 5845 -1845
rect 5845 -1875 5875 -1845
rect 5875 -1875 5876 -1845
rect 5844 -1876 5876 -1875
rect 5844 -1956 5876 -1924
rect 5844 -2005 5876 -2004
rect 5844 -2035 5845 -2005
rect 5845 -2035 5875 -2005
rect 5875 -2035 5876 -2005
rect 5844 -2036 5876 -2035
rect 5844 -2116 5876 -2084
rect 5844 -2165 5876 -2164
rect 5844 -2195 5845 -2165
rect 5845 -2195 5875 -2165
rect 5875 -2195 5876 -2165
rect 5844 -2196 5876 -2195
rect 5844 -2276 5876 -2244
rect 5844 -2325 5876 -2324
rect 5844 -2355 5845 -2325
rect 5845 -2355 5875 -2325
rect 5875 -2355 5876 -2325
rect 5844 -2356 5876 -2355
rect 5844 -2405 5876 -2404
rect 5844 -2435 5845 -2405
rect 5845 -2435 5875 -2405
rect 5875 -2435 5876 -2405
rect 5844 -2436 5876 -2435
rect 5844 -2485 5876 -2484
rect 5844 -2515 5845 -2485
rect 5845 -2515 5875 -2485
rect 5875 -2515 5876 -2485
rect 5844 -2516 5876 -2515
rect 5844 -2565 5876 -2564
rect 5844 -2595 5845 -2565
rect 5845 -2595 5875 -2565
rect 5875 -2595 5876 -2565
rect 5844 -2596 5876 -2595
rect 5844 -2645 5876 -2644
rect 5844 -2675 5845 -2645
rect 5845 -2675 5875 -2645
rect 5875 -2675 5876 -2645
rect 5844 -2676 5876 -2675
rect 5844 -2725 5876 -2724
rect 5844 -2755 5845 -2725
rect 5845 -2755 5875 -2725
rect 5875 -2755 5876 -2725
rect 5844 -2756 5876 -2755
rect 5844 -2836 5876 -2804
rect 5844 -2885 5876 -2884
rect 5844 -2915 5845 -2885
rect 5845 -2915 5875 -2885
rect 5875 -2915 5876 -2885
rect 5844 -2916 5876 -2915
rect 5844 -2996 5876 -2964
rect 5844 -3045 5876 -3044
rect 5844 -3075 5845 -3045
rect 5845 -3075 5875 -3045
rect 5875 -3075 5876 -3045
rect 5844 -3076 5876 -3075
rect 5844 -3156 5876 -3124
rect 5844 -3205 5876 -3204
rect 5844 -3235 5845 -3205
rect 5845 -3235 5875 -3205
rect 5875 -3235 5876 -3205
rect 5844 -3236 5876 -3235
rect 5844 -3285 5876 -3284
rect 5844 -3315 5845 -3285
rect 5845 -3315 5875 -3285
rect 5875 -3315 5876 -3285
rect 5844 -3316 5876 -3315
rect 5844 -3396 5876 -3364
rect 5844 -3476 5876 -3444
rect 5844 -3525 5876 -3524
rect 5844 -3555 5845 -3525
rect 5845 -3555 5875 -3525
rect 5875 -3555 5876 -3525
rect 5844 -3556 5876 -3555
rect 5844 -3605 5876 -3604
rect 5844 -3635 5845 -3605
rect 5845 -3635 5875 -3605
rect 5875 -3635 5876 -3605
rect 5844 -3636 5876 -3635
rect 5844 -3685 5876 -3684
rect 5844 -3715 5845 -3685
rect 5845 -3715 5875 -3685
rect 5875 -3715 5876 -3685
rect 5844 -3716 5876 -3715
rect 5924 1035 5956 1036
rect 5924 1005 5925 1035
rect 5925 1005 5955 1035
rect 5955 1005 5956 1035
rect 5924 1004 5956 1005
rect 5924 955 5956 956
rect 5924 925 5925 955
rect 5925 925 5955 955
rect 5955 925 5956 955
rect 5924 924 5956 925
rect 5924 875 5956 876
rect 5924 845 5925 875
rect 5925 845 5955 875
rect 5955 845 5956 875
rect 5924 844 5956 845
rect 5924 764 5956 796
rect 5924 684 5956 716
rect 5924 635 5956 636
rect 5924 605 5925 635
rect 5925 605 5955 635
rect 5955 605 5956 635
rect 5924 604 5956 605
rect 5924 555 5956 556
rect 5924 525 5925 555
rect 5925 525 5955 555
rect 5955 525 5956 555
rect 5924 524 5956 525
rect 5924 444 5956 476
rect 5924 395 5956 396
rect 5924 365 5925 395
rect 5925 365 5955 395
rect 5955 365 5956 395
rect 5924 364 5956 365
rect 5924 284 5956 316
rect 5924 235 5956 236
rect 5924 205 5925 235
rect 5925 205 5955 235
rect 5955 205 5956 235
rect 5924 204 5956 205
rect 5924 124 5956 156
rect 5924 75 5956 76
rect 5924 45 5925 75
rect 5925 45 5955 75
rect 5955 45 5956 75
rect 5924 44 5956 45
rect 5924 -5 5956 -4
rect 5924 -35 5925 -5
rect 5925 -35 5955 -5
rect 5955 -35 5956 -5
rect 5924 -36 5956 -35
rect 5924 -85 5956 -84
rect 5924 -115 5925 -85
rect 5925 -115 5955 -85
rect 5955 -115 5956 -85
rect 5924 -116 5956 -115
rect 5924 -165 5956 -164
rect 5924 -195 5925 -165
rect 5925 -195 5955 -165
rect 5955 -195 5956 -165
rect 5924 -196 5956 -195
rect 5924 -245 5956 -244
rect 5924 -275 5925 -245
rect 5925 -275 5955 -245
rect 5955 -275 5956 -245
rect 5924 -276 5956 -275
rect 5924 -325 5956 -324
rect 5924 -355 5925 -325
rect 5925 -355 5955 -325
rect 5955 -355 5956 -325
rect 5924 -356 5956 -355
rect 5924 -436 5956 -404
rect 5924 -485 5956 -484
rect 5924 -515 5925 -485
rect 5925 -515 5955 -485
rect 5955 -515 5956 -485
rect 5924 -516 5956 -515
rect 5924 -596 5956 -564
rect 5924 -645 5956 -644
rect 5924 -675 5925 -645
rect 5925 -675 5955 -645
rect 5955 -675 5956 -645
rect 5924 -676 5956 -675
rect 5924 -756 5956 -724
rect 5924 -805 5956 -804
rect 5924 -835 5925 -805
rect 5925 -835 5955 -805
rect 5955 -835 5956 -805
rect 5924 -836 5956 -835
rect 5924 -885 5956 -884
rect 5924 -915 5925 -885
rect 5925 -915 5955 -885
rect 5955 -915 5956 -885
rect 5924 -916 5956 -915
rect 5924 -996 5956 -964
rect 5924 -1076 5956 -1044
rect 5924 -1125 5956 -1124
rect 5924 -1155 5925 -1125
rect 5925 -1155 5955 -1125
rect 5955 -1155 5956 -1125
rect 5924 -1156 5956 -1155
rect 5924 -1205 5956 -1204
rect 5924 -1235 5925 -1205
rect 5925 -1235 5955 -1205
rect 5955 -1235 5956 -1205
rect 5924 -1236 5956 -1235
rect 5924 -1285 5956 -1284
rect 5924 -1315 5925 -1285
rect 5925 -1315 5955 -1285
rect 5955 -1315 5956 -1285
rect 5924 -1316 5956 -1315
rect 5924 -1365 5956 -1364
rect 5924 -1395 5925 -1365
rect 5925 -1395 5955 -1365
rect 5955 -1395 5956 -1365
rect 5924 -1396 5956 -1395
rect 5924 -1445 5956 -1444
rect 5924 -1475 5925 -1445
rect 5925 -1475 5955 -1445
rect 5955 -1475 5956 -1445
rect 5924 -1476 5956 -1475
rect 5924 -1525 5956 -1524
rect 5924 -1555 5925 -1525
rect 5925 -1555 5955 -1525
rect 5955 -1555 5956 -1525
rect 5924 -1556 5956 -1555
rect 5924 -1636 5956 -1604
rect 5924 -1716 5956 -1684
rect 5924 -1765 5956 -1764
rect 5924 -1795 5925 -1765
rect 5925 -1795 5955 -1765
rect 5955 -1795 5956 -1765
rect 5924 -1796 5956 -1795
rect 5924 -1845 5956 -1844
rect 5924 -1875 5925 -1845
rect 5925 -1875 5955 -1845
rect 5955 -1875 5956 -1845
rect 5924 -1876 5956 -1875
rect 5924 -1956 5956 -1924
rect 5924 -2005 5956 -2004
rect 5924 -2035 5925 -2005
rect 5925 -2035 5955 -2005
rect 5955 -2035 5956 -2005
rect 5924 -2036 5956 -2035
rect 5924 -2116 5956 -2084
rect 5924 -2165 5956 -2164
rect 5924 -2195 5925 -2165
rect 5925 -2195 5955 -2165
rect 5955 -2195 5956 -2165
rect 5924 -2196 5956 -2195
rect 5924 -2276 5956 -2244
rect 5924 -2325 5956 -2324
rect 5924 -2355 5925 -2325
rect 5925 -2355 5955 -2325
rect 5955 -2355 5956 -2325
rect 5924 -2356 5956 -2355
rect 5924 -2405 5956 -2404
rect 5924 -2435 5925 -2405
rect 5925 -2435 5955 -2405
rect 5955 -2435 5956 -2405
rect 5924 -2436 5956 -2435
rect 5924 -2485 5956 -2484
rect 5924 -2515 5925 -2485
rect 5925 -2515 5955 -2485
rect 5955 -2515 5956 -2485
rect 5924 -2516 5956 -2515
rect 5924 -2565 5956 -2564
rect 5924 -2595 5925 -2565
rect 5925 -2595 5955 -2565
rect 5955 -2595 5956 -2565
rect 5924 -2596 5956 -2595
rect 5924 -2645 5956 -2644
rect 5924 -2675 5925 -2645
rect 5925 -2675 5955 -2645
rect 5955 -2675 5956 -2645
rect 5924 -2676 5956 -2675
rect 5924 -2725 5956 -2724
rect 5924 -2755 5925 -2725
rect 5925 -2755 5955 -2725
rect 5955 -2755 5956 -2725
rect 5924 -2756 5956 -2755
rect 5924 -2836 5956 -2804
rect 5924 -2885 5956 -2884
rect 5924 -2915 5925 -2885
rect 5925 -2915 5955 -2885
rect 5955 -2915 5956 -2885
rect 5924 -2916 5956 -2915
rect 5924 -2996 5956 -2964
rect 5924 -3045 5956 -3044
rect 5924 -3075 5925 -3045
rect 5925 -3075 5955 -3045
rect 5955 -3075 5956 -3045
rect 5924 -3076 5956 -3075
rect 5924 -3156 5956 -3124
rect 5924 -3205 5956 -3204
rect 5924 -3235 5925 -3205
rect 5925 -3235 5955 -3205
rect 5955 -3235 5956 -3205
rect 5924 -3236 5956 -3235
rect 5924 -3285 5956 -3284
rect 5924 -3315 5925 -3285
rect 5925 -3315 5955 -3285
rect 5955 -3315 5956 -3285
rect 5924 -3316 5956 -3315
rect 5924 -3396 5956 -3364
rect 5924 -3476 5956 -3444
rect 5924 -3525 5956 -3524
rect 5924 -3555 5925 -3525
rect 5925 -3555 5955 -3525
rect 5955 -3555 5956 -3525
rect 5924 -3556 5956 -3555
rect 5924 -3605 5956 -3604
rect 5924 -3635 5925 -3605
rect 5925 -3635 5955 -3605
rect 5955 -3635 5956 -3605
rect 5924 -3636 5956 -3635
rect 5924 -3685 5956 -3684
rect 5924 -3715 5925 -3685
rect 5925 -3715 5955 -3685
rect 5955 -3715 5956 -3685
rect 5924 -3716 5956 -3715
rect 6004 1035 6036 1036
rect 6004 1005 6005 1035
rect 6005 1005 6035 1035
rect 6035 1005 6036 1035
rect 6004 1004 6036 1005
rect 6004 955 6036 956
rect 6004 925 6005 955
rect 6005 925 6035 955
rect 6035 925 6036 955
rect 6004 924 6036 925
rect 6004 875 6036 876
rect 6004 845 6005 875
rect 6005 845 6035 875
rect 6035 845 6036 875
rect 6004 844 6036 845
rect 6004 764 6036 796
rect 6004 684 6036 716
rect 6004 635 6036 636
rect 6004 605 6005 635
rect 6005 605 6035 635
rect 6035 605 6036 635
rect 6004 604 6036 605
rect 6004 555 6036 556
rect 6004 525 6005 555
rect 6005 525 6035 555
rect 6035 525 6036 555
rect 6004 524 6036 525
rect 6004 444 6036 476
rect 6004 395 6036 396
rect 6004 365 6005 395
rect 6005 365 6035 395
rect 6035 365 6036 395
rect 6004 364 6036 365
rect 6004 284 6036 316
rect 6004 235 6036 236
rect 6004 205 6005 235
rect 6005 205 6035 235
rect 6035 205 6036 235
rect 6004 204 6036 205
rect 6004 124 6036 156
rect 6004 75 6036 76
rect 6004 45 6005 75
rect 6005 45 6035 75
rect 6035 45 6036 75
rect 6004 44 6036 45
rect 6004 -5 6036 -4
rect 6004 -35 6005 -5
rect 6005 -35 6035 -5
rect 6035 -35 6036 -5
rect 6004 -36 6036 -35
rect 6004 -85 6036 -84
rect 6004 -115 6005 -85
rect 6005 -115 6035 -85
rect 6035 -115 6036 -85
rect 6004 -116 6036 -115
rect 6004 -165 6036 -164
rect 6004 -195 6005 -165
rect 6005 -195 6035 -165
rect 6035 -195 6036 -165
rect 6004 -196 6036 -195
rect 6004 -245 6036 -244
rect 6004 -275 6005 -245
rect 6005 -275 6035 -245
rect 6035 -275 6036 -245
rect 6004 -276 6036 -275
rect 6004 -325 6036 -324
rect 6004 -355 6005 -325
rect 6005 -355 6035 -325
rect 6035 -355 6036 -325
rect 6004 -356 6036 -355
rect 6004 -436 6036 -404
rect 6004 -485 6036 -484
rect 6004 -515 6005 -485
rect 6005 -515 6035 -485
rect 6035 -515 6036 -485
rect 6004 -516 6036 -515
rect 6004 -596 6036 -564
rect 6004 -645 6036 -644
rect 6004 -675 6005 -645
rect 6005 -675 6035 -645
rect 6035 -675 6036 -645
rect 6004 -676 6036 -675
rect 6004 -756 6036 -724
rect 6004 -805 6036 -804
rect 6004 -835 6005 -805
rect 6005 -835 6035 -805
rect 6035 -835 6036 -805
rect 6004 -836 6036 -835
rect 6004 -885 6036 -884
rect 6004 -915 6005 -885
rect 6005 -915 6035 -885
rect 6035 -915 6036 -885
rect 6004 -916 6036 -915
rect 6004 -996 6036 -964
rect 6004 -1076 6036 -1044
rect 6004 -1125 6036 -1124
rect 6004 -1155 6005 -1125
rect 6005 -1155 6035 -1125
rect 6035 -1155 6036 -1125
rect 6004 -1156 6036 -1155
rect 6004 -1205 6036 -1204
rect 6004 -1235 6005 -1205
rect 6005 -1235 6035 -1205
rect 6035 -1235 6036 -1205
rect 6004 -1236 6036 -1235
rect 6004 -1285 6036 -1284
rect 6004 -1315 6005 -1285
rect 6005 -1315 6035 -1285
rect 6035 -1315 6036 -1285
rect 6004 -1316 6036 -1315
rect 6004 -1365 6036 -1364
rect 6004 -1395 6005 -1365
rect 6005 -1395 6035 -1365
rect 6035 -1395 6036 -1365
rect 6004 -1396 6036 -1395
rect 6004 -1445 6036 -1444
rect 6004 -1475 6005 -1445
rect 6005 -1475 6035 -1445
rect 6035 -1475 6036 -1445
rect 6004 -1476 6036 -1475
rect 6004 -1525 6036 -1524
rect 6004 -1555 6005 -1525
rect 6005 -1555 6035 -1525
rect 6035 -1555 6036 -1525
rect 6004 -1556 6036 -1555
rect 6004 -1636 6036 -1604
rect 6004 -1716 6036 -1684
rect 6004 -1765 6036 -1764
rect 6004 -1795 6005 -1765
rect 6005 -1795 6035 -1765
rect 6035 -1795 6036 -1765
rect 6004 -1796 6036 -1795
rect 6004 -1845 6036 -1844
rect 6004 -1875 6005 -1845
rect 6005 -1875 6035 -1845
rect 6035 -1875 6036 -1845
rect 6004 -1876 6036 -1875
rect 6004 -1956 6036 -1924
rect 6004 -2005 6036 -2004
rect 6004 -2035 6005 -2005
rect 6005 -2035 6035 -2005
rect 6035 -2035 6036 -2005
rect 6004 -2036 6036 -2035
rect 6004 -2116 6036 -2084
rect 6004 -2165 6036 -2164
rect 6004 -2195 6005 -2165
rect 6005 -2195 6035 -2165
rect 6035 -2195 6036 -2165
rect 6004 -2196 6036 -2195
rect 6004 -2276 6036 -2244
rect 6004 -2325 6036 -2324
rect 6004 -2355 6005 -2325
rect 6005 -2355 6035 -2325
rect 6035 -2355 6036 -2325
rect 6004 -2356 6036 -2355
rect 6004 -2405 6036 -2404
rect 6004 -2435 6005 -2405
rect 6005 -2435 6035 -2405
rect 6035 -2435 6036 -2405
rect 6004 -2436 6036 -2435
rect 6004 -2485 6036 -2484
rect 6004 -2515 6005 -2485
rect 6005 -2515 6035 -2485
rect 6035 -2515 6036 -2485
rect 6004 -2516 6036 -2515
rect 6004 -2565 6036 -2564
rect 6004 -2595 6005 -2565
rect 6005 -2595 6035 -2565
rect 6035 -2595 6036 -2565
rect 6004 -2596 6036 -2595
rect 6004 -2645 6036 -2644
rect 6004 -2675 6005 -2645
rect 6005 -2675 6035 -2645
rect 6035 -2675 6036 -2645
rect 6004 -2676 6036 -2675
rect 6004 -2725 6036 -2724
rect 6004 -2755 6005 -2725
rect 6005 -2755 6035 -2725
rect 6035 -2755 6036 -2725
rect 6004 -2756 6036 -2755
rect 6004 -2836 6036 -2804
rect 6004 -2885 6036 -2884
rect 6004 -2915 6005 -2885
rect 6005 -2915 6035 -2885
rect 6035 -2915 6036 -2885
rect 6004 -2916 6036 -2915
rect 6004 -2996 6036 -2964
rect 6004 -3045 6036 -3044
rect 6004 -3075 6005 -3045
rect 6005 -3075 6035 -3045
rect 6035 -3075 6036 -3045
rect 6004 -3076 6036 -3075
rect 6004 -3156 6036 -3124
rect 6004 -3205 6036 -3204
rect 6004 -3235 6005 -3205
rect 6005 -3235 6035 -3205
rect 6035 -3235 6036 -3205
rect 6004 -3236 6036 -3235
rect 6004 -3285 6036 -3284
rect 6004 -3315 6005 -3285
rect 6005 -3315 6035 -3285
rect 6035 -3315 6036 -3285
rect 6004 -3316 6036 -3315
rect 6004 -3396 6036 -3364
rect 6004 -3476 6036 -3444
rect 6004 -3525 6036 -3524
rect 6004 -3555 6005 -3525
rect 6005 -3555 6035 -3525
rect 6035 -3555 6036 -3525
rect 6004 -3556 6036 -3555
rect 6004 -3605 6036 -3604
rect 6004 -3635 6005 -3605
rect 6005 -3635 6035 -3605
rect 6035 -3635 6036 -3605
rect 6004 -3636 6036 -3635
rect 6004 -3685 6036 -3684
rect 6004 -3715 6005 -3685
rect 6005 -3715 6035 -3685
rect 6035 -3715 6036 -3685
rect 6004 -3716 6036 -3715
rect 6084 1035 6116 1036
rect 6084 1005 6085 1035
rect 6085 1005 6115 1035
rect 6115 1005 6116 1035
rect 6084 1004 6116 1005
rect 6084 955 6116 956
rect 6084 925 6085 955
rect 6085 925 6115 955
rect 6115 925 6116 955
rect 6084 924 6116 925
rect 6084 875 6116 876
rect 6084 845 6085 875
rect 6085 845 6115 875
rect 6115 845 6116 875
rect 6084 844 6116 845
rect 6084 764 6116 796
rect 6084 684 6116 716
rect 6084 635 6116 636
rect 6084 605 6085 635
rect 6085 605 6115 635
rect 6115 605 6116 635
rect 6084 604 6116 605
rect 6084 555 6116 556
rect 6084 525 6085 555
rect 6085 525 6115 555
rect 6115 525 6116 555
rect 6084 524 6116 525
rect 6084 444 6116 476
rect 6084 395 6116 396
rect 6084 365 6085 395
rect 6085 365 6115 395
rect 6115 365 6116 395
rect 6084 364 6116 365
rect 6084 284 6116 316
rect 6084 235 6116 236
rect 6084 205 6085 235
rect 6085 205 6115 235
rect 6115 205 6116 235
rect 6084 204 6116 205
rect 6084 124 6116 156
rect 6084 75 6116 76
rect 6084 45 6085 75
rect 6085 45 6115 75
rect 6115 45 6116 75
rect 6084 44 6116 45
rect 6084 -5 6116 -4
rect 6084 -35 6085 -5
rect 6085 -35 6115 -5
rect 6115 -35 6116 -5
rect 6084 -36 6116 -35
rect 6084 -85 6116 -84
rect 6084 -115 6085 -85
rect 6085 -115 6115 -85
rect 6115 -115 6116 -85
rect 6084 -116 6116 -115
rect 6084 -165 6116 -164
rect 6084 -195 6085 -165
rect 6085 -195 6115 -165
rect 6115 -195 6116 -165
rect 6084 -196 6116 -195
rect 6084 -245 6116 -244
rect 6084 -275 6085 -245
rect 6085 -275 6115 -245
rect 6115 -275 6116 -245
rect 6084 -276 6116 -275
rect 6084 -325 6116 -324
rect 6084 -355 6085 -325
rect 6085 -355 6115 -325
rect 6115 -355 6116 -325
rect 6084 -356 6116 -355
rect 6084 -436 6116 -404
rect 6084 -485 6116 -484
rect 6084 -515 6085 -485
rect 6085 -515 6115 -485
rect 6115 -515 6116 -485
rect 6084 -516 6116 -515
rect 6084 -596 6116 -564
rect 6084 -645 6116 -644
rect 6084 -675 6085 -645
rect 6085 -675 6115 -645
rect 6115 -675 6116 -645
rect 6084 -676 6116 -675
rect 6084 -756 6116 -724
rect 6084 -805 6116 -804
rect 6084 -835 6085 -805
rect 6085 -835 6115 -805
rect 6115 -835 6116 -805
rect 6084 -836 6116 -835
rect 6084 -885 6116 -884
rect 6084 -915 6085 -885
rect 6085 -915 6115 -885
rect 6115 -915 6116 -885
rect 6084 -916 6116 -915
rect 6084 -996 6116 -964
rect 6084 -1076 6116 -1044
rect 6084 -1125 6116 -1124
rect 6084 -1155 6085 -1125
rect 6085 -1155 6115 -1125
rect 6115 -1155 6116 -1125
rect 6084 -1156 6116 -1155
rect 6084 -1205 6116 -1204
rect 6084 -1235 6085 -1205
rect 6085 -1235 6115 -1205
rect 6115 -1235 6116 -1205
rect 6084 -1236 6116 -1235
rect 6084 -1285 6116 -1284
rect 6084 -1315 6085 -1285
rect 6085 -1315 6115 -1285
rect 6115 -1315 6116 -1285
rect 6084 -1316 6116 -1315
rect 6084 -1365 6116 -1364
rect 6084 -1395 6085 -1365
rect 6085 -1395 6115 -1365
rect 6115 -1395 6116 -1365
rect 6084 -1396 6116 -1395
rect 6084 -1445 6116 -1444
rect 6084 -1475 6085 -1445
rect 6085 -1475 6115 -1445
rect 6115 -1475 6116 -1445
rect 6084 -1476 6116 -1475
rect 6084 -1525 6116 -1524
rect 6084 -1555 6085 -1525
rect 6085 -1555 6115 -1525
rect 6115 -1555 6116 -1525
rect 6084 -1556 6116 -1555
rect 6084 -1636 6116 -1604
rect 6084 -1716 6116 -1684
rect 6084 -1765 6116 -1764
rect 6084 -1795 6085 -1765
rect 6085 -1795 6115 -1765
rect 6115 -1795 6116 -1765
rect 6084 -1796 6116 -1795
rect 6084 -1845 6116 -1844
rect 6084 -1875 6085 -1845
rect 6085 -1875 6115 -1845
rect 6115 -1875 6116 -1845
rect 6084 -1876 6116 -1875
rect 6084 -1956 6116 -1924
rect 6084 -2005 6116 -2004
rect 6084 -2035 6085 -2005
rect 6085 -2035 6115 -2005
rect 6115 -2035 6116 -2005
rect 6084 -2036 6116 -2035
rect 6084 -2116 6116 -2084
rect 6084 -2165 6116 -2164
rect 6084 -2195 6085 -2165
rect 6085 -2195 6115 -2165
rect 6115 -2195 6116 -2165
rect 6084 -2196 6116 -2195
rect 6084 -2276 6116 -2244
rect 6084 -2325 6116 -2324
rect 6084 -2355 6085 -2325
rect 6085 -2355 6115 -2325
rect 6115 -2355 6116 -2325
rect 6084 -2356 6116 -2355
rect 6084 -2405 6116 -2404
rect 6084 -2435 6085 -2405
rect 6085 -2435 6115 -2405
rect 6115 -2435 6116 -2405
rect 6084 -2436 6116 -2435
rect 6084 -2485 6116 -2484
rect 6084 -2515 6085 -2485
rect 6085 -2515 6115 -2485
rect 6115 -2515 6116 -2485
rect 6084 -2516 6116 -2515
rect 6084 -2565 6116 -2564
rect 6084 -2595 6085 -2565
rect 6085 -2595 6115 -2565
rect 6115 -2595 6116 -2565
rect 6084 -2596 6116 -2595
rect 6084 -2645 6116 -2644
rect 6084 -2675 6085 -2645
rect 6085 -2675 6115 -2645
rect 6115 -2675 6116 -2645
rect 6084 -2676 6116 -2675
rect 6084 -2725 6116 -2724
rect 6084 -2755 6085 -2725
rect 6085 -2755 6115 -2725
rect 6115 -2755 6116 -2725
rect 6084 -2756 6116 -2755
rect 6084 -2836 6116 -2804
rect 6084 -2885 6116 -2884
rect 6084 -2915 6085 -2885
rect 6085 -2915 6115 -2885
rect 6115 -2915 6116 -2885
rect 6084 -2916 6116 -2915
rect 6084 -2996 6116 -2964
rect 6084 -3045 6116 -3044
rect 6084 -3075 6085 -3045
rect 6085 -3075 6115 -3045
rect 6115 -3075 6116 -3045
rect 6084 -3076 6116 -3075
rect 6084 -3156 6116 -3124
rect 6084 -3205 6116 -3204
rect 6084 -3235 6085 -3205
rect 6085 -3235 6115 -3205
rect 6115 -3235 6116 -3205
rect 6084 -3236 6116 -3235
rect 6084 -3285 6116 -3284
rect 6084 -3315 6085 -3285
rect 6085 -3315 6115 -3285
rect 6115 -3315 6116 -3285
rect 6084 -3316 6116 -3315
rect 6084 -3396 6116 -3364
rect 6084 -3476 6116 -3444
rect 6084 -3525 6116 -3524
rect 6084 -3555 6085 -3525
rect 6085 -3555 6115 -3525
rect 6115 -3555 6116 -3525
rect 6084 -3556 6116 -3555
rect 6084 -3605 6116 -3604
rect 6084 -3635 6085 -3605
rect 6085 -3635 6115 -3605
rect 6115 -3635 6116 -3605
rect 6084 -3636 6116 -3635
rect 6084 -3685 6116 -3684
rect 6084 -3715 6085 -3685
rect 6085 -3715 6115 -3685
rect 6115 -3715 6116 -3685
rect 6084 -3716 6116 -3715
rect 6164 1035 6196 1036
rect 6164 1005 6165 1035
rect 6165 1005 6195 1035
rect 6195 1005 6196 1035
rect 6164 1004 6196 1005
rect 6164 955 6196 956
rect 6164 925 6165 955
rect 6165 925 6195 955
rect 6195 925 6196 955
rect 6164 924 6196 925
rect 6164 875 6196 876
rect 6164 845 6165 875
rect 6165 845 6195 875
rect 6195 845 6196 875
rect 6164 844 6196 845
rect 6164 764 6196 796
rect 6164 684 6196 716
rect 6164 635 6196 636
rect 6164 605 6165 635
rect 6165 605 6195 635
rect 6195 605 6196 635
rect 6164 604 6196 605
rect 6164 555 6196 556
rect 6164 525 6165 555
rect 6165 525 6195 555
rect 6195 525 6196 555
rect 6164 524 6196 525
rect 6164 444 6196 476
rect 6164 395 6196 396
rect 6164 365 6165 395
rect 6165 365 6195 395
rect 6195 365 6196 395
rect 6164 364 6196 365
rect 6164 284 6196 316
rect 6164 235 6196 236
rect 6164 205 6165 235
rect 6165 205 6195 235
rect 6195 205 6196 235
rect 6164 204 6196 205
rect 6164 124 6196 156
rect 6164 75 6196 76
rect 6164 45 6165 75
rect 6165 45 6195 75
rect 6195 45 6196 75
rect 6164 44 6196 45
rect 6164 -5 6196 -4
rect 6164 -35 6165 -5
rect 6165 -35 6195 -5
rect 6195 -35 6196 -5
rect 6164 -36 6196 -35
rect 6164 -85 6196 -84
rect 6164 -115 6165 -85
rect 6165 -115 6195 -85
rect 6195 -115 6196 -85
rect 6164 -116 6196 -115
rect 6164 -165 6196 -164
rect 6164 -195 6165 -165
rect 6165 -195 6195 -165
rect 6195 -195 6196 -165
rect 6164 -196 6196 -195
rect 6164 -245 6196 -244
rect 6164 -275 6165 -245
rect 6165 -275 6195 -245
rect 6195 -275 6196 -245
rect 6164 -276 6196 -275
rect 6164 -325 6196 -324
rect 6164 -355 6165 -325
rect 6165 -355 6195 -325
rect 6195 -355 6196 -325
rect 6164 -356 6196 -355
rect 6164 -436 6196 -404
rect 6164 -485 6196 -484
rect 6164 -515 6165 -485
rect 6165 -515 6195 -485
rect 6195 -515 6196 -485
rect 6164 -516 6196 -515
rect 6164 -596 6196 -564
rect 6164 -645 6196 -644
rect 6164 -675 6165 -645
rect 6165 -675 6195 -645
rect 6195 -675 6196 -645
rect 6164 -676 6196 -675
rect 6164 -756 6196 -724
rect 6164 -805 6196 -804
rect 6164 -835 6165 -805
rect 6165 -835 6195 -805
rect 6195 -835 6196 -805
rect 6164 -836 6196 -835
rect 6164 -885 6196 -884
rect 6164 -915 6165 -885
rect 6165 -915 6195 -885
rect 6195 -915 6196 -885
rect 6164 -916 6196 -915
rect 6164 -996 6196 -964
rect 6164 -1076 6196 -1044
rect 6164 -1125 6196 -1124
rect 6164 -1155 6165 -1125
rect 6165 -1155 6195 -1125
rect 6195 -1155 6196 -1125
rect 6164 -1156 6196 -1155
rect 6164 -1205 6196 -1204
rect 6164 -1235 6165 -1205
rect 6165 -1235 6195 -1205
rect 6195 -1235 6196 -1205
rect 6164 -1236 6196 -1235
rect 6164 -1285 6196 -1284
rect 6164 -1315 6165 -1285
rect 6165 -1315 6195 -1285
rect 6195 -1315 6196 -1285
rect 6164 -1316 6196 -1315
rect 6164 -1365 6196 -1364
rect 6164 -1395 6165 -1365
rect 6165 -1395 6195 -1365
rect 6195 -1395 6196 -1365
rect 6164 -1396 6196 -1395
rect 6164 -1445 6196 -1444
rect 6164 -1475 6165 -1445
rect 6165 -1475 6195 -1445
rect 6195 -1475 6196 -1445
rect 6164 -1476 6196 -1475
rect 6164 -1525 6196 -1524
rect 6164 -1555 6165 -1525
rect 6165 -1555 6195 -1525
rect 6195 -1555 6196 -1525
rect 6164 -1556 6196 -1555
rect 6164 -1636 6196 -1604
rect 6164 -1716 6196 -1684
rect 6164 -1765 6196 -1764
rect 6164 -1795 6165 -1765
rect 6165 -1795 6195 -1765
rect 6195 -1795 6196 -1765
rect 6164 -1796 6196 -1795
rect 6164 -1845 6196 -1844
rect 6164 -1875 6165 -1845
rect 6165 -1875 6195 -1845
rect 6195 -1875 6196 -1845
rect 6164 -1876 6196 -1875
rect 6164 -1956 6196 -1924
rect 6164 -2005 6196 -2004
rect 6164 -2035 6165 -2005
rect 6165 -2035 6195 -2005
rect 6195 -2035 6196 -2005
rect 6164 -2036 6196 -2035
rect 6164 -2116 6196 -2084
rect 6164 -2165 6196 -2164
rect 6164 -2195 6165 -2165
rect 6165 -2195 6195 -2165
rect 6195 -2195 6196 -2165
rect 6164 -2196 6196 -2195
rect 6164 -2276 6196 -2244
rect 6164 -2325 6196 -2324
rect 6164 -2355 6165 -2325
rect 6165 -2355 6195 -2325
rect 6195 -2355 6196 -2325
rect 6164 -2356 6196 -2355
rect 6164 -2405 6196 -2404
rect 6164 -2435 6165 -2405
rect 6165 -2435 6195 -2405
rect 6195 -2435 6196 -2405
rect 6164 -2436 6196 -2435
rect 6164 -2485 6196 -2484
rect 6164 -2515 6165 -2485
rect 6165 -2515 6195 -2485
rect 6195 -2515 6196 -2485
rect 6164 -2516 6196 -2515
rect 6164 -2565 6196 -2564
rect 6164 -2595 6165 -2565
rect 6165 -2595 6195 -2565
rect 6195 -2595 6196 -2565
rect 6164 -2596 6196 -2595
rect 6164 -2645 6196 -2644
rect 6164 -2675 6165 -2645
rect 6165 -2675 6195 -2645
rect 6195 -2675 6196 -2645
rect 6164 -2676 6196 -2675
rect 6164 -2725 6196 -2724
rect 6164 -2755 6165 -2725
rect 6165 -2755 6195 -2725
rect 6195 -2755 6196 -2725
rect 6164 -2756 6196 -2755
rect 6164 -2836 6196 -2804
rect 6164 -2885 6196 -2884
rect 6164 -2915 6165 -2885
rect 6165 -2915 6195 -2885
rect 6195 -2915 6196 -2885
rect 6164 -2916 6196 -2915
rect 6164 -2996 6196 -2964
rect 6164 -3045 6196 -3044
rect 6164 -3075 6165 -3045
rect 6165 -3075 6195 -3045
rect 6195 -3075 6196 -3045
rect 6164 -3076 6196 -3075
rect 6164 -3156 6196 -3124
rect 6164 -3205 6196 -3204
rect 6164 -3235 6165 -3205
rect 6165 -3235 6195 -3205
rect 6195 -3235 6196 -3205
rect 6164 -3236 6196 -3235
rect 6164 -3285 6196 -3284
rect 6164 -3315 6165 -3285
rect 6165 -3315 6195 -3285
rect 6195 -3315 6196 -3285
rect 6164 -3316 6196 -3315
rect 6164 -3396 6196 -3364
rect 6164 -3476 6196 -3444
rect 6164 -3525 6196 -3524
rect 6164 -3555 6165 -3525
rect 6165 -3555 6195 -3525
rect 6195 -3555 6196 -3525
rect 6164 -3556 6196 -3555
rect 6164 -3605 6196 -3604
rect 6164 -3635 6165 -3605
rect 6165 -3635 6195 -3605
rect 6195 -3635 6196 -3605
rect 6164 -3636 6196 -3635
rect 6164 -3685 6196 -3684
rect 6164 -3715 6165 -3685
rect 6165 -3715 6195 -3685
rect 6195 -3715 6196 -3685
rect 6164 -3716 6196 -3715
rect 6244 1035 6276 1036
rect 6244 1005 6245 1035
rect 6245 1005 6275 1035
rect 6275 1005 6276 1035
rect 6244 1004 6276 1005
rect 6244 955 6276 956
rect 6244 925 6245 955
rect 6245 925 6275 955
rect 6275 925 6276 955
rect 6244 924 6276 925
rect 6244 875 6276 876
rect 6244 845 6245 875
rect 6245 845 6275 875
rect 6275 845 6276 875
rect 6244 844 6276 845
rect 6244 764 6276 796
rect 6244 684 6276 716
rect 6244 635 6276 636
rect 6244 605 6245 635
rect 6245 605 6275 635
rect 6275 605 6276 635
rect 6244 604 6276 605
rect 6244 555 6276 556
rect 6244 525 6245 555
rect 6245 525 6275 555
rect 6275 525 6276 555
rect 6244 524 6276 525
rect 6244 444 6276 476
rect 6244 395 6276 396
rect 6244 365 6245 395
rect 6245 365 6275 395
rect 6275 365 6276 395
rect 6244 364 6276 365
rect 6244 284 6276 316
rect 6244 235 6276 236
rect 6244 205 6245 235
rect 6245 205 6275 235
rect 6275 205 6276 235
rect 6244 204 6276 205
rect 6244 124 6276 156
rect 6244 75 6276 76
rect 6244 45 6245 75
rect 6245 45 6275 75
rect 6275 45 6276 75
rect 6244 44 6276 45
rect 6244 -5 6276 -4
rect 6244 -35 6245 -5
rect 6245 -35 6275 -5
rect 6275 -35 6276 -5
rect 6244 -36 6276 -35
rect 6244 -85 6276 -84
rect 6244 -115 6245 -85
rect 6245 -115 6275 -85
rect 6275 -115 6276 -85
rect 6244 -116 6276 -115
rect 6244 -165 6276 -164
rect 6244 -195 6245 -165
rect 6245 -195 6275 -165
rect 6275 -195 6276 -165
rect 6244 -196 6276 -195
rect 6244 -245 6276 -244
rect 6244 -275 6245 -245
rect 6245 -275 6275 -245
rect 6275 -275 6276 -245
rect 6244 -276 6276 -275
rect 6244 -325 6276 -324
rect 6244 -355 6245 -325
rect 6245 -355 6275 -325
rect 6275 -355 6276 -325
rect 6244 -356 6276 -355
rect 6244 -436 6276 -404
rect 6244 -485 6276 -484
rect 6244 -515 6245 -485
rect 6245 -515 6275 -485
rect 6275 -515 6276 -485
rect 6244 -516 6276 -515
rect 6244 -596 6276 -564
rect 6244 -645 6276 -644
rect 6244 -675 6245 -645
rect 6245 -675 6275 -645
rect 6275 -675 6276 -645
rect 6244 -676 6276 -675
rect 6244 -756 6276 -724
rect 6244 -805 6276 -804
rect 6244 -835 6245 -805
rect 6245 -835 6275 -805
rect 6275 -835 6276 -805
rect 6244 -836 6276 -835
rect 6244 -885 6276 -884
rect 6244 -915 6245 -885
rect 6245 -915 6275 -885
rect 6275 -915 6276 -885
rect 6244 -916 6276 -915
rect 6244 -996 6276 -964
rect 6244 -1076 6276 -1044
rect 6244 -1125 6276 -1124
rect 6244 -1155 6245 -1125
rect 6245 -1155 6275 -1125
rect 6275 -1155 6276 -1125
rect 6244 -1156 6276 -1155
rect 6244 -1205 6276 -1204
rect 6244 -1235 6245 -1205
rect 6245 -1235 6275 -1205
rect 6275 -1235 6276 -1205
rect 6244 -1236 6276 -1235
rect 6244 -1285 6276 -1284
rect 6244 -1315 6245 -1285
rect 6245 -1315 6275 -1285
rect 6275 -1315 6276 -1285
rect 6244 -1316 6276 -1315
rect 6244 -1365 6276 -1364
rect 6244 -1395 6245 -1365
rect 6245 -1395 6275 -1365
rect 6275 -1395 6276 -1365
rect 6244 -1396 6276 -1395
rect 6244 -1445 6276 -1444
rect 6244 -1475 6245 -1445
rect 6245 -1475 6275 -1445
rect 6275 -1475 6276 -1445
rect 6244 -1476 6276 -1475
rect 6244 -1525 6276 -1524
rect 6244 -1555 6245 -1525
rect 6245 -1555 6275 -1525
rect 6275 -1555 6276 -1525
rect 6244 -1556 6276 -1555
rect 6244 -1636 6276 -1604
rect 6244 -1716 6276 -1684
rect 6244 -1765 6276 -1764
rect 6244 -1795 6245 -1765
rect 6245 -1795 6275 -1765
rect 6275 -1795 6276 -1765
rect 6244 -1796 6276 -1795
rect 6244 -1845 6276 -1844
rect 6244 -1875 6245 -1845
rect 6245 -1875 6275 -1845
rect 6275 -1875 6276 -1845
rect 6244 -1876 6276 -1875
rect 6244 -1956 6276 -1924
rect 6244 -2005 6276 -2004
rect 6244 -2035 6245 -2005
rect 6245 -2035 6275 -2005
rect 6275 -2035 6276 -2005
rect 6244 -2036 6276 -2035
rect 6244 -2116 6276 -2084
rect 6244 -2165 6276 -2164
rect 6244 -2195 6245 -2165
rect 6245 -2195 6275 -2165
rect 6275 -2195 6276 -2165
rect 6244 -2196 6276 -2195
rect 6244 -2276 6276 -2244
rect 6244 -2325 6276 -2324
rect 6244 -2355 6245 -2325
rect 6245 -2355 6275 -2325
rect 6275 -2355 6276 -2325
rect 6244 -2356 6276 -2355
rect 6244 -2405 6276 -2404
rect 6244 -2435 6245 -2405
rect 6245 -2435 6275 -2405
rect 6275 -2435 6276 -2405
rect 6244 -2436 6276 -2435
rect 6244 -2485 6276 -2484
rect 6244 -2515 6245 -2485
rect 6245 -2515 6275 -2485
rect 6275 -2515 6276 -2485
rect 6244 -2516 6276 -2515
rect 6244 -2565 6276 -2564
rect 6244 -2595 6245 -2565
rect 6245 -2595 6275 -2565
rect 6275 -2595 6276 -2565
rect 6244 -2596 6276 -2595
rect 6244 -2645 6276 -2644
rect 6244 -2675 6245 -2645
rect 6245 -2675 6275 -2645
rect 6275 -2675 6276 -2645
rect 6244 -2676 6276 -2675
rect 6244 -2725 6276 -2724
rect 6244 -2755 6245 -2725
rect 6245 -2755 6275 -2725
rect 6275 -2755 6276 -2725
rect 6244 -2756 6276 -2755
rect 6244 -2836 6276 -2804
rect 6244 -2885 6276 -2884
rect 6244 -2915 6245 -2885
rect 6245 -2915 6275 -2885
rect 6275 -2915 6276 -2885
rect 6244 -2916 6276 -2915
rect 6244 -2996 6276 -2964
rect 6244 -3045 6276 -3044
rect 6244 -3075 6245 -3045
rect 6245 -3075 6275 -3045
rect 6275 -3075 6276 -3045
rect 6244 -3076 6276 -3075
rect 6244 -3156 6276 -3124
rect 6244 -3205 6276 -3204
rect 6244 -3235 6245 -3205
rect 6245 -3235 6275 -3205
rect 6275 -3235 6276 -3205
rect 6244 -3236 6276 -3235
rect 6244 -3285 6276 -3284
rect 6244 -3315 6245 -3285
rect 6245 -3315 6275 -3285
rect 6275 -3315 6276 -3285
rect 6244 -3316 6276 -3315
rect 6244 -3396 6276 -3364
rect 6244 -3476 6276 -3444
rect 6244 -3525 6276 -3524
rect 6244 -3555 6245 -3525
rect 6245 -3555 6275 -3525
rect 6275 -3555 6276 -3525
rect 6244 -3556 6276 -3555
rect 6244 -3605 6276 -3604
rect 6244 -3635 6245 -3605
rect 6245 -3635 6275 -3605
rect 6275 -3635 6276 -3605
rect 6244 -3636 6276 -3635
rect 6244 -3685 6276 -3684
rect 6244 -3715 6245 -3685
rect 6245 -3715 6275 -3685
rect 6275 -3715 6276 -3685
rect 6244 -3716 6276 -3715
rect 6324 1035 6356 1036
rect 6324 1005 6325 1035
rect 6325 1005 6355 1035
rect 6355 1005 6356 1035
rect 6324 1004 6356 1005
rect 6324 955 6356 956
rect 6324 925 6325 955
rect 6325 925 6355 955
rect 6355 925 6356 955
rect 6324 924 6356 925
rect 6324 875 6356 876
rect 6324 845 6325 875
rect 6325 845 6355 875
rect 6355 845 6356 875
rect 6324 844 6356 845
rect 6324 764 6356 796
rect 6324 684 6356 716
rect 6324 635 6356 636
rect 6324 605 6325 635
rect 6325 605 6355 635
rect 6355 605 6356 635
rect 6324 604 6356 605
rect 6324 555 6356 556
rect 6324 525 6325 555
rect 6325 525 6355 555
rect 6355 525 6356 555
rect 6324 524 6356 525
rect 6324 444 6356 476
rect 6324 395 6356 396
rect 6324 365 6325 395
rect 6325 365 6355 395
rect 6355 365 6356 395
rect 6324 364 6356 365
rect 6324 284 6356 316
rect 6324 235 6356 236
rect 6324 205 6325 235
rect 6325 205 6355 235
rect 6355 205 6356 235
rect 6324 204 6356 205
rect 6324 124 6356 156
rect 6324 75 6356 76
rect 6324 45 6325 75
rect 6325 45 6355 75
rect 6355 45 6356 75
rect 6324 44 6356 45
rect 6324 -5 6356 -4
rect 6324 -35 6325 -5
rect 6325 -35 6355 -5
rect 6355 -35 6356 -5
rect 6324 -36 6356 -35
rect 6324 -85 6356 -84
rect 6324 -115 6325 -85
rect 6325 -115 6355 -85
rect 6355 -115 6356 -85
rect 6324 -116 6356 -115
rect 6324 -165 6356 -164
rect 6324 -195 6325 -165
rect 6325 -195 6355 -165
rect 6355 -195 6356 -165
rect 6324 -196 6356 -195
rect 6324 -245 6356 -244
rect 6324 -275 6325 -245
rect 6325 -275 6355 -245
rect 6355 -275 6356 -245
rect 6324 -276 6356 -275
rect 6324 -325 6356 -324
rect 6324 -355 6325 -325
rect 6325 -355 6355 -325
rect 6355 -355 6356 -325
rect 6324 -356 6356 -355
rect 6324 -436 6356 -404
rect 6324 -485 6356 -484
rect 6324 -515 6325 -485
rect 6325 -515 6355 -485
rect 6355 -515 6356 -485
rect 6324 -516 6356 -515
rect 6324 -596 6356 -564
rect 6324 -645 6356 -644
rect 6324 -675 6325 -645
rect 6325 -675 6355 -645
rect 6355 -675 6356 -645
rect 6324 -676 6356 -675
rect 6324 -756 6356 -724
rect 6324 -805 6356 -804
rect 6324 -835 6325 -805
rect 6325 -835 6355 -805
rect 6355 -835 6356 -805
rect 6324 -836 6356 -835
rect 6324 -885 6356 -884
rect 6324 -915 6325 -885
rect 6325 -915 6355 -885
rect 6355 -915 6356 -885
rect 6324 -916 6356 -915
rect 6324 -996 6356 -964
rect 6324 -1076 6356 -1044
rect 6324 -1125 6356 -1124
rect 6324 -1155 6325 -1125
rect 6325 -1155 6355 -1125
rect 6355 -1155 6356 -1125
rect 6324 -1156 6356 -1155
rect 6324 -1205 6356 -1204
rect 6324 -1235 6325 -1205
rect 6325 -1235 6355 -1205
rect 6355 -1235 6356 -1205
rect 6324 -1236 6356 -1235
rect 6324 -1285 6356 -1284
rect 6324 -1315 6325 -1285
rect 6325 -1315 6355 -1285
rect 6355 -1315 6356 -1285
rect 6324 -1316 6356 -1315
rect 6324 -1365 6356 -1364
rect 6324 -1395 6325 -1365
rect 6325 -1395 6355 -1365
rect 6355 -1395 6356 -1365
rect 6324 -1396 6356 -1395
rect 6324 -1445 6356 -1444
rect 6324 -1475 6325 -1445
rect 6325 -1475 6355 -1445
rect 6355 -1475 6356 -1445
rect 6324 -1476 6356 -1475
rect 6324 -1525 6356 -1524
rect 6324 -1555 6325 -1525
rect 6325 -1555 6355 -1525
rect 6355 -1555 6356 -1525
rect 6324 -1556 6356 -1555
rect 6324 -1636 6356 -1604
rect 6324 -1716 6356 -1684
rect 6324 -1765 6356 -1764
rect 6324 -1795 6325 -1765
rect 6325 -1795 6355 -1765
rect 6355 -1795 6356 -1765
rect 6324 -1796 6356 -1795
rect 6324 -1845 6356 -1844
rect 6324 -1875 6325 -1845
rect 6325 -1875 6355 -1845
rect 6355 -1875 6356 -1845
rect 6324 -1876 6356 -1875
rect 6324 -1956 6356 -1924
rect 6324 -2005 6356 -2004
rect 6324 -2035 6325 -2005
rect 6325 -2035 6355 -2005
rect 6355 -2035 6356 -2005
rect 6324 -2036 6356 -2035
rect 6324 -2116 6356 -2084
rect 6324 -2165 6356 -2164
rect 6324 -2195 6325 -2165
rect 6325 -2195 6355 -2165
rect 6355 -2195 6356 -2165
rect 6324 -2196 6356 -2195
rect 6324 -2276 6356 -2244
rect 6324 -2325 6356 -2324
rect 6324 -2355 6325 -2325
rect 6325 -2355 6355 -2325
rect 6355 -2355 6356 -2325
rect 6324 -2356 6356 -2355
rect 6324 -2405 6356 -2404
rect 6324 -2435 6325 -2405
rect 6325 -2435 6355 -2405
rect 6355 -2435 6356 -2405
rect 6324 -2436 6356 -2435
rect 6324 -2485 6356 -2484
rect 6324 -2515 6325 -2485
rect 6325 -2515 6355 -2485
rect 6355 -2515 6356 -2485
rect 6324 -2516 6356 -2515
rect 6324 -2565 6356 -2564
rect 6324 -2595 6325 -2565
rect 6325 -2595 6355 -2565
rect 6355 -2595 6356 -2565
rect 6324 -2596 6356 -2595
rect 6324 -2645 6356 -2644
rect 6324 -2675 6325 -2645
rect 6325 -2675 6355 -2645
rect 6355 -2675 6356 -2645
rect 6324 -2676 6356 -2675
rect 6324 -2725 6356 -2724
rect 6324 -2755 6325 -2725
rect 6325 -2755 6355 -2725
rect 6355 -2755 6356 -2725
rect 6324 -2756 6356 -2755
rect 6324 -2836 6356 -2804
rect 6324 -2885 6356 -2884
rect 6324 -2915 6325 -2885
rect 6325 -2915 6355 -2885
rect 6355 -2915 6356 -2885
rect 6324 -2916 6356 -2915
rect 6324 -2996 6356 -2964
rect 6324 -3045 6356 -3044
rect 6324 -3075 6325 -3045
rect 6325 -3075 6355 -3045
rect 6355 -3075 6356 -3045
rect 6324 -3076 6356 -3075
rect 6324 -3156 6356 -3124
rect 6324 -3205 6356 -3204
rect 6324 -3235 6325 -3205
rect 6325 -3235 6355 -3205
rect 6355 -3235 6356 -3205
rect 6324 -3236 6356 -3235
rect 6324 -3285 6356 -3284
rect 6324 -3315 6325 -3285
rect 6325 -3315 6355 -3285
rect 6355 -3315 6356 -3285
rect 6324 -3316 6356 -3315
rect 6324 -3396 6356 -3364
rect 6324 -3476 6356 -3444
rect 6324 -3525 6356 -3524
rect 6324 -3555 6325 -3525
rect 6325 -3555 6355 -3525
rect 6355 -3555 6356 -3525
rect 6324 -3556 6356 -3555
rect 6324 -3605 6356 -3604
rect 6324 -3635 6325 -3605
rect 6325 -3635 6355 -3605
rect 6355 -3635 6356 -3605
rect 6324 -3636 6356 -3635
rect 6324 -3685 6356 -3684
rect 6324 -3715 6325 -3685
rect 6325 -3715 6355 -3685
rect 6355 -3715 6356 -3685
rect 6324 -3716 6356 -3715
rect 6404 1035 6436 1036
rect 6404 1005 6405 1035
rect 6405 1005 6435 1035
rect 6435 1005 6436 1035
rect 6404 1004 6436 1005
rect 6404 955 6436 956
rect 6404 925 6405 955
rect 6405 925 6435 955
rect 6435 925 6436 955
rect 6404 924 6436 925
rect 6404 875 6436 876
rect 6404 845 6405 875
rect 6405 845 6435 875
rect 6435 845 6436 875
rect 6404 844 6436 845
rect 6404 764 6436 796
rect 6404 684 6436 716
rect 6404 635 6436 636
rect 6404 605 6405 635
rect 6405 605 6435 635
rect 6435 605 6436 635
rect 6404 604 6436 605
rect 6404 555 6436 556
rect 6404 525 6405 555
rect 6405 525 6435 555
rect 6435 525 6436 555
rect 6404 524 6436 525
rect 6404 444 6436 476
rect 6404 395 6436 396
rect 6404 365 6405 395
rect 6405 365 6435 395
rect 6435 365 6436 395
rect 6404 364 6436 365
rect 6404 284 6436 316
rect 6404 235 6436 236
rect 6404 205 6405 235
rect 6405 205 6435 235
rect 6435 205 6436 235
rect 6404 204 6436 205
rect 6404 124 6436 156
rect 6404 75 6436 76
rect 6404 45 6405 75
rect 6405 45 6435 75
rect 6435 45 6436 75
rect 6404 44 6436 45
rect 6404 -5 6436 -4
rect 6404 -35 6405 -5
rect 6405 -35 6435 -5
rect 6435 -35 6436 -5
rect 6404 -36 6436 -35
rect 6404 -85 6436 -84
rect 6404 -115 6405 -85
rect 6405 -115 6435 -85
rect 6435 -115 6436 -85
rect 6404 -116 6436 -115
rect 6404 -165 6436 -164
rect 6404 -195 6405 -165
rect 6405 -195 6435 -165
rect 6435 -195 6436 -165
rect 6404 -196 6436 -195
rect 6404 -245 6436 -244
rect 6404 -275 6405 -245
rect 6405 -275 6435 -245
rect 6435 -275 6436 -245
rect 6404 -276 6436 -275
rect 6404 -325 6436 -324
rect 6404 -355 6405 -325
rect 6405 -355 6435 -325
rect 6435 -355 6436 -325
rect 6404 -356 6436 -355
rect 6404 -436 6436 -404
rect 6404 -485 6436 -484
rect 6404 -515 6405 -485
rect 6405 -515 6435 -485
rect 6435 -515 6436 -485
rect 6404 -516 6436 -515
rect 6404 -596 6436 -564
rect 6404 -645 6436 -644
rect 6404 -675 6405 -645
rect 6405 -675 6435 -645
rect 6435 -675 6436 -645
rect 6404 -676 6436 -675
rect 6404 -756 6436 -724
rect 6404 -805 6436 -804
rect 6404 -835 6405 -805
rect 6405 -835 6435 -805
rect 6435 -835 6436 -805
rect 6404 -836 6436 -835
rect 6404 -885 6436 -884
rect 6404 -915 6405 -885
rect 6405 -915 6435 -885
rect 6435 -915 6436 -885
rect 6404 -916 6436 -915
rect 6404 -996 6436 -964
rect 6404 -1076 6436 -1044
rect 6404 -1125 6436 -1124
rect 6404 -1155 6405 -1125
rect 6405 -1155 6435 -1125
rect 6435 -1155 6436 -1125
rect 6404 -1156 6436 -1155
rect 6404 -1205 6436 -1204
rect 6404 -1235 6405 -1205
rect 6405 -1235 6435 -1205
rect 6435 -1235 6436 -1205
rect 6404 -1236 6436 -1235
rect 6404 -1285 6436 -1284
rect 6404 -1315 6405 -1285
rect 6405 -1315 6435 -1285
rect 6435 -1315 6436 -1285
rect 6404 -1316 6436 -1315
rect 6404 -1365 6436 -1364
rect 6404 -1395 6405 -1365
rect 6405 -1395 6435 -1365
rect 6435 -1395 6436 -1365
rect 6404 -1396 6436 -1395
rect 6404 -1445 6436 -1444
rect 6404 -1475 6405 -1445
rect 6405 -1475 6435 -1445
rect 6435 -1475 6436 -1445
rect 6404 -1476 6436 -1475
rect 6404 -1525 6436 -1524
rect 6404 -1555 6405 -1525
rect 6405 -1555 6435 -1525
rect 6435 -1555 6436 -1525
rect 6404 -1556 6436 -1555
rect 6404 -1636 6436 -1604
rect 6404 -1716 6436 -1684
rect 6404 -1765 6436 -1764
rect 6404 -1795 6405 -1765
rect 6405 -1795 6435 -1765
rect 6435 -1795 6436 -1765
rect 6404 -1796 6436 -1795
rect 6404 -1845 6436 -1844
rect 6404 -1875 6405 -1845
rect 6405 -1875 6435 -1845
rect 6435 -1875 6436 -1845
rect 6404 -1876 6436 -1875
rect 6404 -1956 6436 -1924
rect 6404 -2005 6436 -2004
rect 6404 -2035 6405 -2005
rect 6405 -2035 6435 -2005
rect 6435 -2035 6436 -2005
rect 6404 -2036 6436 -2035
rect 6404 -2116 6436 -2084
rect 6404 -2165 6436 -2164
rect 6404 -2195 6405 -2165
rect 6405 -2195 6435 -2165
rect 6435 -2195 6436 -2165
rect 6404 -2196 6436 -2195
rect 6404 -2276 6436 -2244
rect 6404 -2325 6436 -2324
rect 6404 -2355 6405 -2325
rect 6405 -2355 6435 -2325
rect 6435 -2355 6436 -2325
rect 6404 -2356 6436 -2355
rect 6404 -2405 6436 -2404
rect 6404 -2435 6405 -2405
rect 6405 -2435 6435 -2405
rect 6435 -2435 6436 -2405
rect 6404 -2436 6436 -2435
rect 6404 -2485 6436 -2484
rect 6404 -2515 6405 -2485
rect 6405 -2515 6435 -2485
rect 6435 -2515 6436 -2485
rect 6404 -2516 6436 -2515
rect 6404 -2565 6436 -2564
rect 6404 -2595 6405 -2565
rect 6405 -2595 6435 -2565
rect 6435 -2595 6436 -2565
rect 6404 -2596 6436 -2595
rect 6404 -2645 6436 -2644
rect 6404 -2675 6405 -2645
rect 6405 -2675 6435 -2645
rect 6435 -2675 6436 -2645
rect 6404 -2676 6436 -2675
rect 6404 -2725 6436 -2724
rect 6404 -2755 6405 -2725
rect 6405 -2755 6435 -2725
rect 6435 -2755 6436 -2725
rect 6404 -2756 6436 -2755
rect 6404 -2836 6436 -2804
rect 6404 -2885 6436 -2884
rect 6404 -2915 6405 -2885
rect 6405 -2915 6435 -2885
rect 6435 -2915 6436 -2885
rect 6404 -2916 6436 -2915
rect 6404 -2996 6436 -2964
rect 6404 -3045 6436 -3044
rect 6404 -3075 6405 -3045
rect 6405 -3075 6435 -3045
rect 6435 -3075 6436 -3045
rect 6404 -3076 6436 -3075
rect 6404 -3156 6436 -3124
rect 6404 -3205 6436 -3204
rect 6404 -3235 6405 -3205
rect 6405 -3235 6435 -3205
rect 6435 -3235 6436 -3205
rect 6404 -3236 6436 -3235
rect 6404 -3285 6436 -3284
rect 6404 -3315 6405 -3285
rect 6405 -3315 6435 -3285
rect 6435 -3315 6436 -3285
rect 6404 -3316 6436 -3315
rect 6404 -3396 6436 -3364
rect 6404 -3476 6436 -3444
rect 6404 -3525 6436 -3524
rect 6404 -3555 6405 -3525
rect 6405 -3555 6435 -3525
rect 6435 -3555 6436 -3525
rect 6404 -3556 6436 -3555
rect 6404 -3605 6436 -3604
rect 6404 -3635 6405 -3605
rect 6405 -3635 6435 -3605
rect 6435 -3635 6436 -3605
rect 6404 -3636 6436 -3635
rect 6404 -3685 6436 -3684
rect 6404 -3715 6405 -3685
rect 6405 -3715 6435 -3685
rect 6435 -3715 6436 -3685
rect 6404 -3716 6436 -3715
rect 6484 1035 6516 1036
rect 6484 1005 6485 1035
rect 6485 1005 6515 1035
rect 6515 1005 6516 1035
rect 6484 1004 6516 1005
rect 6484 955 6516 956
rect 6484 925 6485 955
rect 6485 925 6515 955
rect 6515 925 6516 955
rect 6484 924 6516 925
rect 6484 875 6516 876
rect 6484 845 6485 875
rect 6485 845 6515 875
rect 6515 845 6516 875
rect 6484 844 6516 845
rect 6484 764 6516 796
rect 6484 684 6516 716
rect 6484 635 6516 636
rect 6484 605 6485 635
rect 6485 605 6515 635
rect 6515 605 6516 635
rect 6484 604 6516 605
rect 6484 555 6516 556
rect 6484 525 6485 555
rect 6485 525 6515 555
rect 6515 525 6516 555
rect 6484 524 6516 525
rect 6484 444 6516 476
rect 6484 395 6516 396
rect 6484 365 6485 395
rect 6485 365 6515 395
rect 6515 365 6516 395
rect 6484 364 6516 365
rect 6484 284 6516 316
rect 6484 235 6516 236
rect 6484 205 6485 235
rect 6485 205 6515 235
rect 6515 205 6516 235
rect 6484 204 6516 205
rect 6484 124 6516 156
rect 6484 75 6516 76
rect 6484 45 6485 75
rect 6485 45 6515 75
rect 6515 45 6516 75
rect 6484 44 6516 45
rect 6484 -5 6516 -4
rect 6484 -35 6485 -5
rect 6485 -35 6515 -5
rect 6515 -35 6516 -5
rect 6484 -36 6516 -35
rect 6484 -85 6516 -84
rect 6484 -115 6485 -85
rect 6485 -115 6515 -85
rect 6515 -115 6516 -85
rect 6484 -116 6516 -115
rect 6484 -165 6516 -164
rect 6484 -195 6485 -165
rect 6485 -195 6515 -165
rect 6515 -195 6516 -165
rect 6484 -196 6516 -195
rect 6484 -245 6516 -244
rect 6484 -275 6485 -245
rect 6485 -275 6515 -245
rect 6515 -275 6516 -245
rect 6484 -276 6516 -275
rect 6484 -325 6516 -324
rect 6484 -355 6485 -325
rect 6485 -355 6515 -325
rect 6515 -355 6516 -325
rect 6484 -356 6516 -355
rect 6484 -436 6516 -404
rect 6484 -485 6516 -484
rect 6484 -515 6485 -485
rect 6485 -515 6515 -485
rect 6515 -515 6516 -485
rect 6484 -516 6516 -515
rect 6484 -596 6516 -564
rect 6484 -645 6516 -644
rect 6484 -675 6485 -645
rect 6485 -675 6515 -645
rect 6515 -675 6516 -645
rect 6484 -676 6516 -675
rect 6484 -756 6516 -724
rect 6484 -805 6516 -804
rect 6484 -835 6485 -805
rect 6485 -835 6515 -805
rect 6515 -835 6516 -805
rect 6484 -836 6516 -835
rect 6484 -885 6516 -884
rect 6484 -915 6485 -885
rect 6485 -915 6515 -885
rect 6515 -915 6516 -885
rect 6484 -916 6516 -915
rect 6484 -996 6516 -964
rect 6484 -1076 6516 -1044
rect 6484 -1125 6516 -1124
rect 6484 -1155 6485 -1125
rect 6485 -1155 6515 -1125
rect 6515 -1155 6516 -1125
rect 6484 -1156 6516 -1155
rect 6484 -1205 6516 -1204
rect 6484 -1235 6485 -1205
rect 6485 -1235 6515 -1205
rect 6515 -1235 6516 -1205
rect 6484 -1236 6516 -1235
rect 6484 -1285 6516 -1284
rect 6484 -1315 6485 -1285
rect 6485 -1315 6515 -1285
rect 6515 -1315 6516 -1285
rect 6484 -1316 6516 -1315
rect 6484 -1365 6516 -1364
rect 6484 -1395 6485 -1365
rect 6485 -1395 6515 -1365
rect 6515 -1395 6516 -1365
rect 6484 -1396 6516 -1395
rect 6484 -1445 6516 -1444
rect 6484 -1475 6485 -1445
rect 6485 -1475 6515 -1445
rect 6515 -1475 6516 -1445
rect 6484 -1476 6516 -1475
rect 6484 -1525 6516 -1524
rect 6484 -1555 6485 -1525
rect 6485 -1555 6515 -1525
rect 6515 -1555 6516 -1525
rect 6484 -1556 6516 -1555
rect 6484 -1636 6516 -1604
rect 6484 -1716 6516 -1684
rect 6484 -1765 6516 -1764
rect 6484 -1795 6485 -1765
rect 6485 -1795 6515 -1765
rect 6515 -1795 6516 -1765
rect 6484 -1796 6516 -1795
rect 6484 -1845 6516 -1844
rect 6484 -1875 6485 -1845
rect 6485 -1875 6515 -1845
rect 6515 -1875 6516 -1845
rect 6484 -1876 6516 -1875
rect 6484 -1956 6516 -1924
rect 6484 -2005 6516 -2004
rect 6484 -2035 6485 -2005
rect 6485 -2035 6515 -2005
rect 6515 -2035 6516 -2005
rect 6484 -2036 6516 -2035
rect 6484 -2116 6516 -2084
rect 6484 -2165 6516 -2164
rect 6484 -2195 6485 -2165
rect 6485 -2195 6515 -2165
rect 6515 -2195 6516 -2165
rect 6484 -2196 6516 -2195
rect 6484 -2276 6516 -2244
rect 6484 -2325 6516 -2324
rect 6484 -2355 6485 -2325
rect 6485 -2355 6515 -2325
rect 6515 -2355 6516 -2325
rect 6484 -2356 6516 -2355
rect 6484 -2405 6516 -2404
rect 6484 -2435 6485 -2405
rect 6485 -2435 6515 -2405
rect 6515 -2435 6516 -2405
rect 6484 -2436 6516 -2435
rect 6484 -2485 6516 -2484
rect 6484 -2515 6485 -2485
rect 6485 -2515 6515 -2485
rect 6515 -2515 6516 -2485
rect 6484 -2516 6516 -2515
rect 6484 -2565 6516 -2564
rect 6484 -2595 6485 -2565
rect 6485 -2595 6515 -2565
rect 6515 -2595 6516 -2565
rect 6484 -2596 6516 -2595
rect 6484 -2645 6516 -2644
rect 6484 -2675 6485 -2645
rect 6485 -2675 6515 -2645
rect 6515 -2675 6516 -2645
rect 6484 -2676 6516 -2675
rect 6484 -2725 6516 -2724
rect 6484 -2755 6485 -2725
rect 6485 -2755 6515 -2725
rect 6515 -2755 6516 -2725
rect 6484 -2756 6516 -2755
rect 6484 -2836 6516 -2804
rect 6484 -2885 6516 -2884
rect 6484 -2915 6485 -2885
rect 6485 -2915 6515 -2885
rect 6515 -2915 6516 -2885
rect 6484 -2916 6516 -2915
rect 6484 -2996 6516 -2964
rect 6484 -3045 6516 -3044
rect 6484 -3075 6485 -3045
rect 6485 -3075 6515 -3045
rect 6515 -3075 6516 -3045
rect 6484 -3076 6516 -3075
rect 6484 -3156 6516 -3124
rect 6484 -3205 6516 -3204
rect 6484 -3235 6485 -3205
rect 6485 -3235 6515 -3205
rect 6515 -3235 6516 -3205
rect 6484 -3236 6516 -3235
rect 6484 -3285 6516 -3284
rect 6484 -3315 6485 -3285
rect 6485 -3315 6515 -3285
rect 6515 -3315 6516 -3285
rect 6484 -3316 6516 -3315
rect 6484 -3396 6516 -3364
rect 6484 -3476 6516 -3444
rect 6484 -3525 6516 -3524
rect 6484 -3555 6485 -3525
rect 6485 -3555 6515 -3525
rect 6515 -3555 6516 -3525
rect 6484 -3556 6516 -3555
rect 6484 -3605 6516 -3604
rect 6484 -3635 6485 -3605
rect 6485 -3635 6515 -3605
rect 6515 -3635 6516 -3605
rect 6484 -3636 6516 -3635
rect 6484 -3685 6516 -3684
rect 6484 -3715 6485 -3685
rect 6485 -3715 6515 -3685
rect 6515 -3715 6516 -3685
rect 6484 -3716 6516 -3715
rect 6564 1035 6596 1036
rect 6564 1005 6565 1035
rect 6565 1005 6595 1035
rect 6595 1005 6596 1035
rect 6564 1004 6596 1005
rect 6564 955 6596 956
rect 6564 925 6565 955
rect 6565 925 6595 955
rect 6595 925 6596 955
rect 6564 924 6596 925
rect 6564 875 6596 876
rect 6564 845 6565 875
rect 6565 845 6595 875
rect 6595 845 6596 875
rect 6564 844 6596 845
rect 6564 764 6596 796
rect 6564 684 6596 716
rect 6564 635 6596 636
rect 6564 605 6565 635
rect 6565 605 6595 635
rect 6595 605 6596 635
rect 6564 604 6596 605
rect 6564 555 6596 556
rect 6564 525 6565 555
rect 6565 525 6595 555
rect 6595 525 6596 555
rect 6564 524 6596 525
rect 6564 444 6596 476
rect 6564 395 6596 396
rect 6564 365 6565 395
rect 6565 365 6595 395
rect 6595 365 6596 395
rect 6564 364 6596 365
rect 6564 284 6596 316
rect 6564 235 6596 236
rect 6564 205 6565 235
rect 6565 205 6595 235
rect 6595 205 6596 235
rect 6564 204 6596 205
rect 6564 124 6596 156
rect 6564 75 6596 76
rect 6564 45 6565 75
rect 6565 45 6595 75
rect 6595 45 6596 75
rect 6564 44 6596 45
rect 6564 -5 6596 -4
rect 6564 -35 6565 -5
rect 6565 -35 6595 -5
rect 6595 -35 6596 -5
rect 6564 -36 6596 -35
rect 6564 -85 6596 -84
rect 6564 -115 6565 -85
rect 6565 -115 6595 -85
rect 6595 -115 6596 -85
rect 6564 -116 6596 -115
rect 6564 -165 6596 -164
rect 6564 -195 6565 -165
rect 6565 -195 6595 -165
rect 6595 -195 6596 -165
rect 6564 -196 6596 -195
rect 6564 -245 6596 -244
rect 6564 -275 6565 -245
rect 6565 -275 6595 -245
rect 6595 -275 6596 -245
rect 6564 -276 6596 -275
rect 6564 -325 6596 -324
rect 6564 -355 6565 -325
rect 6565 -355 6595 -325
rect 6595 -355 6596 -325
rect 6564 -356 6596 -355
rect 6564 -436 6596 -404
rect 6564 -485 6596 -484
rect 6564 -515 6565 -485
rect 6565 -515 6595 -485
rect 6595 -515 6596 -485
rect 6564 -516 6596 -515
rect 6564 -596 6596 -564
rect 6564 -645 6596 -644
rect 6564 -675 6565 -645
rect 6565 -675 6595 -645
rect 6595 -675 6596 -645
rect 6564 -676 6596 -675
rect 6564 -756 6596 -724
rect 6564 -805 6596 -804
rect 6564 -835 6565 -805
rect 6565 -835 6595 -805
rect 6595 -835 6596 -805
rect 6564 -836 6596 -835
rect 6564 -885 6596 -884
rect 6564 -915 6565 -885
rect 6565 -915 6595 -885
rect 6595 -915 6596 -885
rect 6564 -916 6596 -915
rect 6564 -996 6596 -964
rect 6564 -1076 6596 -1044
rect 6564 -1125 6596 -1124
rect 6564 -1155 6565 -1125
rect 6565 -1155 6595 -1125
rect 6595 -1155 6596 -1125
rect 6564 -1156 6596 -1155
rect 6564 -1205 6596 -1204
rect 6564 -1235 6565 -1205
rect 6565 -1235 6595 -1205
rect 6595 -1235 6596 -1205
rect 6564 -1236 6596 -1235
rect 6564 -1285 6596 -1284
rect 6564 -1315 6565 -1285
rect 6565 -1315 6595 -1285
rect 6595 -1315 6596 -1285
rect 6564 -1316 6596 -1315
rect 6564 -1365 6596 -1364
rect 6564 -1395 6565 -1365
rect 6565 -1395 6595 -1365
rect 6595 -1395 6596 -1365
rect 6564 -1396 6596 -1395
rect 6564 -1445 6596 -1444
rect 6564 -1475 6565 -1445
rect 6565 -1475 6595 -1445
rect 6595 -1475 6596 -1445
rect 6564 -1476 6596 -1475
rect 6564 -1525 6596 -1524
rect 6564 -1555 6565 -1525
rect 6565 -1555 6595 -1525
rect 6595 -1555 6596 -1525
rect 6564 -1556 6596 -1555
rect 6564 -1636 6596 -1604
rect 6564 -1716 6596 -1684
rect 6564 -1765 6596 -1764
rect 6564 -1795 6565 -1765
rect 6565 -1795 6595 -1765
rect 6595 -1795 6596 -1765
rect 6564 -1796 6596 -1795
rect 6564 -1845 6596 -1844
rect 6564 -1875 6565 -1845
rect 6565 -1875 6595 -1845
rect 6595 -1875 6596 -1845
rect 6564 -1876 6596 -1875
rect 6564 -1956 6596 -1924
rect 6564 -2005 6596 -2004
rect 6564 -2035 6565 -2005
rect 6565 -2035 6595 -2005
rect 6595 -2035 6596 -2005
rect 6564 -2036 6596 -2035
rect 6564 -2116 6596 -2084
rect 6564 -2165 6596 -2164
rect 6564 -2195 6565 -2165
rect 6565 -2195 6595 -2165
rect 6595 -2195 6596 -2165
rect 6564 -2196 6596 -2195
rect 6564 -2276 6596 -2244
rect 6564 -2325 6596 -2324
rect 6564 -2355 6565 -2325
rect 6565 -2355 6595 -2325
rect 6595 -2355 6596 -2325
rect 6564 -2356 6596 -2355
rect 6564 -2405 6596 -2404
rect 6564 -2435 6565 -2405
rect 6565 -2435 6595 -2405
rect 6595 -2435 6596 -2405
rect 6564 -2436 6596 -2435
rect 6564 -2485 6596 -2484
rect 6564 -2515 6565 -2485
rect 6565 -2515 6595 -2485
rect 6595 -2515 6596 -2485
rect 6564 -2516 6596 -2515
rect 6564 -2565 6596 -2564
rect 6564 -2595 6565 -2565
rect 6565 -2595 6595 -2565
rect 6595 -2595 6596 -2565
rect 6564 -2596 6596 -2595
rect 6564 -2645 6596 -2644
rect 6564 -2675 6565 -2645
rect 6565 -2675 6595 -2645
rect 6595 -2675 6596 -2645
rect 6564 -2676 6596 -2675
rect 6564 -2725 6596 -2724
rect 6564 -2755 6565 -2725
rect 6565 -2755 6595 -2725
rect 6595 -2755 6596 -2725
rect 6564 -2756 6596 -2755
rect 6564 -2836 6596 -2804
rect 6564 -2885 6596 -2884
rect 6564 -2915 6565 -2885
rect 6565 -2915 6595 -2885
rect 6595 -2915 6596 -2885
rect 6564 -2916 6596 -2915
rect 6564 -2996 6596 -2964
rect 6564 -3045 6596 -3044
rect 6564 -3075 6565 -3045
rect 6565 -3075 6595 -3045
rect 6595 -3075 6596 -3045
rect 6564 -3076 6596 -3075
rect 6564 -3156 6596 -3124
rect 6564 -3205 6596 -3204
rect 6564 -3235 6565 -3205
rect 6565 -3235 6595 -3205
rect 6595 -3235 6596 -3205
rect 6564 -3236 6596 -3235
rect 6564 -3285 6596 -3284
rect 6564 -3315 6565 -3285
rect 6565 -3315 6595 -3285
rect 6595 -3315 6596 -3285
rect 6564 -3316 6596 -3315
rect 6564 -3396 6596 -3364
rect 6564 -3476 6596 -3444
rect 6564 -3525 6596 -3524
rect 6564 -3555 6565 -3525
rect 6565 -3555 6595 -3525
rect 6595 -3555 6596 -3525
rect 6564 -3556 6596 -3555
rect 6564 -3605 6596 -3604
rect 6564 -3635 6565 -3605
rect 6565 -3635 6595 -3605
rect 6595 -3635 6596 -3605
rect 6564 -3636 6596 -3635
rect 6564 -3685 6596 -3684
rect 6564 -3715 6565 -3685
rect 6565 -3715 6595 -3685
rect 6595 -3715 6596 -3685
rect 6564 -3716 6596 -3715
rect 6644 1035 6676 1036
rect 6644 1005 6645 1035
rect 6645 1005 6675 1035
rect 6675 1005 6676 1035
rect 6644 1004 6676 1005
rect 6644 955 6676 956
rect 6644 925 6645 955
rect 6645 925 6675 955
rect 6675 925 6676 955
rect 6644 924 6676 925
rect 6644 875 6676 876
rect 6644 845 6645 875
rect 6645 845 6675 875
rect 6675 845 6676 875
rect 6644 844 6676 845
rect 6644 764 6676 796
rect 6644 684 6676 716
rect 6644 635 6676 636
rect 6644 605 6645 635
rect 6645 605 6675 635
rect 6675 605 6676 635
rect 6644 604 6676 605
rect 6644 555 6676 556
rect 6644 525 6645 555
rect 6645 525 6675 555
rect 6675 525 6676 555
rect 6644 524 6676 525
rect 6644 444 6676 476
rect 6644 395 6676 396
rect 6644 365 6645 395
rect 6645 365 6675 395
rect 6675 365 6676 395
rect 6644 364 6676 365
rect 6644 284 6676 316
rect 6644 235 6676 236
rect 6644 205 6645 235
rect 6645 205 6675 235
rect 6675 205 6676 235
rect 6644 204 6676 205
rect 6644 124 6676 156
rect 6644 75 6676 76
rect 6644 45 6645 75
rect 6645 45 6675 75
rect 6675 45 6676 75
rect 6644 44 6676 45
rect 6644 -5 6676 -4
rect 6644 -35 6645 -5
rect 6645 -35 6675 -5
rect 6675 -35 6676 -5
rect 6644 -36 6676 -35
rect 6644 -85 6676 -84
rect 6644 -115 6645 -85
rect 6645 -115 6675 -85
rect 6675 -115 6676 -85
rect 6644 -116 6676 -115
rect 6644 -165 6676 -164
rect 6644 -195 6645 -165
rect 6645 -195 6675 -165
rect 6675 -195 6676 -165
rect 6644 -196 6676 -195
rect 6644 -245 6676 -244
rect 6644 -275 6645 -245
rect 6645 -275 6675 -245
rect 6675 -275 6676 -245
rect 6644 -276 6676 -275
rect 6644 -325 6676 -324
rect 6644 -355 6645 -325
rect 6645 -355 6675 -325
rect 6675 -355 6676 -325
rect 6644 -356 6676 -355
rect 6644 -436 6676 -404
rect 6644 -485 6676 -484
rect 6644 -515 6645 -485
rect 6645 -515 6675 -485
rect 6675 -515 6676 -485
rect 6644 -516 6676 -515
rect 6644 -596 6676 -564
rect 6644 -645 6676 -644
rect 6644 -675 6645 -645
rect 6645 -675 6675 -645
rect 6675 -675 6676 -645
rect 6644 -676 6676 -675
rect 6644 -756 6676 -724
rect 6644 -805 6676 -804
rect 6644 -835 6645 -805
rect 6645 -835 6675 -805
rect 6675 -835 6676 -805
rect 6644 -836 6676 -835
rect 6644 -885 6676 -884
rect 6644 -915 6645 -885
rect 6645 -915 6675 -885
rect 6675 -915 6676 -885
rect 6644 -916 6676 -915
rect 6644 -996 6676 -964
rect 6644 -1076 6676 -1044
rect 6644 -1125 6676 -1124
rect 6644 -1155 6645 -1125
rect 6645 -1155 6675 -1125
rect 6675 -1155 6676 -1125
rect 6644 -1156 6676 -1155
rect 6644 -1205 6676 -1204
rect 6644 -1235 6645 -1205
rect 6645 -1235 6675 -1205
rect 6675 -1235 6676 -1205
rect 6644 -1236 6676 -1235
rect 6644 -1285 6676 -1284
rect 6644 -1315 6645 -1285
rect 6645 -1315 6675 -1285
rect 6675 -1315 6676 -1285
rect 6644 -1316 6676 -1315
rect 6644 -1365 6676 -1364
rect 6644 -1395 6645 -1365
rect 6645 -1395 6675 -1365
rect 6675 -1395 6676 -1365
rect 6644 -1396 6676 -1395
rect 6644 -1445 6676 -1444
rect 6644 -1475 6645 -1445
rect 6645 -1475 6675 -1445
rect 6675 -1475 6676 -1445
rect 6644 -1476 6676 -1475
rect 6644 -1525 6676 -1524
rect 6644 -1555 6645 -1525
rect 6645 -1555 6675 -1525
rect 6675 -1555 6676 -1525
rect 6644 -1556 6676 -1555
rect 6644 -1636 6676 -1604
rect 6644 -1716 6676 -1684
rect 6644 -1765 6676 -1764
rect 6644 -1795 6645 -1765
rect 6645 -1795 6675 -1765
rect 6675 -1795 6676 -1765
rect 6644 -1796 6676 -1795
rect 6644 -1845 6676 -1844
rect 6644 -1875 6645 -1845
rect 6645 -1875 6675 -1845
rect 6675 -1875 6676 -1845
rect 6644 -1876 6676 -1875
rect 6644 -1956 6676 -1924
rect 6644 -2005 6676 -2004
rect 6644 -2035 6645 -2005
rect 6645 -2035 6675 -2005
rect 6675 -2035 6676 -2005
rect 6644 -2036 6676 -2035
rect 6644 -2116 6676 -2084
rect 6644 -2165 6676 -2164
rect 6644 -2195 6645 -2165
rect 6645 -2195 6675 -2165
rect 6675 -2195 6676 -2165
rect 6644 -2196 6676 -2195
rect 6644 -2276 6676 -2244
rect 6644 -2325 6676 -2324
rect 6644 -2355 6645 -2325
rect 6645 -2355 6675 -2325
rect 6675 -2355 6676 -2325
rect 6644 -2356 6676 -2355
rect 6644 -2405 6676 -2404
rect 6644 -2435 6645 -2405
rect 6645 -2435 6675 -2405
rect 6675 -2435 6676 -2405
rect 6644 -2436 6676 -2435
rect 6644 -2485 6676 -2484
rect 6644 -2515 6645 -2485
rect 6645 -2515 6675 -2485
rect 6675 -2515 6676 -2485
rect 6644 -2516 6676 -2515
rect 6644 -2565 6676 -2564
rect 6644 -2595 6645 -2565
rect 6645 -2595 6675 -2565
rect 6675 -2595 6676 -2565
rect 6644 -2596 6676 -2595
rect 6644 -2645 6676 -2644
rect 6644 -2675 6645 -2645
rect 6645 -2675 6675 -2645
rect 6675 -2675 6676 -2645
rect 6644 -2676 6676 -2675
rect 6644 -2725 6676 -2724
rect 6644 -2755 6645 -2725
rect 6645 -2755 6675 -2725
rect 6675 -2755 6676 -2725
rect 6644 -2756 6676 -2755
rect 6644 -2836 6676 -2804
rect 6644 -2885 6676 -2884
rect 6644 -2915 6645 -2885
rect 6645 -2915 6675 -2885
rect 6675 -2915 6676 -2885
rect 6644 -2916 6676 -2915
rect 6644 -2996 6676 -2964
rect 6644 -3045 6676 -3044
rect 6644 -3075 6645 -3045
rect 6645 -3075 6675 -3045
rect 6675 -3075 6676 -3045
rect 6644 -3076 6676 -3075
rect 6644 -3156 6676 -3124
rect 6644 -3205 6676 -3204
rect 6644 -3235 6645 -3205
rect 6645 -3235 6675 -3205
rect 6675 -3235 6676 -3205
rect 6644 -3236 6676 -3235
rect 6644 -3285 6676 -3284
rect 6644 -3315 6645 -3285
rect 6645 -3315 6675 -3285
rect 6675 -3315 6676 -3285
rect 6644 -3316 6676 -3315
rect 6644 -3396 6676 -3364
rect 6644 -3476 6676 -3444
rect 6644 -3525 6676 -3524
rect 6644 -3555 6645 -3525
rect 6645 -3555 6675 -3525
rect 6675 -3555 6676 -3525
rect 6644 -3556 6676 -3555
rect 6644 -3605 6676 -3604
rect 6644 -3635 6645 -3605
rect 6645 -3635 6675 -3605
rect 6675 -3635 6676 -3605
rect 6644 -3636 6676 -3635
rect 6644 -3685 6676 -3684
rect 6644 -3715 6645 -3685
rect 6645 -3715 6675 -3685
rect 6675 -3715 6676 -3685
rect 6644 -3716 6676 -3715
rect 6724 1035 6756 1036
rect 6724 1005 6725 1035
rect 6725 1005 6755 1035
rect 6755 1005 6756 1035
rect 6724 1004 6756 1005
rect 6724 955 6756 956
rect 6724 925 6725 955
rect 6725 925 6755 955
rect 6755 925 6756 955
rect 6724 924 6756 925
rect 6724 875 6756 876
rect 6724 845 6725 875
rect 6725 845 6755 875
rect 6755 845 6756 875
rect 6724 844 6756 845
rect 6724 764 6756 796
rect 6724 684 6756 716
rect 6724 635 6756 636
rect 6724 605 6725 635
rect 6725 605 6755 635
rect 6755 605 6756 635
rect 6724 604 6756 605
rect 6724 555 6756 556
rect 6724 525 6725 555
rect 6725 525 6755 555
rect 6755 525 6756 555
rect 6724 524 6756 525
rect 6724 444 6756 476
rect 6724 395 6756 396
rect 6724 365 6725 395
rect 6725 365 6755 395
rect 6755 365 6756 395
rect 6724 364 6756 365
rect 6724 284 6756 316
rect 6724 235 6756 236
rect 6724 205 6725 235
rect 6725 205 6755 235
rect 6755 205 6756 235
rect 6724 204 6756 205
rect 6724 124 6756 156
rect 6724 75 6756 76
rect 6724 45 6725 75
rect 6725 45 6755 75
rect 6755 45 6756 75
rect 6724 44 6756 45
rect 6724 -5 6756 -4
rect 6724 -35 6725 -5
rect 6725 -35 6755 -5
rect 6755 -35 6756 -5
rect 6724 -36 6756 -35
rect 6724 -85 6756 -84
rect 6724 -115 6725 -85
rect 6725 -115 6755 -85
rect 6755 -115 6756 -85
rect 6724 -116 6756 -115
rect 6724 -165 6756 -164
rect 6724 -195 6725 -165
rect 6725 -195 6755 -165
rect 6755 -195 6756 -165
rect 6724 -196 6756 -195
rect 6724 -245 6756 -244
rect 6724 -275 6725 -245
rect 6725 -275 6755 -245
rect 6755 -275 6756 -245
rect 6724 -276 6756 -275
rect 6724 -325 6756 -324
rect 6724 -355 6725 -325
rect 6725 -355 6755 -325
rect 6755 -355 6756 -325
rect 6724 -356 6756 -355
rect 6724 -436 6756 -404
rect 6724 -485 6756 -484
rect 6724 -515 6725 -485
rect 6725 -515 6755 -485
rect 6755 -515 6756 -485
rect 6724 -516 6756 -515
rect 6724 -596 6756 -564
rect 6724 -645 6756 -644
rect 6724 -675 6725 -645
rect 6725 -675 6755 -645
rect 6755 -675 6756 -645
rect 6724 -676 6756 -675
rect 6724 -756 6756 -724
rect 6724 -805 6756 -804
rect 6724 -835 6725 -805
rect 6725 -835 6755 -805
rect 6755 -835 6756 -805
rect 6724 -836 6756 -835
rect 6724 -885 6756 -884
rect 6724 -915 6725 -885
rect 6725 -915 6755 -885
rect 6755 -915 6756 -885
rect 6724 -916 6756 -915
rect 6724 -996 6756 -964
rect 6724 -1076 6756 -1044
rect 6724 -1125 6756 -1124
rect 6724 -1155 6725 -1125
rect 6725 -1155 6755 -1125
rect 6755 -1155 6756 -1125
rect 6724 -1156 6756 -1155
rect 6724 -1205 6756 -1204
rect 6724 -1235 6725 -1205
rect 6725 -1235 6755 -1205
rect 6755 -1235 6756 -1205
rect 6724 -1236 6756 -1235
rect 6724 -1285 6756 -1284
rect 6724 -1315 6725 -1285
rect 6725 -1315 6755 -1285
rect 6755 -1315 6756 -1285
rect 6724 -1316 6756 -1315
rect 6724 -1365 6756 -1364
rect 6724 -1395 6725 -1365
rect 6725 -1395 6755 -1365
rect 6755 -1395 6756 -1365
rect 6724 -1396 6756 -1395
rect 6724 -1445 6756 -1444
rect 6724 -1475 6725 -1445
rect 6725 -1475 6755 -1445
rect 6755 -1475 6756 -1445
rect 6724 -1476 6756 -1475
rect 6724 -1525 6756 -1524
rect 6724 -1555 6725 -1525
rect 6725 -1555 6755 -1525
rect 6755 -1555 6756 -1525
rect 6724 -1556 6756 -1555
rect 6724 -1636 6756 -1604
rect 6724 -1716 6756 -1684
rect 6724 -1765 6756 -1764
rect 6724 -1795 6725 -1765
rect 6725 -1795 6755 -1765
rect 6755 -1795 6756 -1765
rect 6724 -1796 6756 -1795
rect 6724 -1845 6756 -1844
rect 6724 -1875 6725 -1845
rect 6725 -1875 6755 -1845
rect 6755 -1875 6756 -1845
rect 6724 -1876 6756 -1875
rect 6724 -1956 6756 -1924
rect 6724 -2005 6756 -2004
rect 6724 -2035 6725 -2005
rect 6725 -2035 6755 -2005
rect 6755 -2035 6756 -2005
rect 6724 -2036 6756 -2035
rect 6724 -2116 6756 -2084
rect 6724 -2165 6756 -2164
rect 6724 -2195 6725 -2165
rect 6725 -2195 6755 -2165
rect 6755 -2195 6756 -2165
rect 6724 -2196 6756 -2195
rect 6724 -2276 6756 -2244
rect 6724 -2325 6756 -2324
rect 6724 -2355 6725 -2325
rect 6725 -2355 6755 -2325
rect 6755 -2355 6756 -2325
rect 6724 -2356 6756 -2355
rect 6724 -2405 6756 -2404
rect 6724 -2435 6725 -2405
rect 6725 -2435 6755 -2405
rect 6755 -2435 6756 -2405
rect 6724 -2436 6756 -2435
rect 6724 -2485 6756 -2484
rect 6724 -2515 6725 -2485
rect 6725 -2515 6755 -2485
rect 6755 -2515 6756 -2485
rect 6724 -2516 6756 -2515
rect 6724 -2565 6756 -2564
rect 6724 -2595 6725 -2565
rect 6725 -2595 6755 -2565
rect 6755 -2595 6756 -2565
rect 6724 -2596 6756 -2595
rect 6724 -2645 6756 -2644
rect 6724 -2675 6725 -2645
rect 6725 -2675 6755 -2645
rect 6755 -2675 6756 -2645
rect 6724 -2676 6756 -2675
rect 6724 -2725 6756 -2724
rect 6724 -2755 6725 -2725
rect 6725 -2755 6755 -2725
rect 6755 -2755 6756 -2725
rect 6724 -2756 6756 -2755
rect 6724 -2836 6756 -2804
rect 6724 -2885 6756 -2884
rect 6724 -2915 6725 -2885
rect 6725 -2915 6755 -2885
rect 6755 -2915 6756 -2885
rect 6724 -2916 6756 -2915
rect 6724 -2996 6756 -2964
rect 6724 -3045 6756 -3044
rect 6724 -3075 6725 -3045
rect 6725 -3075 6755 -3045
rect 6755 -3075 6756 -3045
rect 6724 -3076 6756 -3075
rect 6724 -3156 6756 -3124
rect 6724 -3205 6756 -3204
rect 6724 -3235 6725 -3205
rect 6725 -3235 6755 -3205
rect 6755 -3235 6756 -3205
rect 6724 -3236 6756 -3235
rect 6724 -3285 6756 -3284
rect 6724 -3315 6725 -3285
rect 6725 -3315 6755 -3285
rect 6755 -3315 6756 -3285
rect 6724 -3316 6756 -3315
rect 6724 -3396 6756 -3364
rect 6724 -3476 6756 -3444
rect 6724 -3525 6756 -3524
rect 6724 -3555 6725 -3525
rect 6725 -3555 6755 -3525
rect 6755 -3555 6756 -3525
rect 6724 -3556 6756 -3555
rect 6724 -3605 6756 -3604
rect 6724 -3635 6725 -3605
rect 6725 -3635 6755 -3605
rect 6755 -3635 6756 -3605
rect 6724 -3636 6756 -3635
rect 6724 -3685 6756 -3684
rect 6724 -3715 6725 -3685
rect 6725 -3715 6755 -3685
rect 6755 -3715 6756 -3685
rect 6724 -3716 6756 -3715
rect 6804 1035 6836 1036
rect 6804 1005 6805 1035
rect 6805 1005 6835 1035
rect 6835 1005 6836 1035
rect 6804 1004 6836 1005
rect 6804 955 6836 956
rect 6804 925 6805 955
rect 6805 925 6835 955
rect 6835 925 6836 955
rect 6804 924 6836 925
rect 6804 875 6836 876
rect 6804 845 6805 875
rect 6805 845 6835 875
rect 6835 845 6836 875
rect 6804 844 6836 845
rect 6804 764 6836 796
rect 6804 684 6836 716
rect 6804 635 6836 636
rect 6804 605 6805 635
rect 6805 605 6835 635
rect 6835 605 6836 635
rect 6804 604 6836 605
rect 6804 555 6836 556
rect 6804 525 6805 555
rect 6805 525 6835 555
rect 6835 525 6836 555
rect 6804 524 6836 525
rect 6804 444 6836 476
rect 6804 395 6836 396
rect 6804 365 6805 395
rect 6805 365 6835 395
rect 6835 365 6836 395
rect 6804 364 6836 365
rect 6804 284 6836 316
rect 6804 235 6836 236
rect 6804 205 6805 235
rect 6805 205 6835 235
rect 6835 205 6836 235
rect 6804 204 6836 205
rect 6804 124 6836 156
rect 6804 75 6836 76
rect 6804 45 6805 75
rect 6805 45 6835 75
rect 6835 45 6836 75
rect 6804 44 6836 45
rect 6804 -5 6836 -4
rect 6804 -35 6805 -5
rect 6805 -35 6835 -5
rect 6835 -35 6836 -5
rect 6804 -36 6836 -35
rect 6804 -85 6836 -84
rect 6804 -115 6805 -85
rect 6805 -115 6835 -85
rect 6835 -115 6836 -85
rect 6804 -116 6836 -115
rect 6804 -165 6836 -164
rect 6804 -195 6805 -165
rect 6805 -195 6835 -165
rect 6835 -195 6836 -165
rect 6804 -196 6836 -195
rect 6804 -245 6836 -244
rect 6804 -275 6805 -245
rect 6805 -275 6835 -245
rect 6835 -275 6836 -245
rect 6804 -276 6836 -275
rect 6804 -325 6836 -324
rect 6804 -355 6805 -325
rect 6805 -355 6835 -325
rect 6835 -355 6836 -325
rect 6804 -356 6836 -355
rect 6804 -436 6836 -404
rect 6804 -485 6836 -484
rect 6804 -515 6805 -485
rect 6805 -515 6835 -485
rect 6835 -515 6836 -485
rect 6804 -516 6836 -515
rect 6804 -596 6836 -564
rect 6804 -645 6836 -644
rect 6804 -675 6805 -645
rect 6805 -675 6835 -645
rect 6835 -675 6836 -645
rect 6804 -676 6836 -675
rect 6804 -756 6836 -724
rect 6804 -805 6836 -804
rect 6804 -835 6805 -805
rect 6805 -835 6835 -805
rect 6835 -835 6836 -805
rect 6804 -836 6836 -835
rect 6804 -885 6836 -884
rect 6804 -915 6805 -885
rect 6805 -915 6835 -885
rect 6835 -915 6836 -885
rect 6804 -916 6836 -915
rect 6804 -996 6836 -964
rect 6804 -1076 6836 -1044
rect 6804 -1125 6836 -1124
rect 6804 -1155 6805 -1125
rect 6805 -1155 6835 -1125
rect 6835 -1155 6836 -1125
rect 6804 -1156 6836 -1155
rect 6804 -1205 6836 -1204
rect 6804 -1235 6805 -1205
rect 6805 -1235 6835 -1205
rect 6835 -1235 6836 -1205
rect 6804 -1236 6836 -1235
rect 6804 -1285 6836 -1284
rect 6804 -1315 6805 -1285
rect 6805 -1315 6835 -1285
rect 6835 -1315 6836 -1285
rect 6804 -1316 6836 -1315
rect 6804 -1365 6836 -1364
rect 6804 -1395 6805 -1365
rect 6805 -1395 6835 -1365
rect 6835 -1395 6836 -1365
rect 6804 -1396 6836 -1395
rect 6804 -1445 6836 -1444
rect 6804 -1475 6805 -1445
rect 6805 -1475 6835 -1445
rect 6835 -1475 6836 -1445
rect 6804 -1476 6836 -1475
rect 6804 -1525 6836 -1524
rect 6804 -1555 6805 -1525
rect 6805 -1555 6835 -1525
rect 6835 -1555 6836 -1525
rect 6804 -1556 6836 -1555
rect 6804 -1636 6836 -1604
rect 6804 -1716 6836 -1684
rect 6804 -1765 6836 -1764
rect 6804 -1795 6805 -1765
rect 6805 -1795 6835 -1765
rect 6835 -1795 6836 -1765
rect 6804 -1796 6836 -1795
rect 6804 -1845 6836 -1844
rect 6804 -1875 6805 -1845
rect 6805 -1875 6835 -1845
rect 6835 -1875 6836 -1845
rect 6804 -1876 6836 -1875
rect 6804 -1956 6836 -1924
rect 6804 -2005 6836 -2004
rect 6804 -2035 6805 -2005
rect 6805 -2035 6835 -2005
rect 6835 -2035 6836 -2005
rect 6804 -2036 6836 -2035
rect 6804 -2116 6836 -2084
rect 6804 -2165 6836 -2164
rect 6804 -2195 6805 -2165
rect 6805 -2195 6835 -2165
rect 6835 -2195 6836 -2165
rect 6804 -2196 6836 -2195
rect 6804 -2276 6836 -2244
rect 6804 -2325 6836 -2324
rect 6804 -2355 6805 -2325
rect 6805 -2355 6835 -2325
rect 6835 -2355 6836 -2325
rect 6804 -2356 6836 -2355
rect 6804 -2405 6836 -2404
rect 6804 -2435 6805 -2405
rect 6805 -2435 6835 -2405
rect 6835 -2435 6836 -2405
rect 6804 -2436 6836 -2435
rect 6804 -2485 6836 -2484
rect 6804 -2515 6805 -2485
rect 6805 -2515 6835 -2485
rect 6835 -2515 6836 -2485
rect 6804 -2516 6836 -2515
rect 6804 -2565 6836 -2564
rect 6804 -2595 6805 -2565
rect 6805 -2595 6835 -2565
rect 6835 -2595 6836 -2565
rect 6804 -2596 6836 -2595
rect 6804 -2645 6836 -2644
rect 6804 -2675 6805 -2645
rect 6805 -2675 6835 -2645
rect 6835 -2675 6836 -2645
rect 6804 -2676 6836 -2675
rect 6804 -2725 6836 -2724
rect 6804 -2755 6805 -2725
rect 6805 -2755 6835 -2725
rect 6835 -2755 6836 -2725
rect 6804 -2756 6836 -2755
rect 6804 -2836 6836 -2804
rect 6804 -2885 6836 -2884
rect 6804 -2915 6805 -2885
rect 6805 -2915 6835 -2885
rect 6835 -2915 6836 -2885
rect 6804 -2916 6836 -2915
rect 6804 -2996 6836 -2964
rect 6804 -3045 6836 -3044
rect 6804 -3075 6805 -3045
rect 6805 -3075 6835 -3045
rect 6835 -3075 6836 -3045
rect 6804 -3076 6836 -3075
rect 6804 -3156 6836 -3124
rect 6804 -3205 6836 -3204
rect 6804 -3235 6805 -3205
rect 6805 -3235 6835 -3205
rect 6835 -3235 6836 -3205
rect 6804 -3236 6836 -3235
rect 6804 -3285 6836 -3284
rect 6804 -3315 6805 -3285
rect 6805 -3315 6835 -3285
rect 6835 -3315 6836 -3285
rect 6804 -3316 6836 -3315
rect 6804 -3396 6836 -3364
rect 6804 -3476 6836 -3444
rect 6804 -3525 6836 -3524
rect 6804 -3555 6805 -3525
rect 6805 -3555 6835 -3525
rect 6835 -3555 6836 -3525
rect 6804 -3556 6836 -3555
rect 6804 -3605 6836 -3604
rect 6804 -3635 6805 -3605
rect 6805 -3635 6835 -3605
rect 6835 -3635 6836 -3605
rect 6804 -3636 6836 -3635
rect 6804 -3685 6836 -3684
rect 6804 -3715 6805 -3685
rect 6805 -3715 6835 -3685
rect 6835 -3715 6836 -3685
rect 6804 -3716 6836 -3715
rect 6884 1035 6916 1036
rect 6884 1005 6885 1035
rect 6885 1005 6915 1035
rect 6915 1005 6916 1035
rect 6884 1004 6916 1005
rect 6884 955 6916 956
rect 6884 925 6885 955
rect 6885 925 6915 955
rect 6915 925 6916 955
rect 6884 924 6916 925
rect 6884 875 6916 876
rect 6884 845 6885 875
rect 6885 845 6915 875
rect 6915 845 6916 875
rect 6884 844 6916 845
rect 6884 764 6916 796
rect 6884 684 6916 716
rect 6884 635 6916 636
rect 6884 605 6885 635
rect 6885 605 6915 635
rect 6915 605 6916 635
rect 6884 604 6916 605
rect 6884 555 6916 556
rect 6884 525 6885 555
rect 6885 525 6915 555
rect 6915 525 6916 555
rect 6884 524 6916 525
rect 6884 444 6916 476
rect 6884 395 6916 396
rect 6884 365 6885 395
rect 6885 365 6915 395
rect 6915 365 6916 395
rect 6884 364 6916 365
rect 6884 284 6916 316
rect 6884 235 6916 236
rect 6884 205 6885 235
rect 6885 205 6915 235
rect 6915 205 6916 235
rect 6884 204 6916 205
rect 6884 124 6916 156
rect 6884 75 6916 76
rect 6884 45 6885 75
rect 6885 45 6915 75
rect 6915 45 6916 75
rect 6884 44 6916 45
rect 6884 -5 6916 -4
rect 6884 -35 6885 -5
rect 6885 -35 6915 -5
rect 6915 -35 6916 -5
rect 6884 -36 6916 -35
rect 6884 -85 6916 -84
rect 6884 -115 6885 -85
rect 6885 -115 6915 -85
rect 6915 -115 6916 -85
rect 6884 -116 6916 -115
rect 6884 -165 6916 -164
rect 6884 -195 6885 -165
rect 6885 -195 6915 -165
rect 6915 -195 6916 -165
rect 6884 -196 6916 -195
rect 6884 -245 6916 -244
rect 6884 -275 6885 -245
rect 6885 -275 6915 -245
rect 6915 -275 6916 -245
rect 6884 -276 6916 -275
rect 6884 -325 6916 -324
rect 6884 -355 6885 -325
rect 6885 -355 6915 -325
rect 6915 -355 6916 -325
rect 6884 -356 6916 -355
rect 6884 -436 6916 -404
rect 6884 -485 6916 -484
rect 6884 -515 6885 -485
rect 6885 -515 6915 -485
rect 6915 -515 6916 -485
rect 6884 -516 6916 -515
rect 6884 -596 6916 -564
rect 6884 -645 6916 -644
rect 6884 -675 6885 -645
rect 6885 -675 6915 -645
rect 6915 -675 6916 -645
rect 6884 -676 6916 -675
rect 6884 -756 6916 -724
rect 6884 -805 6916 -804
rect 6884 -835 6885 -805
rect 6885 -835 6915 -805
rect 6915 -835 6916 -805
rect 6884 -836 6916 -835
rect 6884 -885 6916 -884
rect 6884 -915 6885 -885
rect 6885 -915 6915 -885
rect 6915 -915 6916 -885
rect 6884 -916 6916 -915
rect 6884 -996 6916 -964
rect 6884 -1076 6916 -1044
rect 6884 -1125 6916 -1124
rect 6884 -1155 6885 -1125
rect 6885 -1155 6915 -1125
rect 6915 -1155 6916 -1125
rect 6884 -1156 6916 -1155
rect 6884 -1205 6916 -1204
rect 6884 -1235 6885 -1205
rect 6885 -1235 6915 -1205
rect 6915 -1235 6916 -1205
rect 6884 -1236 6916 -1235
rect 6884 -1285 6916 -1284
rect 6884 -1315 6885 -1285
rect 6885 -1315 6915 -1285
rect 6915 -1315 6916 -1285
rect 6884 -1316 6916 -1315
rect 6884 -1365 6916 -1364
rect 6884 -1395 6885 -1365
rect 6885 -1395 6915 -1365
rect 6915 -1395 6916 -1365
rect 6884 -1396 6916 -1395
rect 6884 -1445 6916 -1444
rect 6884 -1475 6885 -1445
rect 6885 -1475 6915 -1445
rect 6915 -1475 6916 -1445
rect 6884 -1476 6916 -1475
rect 6884 -1525 6916 -1524
rect 6884 -1555 6885 -1525
rect 6885 -1555 6915 -1525
rect 6915 -1555 6916 -1525
rect 6884 -1556 6916 -1555
rect 6884 -1636 6916 -1604
rect 6884 -1716 6916 -1684
rect 6884 -1765 6916 -1764
rect 6884 -1795 6885 -1765
rect 6885 -1795 6915 -1765
rect 6915 -1795 6916 -1765
rect 6884 -1796 6916 -1795
rect 6884 -1845 6916 -1844
rect 6884 -1875 6885 -1845
rect 6885 -1875 6915 -1845
rect 6915 -1875 6916 -1845
rect 6884 -1876 6916 -1875
rect 6884 -1956 6916 -1924
rect 6884 -2005 6916 -2004
rect 6884 -2035 6885 -2005
rect 6885 -2035 6915 -2005
rect 6915 -2035 6916 -2005
rect 6884 -2036 6916 -2035
rect 6884 -2116 6916 -2084
rect 6884 -2165 6916 -2164
rect 6884 -2195 6885 -2165
rect 6885 -2195 6915 -2165
rect 6915 -2195 6916 -2165
rect 6884 -2196 6916 -2195
rect 6884 -2276 6916 -2244
rect 6884 -2325 6916 -2324
rect 6884 -2355 6885 -2325
rect 6885 -2355 6915 -2325
rect 6915 -2355 6916 -2325
rect 6884 -2356 6916 -2355
rect 6884 -2405 6916 -2404
rect 6884 -2435 6885 -2405
rect 6885 -2435 6915 -2405
rect 6915 -2435 6916 -2405
rect 6884 -2436 6916 -2435
rect 6884 -2485 6916 -2484
rect 6884 -2515 6885 -2485
rect 6885 -2515 6915 -2485
rect 6915 -2515 6916 -2485
rect 6884 -2516 6916 -2515
rect 6884 -2565 6916 -2564
rect 6884 -2595 6885 -2565
rect 6885 -2595 6915 -2565
rect 6915 -2595 6916 -2565
rect 6884 -2596 6916 -2595
rect 6884 -2645 6916 -2644
rect 6884 -2675 6885 -2645
rect 6885 -2675 6915 -2645
rect 6915 -2675 6916 -2645
rect 6884 -2676 6916 -2675
rect 6884 -2725 6916 -2724
rect 6884 -2755 6885 -2725
rect 6885 -2755 6915 -2725
rect 6915 -2755 6916 -2725
rect 6884 -2756 6916 -2755
rect 6884 -2836 6916 -2804
rect 6884 -2885 6916 -2884
rect 6884 -2915 6885 -2885
rect 6885 -2915 6915 -2885
rect 6915 -2915 6916 -2885
rect 6884 -2916 6916 -2915
rect 6884 -2996 6916 -2964
rect 6884 -3045 6916 -3044
rect 6884 -3075 6885 -3045
rect 6885 -3075 6915 -3045
rect 6915 -3075 6916 -3045
rect 6884 -3076 6916 -3075
rect 6884 -3156 6916 -3124
rect 6884 -3205 6916 -3204
rect 6884 -3235 6885 -3205
rect 6885 -3235 6915 -3205
rect 6915 -3235 6916 -3205
rect 6884 -3236 6916 -3235
rect 6884 -3285 6916 -3284
rect 6884 -3315 6885 -3285
rect 6885 -3315 6915 -3285
rect 6915 -3315 6916 -3285
rect 6884 -3316 6916 -3315
rect 6884 -3396 6916 -3364
rect 6884 -3476 6916 -3444
rect 6884 -3525 6916 -3524
rect 6884 -3555 6885 -3525
rect 6885 -3555 6915 -3525
rect 6915 -3555 6916 -3525
rect 6884 -3556 6916 -3555
rect 6884 -3605 6916 -3604
rect 6884 -3635 6885 -3605
rect 6885 -3635 6915 -3605
rect 6915 -3635 6916 -3605
rect 6884 -3636 6916 -3635
rect 6884 -3685 6916 -3684
rect 6884 -3715 6885 -3685
rect 6885 -3715 6915 -3685
rect 6915 -3715 6916 -3685
rect 6884 -3716 6916 -3715
rect 6964 1035 6996 1036
rect 6964 1005 6965 1035
rect 6965 1005 6995 1035
rect 6995 1005 6996 1035
rect 6964 1004 6996 1005
rect 6964 955 6996 956
rect 6964 925 6965 955
rect 6965 925 6995 955
rect 6995 925 6996 955
rect 6964 924 6996 925
rect 6964 875 6996 876
rect 6964 845 6965 875
rect 6965 845 6995 875
rect 6995 845 6996 875
rect 6964 844 6996 845
rect 6964 764 6996 796
rect 6964 684 6996 716
rect 6964 635 6996 636
rect 6964 605 6965 635
rect 6965 605 6995 635
rect 6995 605 6996 635
rect 6964 604 6996 605
rect 6964 555 6996 556
rect 6964 525 6965 555
rect 6965 525 6995 555
rect 6995 525 6996 555
rect 6964 524 6996 525
rect 6964 444 6996 476
rect 6964 395 6996 396
rect 6964 365 6965 395
rect 6965 365 6995 395
rect 6995 365 6996 395
rect 6964 364 6996 365
rect 6964 284 6996 316
rect 6964 235 6996 236
rect 6964 205 6965 235
rect 6965 205 6995 235
rect 6995 205 6996 235
rect 6964 204 6996 205
rect 6964 124 6996 156
rect 6964 75 6996 76
rect 6964 45 6965 75
rect 6965 45 6995 75
rect 6995 45 6996 75
rect 6964 44 6996 45
rect 6964 -5 6996 -4
rect 6964 -35 6965 -5
rect 6965 -35 6995 -5
rect 6995 -35 6996 -5
rect 6964 -36 6996 -35
rect 6964 -85 6996 -84
rect 6964 -115 6965 -85
rect 6965 -115 6995 -85
rect 6995 -115 6996 -85
rect 6964 -116 6996 -115
rect 6964 -165 6996 -164
rect 6964 -195 6965 -165
rect 6965 -195 6995 -165
rect 6995 -195 6996 -165
rect 6964 -196 6996 -195
rect 6964 -245 6996 -244
rect 6964 -275 6965 -245
rect 6965 -275 6995 -245
rect 6995 -275 6996 -245
rect 6964 -276 6996 -275
rect 6964 -325 6996 -324
rect 6964 -355 6965 -325
rect 6965 -355 6995 -325
rect 6995 -355 6996 -325
rect 6964 -356 6996 -355
rect 6964 -436 6996 -404
rect 6964 -485 6996 -484
rect 6964 -515 6965 -485
rect 6965 -515 6995 -485
rect 6995 -515 6996 -485
rect 6964 -516 6996 -515
rect 6964 -596 6996 -564
rect 6964 -645 6996 -644
rect 6964 -675 6965 -645
rect 6965 -675 6995 -645
rect 6995 -675 6996 -645
rect 6964 -676 6996 -675
rect 6964 -756 6996 -724
rect 6964 -805 6996 -804
rect 6964 -835 6965 -805
rect 6965 -835 6995 -805
rect 6995 -835 6996 -805
rect 6964 -836 6996 -835
rect 6964 -885 6996 -884
rect 6964 -915 6965 -885
rect 6965 -915 6995 -885
rect 6995 -915 6996 -885
rect 6964 -916 6996 -915
rect 6964 -996 6996 -964
rect 6964 -1076 6996 -1044
rect 6964 -1125 6996 -1124
rect 6964 -1155 6965 -1125
rect 6965 -1155 6995 -1125
rect 6995 -1155 6996 -1125
rect 6964 -1156 6996 -1155
rect 6964 -1205 6996 -1204
rect 6964 -1235 6965 -1205
rect 6965 -1235 6995 -1205
rect 6995 -1235 6996 -1205
rect 6964 -1236 6996 -1235
rect 6964 -1285 6996 -1284
rect 6964 -1315 6965 -1285
rect 6965 -1315 6995 -1285
rect 6995 -1315 6996 -1285
rect 6964 -1316 6996 -1315
rect 6964 -1365 6996 -1364
rect 6964 -1395 6965 -1365
rect 6965 -1395 6995 -1365
rect 6995 -1395 6996 -1365
rect 6964 -1396 6996 -1395
rect 6964 -1445 6996 -1444
rect 6964 -1475 6965 -1445
rect 6965 -1475 6995 -1445
rect 6995 -1475 6996 -1445
rect 6964 -1476 6996 -1475
rect 6964 -1525 6996 -1524
rect 6964 -1555 6965 -1525
rect 6965 -1555 6995 -1525
rect 6995 -1555 6996 -1525
rect 6964 -1556 6996 -1555
rect 6964 -1636 6996 -1604
rect 6964 -1716 6996 -1684
rect 6964 -1765 6996 -1764
rect 6964 -1795 6965 -1765
rect 6965 -1795 6995 -1765
rect 6995 -1795 6996 -1765
rect 6964 -1796 6996 -1795
rect 6964 -1845 6996 -1844
rect 6964 -1875 6965 -1845
rect 6965 -1875 6995 -1845
rect 6995 -1875 6996 -1845
rect 6964 -1876 6996 -1875
rect 6964 -1956 6996 -1924
rect 6964 -2005 6996 -2004
rect 6964 -2035 6965 -2005
rect 6965 -2035 6995 -2005
rect 6995 -2035 6996 -2005
rect 6964 -2036 6996 -2035
rect 6964 -2116 6996 -2084
rect 6964 -2165 6996 -2164
rect 6964 -2195 6965 -2165
rect 6965 -2195 6995 -2165
rect 6995 -2195 6996 -2165
rect 6964 -2196 6996 -2195
rect 6964 -2276 6996 -2244
rect 6964 -2325 6996 -2324
rect 6964 -2355 6965 -2325
rect 6965 -2355 6995 -2325
rect 6995 -2355 6996 -2325
rect 6964 -2356 6996 -2355
rect 6964 -2405 6996 -2404
rect 6964 -2435 6965 -2405
rect 6965 -2435 6995 -2405
rect 6995 -2435 6996 -2405
rect 6964 -2436 6996 -2435
rect 6964 -2485 6996 -2484
rect 6964 -2515 6965 -2485
rect 6965 -2515 6995 -2485
rect 6995 -2515 6996 -2485
rect 6964 -2516 6996 -2515
rect 6964 -2565 6996 -2564
rect 6964 -2595 6965 -2565
rect 6965 -2595 6995 -2565
rect 6995 -2595 6996 -2565
rect 6964 -2596 6996 -2595
rect 6964 -2645 6996 -2644
rect 6964 -2675 6965 -2645
rect 6965 -2675 6995 -2645
rect 6995 -2675 6996 -2645
rect 6964 -2676 6996 -2675
rect 6964 -2725 6996 -2724
rect 6964 -2755 6965 -2725
rect 6965 -2755 6995 -2725
rect 6995 -2755 6996 -2725
rect 6964 -2756 6996 -2755
rect 6964 -2836 6996 -2804
rect 6964 -2885 6996 -2884
rect 6964 -2915 6965 -2885
rect 6965 -2915 6995 -2885
rect 6995 -2915 6996 -2885
rect 6964 -2916 6996 -2915
rect 6964 -2996 6996 -2964
rect 6964 -3045 6996 -3044
rect 6964 -3075 6965 -3045
rect 6965 -3075 6995 -3045
rect 6995 -3075 6996 -3045
rect 6964 -3076 6996 -3075
rect 6964 -3156 6996 -3124
rect 6964 -3205 6996 -3204
rect 6964 -3235 6965 -3205
rect 6965 -3235 6995 -3205
rect 6995 -3235 6996 -3205
rect 6964 -3236 6996 -3235
rect 6964 -3285 6996 -3284
rect 6964 -3315 6965 -3285
rect 6965 -3315 6995 -3285
rect 6995 -3315 6996 -3285
rect 6964 -3316 6996 -3315
rect 6964 -3396 6996 -3364
rect 6964 -3476 6996 -3444
rect 6964 -3525 6996 -3524
rect 6964 -3555 6965 -3525
rect 6965 -3555 6995 -3525
rect 6995 -3555 6996 -3525
rect 6964 -3556 6996 -3555
rect 6964 -3605 6996 -3604
rect 6964 -3635 6965 -3605
rect 6965 -3635 6995 -3605
rect 6995 -3635 6996 -3605
rect 6964 -3636 6996 -3635
rect 6964 -3685 6996 -3684
rect 6964 -3715 6965 -3685
rect 6965 -3715 6995 -3685
rect 6995 -3715 6996 -3685
rect 6964 -3716 6996 -3715
rect 7044 1035 7076 1036
rect 7044 1005 7045 1035
rect 7045 1005 7075 1035
rect 7075 1005 7076 1035
rect 7044 1004 7076 1005
rect 7044 955 7076 956
rect 7044 925 7045 955
rect 7045 925 7075 955
rect 7075 925 7076 955
rect 7044 924 7076 925
rect 7044 875 7076 876
rect 7044 845 7045 875
rect 7045 845 7075 875
rect 7075 845 7076 875
rect 7044 844 7076 845
rect 7044 764 7076 796
rect 7044 684 7076 716
rect 7044 635 7076 636
rect 7044 605 7045 635
rect 7045 605 7075 635
rect 7075 605 7076 635
rect 7044 604 7076 605
rect 7044 555 7076 556
rect 7044 525 7045 555
rect 7045 525 7075 555
rect 7075 525 7076 555
rect 7044 524 7076 525
rect 7044 444 7076 476
rect 7044 395 7076 396
rect 7044 365 7045 395
rect 7045 365 7075 395
rect 7075 365 7076 395
rect 7044 364 7076 365
rect 7044 284 7076 316
rect 7044 235 7076 236
rect 7044 205 7045 235
rect 7045 205 7075 235
rect 7075 205 7076 235
rect 7044 204 7076 205
rect 7044 124 7076 156
rect 7044 75 7076 76
rect 7044 45 7045 75
rect 7045 45 7075 75
rect 7075 45 7076 75
rect 7044 44 7076 45
rect 7044 -5 7076 -4
rect 7044 -35 7045 -5
rect 7045 -35 7075 -5
rect 7075 -35 7076 -5
rect 7044 -36 7076 -35
rect 7044 -85 7076 -84
rect 7044 -115 7045 -85
rect 7045 -115 7075 -85
rect 7075 -115 7076 -85
rect 7044 -116 7076 -115
rect 7044 -165 7076 -164
rect 7044 -195 7045 -165
rect 7045 -195 7075 -165
rect 7075 -195 7076 -165
rect 7044 -196 7076 -195
rect 7044 -245 7076 -244
rect 7044 -275 7045 -245
rect 7045 -275 7075 -245
rect 7075 -275 7076 -245
rect 7044 -276 7076 -275
rect 7044 -325 7076 -324
rect 7044 -355 7045 -325
rect 7045 -355 7075 -325
rect 7075 -355 7076 -325
rect 7044 -356 7076 -355
rect 7044 -436 7076 -404
rect 7044 -485 7076 -484
rect 7044 -515 7045 -485
rect 7045 -515 7075 -485
rect 7075 -515 7076 -485
rect 7044 -516 7076 -515
rect 7044 -596 7076 -564
rect 7044 -645 7076 -644
rect 7044 -675 7045 -645
rect 7045 -675 7075 -645
rect 7075 -675 7076 -645
rect 7044 -676 7076 -675
rect 7044 -756 7076 -724
rect 7044 -805 7076 -804
rect 7044 -835 7045 -805
rect 7045 -835 7075 -805
rect 7075 -835 7076 -805
rect 7044 -836 7076 -835
rect 7044 -885 7076 -884
rect 7044 -915 7045 -885
rect 7045 -915 7075 -885
rect 7075 -915 7076 -885
rect 7044 -916 7076 -915
rect 7044 -996 7076 -964
rect 7044 -1076 7076 -1044
rect 7044 -1125 7076 -1124
rect 7044 -1155 7045 -1125
rect 7045 -1155 7075 -1125
rect 7075 -1155 7076 -1125
rect 7044 -1156 7076 -1155
rect 7044 -1205 7076 -1204
rect 7044 -1235 7045 -1205
rect 7045 -1235 7075 -1205
rect 7075 -1235 7076 -1205
rect 7044 -1236 7076 -1235
rect 7044 -1285 7076 -1284
rect 7044 -1315 7045 -1285
rect 7045 -1315 7075 -1285
rect 7075 -1315 7076 -1285
rect 7044 -1316 7076 -1315
rect 7044 -1365 7076 -1364
rect 7044 -1395 7045 -1365
rect 7045 -1395 7075 -1365
rect 7075 -1395 7076 -1365
rect 7044 -1396 7076 -1395
rect 7044 -1445 7076 -1444
rect 7044 -1475 7045 -1445
rect 7045 -1475 7075 -1445
rect 7075 -1475 7076 -1445
rect 7044 -1476 7076 -1475
rect 7044 -1525 7076 -1524
rect 7044 -1555 7045 -1525
rect 7045 -1555 7075 -1525
rect 7075 -1555 7076 -1525
rect 7044 -1556 7076 -1555
rect 7044 -1636 7076 -1604
rect 7044 -1716 7076 -1684
rect 7044 -1765 7076 -1764
rect 7044 -1795 7045 -1765
rect 7045 -1795 7075 -1765
rect 7075 -1795 7076 -1765
rect 7044 -1796 7076 -1795
rect 7044 -1845 7076 -1844
rect 7044 -1875 7045 -1845
rect 7045 -1875 7075 -1845
rect 7075 -1875 7076 -1845
rect 7044 -1876 7076 -1875
rect 7044 -1956 7076 -1924
rect 7044 -2005 7076 -2004
rect 7044 -2035 7045 -2005
rect 7045 -2035 7075 -2005
rect 7075 -2035 7076 -2005
rect 7044 -2036 7076 -2035
rect 7044 -2116 7076 -2084
rect 7044 -2165 7076 -2164
rect 7044 -2195 7045 -2165
rect 7045 -2195 7075 -2165
rect 7075 -2195 7076 -2165
rect 7044 -2196 7076 -2195
rect 7044 -2276 7076 -2244
rect 7044 -2325 7076 -2324
rect 7044 -2355 7045 -2325
rect 7045 -2355 7075 -2325
rect 7075 -2355 7076 -2325
rect 7044 -2356 7076 -2355
rect 7044 -2405 7076 -2404
rect 7044 -2435 7045 -2405
rect 7045 -2435 7075 -2405
rect 7075 -2435 7076 -2405
rect 7044 -2436 7076 -2435
rect 7044 -2485 7076 -2484
rect 7044 -2515 7045 -2485
rect 7045 -2515 7075 -2485
rect 7075 -2515 7076 -2485
rect 7044 -2516 7076 -2515
rect 7044 -2565 7076 -2564
rect 7044 -2595 7045 -2565
rect 7045 -2595 7075 -2565
rect 7075 -2595 7076 -2565
rect 7044 -2596 7076 -2595
rect 7044 -2645 7076 -2644
rect 7044 -2675 7045 -2645
rect 7045 -2675 7075 -2645
rect 7075 -2675 7076 -2645
rect 7044 -2676 7076 -2675
rect 7044 -2725 7076 -2724
rect 7044 -2755 7045 -2725
rect 7045 -2755 7075 -2725
rect 7075 -2755 7076 -2725
rect 7044 -2756 7076 -2755
rect 7044 -2836 7076 -2804
rect 7044 -2885 7076 -2884
rect 7044 -2915 7045 -2885
rect 7045 -2915 7075 -2885
rect 7075 -2915 7076 -2885
rect 7044 -2916 7076 -2915
rect 7044 -2996 7076 -2964
rect 7044 -3045 7076 -3044
rect 7044 -3075 7045 -3045
rect 7045 -3075 7075 -3045
rect 7075 -3075 7076 -3045
rect 7044 -3076 7076 -3075
rect 7044 -3156 7076 -3124
rect 7044 -3205 7076 -3204
rect 7044 -3235 7045 -3205
rect 7045 -3235 7075 -3205
rect 7075 -3235 7076 -3205
rect 7044 -3236 7076 -3235
rect 7044 -3285 7076 -3284
rect 7044 -3315 7045 -3285
rect 7045 -3315 7075 -3285
rect 7075 -3315 7076 -3285
rect 7044 -3316 7076 -3315
rect 7044 -3396 7076 -3364
rect 7044 -3476 7076 -3444
rect 7044 -3525 7076 -3524
rect 7044 -3555 7045 -3525
rect 7045 -3555 7075 -3525
rect 7075 -3555 7076 -3525
rect 7044 -3556 7076 -3555
rect 7044 -3605 7076 -3604
rect 7044 -3635 7045 -3605
rect 7045 -3635 7075 -3605
rect 7075 -3635 7076 -3605
rect 7044 -3636 7076 -3635
rect 7044 -3685 7076 -3684
rect 7044 -3715 7045 -3685
rect 7045 -3715 7075 -3685
rect 7075 -3715 7076 -3685
rect 7044 -3716 7076 -3715
rect 7124 1035 7156 1036
rect 7124 1005 7125 1035
rect 7125 1005 7155 1035
rect 7155 1005 7156 1035
rect 7124 1004 7156 1005
rect 7124 955 7156 956
rect 7124 925 7125 955
rect 7125 925 7155 955
rect 7155 925 7156 955
rect 7124 924 7156 925
rect 7124 875 7156 876
rect 7124 845 7125 875
rect 7125 845 7155 875
rect 7155 845 7156 875
rect 7124 844 7156 845
rect 7124 764 7156 796
rect 7124 684 7156 716
rect 7124 635 7156 636
rect 7124 605 7125 635
rect 7125 605 7155 635
rect 7155 605 7156 635
rect 7124 604 7156 605
rect 7124 555 7156 556
rect 7124 525 7125 555
rect 7125 525 7155 555
rect 7155 525 7156 555
rect 7124 524 7156 525
rect 7124 444 7156 476
rect 7124 395 7156 396
rect 7124 365 7125 395
rect 7125 365 7155 395
rect 7155 365 7156 395
rect 7124 364 7156 365
rect 7124 284 7156 316
rect 7124 235 7156 236
rect 7124 205 7125 235
rect 7125 205 7155 235
rect 7155 205 7156 235
rect 7124 204 7156 205
rect 7124 124 7156 156
rect 7124 75 7156 76
rect 7124 45 7125 75
rect 7125 45 7155 75
rect 7155 45 7156 75
rect 7124 44 7156 45
rect 7124 -5 7156 -4
rect 7124 -35 7125 -5
rect 7125 -35 7155 -5
rect 7155 -35 7156 -5
rect 7124 -36 7156 -35
rect 7124 -85 7156 -84
rect 7124 -115 7125 -85
rect 7125 -115 7155 -85
rect 7155 -115 7156 -85
rect 7124 -116 7156 -115
rect 7124 -165 7156 -164
rect 7124 -195 7125 -165
rect 7125 -195 7155 -165
rect 7155 -195 7156 -165
rect 7124 -196 7156 -195
rect 7124 -245 7156 -244
rect 7124 -275 7125 -245
rect 7125 -275 7155 -245
rect 7155 -275 7156 -245
rect 7124 -276 7156 -275
rect 7124 -325 7156 -324
rect 7124 -355 7125 -325
rect 7125 -355 7155 -325
rect 7155 -355 7156 -325
rect 7124 -356 7156 -355
rect 7124 -436 7156 -404
rect 7124 -485 7156 -484
rect 7124 -515 7125 -485
rect 7125 -515 7155 -485
rect 7155 -515 7156 -485
rect 7124 -516 7156 -515
rect 7124 -596 7156 -564
rect 7124 -645 7156 -644
rect 7124 -675 7125 -645
rect 7125 -675 7155 -645
rect 7155 -675 7156 -645
rect 7124 -676 7156 -675
rect 7124 -756 7156 -724
rect 7124 -805 7156 -804
rect 7124 -835 7125 -805
rect 7125 -835 7155 -805
rect 7155 -835 7156 -805
rect 7124 -836 7156 -835
rect 7124 -885 7156 -884
rect 7124 -915 7125 -885
rect 7125 -915 7155 -885
rect 7155 -915 7156 -885
rect 7124 -916 7156 -915
rect 7124 -996 7156 -964
rect 7124 -1076 7156 -1044
rect 7124 -1125 7156 -1124
rect 7124 -1155 7125 -1125
rect 7125 -1155 7155 -1125
rect 7155 -1155 7156 -1125
rect 7124 -1156 7156 -1155
rect 7124 -1205 7156 -1204
rect 7124 -1235 7125 -1205
rect 7125 -1235 7155 -1205
rect 7155 -1235 7156 -1205
rect 7124 -1236 7156 -1235
rect 7124 -1285 7156 -1284
rect 7124 -1315 7125 -1285
rect 7125 -1315 7155 -1285
rect 7155 -1315 7156 -1285
rect 7124 -1316 7156 -1315
rect 7124 -1365 7156 -1364
rect 7124 -1395 7125 -1365
rect 7125 -1395 7155 -1365
rect 7155 -1395 7156 -1365
rect 7124 -1396 7156 -1395
rect 7124 -1445 7156 -1444
rect 7124 -1475 7125 -1445
rect 7125 -1475 7155 -1445
rect 7155 -1475 7156 -1445
rect 7124 -1476 7156 -1475
rect 7124 -1525 7156 -1524
rect 7124 -1555 7125 -1525
rect 7125 -1555 7155 -1525
rect 7155 -1555 7156 -1525
rect 7124 -1556 7156 -1555
rect 7124 -1636 7156 -1604
rect 7124 -1716 7156 -1684
rect 7124 -1765 7156 -1764
rect 7124 -1795 7125 -1765
rect 7125 -1795 7155 -1765
rect 7155 -1795 7156 -1765
rect 7124 -1796 7156 -1795
rect 7124 -1845 7156 -1844
rect 7124 -1875 7125 -1845
rect 7125 -1875 7155 -1845
rect 7155 -1875 7156 -1845
rect 7124 -1876 7156 -1875
rect 7124 -1956 7156 -1924
rect 7124 -2005 7156 -2004
rect 7124 -2035 7125 -2005
rect 7125 -2035 7155 -2005
rect 7155 -2035 7156 -2005
rect 7124 -2036 7156 -2035
rect 7124 -2116 7156 -2084
rect 7124 -2165 7156 -2164
rect 7124 -2195 7125 -2165
rect 7125 -2195 7155 -2165
rect 7155 -2195 7156 -2165
rect 7124 -2196 7156 -2195
rect 7124 -2276 7156 -2244
rect 7124 -2325 7156 -2324
rect 7124 -2355 7125 -2325
rect 7125 -2355 7155 -2325
rect 7155 -2355 7156 -2325
rect 7124 -2356 7156 -2355
rect 7124 -2405 7156 -2404
rect 7124 -2435 7125 -2405
rect 7125 -2435 7155 -2405
rect 7155 -2435 7156 -2405
rect 7124 -2436 7156 -2435
rect 7124 -2485 7156 -2484
rect 7124 -2515 7125 -2485
rect 7125 -2515 7155 -2485
rect 7155 -2515 7156 -2485
rect 7124 -2516 7156 -2515
rect 7124 -2565 7156 -2564
rect 7124 -2595 7125 -2565
rect 7125 -2595 7155 -2565
rect 7155 -2595 7156 -2565
rect 7124 -2596 7156 -2595
rect 7124 -2645 7156 -2644
rect 7124 -2675 7125 -2645
rect 7125 -2675 7155 -2645
rect 7155 -2675 7156 -2645
rect 7124 -2676 7156 -2675
rect 7124 -2725 7156 -2724
rect 7124 -2755 7125 -2725
rect 7125 -2755 7155 -2725
rect 7155 -2755 7156 -2725
rect 7124 -2756 7156 -2755
rect 7124 -2836 7156 -2804
rect 7124 -2885 7156 -2884
rect 7124 -2915 7125 -2885
rect 7125 -2915 7155 -2885
rect 7155 -2915 7156 -2885
rect 7124 -2916 7156 -2915
rect 7124 -2996 7156 -2964
rect 7124 -3045 7156 -3044
rect 7124 -3075 7125 -3045
rect 7125 -3075 7155 -3045
rect 7155 -3075 7156 -3045
rect 7124 -3076 7156 -3075
rect 7124 -3156 7156 -3124
rect 7124 -3205 7156 -3204
rect 7124 -3235 7125 -3205
rect 7125 -3235 7155 -3205
rect 7155 -3235 7156 -3205
rect 7124 -3236 7156 -3235
rect 7124 -3285 7156 -3284
rect 7124 -3315 7125 -3285
rect 7125 -3315 7155 -3285
rect 7155 -3315 7156 -3285
rect 7124 -3316 7156 -3315
rect 7124 -3396 7156 -3364
rect 7124 -3476 7156 -3444
rect 7124 -3525 7156 -3524
rect 7124 -3555 7125 -3525
rect 7125 -3555 7155 -3525
rect 7155 -3555 7156 -3525
rect 7124 -3556 7156 -3555
rect 7124 -3605 7156 -3604
rect 7124 -3635 7125 -3605
rect 7125 -3635 7155 -3605
rect 7155 -3635 7156 -3605
rect 7124 -3636 7156 -3635
rect 7124 -3685 7156 -3684
rect 7124 -3715 7125 -3685
rect 7125 -3715 7155 -3685
rect 7155 -3715 7156 -3685
rect 7124 -3716 7156 -3715
rect 7204 1035 7236 1036
rect 7204 1005 7205 1035
rect 7205 1005 7235 1035
rect 7235 1005 7236 1035
rect 7204 1004 7236 1005
rect 7204 955 7236 956
rect 7204 925 7205 955
rect 7205 925 7235 955
rect 7235 925 7236 955
rect 7204 924 7236 925
rect 7204 875 7236 876
rect 7204 845 7205 875
rect 7205 845 7235 875
rect 7235 845 7236 875
rect 7204 844 7236 845
rect 7204 764 7236 796
rect 7204 684 7236 716
rect 7204 635 7236 636
rect 7204 605 7205 635
rect 7205 605 7235 635
rect 7235 605 7236 635
rect 7204 604 7236 605
rect 7204 555 7236 556
rect 7204 525 7205 555
rect 7205 525 7235 555
rect 7235 525 7236 555
rect 7204 524 7236 525
rect 7204 444 7236 476
rect 7204 395 7236 396
rect 7204 365 7205 395
rect 7205 365 7235 395
rect 7235 365 7236 395
rect 7204 364 7236 365
rect 7204 284 7236 316
rect 7204 235 7236 236
rect 7204 205 7205 235
rect 7205 205 7235 235
rect 7235 205 7236 235
rect 7204 204 7236 205
rect 7204 124 7236 156
rect 7204 75 7236 76
rect 7204 45 7205 75
rect 7205 45 7235 75
rect 7235 45 7236 75
rect 7204 44 7236 45
rect 7204 -5 7236 -4
rect 7204 -35 7205 -5
rect 7205 -35 7235 -5
rect 7235 -35 7236 -5
rect 7204 -36 7236 -35
rect 7204 -85 7236 -84
rect 7204 -115 7205 -85
rect 7205 -115 7235 -85
rect 7235 -115 7236 -85
rect 7204 -116 7236 -115
rect 7204 -165 7236 -164
rect 7204 -195 7205 -165
rect 7205 -195 7235 -165
rect 7235 -195 7236 -165
rect 7204 -196 7236 -195
rect 7204 -245 7236 -244
rect 7204 -275 7205 -245
rect 7205 -275 7235 -245
rect 7235 -275 7236 -245
rect 7204 -276 7236 -275
rect 7204 -325 7236 -324
rect 7204 -355 7205 -325
rect 7205 -355 7235 -325
rect 7235 -355 7236 -325
rect 7204 -356 7236 -355
rect 7204 -436 7236 -404
rect 7204 -485 7236 -484
rect 7204 -515 7205 -485
rect 7205 -515 7235 -485
rect 7235 -515 7236 -485
rect 7204 -516 7236 -515
rect 7204 -596 7236 -564
rect 7204 -645 7236 -644
rect 7204 -675 7205 -645
rect 7205 -675 7235 -645
rect 7235 -675 7236 -645
rect 7204 -676 7236 -675
rect 7204 -756 7236 -724
rect 7204 -805 7236 -804
rect 7204 -835 7205 -805
rect 7205 -835 7235 -805
rect 7235 -835 7236 -805
rect 7204 -836 7236 -835
rect 7204 -885 7236 -884
rect 7204 -915 7205 -885
rect 7205 -915 7235 -885
rect 7235 -915 7236 -885
rect 7204 -916 7236 -915
rect 7204 -996 7236 -964
rect 7204 -1076 7236 -1044
rect 7204 -1125 7236 -1124
rect 7204 -1155 7205 -1125
rect 7205 -1155 7235 -1125
rect 7235 -1155 7236 -1125
rect 7204 -1156 7236 -1155
rect 7204 -1205 7236 -1204
rect 7204 -1235 7205 -1205
rect 7205 -1235 7235 -1205
rect 7235 -1235 7236 -1205
rect 7204 -1236 7236 -1235
rect 7204 -1285 7236 -1284
rect 7204 -1315 7205 -1285
rect 7205 -1315 7235 -1285
rect 7235 -1315 7236 -1285
rect 7204 -1316 7236 -1315
rect 7204 -1365 7236 -1364
rect 7204 -1395 7205 -1365
rect 7205 -1395 7235 -1365
rect 7235 -1395 7236 -1365
rect 7204 -1396 7236 -1395
rect 7204 -1445 7236 -1444
rect 7204 -1475 7205 -1445
rect 7205 -1475 7235 -1445
rect 7235 -1475 7236 -1445
rect 7204 -1476 7236 -1475
rect 7204 -1525 7236 -1524
rect 7204 -1555 7205 -1525
rect 7205 -1555 7235 -1525
rect 7235 -1555 7236 -1525
rect 7204 -1556 7236 -1555
rect 7204 -1636 7236 -1604
rect 7204 -1716 7236 -1684
rect 7204 -1765 7236 -1764
rect 7204 -1795 7205 -1765
rect 7205 -1795 7235 -1765
rect 7235 -1795 7236 -1765
rect 7204 -1796 7236 -1795
rect 7204 -1845 7236 -1844
rect 7204 -1875 7205 -1845
rect 7205 -1875 7235 -1845
rect 7235 -1875 7236 -1845
rect 7204 -1876 7236 -1875
rect 7204 -1956 7236 -1924
rect 7204 -2005 7236 -2004
rect 7204 -2035 7205 -2005
rect 7205 -2035 7235 -2005
rect 7235 -2035 7236 -2005
rect 7204 -2036 7236 -2035
rect 7204 -2116 7236 -2084
rect 7204 -2165 7236 -2164
rect 7204 -2195 7205 -2165
rect 7205 -2195 7235 -2165
rect 7235 -2195 7236 -2165
rect 7204 -2196 7236 -2195
rect 7204 -2276 7236 -2244
rect 7204 -2325 7236 -2324
rect 7204 -2355 7205 -2325
rect 7205 -2355 7235 -2325
rect 7235 -2355 7236 -2325
rect 7204 -2356 7236 -2355
rect 7204 -2405 7236 -2404
rect 7204 -2435 7205 -2405
rect 7205 -2435 7235 -2405
rect 7235 -2435 7236 -2405
rect 7204 -2436 7236 -2435
rect 7204 -2485 7236 -2484
rect 7204 -2515 7205 -2485
rect 7205 -2515 7235 -2485
rect 7235 -2515 7236 -2485
rect 7204 -2516 7236 -2515
rect 7204 -2565 7236 -2564
rect 7204 -2595 7205 -2565
rect 7205 -2595 7235 -2565
rect 7235 -2595 7236 -2565
rect 7204 -2596 7236 -2595
rect 7204 -2645 7236 -2644
rect 7204 -2675 7205 -2645
rect 7205 -2675 7235 -2645
rect 7235 -2675 7236 -2645
rect 7204 -2676 7236 -2675
rect 7204 -2725 7236 -2724
rect 7204 -2755 7205 -2725
rect 7205 -2755 7235 -2725
rect 7235 -2755 7236 -2725
rect 7204 -2756 7236 -2755
rect 7204 -2836 7236 -2804
rect 7204 -2885 7236 -2884
rect 7204 -2915 7205 -2885
rect 7205 -2915 7235 -2885
rect 7235 -2915 7236 -2885
rect 7204 -2916 7236 -2915
rect 7204 -2996 7236 -2964
rect 7204 -3045 7236 -3044
rect 7204 -3075 7205 -3045
rect 7205 -3075 7235 -3045
rect 7235 -3075 7236 -3045
rect 7204 -3076 7236 -3075
rect 7204 -3156 7236 -3124
rect 7204 -3205 7236 -3204
rect 7204 -3235 7205 -3205
rect 7205 -3235 7235 -3205
rect 7235 -3235 7236 -3205
rect 7204 -3236 7236 -3235
rect 7204 -3285 7236 -3284
rect 7204 -3315 7205 -3285
rect 7205 -3315 7235 -3285
rect 7235 -3315 7236 -3285
rect 7204 -3316 7236 -3315
rect 7204 -3396 7236 -3364
rect 7204 -3476 7236 -3444
rect 7204 -3525 7236 -3524
rect 7204 -3555 7205 -3525
rect 7205 -3555 7235 -3525
rect 7235 -3555 7236 -3525
rect 7204 -3556 7236 -3555
rect 7204 -3605 7236 -3604
rect 7204 -3635 7205 -3605
rect 7205 -3635 7235 -3605
rect 7235 -3635 7236 -3605
rect 7204 -3636 7236 -3635
rect 7204 -3685 7236 -3684
rect 7204 -3715 7205 -3685
rect 7205 -3715 7235 -3685
rect 7235 -3715 7236 -3685
rect 7204 -3716 7236 -3715
rect 7284 1035 7316 1036
rect 7284 1005 7285 1035
rect 7285 1005 7315 1035
rect 7315 1005 7316 1035
rect 7284 1004 7316 1005
rect 7284 955 7316 956
rect 7284 925 7285 955
rect 7285 925 7315 955
rect 7315 925 7316 955
rect 7284 924 7316 925
rect 7284 875 7316 876
rect 7284 845 7285 875
rect 7285 845 7315 875
rect 7315 845 7316 875
rect 7284 844 7316 845
rect 7284 764 7316 796
rect 7284 684 7316 716
rect 7284 635 7316 636
rect 7284 605 7285 635
rect 7285 605 7315 635
rect 7315 605 7316 635
rect 7284 604 7316 605
rect 7284 555 7316 556
rect 7284 525 7285 555
rect 7285 525 7315 555
rect 7315 525 7316 555
rect 7284 524 7316 525
rect 7284 444 7316 476
rect 7284 395 7316 396
rect 7284 365 7285 395
rect 7285 365 7315 395
rect 7315 365 7316 395
rect 7284 364 7316 365
rect 7284 284 7316 316
rect 7284 235 7316 236
rect 7284 205 7285 235
rect 7285 205 7315 235
rect 7315 205 7316 235
rect 7284 204 7316 205
rect 7284 124 7316 156
rect 7284 75 7316 76
rect 7284 45 7285 75
rect 7285 45 7315 75
rect 7315 45 7316 75
rect 7284 44 7316 45
rect 7284 -5 7316 -4
rect 7284 -35 7285 -5
rect 7285 -35 7315 -5
rect 7315 -35 7316 -5
rect 7284 -36 7316 -35
rect 7284 -85 7316 -84
rect 7284 -115 7285 -85
rect 7285 -115 7315 -85
rect 7315 -115 7316 -85
rect 7284 -116 7316 -115
rect 7284 -165 7316 -164
rect 7284 -195 7285 -165
rect 7285 -195 7315 -165
rect 7315 -195 7316 -165
rect 7284 -196 7316 -195
rect 7284 -245 7316 -244
rect 7284 -275 7285 -245
rect 7285 -275 7315 -245
rect 7315 -275 7316 -245
rect 7284 -276 7316 -275
rect 7284 -325 7316 -324
rect 7284 -355 7285 -325
rect 7285 -355 7315 -325
rect 7315 -355 7316 -325
rect 7284 -356 7316 -355
rect 7284 -436 7316 -404
rect 7284 -485 7316 -484
rect 7284 -515 7285 -485
rect 7285 -515 7315 -485
rect 7315 -515 7316 -485
rect 7284 -516 7316 -515
rect 7284 -596 7316 -564
rect 7284 -645 7316 -644
rect 7284 -675 7285 -645
rect 7285 -675 7315 -645
rect 7315 -675 7316 -645
rect 7284 -676 7316 -675
rect 7284 -756 7316 -724
rect 7284 -805 7316 -804
rect 7284 -835 7285 -805
rect 7285 -835 7315 -805
rect 7315 -835 7316 -805
rect 7284 -836 7316 -835
rect 7284 -885 7316 -884
rect 7284 -915 7285 -885
rect 7285 -915 7315 -885
rect 7315 -915 7316 -885
rect 7284 -916 7316 -915
rect 7284 -996 7316 -964
rect 7284 -1076 7316 -1044
rect 7284 -1125 7316 -1124
rect 7284 -1155 7285 -1125
rect 7285 -1155 7315 -1125
rect 7315 -1155 7316 -1125
rect 7284 -1156 7316 -1155
rect 7284 -1205 7316 -1204
rect 7284 -1235 7285 -1205
rect 7285 -1235 7315 -1205
rect 7315 -1235 7316 -1205
rect 7284 -1236 7316 -1235
rect 7284 -1285 7316 -1284
rect 7284 -1315 7285 -1285
rect 7285 -1315 7315 -1285
rect 7315 -1315 7316 -1285
rect 7284 -1316 7316 -1315
rect 7284 -1365 7316 -1364
rect 7284 -1395 7285 -1365
rect 7285 -1395 7315 -1365
rect 7315 -1395 7316 -1365
rect 7284 -1396 7316 -1395
rect 7284 -1445 7316 -1444
rect 7284 -1475 7285 -1445
rect 7285 -1475 7315 -1445
rect 7315 -1475 7316 -1445
rect 7284 -1476 7316 -1475
rect 7284 -1525 7316 -1524
rect 7284 -1555 7285 -1525
rect 7285 -1555 7315 -1525
rect 7315 -1555 7316 -1525
rect 7284 -1556 7316 -1555
rect 7284 -1636 7316 -1604
rect 7284 -1716 7316 -1684
rect 7284 -1765 7316 -1764
rect 7284 -1795 7285 -1765
rect 7285 -1795 7315 -1765
rect 7315 -1795 7316 -1765
rect 7284 -1796 7316 -1795
rect 7284 -1845 7316 -1844
rect 7284 -1875 7285 -1845
rect 7285 -1875 7315 -1845
rect 7315 -1875 7316 -1845
rect 7284 -1876 7316 -1875
rect 7284 -1956 7316 -1924
rect 7284 -2005 7316 -2004
rect 7284 -2035 7285 -2005
rect 7285 -2035 7315 -2005
rect 7315 -2035 7316 -2005
rect 7284 -2036 7316 -2035
rect 7284 -2116 7316 -2084
rect 7284 -2165 7316 -2164
rect 7284 -2195 7285 -2165
rect 7285 -2195 7315 -2165
rect 7315 -2195 7316 -2165
rect 7284 -2196 7316 -2195
rect 7284 -2276 7316 -2244
rect 7284 -2325 7316 -2324
rect 7284 -2355 7285 -2325
rect 7285 -2355 7315 -2325
rect 7315 -2355 7316 -2325
rect 7284 -2356 7316 -2355
rect 7284 -2405 7316 -2404
rect 7284 -2435 7285 -2405
rect 7285 -2435 7315 -2405
rect 7315 -2435 7316 -2405
rect 7284 -2436 7316 -2435
rect 7284 -2485 7316 -2484
rect 7284 -2515 7285 -2485
rect 7285 -2515 7315 -2485
rect 7315 -2515 7316 -2485
rect 7284 -2516 7316 -2515
rect 7284 -2565 7316 -2564
rect 7284 -2595 7285 -2565
rect 7285 -2595 7315 -2565
rect 7315 -2595 7316 -2565
rect 7284 -2596 7316 -2595
rect 7284 -2645 7316 -2644
rect 7284 -2675 7285 -2645
rect 7285 -2675 7315 -2645
rect 7315 -2675 7316 -2645
rect 7284 -2676 7316 -2675
rect 7284 -2725 7316 -2724
rect 7284 -2755 7285 -2725
rect 7285 -2755 7315 -2725
rect 7315 -2755 7316 -2725
rect 7284 -2756 7316 -2755
rect 7284 -2836 7316 -2804
rect 7284 -2885 7316 -2884
rect 7284 -2915 7285 -2885
rect 7285 -2915 7315 -2885
rect 7315 -2915 7316 -2885
rect 7284 -2916 7316 -2915
rect 7284 -2996 7316 -2964
rect 7284 -3045 7316 -3044
rect 7284 -3075 7285 -3045
rect 7285 -3075 7315 -3045
rect 7315 -3075 7316 -3045
rect 7284 -3076 7316 -3075
rect 7284 -3156 7316 -3124
rect 7284 -3205 7316 -3204
rect 7284 -3235 7285 -3205
rect 7285 -3235 7315 -3205
rect 7315 -3235 7316 -3205
rect 7284 -3236 7316 -3235
rect 7284 -3285 7316 -3284
rect 7284 -3315 7285 -3285
rect 7285 -3315 7315 -3285
rect 7315 -3315 7316 -3285
rect 7284 -3316 7316 -3315
rect 7284 -3396 7316 -3364
rect 7284 -3476 7316 -3444
rect 7284 -3525 7316 -3524
rect 7284 -3555 7285 -3525
rect 7285 -3555 7315 -3525
rect 7315 -3555 7316 -3525
rect 7284 -3556 7316 -3555
rect 7284 -3605 7316 -3604
rect 7284 -3635 7285 -3605
rect 7285 -3635 7315 -3605
rect 7315 -3635 7316 -3605
rect 7284 -3636 7316 -3635
rect 7284 -3685 7316 -3684
rect 7284 -3715 7285 -3685
rect 7285 -3715 7315 -3685
rect 7315 -3715 7316 -3685
rect 7284 -3716 7316 -3715
rect 7364 1035 7396 1036
rect 7364 1005 7365 1035
rect 7365 1005 7395 1035
rect 7395 1005 7396 1035
rect 7364 1004 7396 1005
rect 7364 955 7396 956
rect 7364 925 7365 955
rect 7365 925 7395 955
rect 7395 925 7396 955
rect 7364 924 7396 925
rect 7364 875 7396 876
rect 7364 845 7365 875
rect 7365 845 7395 875
rect 7395 845 7396 875
rect 7364 844 7396 845
rect 7364 764 7396 796
rect 7364 684 7396 716
rect 7364 635 7396 636
rect 7364 605 7365 635
rect 7365 605 7395 635
rect 7395 605 7396 635
rect 7364 604 7396 605
rect 7364 555 7396 556
rect 7364 525 7365 555
rect 7365 525 7395 555
rect 7395 525 7396 555
rect 7364 524 7396 525
rect 7364 444 7396 476
rect 7364 395 7396 396
rect 7364 365 7365 395
rect 7365 365 7395 395
rect 7395 365 7396 395
rect 7364 364 7396 365
rect 7364 284 7396 316
rect 7364 235 7396 236
rect 7364 205 7365 235
rect 7365 205 7395 235
rect 7395 205 7396 235
rect 7364 204 7396 205
rect 7364 124 7396 156
rect 7364 75 7396 76
rect 7364 45 7365 75
rect 7365 45 7395 75
rect 7395 45 7396 75
rect 7364 44 7396 45
rect 7364 -5 7396 -4
rect 7364 -35 7365 -5
rect 7365 -35 7395 -5
rect 7395 -35 7396 -5
rect 7364 -36 7396 -35
rect 7364 -85 7396 -84
rect 7364 -115 7365 -85
rect 7365 -115 7395 -85
rect 7395 -115 7396 -85
rect 7364 -116 7396 -115
rect 7364 -165 7396 -164
rect 7364 -195 7365 -165
rect 7365 -195 7395 -165
rect 7395 -195 7396 -165
rect 7364 -196 7396 -195
rect 7364 -245 7396 -244
rect 7364 -275 7365 -245
rect 7365 -275 7395 -245
rect 7395 -275 7396 -245
rect 7364 -276 7396 -275
rect 7364 -325 7396 -324
rect 7364 -355 7365 -325
rect 7365 -355 7395 -325
rect 7395 -355 7396 -325
rect 7364 -356 7396 -355
rect 7364 -436 7396 -404
rect 7364 -485 7396 -484
rect 7364 -515 7365 -485
rect 7365 -515 7395 -485
rect 7395 -515 7396 -485
rect 7364 -516 7396 -515
rect 7364 -596 7396 -564
rect 7364 -645 7396 -644
rect 7364 -675 7365 -645
rect 7365 -675 7395 -645
rect 7395 -675 7396 -645
rect 7364 -676 7396 -675
rect 7364 -756 7396 -724
rect 7364 -805 7396 -804
rect 7364 -835 7365 -805
rect 7365 -835 7395 -805
rect 7395 -835 7396 -805
rect 7364 -836 7396 -835
rect 7364 -885 7396 -884
rect 7364 -915 7365 -885
rect 7365 -915 7395 -885
rect 7395 -915 7396 -885
rect 7364 -916 7396 -915
rect 7364 -996 7396 -964
rect 7364 -1076 7396 -1044
rect 7364 -1125 7396 -1124
rect 7364 -1155 7365 -1125
rect 7365 -1155 7395 -1125
rect 7395 -1155 7396 -1125
rect 7364 -1156 7396 -1155
rect 7364 -1205 7396 -1204
rect 7364 -1235 7365 -1205
rect 7365 -1235 7395 -1205
rect 7395 -1235 7396 -1205
rect 7364 -1236 7396 -1235
rect 7364 -1285 7396 -1284
rect 7364 -1315 7365 -1285
rect 7365 -1315 7395 -1285
rect 7395 -1315 7396 -1285
rect 7364 -1316 7396 -1315
rect 7364 -1365 7396 -1364
rect 7364 -1395 7365 -1365
rect 7365 -1395 7395 -1365
rect 7395 -1395 7396 -1365
rect 7364 -1396 7396 -1395
rect 7364 -1445 7396 -1444
rect 7364 -1475 7365 -1445
rect 7365 -1475 7395 -1445
rect 7395 -1475 7396 -1445
rect 7364 -1476 7396 -1475
rect 7364 -1525 7396 -1524
rect 7364 -1555 7365 -1525
rect 7365 -1555 7395 -1525
rect 7395 -1555 7396 -1525
rect 7364 -1556 7396 -1555
rect 7364 -1636 7396 -1604
rect 7364 -1716 7396 -1684
rect 7364 -1765 7396 -1764
rect 7364 -1795 7365 -1765
rect 7365 -1795 7395 -1765
rect 7395 -1795 7396 -1765
rect 7364 -1796 7396 -1795
rect 7364 -1845 7396 -1844
rect 7364 -1875 7365 -1845
rect 7365 -1875 7395 -1845
rect 7395 -1875 7396 -1845
rect 7364 -1876 7396 -1875
rect 7364 -1956 7396 -1924
rect 7364 -2005 7396 -2004
rect 7364 -2035 7365 -2005
rect 7365 -2035 7395 -2005
rect 7395 -2035 7396 -2005
rect 7364 -2036 7396 -2035
rect 7364 -2116 7396 -2084
rect 7364 -2165 7396 -2164
rect 7364 -2195 7365 -2165
rect 7365 -2195 7395 -2165
rect 7395 -2195 7396 -2165
rect 7364 -2196 7396 -2195
rect 7364 -2276 7396 -2244
rect 7364 -2325 7396 -2324
rect 7364 -2355 7365 -2325
rect 7365 -2355 7395 -2325
rect 7395 -2355 7396 -2325
rect 7364 -2356 7396 -2355
rect 7364 -2405 7396 -2404
rect 7364 -2435 7365 -2405
rect 7365 -2435 7395 -2405
rect 7395 -2435 7396 -2405
rect 7364 -2436 7396 -2435
rect 7364 -2485 7396 -2484
rect 7364 -2515 7365 -2485
rect 7365 -2515 7395 -2485
rect 7395 -2515 7396 -2485
rect 7364 -2516 7396 -2515
rect 7364 -2565 7396 -2564
rect 7364 -2595 7365 -2565
rect 7365 -2595 7395 -2565
rect 7395 -2595 7396 -2565
rect 7364 -2596 7396 -2595
rect 7364 -2645 7396 -2644
rect 7364 -2675 7365 -2645
rect 7365 -2675 7395 -2645
rect 7395 -2675 7396 -2645
rect 7364 -2676 7396 -2675
rect 7364 -2725 7396 -2724
rect 7364 -2755 7365 -2725
rect 7365 -2755 7395 -2725
rect 7395 -2755 7396 -2725
rect 7364 -2756 7396 -2755
rect 7364 -2836 7396 -2804
rect 7364 -2885 7396 -2884
rect 7364 -2915 7365 -2885
rect 7365 -2915 7395 -2885
rect 7395 -2915 7396 -2885
rect 7364 -2916 7396 -2915
rect 7364 -2996 7396 -2964
rect 7364 -3045 7396 -3044
rect 7364 -3075 7365 -3045
rect 7365 -3075 7395 -3045
rect 7395 -3075 7396 -3045
rect 7364 -3076 7396 -3075
rect 7364 -3156 7396 -3124
rect 7364 -3205 7396 -3204
rect 7364 -3235 7365 -3205
rect 7365 -3235 7395 -3205
rect 7395 -3235 7396 -3205
rect 7364 -3236 7396 -3235
rect 7364 -3285 7396 -3284
rect 7364 -3315 7365 -3285
rect 7365 -3315 7395 -3285
rect 7395 -3315 7396 -3285
rect 7364 -3316 7396 -3315
rect 7364 -3396 7396 -3364
rect 7364 -3476 7396 -3444
rect 7364 -3525 7396 -3524
rect 7364 -3555 7365 -3525
rect 7365 -3555 7395 -3525
rect 7395 -3555 7396 -3525
rect 7364 -3556 7396 -3555
rect 7364 -3605 7396 -3604
rect 7364 -3635 7365 -3605
rect 7365 -3635 7395 -3605
rect 7395 -3635 7396 -3605
rect 7364 -3636 7396 -3635
rect 7364 -3685 7396 -3684
rect 7364 -3715 7365 -3685
rect 7365 -3715 7395 -3685
rect 7395 -3715 7396 -3685
rect 7364 -3716 7396 -3715
rect 7444 1035 7476 1036
rect 7444 1005 7445 1035
rect 7445 1005 7475 1035
rect 7475 1005 7476 1035
rect 7444 1004 7476 1005
rect 7444 955 7476 956
rect 7444 925 7445 955
rect 7445 925 7475 955
rect 7475 925 7476 955
rect 7444 924 7476 925
rect 7444 875 7476 876
rect 7444 845 7445 875
rect 7445 845 7475 875
rect 7475 845 7476 875
rect 7444 844 7476 845
rect 7444 764 7476 796
rect 7444 684 7476 716
rect 7444 635 7476 636
rect 7444 605 7445 635
rect 7445 605 7475 635
rect 7475 605 7476 635
rect 7444 604 7476 605
rect 7444 555 7476 556
rect 7444 525 7445 555
rect 7445 525 7475 555
rect 7475 525 7476 555
rect 7444 524 7476 525
rect 7444 444 7476 476
rect 7444 395 7476 396
rect 7444 365 7445 395
rect 7445 365 7475 395
rect 7475 365 7476 395
rect 7444 364 7476 365
rect 7444 284 7476 316
rect 7444 235 7476 236
rect 7444 205 7445 235
rect 7445 205 7475 235
rect 7475 205 7476 235
rect 7444 204 7476 205
rect 7444 124 7476 156
rect 7444 75 7476 76
rect 7444 45 7445 75
rect 7445 45 7475 75
rect 7475 45 7476 75
rect 7444 44 7476 45
rect 7444 -5 7476 -4
rect 7444 -35 7445 -5
rect 7445 -35 7475 -5
rect 7475 -35 7476 -5
rect 7444 -36 7476 -35
rect 7444 -85 7476 -84
rect 7444 -115 7445 -85
rect 7445 -115 7475 -85
rect 7475 -115 7476 -85
rect 7444 -116 7476 -115
rect 7444 -165 7476 -164
rect 7444 -195 7445 -165
rect 7445 -195 7475 -165
rect 7475 -195 7476 -165
rect 7444 -196 7476 -195
rect 7444 -245 7476 -244
rect 7444 -275 7445 -245
rect 7445 -275 7475 -245
rect 7475 -275 7476 -245
rect 7444 -276 7476 -275
rect 7444 -325 7476 -324
rect 7444 -355 7445 -325
rect 7445 -355 7475 -325
rect 7475 -355 7476 -325
rect 7444 -356 7476 -355
rect 7444 -436 7476 -404
rect 7444 -485 7476 -484
rect 7444 -515 7445 -485
rect 7445 -515 7475 -485
rect 7475 -515 7476 -485
rect 7444 -516 7476 -515
rect 7444 -596 7476 -564
rect 7444 -645 7476 -644
rect 7444 -675 7445 -645
rect 7445 -675 7475 -645
rect 7475 -675 7476 -645
rect 7444 -676 7476 -675
rect 7444 -756 7476 -724
rect 7444 -805 7476 -804
rect 7444 -835 7445 -805
rect 7445 -835 7475 -805
rect 7475 -835 7476 -805
rect 7444 -836 7476 -835
rect 7444 -885 7476 -884
rect 7444 -915 7445 -885
rect 7445 -915 7475 -885
rect 7475 -915 7476 -885
rect 7444 -916 7476 -915
rect 7444 -996 7476 -964
rect 7444 -1076 7476 -1044
rect 7444 -1125 7476 -1124
rect 7444 -1155 7445 -1125
rect 7445 -1155 7475 -1125
rect 7475 -1155 7476 -1125
rect 7444 -1156 7476 -1155
rect 7444 -1205 7476 -1204
rect 7444 -1235 7445 -1205
rect 7445 -1235 7475 -1205
rect 7475 -1235 7476 -1205
rect 7444 -1236 7476 -1235
rect 7444 -1285 7476 -1284
rect 7444 -1315 7445 -1285
rect 7445 -1315 7475 -1285
rect 7475 -1315 7476 -1285
rect 7444 -1316 7476 -1315
rect 7444 -1365 7476 -1364
rect 7444 -1395 7445 -1365
rect 7445 -1395 7475 -1365
rect 7475 -1395 7476 -1365
rect 7444 -1396 7476 -1395
rect 7444 -1445 7476 -1444
rect 7444 -1475 7445 -1445
rect 7445 -1475 7475 -1445
rect 7475 -1475 7476 -1445
rect 7444 -1476 7476 -1475
rect 7444 -1525 7476 -1524
rect 7444 -1555 7445 -1525
rect 7445 -1555 7475 -1525
rect 7475 -1555 7476 -1525
rect 7444 -1556 7476 -1555
rect 7444 -1636 7476 -1604
rect 7444 -1716 7476 -1684
rect 7444 -1765 7476 -1764
rect 7444 -1795 7445 -1765
rect 7445 -1795 7475 -1765
rect 7475 -1795 7476 -1765
rect 7444 -1796 7476 -1795
rect 7444 -1845 7476 -1844
rect 7444 -1875 7445 -1845
rect 7445 -1875 7475 -1845
rect 7475 -1875 7476 -1845
rect 7444 -1876 7476 -1875
rect 7444 -1956 7476 -1924
rect 7444 -2005 7476 -2004
rect 7444 -2035 7445 -2005
rect 7445 -2035 7475 -2005
rect 7475 -2035 7476 -2005
rect 7444 -2036 7476 -2035
rect 7444 -2116 7476 -2084
rect 7444 -2165 7476 -2164
rect 7444 -2195 7445 -2165
rect 7445 -2195 7475 -2165
rect 7475 -2195 7476 -2165
rect 7444 -2196 7476 -2195
rect 7444 -2276 7476 -2244
rect 7444 -2325 7476 -2324
rect 7444 -2355 7445 -2325
rect 7445 -2355 7475 -2325
rect 7475 -2355 7476 -2325
rect 7444 -2356 7476 -2355
rect 7444 -2405 7476 -2404
rect 7444 -2435 7445 -2405
rect 7445 -2435 7475 -2405
rect 7475 -2435 7476 -2405
rect 7444 -2436 7476 -2435
rect 7444 -2485 7476 -2484
rect 7444 -2515 7445 -2485
rect 7445 -2515 7475 -2485
rect 7475 -2515 7476 -2485
rect 7444 -2516 7476 -2515
rect 7444 -2565 7476 -2564
rect 7444 -2595 7445 -2565
rect 7445 -2595 7475 -2565
rect 7475 -2595 7476 -2565
rect 7444 -2596 7476 -2595
rect 7444 -2645 7476 -2644
rect 7444 -2675 7445 -2645
rect 7445 -2675 7475 -2645
rect 7475 -2675 7476 -2645
rect 7444 -2676 7476 -2675
rect 7444 -2725 7476 -2724
rect 7444 -2755 7445 -2725
rect 7445 -2755 7475 -2725
rect 7475 -2755 7476 -2725
rect 7444 -2756 7476 -2755
rect 7444 -2836 7476 -2804
rect 7444 -2885 7476 -2884
rect 7444 -2915 7445 -2885
rect 7445 -2915 7475 -2885
rect 7475 -2915 7476 -2885
rect 7444 -2916 7476 -2915
rect 7444 -2996 7476 -2964
rect 7444 -3045 7476 -3044
rect 7444 -3075 7445 -3045
rect 7445 -3075 7475 -3045
rect 7475 -3075 7476 -3045
rect 7444 -3076 7476 -3075
rect 7444 -3156 7476 -3124
rect 7444 -3205 7476 -3204
rect 7444 -3235 7445 -3205
rect 7445 -3235 7475 -3205
rect 7475 -3235 7476 -3205
rect 7444 -3236 7476 -3235
rect 7444 -3285 7476 -3284
rect 7444 -3315 7445 -3285
rect 7445 -3315 7475 -3285
rect 7475 -3315 7476 -3285
rect 7444 -3316 7476 -3315
rect 7444 -3396 7476 -3364
rect 7444 -3476 7476 -3444
rect 7444 -3525 7476 -3524
rect 7444 -3555 7445 -3525
rect 7445 -3555 7475 -3525
rect 7475 -3555 7476 -3525
rect 7444 -3556 7476 -3555
rect 7444 -3605 7476 -3604
rect 7444 -3635 7445 -3605
rect 7445 -3635 7475 -3605
rect 7475 -3635 7476 -3605
rect 7444 -3636 7476 -3635
rect 7444 -3685 7476 -3684
rect 7444 -3715 7445 -3685
rect 7445 -3715 7475 -3685
rect 7475 -3715 7476 -3685
rect 7444 -3716 7476 -3715
rect 7524 1035 7556 1036
rect 7524 1005 7525 1035
rect 7525 1005 7555 1035
rect 7555 1005 7556 1035
rect 7524 1004 7556 1005
rect 7524 955 7556 956
rect 7524 925 7525 955
rect 7525 925 7555 955
rect 7555 925 7556 955
rect 7524 924 7556 925
rect 7524 875 7556 876
rect 7524 845 7525 875
rect 7525 845 7555 875
rect 7555 845 7556 875
rect 7524 844 7556 845
rect 7524 764 7556 796
rect 7524 684 7556 716
rect 7524 635 7556 636
rect 7524 605 7525 635
rect 7525 605 7555 635
rect 7555 605 7556 635
rect 7524 604 7556 605
rect 7524 555 7556 556
rect 7524 525 7525 555
rect 7525 525 7555 555
rect 7555 525 7556 555
rect 7524 524 7556 525
rect 7524 444 7556 476
rect 7524 395 7556 396
rect 7524 365 7525 395
rect 7525 365 7555 395
rect 7555 365 7556 395
rect 7524 364 7556 365
rect 7524 284 7556 316
rect 7524 235 7556 236
rect 7524 205 7525 235
rect 7525 205 7555 235
rect 7555 205 7556 235
rect 7524 204 7556 205
rect 7524 124 7556 156
rect 7524 75 7556 76
rect 7524 45 7525 75
rect 7525 45 7555 75
rect 7555 45 7556 75
rect 7524 44 7556 45
rect 7524 -5 7556 -4
rect 7524 -35 7525 -5
rect 7525 -35 7555 -5
rect 7555 -35 7556 -5
rect 7524 -36 7556 -35
rect 7524 -85 7556 -84
rect 7524 -115 7525 -85
rect 7525 -115 7555 -85
rect 7555 -115 7556 -85
rect 7524 -116 7556 -115
rect 7524 -165 7556 -164
rect 7524 -195 7525 -165
rect 7525 -195 7555 -165
rect 7555 -195 7556 -165
rect 7524 -196 7556 -195
rect 7524 -245 7556 -244
rect 7524 -275 7525 -245
rect 7525 -275 7555 -245
rect 7555 -275 7556 -245
rect 7524 -276 7556 -275
rect 7524 -325 7556 -324
rect 7524 -355 7525 -325
rect 7525 -355 7555 -325
rect 7555 -355 7556 -325
rect 7524 -356 7556 -355
rect 7524 -436 7556 -404
rect 7524 -485 7556 -484
rect 7524 -515 7525 -485
rect 7525 -515 7555 -485
rect 7555 -515 7556 -485
rect 7524 -516 7556 -515
rect 7524 -596 7556 -564
rect 7524 -645 7556 -644
rect 7524 -675 7525 -645
rect 7525 -675 7555 -645
rect 7555 -675 7556 -645
rect 7524 -676 7556 -675
rect 7524 -756 7556 -724
rect 7524 -805 7556 -804
rect 7524 -835 7525 -805
rect 7525 -835 7555 -805
rect 7555 -835 7556 -805
rect 7524 -836 7556 -835
rect 7524 -885 7556 -884
rect 7524 -915 7525 -885
rect 7525 -915 7555 -885
rect 7555 -915 7556 -885
rect 7524 -916 7556 -915
rect 7524 -996 7556 -964
rect 7524 -1076 7556 -1044
rect 7524 -1125 7556 -1124
rect 7524 -1155 7525 -1125
rect 7525 -1155 7555 -1125
rect 7555 -1155 7556 -1125
rect 7524 -1156 7556 -1155
rect 7524 -1205 7556 -1204
rect 7524 -1235 7525 -1205
rect 7525 -1235 7555 -1205
rect 7555 -1235 7556 -1205
rect 7524 -1236 7556 -1235
rect 7524 -1285 7556 -1284
rect 7524 -1315 7525 -1285
rect 7525 -1315 7555 -1285
rect 7555 -1315 7556 -1285
rect 7524 -1316 7556 -1315
rect 7524 -1365 7556 -1364
rect 7524 -1395 7525 -1365
rect 7525 -1395 7555 -1365
rect 7555 -1395 7556 -1365
rect 7524 -1396 7556 -1395
rect 7524 -1445 7556 -1444
rect 7524 -1475 7525 -1445
rect 7525 -1475 7555 -1445
rect 7555 -1475 7556 -1445
rect 7524 -1476 7556 -1475
rect 7524 -1525 7556 -1524
rect 7524 -1555 7525 -1525
rect 7525 -1555 7555 -1525
rect 7555 -1555 7556 -1525
rect 7524 -1556 7556 -1555
rect 7524 -1636 7556 -1604
rect 7524 -1716 7556 -1684
rect 7524 -1765 7556 -1764
rect 7524 -1795 7525 -1765
rect 7525 -1795 7555 -1765
rect 7555 -1795 7556 -1765
rect 7524 -1796 7556 -1795
rect 7524 -1845 7556 -1844
rect 7524 -1875 7525 -1845
rect 7525 -1875 7555 -1845
rect 7555 -1875 7556 -1845
rect 7524 -1876 7556 -1875
rect 7524 -1956 7556 -1924
rect 7524 -2005 7556 -2004
rect 7524 -2035 7525 -2005
rect 7525 -2035 7555 -2005
rect 7555 -2035 7556 -2005
rect 7524 -2036 7556 -2035
rect 7524 -2116 7556 -2084
rect 7524 -2165 7556 -2164
rect 7524 -2195 7525 -2165
rect 7525 -2195 7555 -2165
rect 7555 -2195 7556 -2165
rect 7524 -2196 7556 -2195
rect 7524 -2276 7556 -2244
rect 7524 -2325 7556 -2324
rect 7524 -2355 7525 -2325
rect 7525 -2355 7555 -2325
rect 7555 -2355 7556 -2325
rect 7524 -2356 7556 -2355
rect 7524 -2405 7556 -2404
rect 7524 -2435 7525 -2405
rect 7525 -2435 7555 -2405
rect 7555 -2435 7556 -2405
rect 7524 -2436 7556 -2435
rect 7524 -2485 7556 -2484
rect 7524 -2515 7525 -2485
rect 7525 -2515 7555 -2485
rect 7555 -2515 7556 -2485
rect 7524 -2516 7556 -2515
rect 7524 -2565 7556 -2564
rect 7524 -2595 7525 -2565
rect 7525 -2595 7555 -2565
rect 7555 -2595 7556 -2565
rect 7524 -2596 7556 -2595
rect 7524 -2645 7556 -2644
rect 7524 -2675 7525 -2645
rect 7525 -2675 7555 -2645
rect 7555 -2675 7556 -2645
rect 7524 -2676 7556 -2675
rect 7524 -2725 7556 -2724
rect 7524 -2755 7525 -2725
rect 7525 -2755 7555 -2725
rect 7555 -2755 7556 -2725
rect 7524 -2756 7556 -2755
rect 7524 -2836 7556 -2804
rect 7524 -2885 7556 -2884
rect 7524 -2915 7525 -2885
rect 7525 -2915 7555 -2885
rect 7555 -2915 7556 -2885
rect 7524 -2916 7556 -2915
rect 7524 -2996 7556 -2964
rect 7524 -3045 7556 -3044
rect 7524 -3075 7525 -3045
rect 7525 -3075 7555 -3045
rect 7555 -3075 7556 -3045
rect 7524 -3076 7556 -3075
rect 7524 -3156 7556 -3124
rect 7524 -3205 7556 -3204
rect 7524 -3235 7525 -3205
rect 7525 -3235 7555 -3205
rect 7555 -3235 7556 -3205
rect 7524 -3236 7556 -3235
rect 7524 -3285 7556 -3284
rect 7524 -3315 7525 -3285
rect 7525 -3315 7555 -3285
rect 7555 -3315 7556 -3285
rect 7524 -3316 7556 -3315
rect 7524 -3396 7556 -3364
rect 7524 -3476 7556 -3444
rect 7524 -3525 7556 -3524
rect 7524 -3555 7525 -3525
rect 7525 -3555 7555 -3525
rect 7555 -3555 7556 -3525
rect 7524 -3556 7556 -3555
rect 7524 -3605 7556 -3604
rect 7524 -3635 7525 -3605
rect 7525 -3635 7555 -3605
rect 7555 -3635 7556 -3605
rect 7524 -3636 7556 -3635
rect 7524 -3685 7556 -3684
rect 7524 -3715 7525 -3685
rect 7525 -3715 7555 -3685
rect 7555 -3715 7556 -3685
rect 7524 -3716 7556 -3715
rect 7604 1035 7636 1036
rect 7604 1005 7605 1035
rect 7605 1005 7635 1035
rect 7635 1005 7636 1035
rect 7604 1004 7636 1005
rect 7604 955 7636 956
rect 7604 925 7605 955
rect 7605 925 7635 955
rect 7635 925 7636 955
rect 7604 924 7636 925
rect 7604 875 7636 876
rect 7604 845 7605 875
rect 7605 845 7635 875
rect 7635 845 7636 875
rect 7604 844 7636 845
rect 7604 764 7636 796
rect 7604 684 7636 716
rect 7604 635 7636 636
rect 7604 605 7605 635
rect 7605 605 7635 635
rect 7635 605 7636 635
rect 7604 604 7636 605
rect 7604 555 7636 556
rect 7604 525 7605 555
rect 7605 525 7635 555
rect 7635 525 7636 555
rect 7604 524 7636 525
rect 7604 444 7636 476
rect 7604 395 7636 396
rect 7604 365 7605 395
rect 7605 365 7635 395
rect 7635 365 7636 395
rect 7604 364 7636 365
rect 7604 284 7636 316
rect 7604 235 7636 236
rect 7604 205 7605 235
rect 7605 205 7635 235
rect 7635 205 7636 235
rect 7604 204 7636 205
rect 7604 124 7636 156
rect 7604 75 7636 76
rect 7604 45 7605 75
rect 7605 45 7635 75
rect 7635 45 7636 75
rect 7604 44 7636 45
rect 7604 -5 7636 -4
rect 7604 -35 7605 -5
rect 7605 -35 7635 -5
rect 7635 -35 7636 -5
rect 7604 -36 7636 -35
rect 7604 -85 7636 -84
rect 7604 -115 7605 -85
rect 7605 -115 7635 -85
rect 7635 -115 7636 -85
rect 7604 -116 7636 -115
rect 7604 -165 7636 -164
rect 7604 -195 7605 -165
rect 7605 -195 7635 -165
rect 7635 -195 7636 -165
rect 7604 -196 7636 -195
rect 7604 -245 7636 -244
rect 7604 -275 7605 -245
rect 7605 -275 7635 -245
rect 7635 -275 7636 -245
rect 7604 -276 7636 -275
rect 7604 -325 7636 -324
rect 7604 -355 7605 -325
rect 7605 -355 7635 -325
rect 7635 -355 7636 -325
rect 7604 -356 7636 -355
rect 7604 -436 7636 -404
rect 7604 -485 7636 -484
rect 7604 -515 7605 -485
rect 7605 -515 7635 -485
rect 7635 -515 7636 -485
rect 7604 -516 7636 -515
rect 7604 -596 7636 -564
rect 7604 -645 7636 -644
rect 7604 -675 7605 -645
rect 7605 -675 7635 -645
rect 7635 -675 7636 -645
rect 7604 -676 7636 -675
rect 7604 -756 7636 -724
rect 7604 -805 7636 -804
rect 7604 -835 7605 -805
rect 7605 -835 7635 -805
rect 7635 -835 7636 -805
rect 7604 -836 7636 -835
rect 7604 -885 7636 -884
rect 7604 -915 7605 -885
rect 7605 -915 7635 -885
rect 7635 -915 7636 -885
rect 7604 -916 7636 -915
rect 7604 -996 7636 -964
rect 7604 -1076 7636 -1044
rect 7604 -1125 7636 -1124
rect 7604 -1155 7605 -1125
rect 7605 -1155 7635 -1125
rect 7635 -1155 7636 -1125
rect 7604 -1156 7636 -1155
rect 7604 -1205 7636 -1204
rect 7604 -1235 7605 -1205
rect 7605 -1235 7635 -1205
rect 7635 -1235 7636 -1205
rect 7604 -1236 7636 -1235
rect 7604 -1285 7636 -1284
rect 7604 -1315 7605 -1285
rect 7605 -1315 7635 -1285
rect 7635 -1315 7636 -1285
rect 7604 -1316 7636 -1315
rect 7604 -1365 7636 -1364
rect 7604 -1395 7605 -1365
rect 7605 -1395 7635 -1365
rect 7635 -1395 7636 -1365
rect 7604 -1396 7636 -1395
rect 7604 -1445 7636 -1444
rect 7604 -1475 7605 -1445
rect 7605 -1475 7635 -1445
rect 7635 -1475 7636 -1445
rect 7604 -1476 7636 -1475
rect 7604 -1525 7636 -1524
rect 7604 -1555 7605 -1525
rect 7605 -1555 7635 -1525
rect 7635 -1555 7636 -1525
rect 7604 -1556 7636 -1555
rect 7604 -1636 7636 -1604
rect 7604 -1716 7636 -1684
rect 7604 -1765 7636 -1764
rect 7604 -1795 7605 -1765
rect 7605 -1795 7635 -1765
rect 7635 -1795 7636 -1765
rect 7604 -1796 7636 -1795
rect 7604 -1845 7636 -1844
rect 7604 -1875 7605 -1845
rect 7605 -1875 7635 -1845
rect 7635 -1875 7636 -1845
rect 7604 -1876 7636 -1875
rect 7604 -1956 7636 -1924
rect 7604 -2005 7636 -2004
rect 7604 -2035 7605 -2005
rect 7605 -2035 7635 -2005
rect 7635 -2035 7636 -2005
rect 7604 -2036 7636 -2035
rect 7604 -2116 7636 -2084
rect 7604 -2165 7636 -2164
rect 7604 -2195 7605 -2165
rect 7605 -2195 7635 -2165
rect 7635 -2195 7636 -2165
rect 7604 -2196 7636 -2195
rect 7604 -2276 7636 -2244
rect 7604 -2325 7636 -2324
rect 7604 -2355 7605 -2325
rect 7605 -2355 7635 -2325
rect 7635 -2355 7636 -2325
rect 7604 -2356 7636 -2355
rect 7604 -2405 7636 -2404
rect 7604 -2435 7605 -2405
rect 7605 -2435 7635 -2405
rect 7635 -2435 7636 -2405
rect 7604 -2436 7636 -2435
rect 7604 -2485 7636 -2484
rect 7604 -2515 7605 -2485
rect 7605 -2515 7635 -2485
rect 7635 -2515 7636 -2485
rect 7604 -2516 7636 -2515
rect 7604 -2565 7636 -2564
rect 7604 -2595 7605 -2565
rect 7605 -2595 7635 -2565
rect 7635 -2595 7636 -2565
rect 7604 -2596 7636 -2595
rect 7604 -2645 7636 -2644
rect 7604 -2675 7605 -2645
rect 7605 -2675 7635 -2645
rect 7635 -2675 7636 -2645
rect 7604 -2676 7636 -2675
rect 7604 -2725 7636 -2724
rect 7604 -2755 7605 -2725
rect 7605 -2755 7635 -2725
rect 7635 -2755 7636 -2725
rect 7604 -2756 7636 -2755
rect 7604 -2836 7636 -2804
rect 7604 -2885 7636 -2884
rect 7604 -2915 7605 -2885
rect 7605 -2915 7635 -2885
rect 7635 -2915 7636 -2885
rect 7604 -2916 7636 -2915
rect 7604 -2996 7636 -2964
rect 7604 -3045 7636 -3044
rect 7604 -3075 7605 -3045
rect 7605 -3075 7635 -3045
rect 7635 -3075 7636 -3045
rect 7604 -3076 7636 -3075
rect 7604 -3156 7636 -3124
rect 7604 -3205 7636 -3204
rect 7604 -3235 7605 -3205
rect 7605 -3235 7635 -3205
rect 7635 -3235 7636 -3205
rect 7604 -3236 7636 -3235
rect 7604 -3285 7636 -3284
rect 7604 -3315 7605 -3285
rect 7605 -3315 7635 -3285
rect 7635 -3315 7636 -3285
rect 7604 -3316 7636 -3315
rect 7604 -3396 7636 -3364
rect 7604 -3476 7636 -3444
rect 7604 -3525 7636 -3524
rect 7604 -3555 7605 -3525
rect 7605 -3555 7635 -3525
rect 7635 -3555 7636 -3525
rect 7604 -3556 7636 -3555
rect 7604 -3605 7636 -3604
rect 7604 -3635 7605 -3605
rect 7605 -3635 7635 -3605
rect 7635 -3635 7636 -3605
rect 7604 -3636 7636 -3635
rect 7604 -3685 7636 -3684
rect 7604 -3715 7605 -3685
rect 7605 -3715 7635 -3685
rect 7635 -3715 7636 -3685
rect 7604 -3716 7636 -3715
rect 7684 1035 7716 1036
rect 7684 1005 7685 1035
rect 7685 1005 7715 1035
rect 7715 1005 7716 1035
rect 7684 1004 7716 1005
rect 7684 955 7716 956
rect 7684 925 7685 955
rect 7685 925 7715 955
rect 7715 925 7716 955
rect 7684 924 7716 925
rect 7684 875 7716 876
rect 7684 845 7685 875
rect 7685 845 7715 875
rect 7715 845 7716 875
rect 7684 844 7716 845
rect 7684 764 7716 796
rect 7684 684 7716 716
rect 7684 635 7716 636
rect 7684 605 7685 635
rect 7685 605 7715 635
rect 7715 605 7716 635
rect 7684 604 7716 605
rect 7684 555 7716 556
rect 7684 525 7685 555
rect 7685 525 7715 555
rect 7715 525 7716 555
rect 7684 524 7716 525
rect 7684 444 7716 476
rect 7684 395 7716 396
rect 7684 365 7685 395
rect 7685 365 7715 395
rect 7715 365 7716 395
rect 7684 364 7716 365
rect 7684 284 7716 316
rect 7684 235 7716 236
rect 7684 205 7685 235
rect 7685 205 7715 235
rect 7715 205 7716 235
rect 7684 204 7716 205
rect 7684 124 7716 156
rect 7684 75 7716 76
rect 7684 45 7685 75
rect 7685 45 7715 75
rect 7715 45 7716 75
rect 7684 44 7716 45
rect 7684 -5 7716 -4
rect 7684 -35 7685 -5
rect 7685 -35 7715 -5
rect 7715 -35 7716 -5
rect 7684 -36 7716 -35
rect 7684 -85 7716 -84
rect 7684 -115 7685 -85
rect 7685 -115 7715 -85
rect 7715 -115 7716 -85
rect 7684 -116 7716 -115
rect 7684 -165 7716 -164
rect 7684 -195 7685 -165
rect 7685 -195 7715 -165
rect 7715 -195 7716 -165
rect 7684 -196 7716 -195
rect 7684 -245 7716 -244
rect 7684 -275 7685 -245
rect 7685 -275 7715 -245
rect 7715 -275 7716 -245
rect 7684 -276 7716 -275
rect 7684 -325 7716 -324
rect 7684 -355 7685 -325
rect 7685 -355 7715 -325
rect 7715 -355 7716 -325
rect 7684 -356 7716 -355
rect 7684 -436 7716 -404
rect 7684 -485 7716 -484
rect 7684 -515 7685 -485
rect 7685 -515 7715 -485
rect 7715 -515 7716 -485
rect 7684 -516 7716 -515
rect 7684 -596 7716 -564
rect 7684 -645 7716 -644
rect 7684 -675 7685 -645
rect 7685 -675 7715 -645
rect 7715 -675 7716 -645
rect 7684 -676 7716 -675
rect 7684 -756 7716 -724
rect 7684 -805 7716 -804
rect 7684 -835 7685 -805
rect 7685 -835 7715 -805
rect 7715 -835 7716 -805
rect 7684 -836 7716 -835
rect 7684 -885 7716 -884
rect 7684 -915 7685 -885
rect 7685 -915 7715 -885
rect 7715 -915 7716 -885
rect 7684 -916 7716 -915
rect 7684 -996 7716 -964
rect 7684 -1076 7716 -1044
rect 7684 -1125 7716 -1124
rect 7684 -1155 7685 -1125
rect 7685 -1155 7715 -1125
rect 7715 -1155 7716 -1125
rect 7684 -1156 7716 -1155
rect 7684 -1205 7716 -1204
rect 7684 -1235 7685 -1205
rect 7685 -1235 7715 -1205
rect 7715 -1235 7716 -1205
rect 7684 -1236 7716 -1235
rect 7684 -1285 7716 -1284
rect 7684 -1315 7685 -1285
rect 7685 -1315 7715 -1285
rect 7715 -1315 7716 -1285
rect 7684 -1316 7716 -1315
rect 7684 -1365 7716 -1364
rect 7684 -1395 7685 -1365
rect 7685 -1395 7715 -1365
rect 7715 -1395 7716 -1365
rect 7684 -1396 7716 -1395
rect 7684 -1445 7716 -1444
rect 7684 -1475 7685 -1445
rect 7685 -1475 7715 -1445
rect 7715 -1475 7716 -1445
rect 7684 -1476 7716 -1475
rect 7684 -1525 7716 -1524
rect 7684 -1555 7685 -1525
rect 7685 -1555 7715 -1525
rect 7715 -1555 7716 -1525
rect 7684 -1556 7716 -1555
rect 7684 -1636 7716 -1604
rect 7684 -1716 7716 -1684
rect 7684 -1765 7716 -1764
rect 7684 -1795 7685 -1765
rect 7685 -1795 7715 -1765
rect 7715 -1795 7716 -1765
rect 7684 -1796 7716 -1795
rect 7684 -1845 7716 -1844
rect 7684 -1875 7685 -1845
rect 7685 -1875 7715 -1845
rect 7715 -1875 7716 -1845
rect 7684 -1876 7716 -1875
rect 7684 -1956 7716 -1924
rect 7684 -2005 7716 -2004
rect 7684 -2035 7685 -2005
rect 7685 -2035 7715 -2005
rect 7715 -2035 7716 -2005
rect 7684 -2036 7716 -2035
rect 7684 -2116 7716 -2084
rect 7684 -2165 7716 -2164
rect 7684 -2195 7685 -2165
rect 7685 -2195 7715 -2165
rect 7715 -2195 7716 -2165
rect 7684 -2196 7716 -2195
rect 7684 -2276 7716 -2244
rect 7684 -2325 7716 -2324
rect 7684 -2355 7685 -2325
rect 7685 -2355 7715 -2325
rect 7715 -2355 7716 -2325
rect 7684 -2356 7716 -2355
rect 7684 -2405 7716 -2404
rect 7684 -2435 7685 -2405
rect 7685 -2435 7715 -2405
rect 7715 -2435 7716 -2405
rect 7684 -2436 7716 -2435
rect 7684 -2485 7716 -2484
rect 7684 -2515 7685 -2485
rect 7685 -2515 7715 -2485
rect 7715 -2515 7716 -2485
rect 7684 -2516 7716 -2515
rect 7684 -2565 7716 -2564
rect 7684 -2595 7685 -2565
rect 7685 -2595 7715 -2565
rect 7715 -2595 7716 -2565
rect 7684 -2596 7716 -2595
rect 7684 -2645 7716 -2644
rect 7684 -2675 7685 -2645
rect 7685 -2675 7715 -2645
rect 7715 -2675 7716 -2645
rect 7684 -2676 7716 -2675
rect 7684 -2725 7716 -2724
rect 7684 -2755 7685 -2725
rect 7685 -2755 7715 -2725
rect 7715 -2755 7716 -2725
rect 7684 -2756 7716 -2755
rect 7684 -2836 7716 -2804
rect 7684 -2885 7716 -2884
rect 7684 -2915 7685 -2885
rect 7685 -2915 7715 -2885
rect 7715 -2915 7716 -2885
rect 7684 -2916 7716 -2915
rect 7684 -2996 7716 -2964
rect 7684 -3045 7716 -3044
rect 7684 -3075 7685 -3045
rect 7685 -3075 7715 -3045
rect 7715 -3075 7716 -3045
rect 7684 -3076 7716 -3075
rect 7684 -3156 7716 -3124
rect 7684 -3205 7716 -3204
rect 7684 -3235 7685 -3205
rect 7685 -3235 7715 -3205
rect 7715 -3235 7716 -3205
rect 7684 -3236 7716 -3235
rect 7684 -3285 7716 -3284
rect 7684 -3315 7685 -3285
rect 7685 -3315 7715 -3285
rect 7715 -3315 7716 -3285
rect 7684 -3316 7716 -3315
rect 7684 -3396 7716 -3364
rect 7684 -3476 7716 -3444
rect 7684 -3525 7716 -3524
rect 7684 -3555 7685 -3525
rect 7685 -3555 7715 -3525
rect 7715 -3555 7716 -3525
rect 7684 -3556 7716 -3555
rect 7684 -3605 7716 -3604
rect 7684 -3635 7685 -3605
rect 7685 -3635 7715 -3605
rect 7715 -3635 7716 -3605
rect 7684 -3636 7716 -3635
rect 7684 -3685 7716 -3684
rect 7684 -3715 7685 -3685
rect 7685 -3715 7715 -3685
rect 7715 -3715 7716 -3685
rect 7684 -3716 7716 -3715
rect 7764 1035 7796 1036
rect 7764 1005 7765 1035
rect 7765 1005 7795 1035
rect 7795 1005 7796 1035
rect 7764 1004 7796 1005
rect 7764 955 7796 956
rect 7764 925 7765 955
rect 7765 925 7795 955
rect 7795 925 7796 955
rect 7764 924 7796 925
rect 7764 875 7796 876
rect 7764 845 7765 875
rect 7765 845 7795 875
rect 7795 845 7796 875
rect 7764 844 7796 845
rect 7764 764 7796 796
rect 7764 684 7796 716
rect 7764 635 7796 636
rect 7764 605 7765 635
rect 7765 605 7795 635
rect 7795 605 7796 635
rect 7764 604 7796 605
rect 7764 555 7796 556
rect 7764 525 7765 555
rect 7765 525 7795 555
rect 7795 525 7796 555
rect 7764 524 7796 525
rect 7764 444 7796 476
rect 7764 395 7796 396
rect 7764 365 7765 395
rect 7765 365 7795 395
rect 7795 365 7796 395
rect 7764 364 7796 365
rect 7764 284 7796 316
rect 7764 235 7796 236
rect 7764 205 7765 235
rect 7765 205 7795 235
rect 7795 205 7796 235
rect 7764 204 7796 205
rect 7764 124 7796 156
rect 7764 75 7796 76
rect 7764 45 7765 75
rect 7765 45 7795 75
rect 7795 45 7796 75
rect 7764 44 7796 45
rect 7764 -5 7796 -4
rect 7764 -35 7765 -5
rect 7765 -35 7795 -5
rect 7795 -35 7796 -5
rect 7764 -36 7796 -35
rect 7764 -85 7796 -84
rect 7764 -115 7765 -85
rect 7765 -115 7795 -85
rect 7795 -115 7796 -85
rect 7764 -116 7796 -115
rect 7764 -165 7796 -164
rect 7764 -195 7765 -165
rect 7765 -195 7795 -165
rect 7795 -195 7796 -165
rect 7764 -196 7796 -195
rect 7764 -245 7796 -244
rect 7764 -275 7765 -245
rect 7765 -275 7795 -245
rect 7795 -275 7796 -245
rect 7764 -276 7796 -275
rect 7764 -325 7796 -324
rect 7764 -355 7765 -325
rect 7765 -355 7795 -325
rect 7795 -355 7796 -325
rect 7764 -356 7796 -355
rect 7764 -436 7796 -404
rect 7764 -485 7796 -484
rect 7764 -515 7765 -485
rect 7765 -515 7795 -485
rect 7795 -515 7796 -485
rect 7764 -516 7796 -515
rect 7764 -596 7796 -564
rect 7764 -645 7796 -644
rect 7764 -675 7765 -645
rect 7765 -675 7795 -645
rect 7795 -675 7796 -645
rect 7764 -676 7796 -675
rect 7764 -756 7796 -724
rect 7764 -805 7796 -804
rect 7764 -835 7765 -805
rect 7765 -835 7795 -805
rect 7795 -835 7796 -805
rect 7764 -836 7796 -835
rect 7764 -885 7796 -884
rect 7764 -915 7765 -885
rect 7765 -915 7795 -885
rect 7795 -915 7796 -885
rect 7764 -916 7796 -915
rect 7764 -996 7796 -964
rect 7764 -1076 7796 -1044
rect 7764 -1125 7796 -1124
rect 7764 -1155 7765 -1125
rect 7765 -1155 7795 -1125
rect 7795 -1155 7796 -1125
rect 7764 -1156 7796 -1155
rect 7764 -1205 7796 -1204
rect 7764 -1235 7765 -1205
rect 7765 -1235 7795 -1205
rect 7795 -1235 7796 -1205
rect 7764 -1236 7796 -1235
rect 7764 -1285 7796 -1284
rect 7764 -1315 7765 -1285
rect 7765 -1315 7795 -1285
rect 7795 -1315 7796 -1285
rect 7764 -1316 7796 -1315
rect 7764 -1365 7796 -1364
rect 7764 -1395 7765 -1365
rect 7765 -1395 7795 -1365
rect 7795 -1395 7796 -1365
rect 7764 -1396 7796 -1395
rect 7764 -1445 7796 -1444
rect 7764 -1475 7765 -1445
rect 7765 -1475 7795 -1445
rect 7795 -1475 7796 -1445
rect 7764 -1476 7796 -1475
rect 7764 -1525 7796 -1524
rect 7764 -1555 7765 -1525
rect 7765 -1555 7795 -1525
rect 7795 -1555 7796 -1525
rect 7764 -1556 7796 -1555
rect 7764 -1636 7796 -1604
rect 7764 -1716 7796 -1684
rect 7764 -1765 7796 -1764
rect 7764 -1795 7765 -1765
rect 7765 -1795 7795 -1765
rect 7795 -1795 7796 -1765
rect 7764 -1796 7796 -1795
rect 7764 -1845 7796 -1844
rect 7764 -1875 7765 -1845
rect 7765 -1875 7795 -1845
rect 7795 -1875 7796 -1845
rect 7764 -1876 7796 -1875
rect 7764 -1956 7796 -1924
rect 7764 -2005 7796 -2004
rect 7764 -2035 7765 -2005
rect 7765 -2035 7795 -2005
rect 7795 -2035 7796 -2005
rect 7764 -2036 7796 -2035
rect 7764 -2116 7796 -2084
rect 7764 -2165 7796 -2164
rect 7764 -2195 7765 -2165
rect 7765 -2195 7795 -2165
rect 7795 -2195 7796 -2165
rect 7764 -2196 7796 -2195
rect 7764 -2276 7796 -2244
rect 7764 -2325 7796 -2324
rect 7764 -2355 7765 -2325
rect 7765 -2355 7795 -2325
rect 7795 -2355 7796 -2325
rect 7764 -2356 7796 -2355
rect 7764 -2405 7796 -2404
rect 7764 -2435 7765 -2405
rect 7765 -2435 7795 -2405
rect 7795 -2435 7796 -2405
rect 7764 -2436 7796 -2435
rect 7764 -2485 7796 -2484
rect 7764 -2515 7765 -2485
rect 7765 -2515 7795 -2485
rect 7795 -2515 7796 -2485
rect 7764 -2516 7796 -2515
rect 7764 -2565 7796 -2564
rect 7764 -2595 7765 -2565
rect 7765 -2595 7795 -2565
rect 7795 -2595 7796 -2565
rect 7764 -2596 7796 -2595
rect 7764 -2645 7796 -2644
rect 7764 -2675 7765 -2645
rect 7765 -2675 7795 -2645
rect 7795 -2675 7796 -2645
rect 7764 -2676 7796 -2675
rect 7764 -2725 7796 -2724
rect 7764 -2755 7765 -2725
rect 7765 -2755 7795 -2725
rect 7795 -2755 7796 -2725
rect 7764 -2756 7796 -2755
rect 7764 -2836 7796 -2804
rect 7764 -2885 7796 -2884
rect 7764 -2915 7765 -2885
rect 7765 -2915 7795 -2885
rect 7795 -2915 7796 -2885
rect 7764 -2916 7796 -2915
rect 7764 -2996 7796 -2964
rect 7764 -3045 7796 -3044
rect 7764 -3075 7765 -3045
rect 7765 -3075 7795 -3045
rect 7795 -3075 7796 -3045
rect 7764 -3076 7796 -3075
rect 7764 -3156 7796 -3124
rect 7764 -3205 7796 -3204
rect 7764 -3235 7765 -3205
rect 7765 -3235 7795 -3205
rect 7795 -3235 7796 -3205
rect 7764 -3236 7796 -3235
rect 7764 -3285 7796 -3284
rect 7764 -3315 7765 -3285
rect 7765 -3315 7795 -3285
rect 7795 -3315 7796 -3285
rect 7764 -3316 7796 -3315
rect 7764 -3396 7796 -3364
rect 7764 -3476 7796 -3444
rect 7764 -3525 7796 -3524
rect 7764 -3555 7765 -3525
rect 7765 -3555 7795 -3525
rect 7795 -3555 7796 -3525
rect 7764 -3556 7796 -3555
rect 7764 -3605 7796 -3604
rect 7764 -3635 7765 -3605
rect 7765 -3635 7795 -3605
rect 7795 -3635 7796 -3605
rect 7764 -3636 7796 -3635
rect 7764 -3685 7796 -3684
rect 7764 -3715 7765 -3685
rect 7765 -3715 7795 -3685
rect 7795 -3715 7796 -3685
rect 7764 -3716 7796 -3715
rect 7844 1035 7876 1036
rect 7844 1005 7845 1035
rect 7845 1005 7875 1035
rect 7875 1005 7876 1035
rect 7844 1004 7876 1005
rect 7844 955 7876 956
rect 7844 925 7845 955
rect 7845 925 7875 955
rect 7875 925 7876 955
rect 7844 924 7876 925
rect 7844 875 7876 876
rect 7844 845 7845 875
rect 7845 845 7875 875
rect 7875 845 7876 875
rect 7844 844 7876 845
rect 7844 764 7876 796
rect 7844 684 7876 716
rect 7844 635 7876 636
rect 7844 605 7845 635
rect 7845 605 7875 635
rect 7875 605 7876 635
rect 7844 604 7876 605
rect 7844 555 7876 556
rect 7844 525 7845 555
rect 7845 525 7875 555
rect 7875 525 7876 555
rect 7844 524 7876 525
rect 7844 444 7876 476
rect 7844 395 7876 396
rect 7844 365 7845 395
rect 7845 365 7875 395
rect 7875 365 7876 395
rect 7844 364 7876 365
rect 7844 284 7876 316
rect 7844 235 7876 236
rect 7844 205 7845 235
rect 7845 205 7875 235
rect 7875 205 7876 235
rect 7844 204 7876 205
rect 7844 124 7876 156
rect 7844 75 7876 76
rect 7844 45 7845 75
rect 7845 45 7875 75
rect 7875 45 7876 75
rect 7844 44 7876 45
rect 7844 -5 7876 -4
rect 7844 -35 7845 -5
rect 7845 -35 7875 -5
rect 7875 -35 7876 -5
rect 7844 -36 7876 -35
rect 7844 -85 7876 -84
rect 7844 -115 7845 -85
rect 7845 -115 7875 -85
rect 7875 -115 7876 -85
rect 7844 -116 7876 -115
rect 7844 -165 7876 -164
rect 7844 -195 7845 -165
rect 7845 -195 7875 -165
rect 7875 -195 7876 -165
rect 7844 -196 7876 -195
rect 7844 -245 7876 -244
rect 7844 -275 7845 -245
rect 7845 -275 7875 -245
rect 7875 -275 7876 -245
rect 7844 -276 7876 -275
rect 7844 -325 7876 -324
rect 7844 -355 7845 -325
rect 7845 -355 7875 -325
rect 7875 -355 7876 -325
rect 7844 -356 7876 -355
rect 7844 -436 7876 -404
rect 7844 -485 7876 -484
rect 7844 -515 7845 -485
rect 7845 -515 7875 -485
rect 7875 -515 7876 -485
rect 7844 -516 7876 -515
rect 7844 -596 7876 -564
rect 7844 -645 7876 -644
rect 7844 -675 7845 -645
rect 7845 -675 7875 -645
rect 7875 -675 7876 -645
rect 7844 -676 7876 -675
rect 7844 -756 7876 -724
rect 7844 -805 7876 -804
rect 7844 -835 7845 -805
rect 7845 -835 7875 -805
rect 7875 -835 7876 -805
rect 7844 -836 7876 -835
rect 7844 -885 7876 -884
rect 7844 -915 7845 -885
rect 7845 -915 7875 -885
rect 7875 -915 7876 -885
rect 7844 -916 7876 -915
rect 7844 -996 7876 -964
rect 7844 -1076 7876 -1044
rect 7844 -1125 7876 -1124
rect 7844 -1155 7845 -1125
rect 7845 -1155 7875 -1125
rect 7875 -1155 7876 -1125
rect 7844 -1156 7876 -1155
rect 7844 -1205 7876 -1204
rect 7844 -1235 7845 -1205
rect 7845 -1235 7875 -1205
rect 7875 -1235 7876 -1205
rect 7844 -1236 7876 -1235
rect 7844 -1285 7876 -1284
rect 7844 -1315 7845 -1285
rect 7845 -1315 7875 -1285
rect 7875 -1315 7876 -1285
rect 7844 -1316 7876 -1315
rect 7844 -1365 7876 -1364
rect 7844 -1395 7845 -1365
rect 7845 -1395 7875 -1365
rect 7875 -1395 7876 -1365
rect 7844 -1396 7876 -1395
rect 7844 -1445 7876 -1444
rect 7844 -1475 7845 -1445
rect 7845 -1475 7875 -1445
rect 7875 -1475 7876 -1445
rect 7844 -1476 7876 -1475
rect 7844 -1525 7876 -1524
rect 7844 -1555 7845 -1525
rect 7845 -1555 7875 -1525
rect 7875 -1555 7876 -1525
rect 7844 -1556 7876 -1555
rect 7844 -1636 7876 -1604
rect 7844 -1716 7876 -1684
rect 7844 -1765 7876 -1764
rect 7844 -1795 7845 -1765
rect 7845 -1795 7875 -1765
rect 7875 -1795 7876 -1765
rect 7844 -1796 7876 -1795
rect 7844 -1845 7876 -1844
rect 7844 -1875 7845 -1845
rect 7845 -1875 7875 -1845
rect 7875 -1875 7876 -1845
rect 7844 -1876 7876 -1875
rect 7844 -1956 7876 -1924
rect 7844 -2005 7876 -2004
rect 7844 -2035 7845 -2005
rect 7845 -2035 7875 -2005
rect 7875 -2035 7876 -2005
rect 7844 -2036 7876 -2035
rect 7844 -2116 7876 -2084
rect 7844 -2165 7876 -2164
rect 7844 -2195 7845 -2165
rect 7845 -2195 7875 -2165
rect 7875 -2195 7876 -2165
rect 7844 -2196 7876 -2195
rect 7844 -2276 7876 -2244
rect 7844 -2325 7876 -2324
rect 7844 -2355 7845 -2325
rect 7845 -2355 7875 -2325
rect 7875 -2355 7876 -2325
rect 7844 -2356 7876 -2355
rect 7844 -2405 7876 -2404
rect 7844 -2435 7845 -2405
rect 7845 -2435 7875 -2405
rect 7875 -2435 7876 -2405
rect 7844 -2436 7876 -2435
rect 7844 -2485 7876 -2484
rect 7844 -2515 7845 -2485
rect 7845 -2515 7875 -2485
rect 7875 -2515 7876 -2485
rect 7844 -2516 7876 -2515
rect 7844 -2565 7876 -2564
rect 7844 -2595 7845 -2565
rect 7845 -2595 7875 -2565
rect 7875 -2595 7876 -2565
rect 7844 -2596 7876 -2595
rect 7844 -2645 7876 -2644
rect 7844 -2675 7845 -2645
rect 7845 -2675 7875 -2645
rect 7875 -2675 7876 -2645
rect 7844 -2676 7876 -2675
rect 7844 -2725 7876 -2724
rect 7844 -2755 7845 -2725
rect 7845 -2755 7875 -2725
rect 7875 -2755 7876 -2725
rect 7844 -2756 7876 -2755
rect 7844 -2836 7876 -2804
rect 7844 -2885 7876 -2884
rect 7844 -2915 7845 -2885
rect 7845 -2915 7875 -2885
rect 7875 -2915 7876 -2885
rect 7844 -2916 7876 -2915
rect 7844 -2996 7876 -2964
rect 7844 -3045 7876 -3044
rect 7844 -3075 7845 -3045
rect 7845 -3075 7875 -3045
rect 7875 -3075 7876 -3045
rect 7844 -3076 7876 -3075
rect 7844 -3156 7876 -3124
rect 7844 -3205 7876 -3204
rect 7844 -3235 7845 -3205
rect 7845 -3235 7875 -3205
rect 7875 -3235 7876 -3205
rect 7844 -3236 7876 -3235
rect 7844 -3285 7876 -3284
rect 7844 -3315 7845 -3285
rect 7845 -3315 7875 -3285
rect 7875 -3315 7876 -3285
rect 7844 -3316 7876 -3315
rect 7844 -3396 7876 -3364
rect 7844 -3476 7876 -3444
rect 7844 -3525 7876 -3524
rect 7844 -3555 7845 -3525
rect 7845 -3555 7875 -3525
rect 7875 -3555 7876 -3525
rect 7844 -3556 7876 -3555
rect 7844 -3605 7876 -3604
rect 7844 -3635 7845 -3605
rect 7845 -3635 7875 -3605
rect 7875 -3635 7876 -3605
rect 7844 -3636 7876 -3635
rect 7844 -3685 7876 -3684
rect 7844 -3715 7845 -3685
rect 7845 -3715 7875 -3685
rect 7875 -3715 7876 -3685
rect 7844 -3716 7876 -3715
rect 7924 1035 7956 1036
rect 7924 1005 7925 1035
rect 7925 1005 7955 1035
rect 7955 1005 7956 1035
rect 7924 1004 7956 1005
rect 7924 955 7956 956
rect 7924 925 7925 955
rect 7925 925 7955 955
rect 7955 925 7956 955
rect 7924 924 7956 925
rect 7924 875 7956 876
rect 7924 845 7925 875
rect 7925 845 7955 875
rect 7955 845 7956 875
rect 7924 844 7956 845
rect 7924 764 7956 796
rect 7924 684 7956 716
rect 7924 635 7956 636
rect 7924 605 7925 635
rect 7925 605 7955 635
rect 7955 605 7956 635
rect 7924 604 7956 605
rect 7924 555 7956 556
rect 7924 525 7925 555
rect 7925 525 7955 555
rect 7955 525 7956 555
rect 7924 524 7956 525
rect 7924 444 7956 476
rect 7924 395 7956 396
rect 7924 365 7925 395
rect 7925 365 7955 395
rect 7955 365 7956 395
rect 7924 364 7956 365
rect 7924 284 7956 316
rect 7924 235 7956 236
rect 7924 205 7925 235
rect 7925 205 7955 235
rect 7955 205 7956 235
rect 7924 204 7956 205
rect 7924 124 7956 156
rect 7924 75 7956 76
rect 7924 45 7925 75
rect 7925 45 7955 75
rect 7955 45 7956 75
rect 7924 44 7956 45
rect 7924 -5 7956 -4
rect 7924 -35 7925 -5
rect 7925 -35 7955 -5
rect 7955 -35 7956 -5
rect 7924 -36 7956 -35
rect 7924 -85 7956 -84
rect 7924 -115 7925 -85
rect 7925 -115 7955 -85
rect 7955 -115 7956 -85
rect 7924 -116 7956 -115
rect 7924 -165 7956 -164
rect 7924 -195 7925 -165
rect 7925 -195 7955 -165
rect 7955 -195 7956 -165
rect 7924 -196 7956 -195
rect 7924 -245 7956 -244
rect 7924 -275 7925 -245
rect 7925 -275 7955 -245
rect 7955 -275 7956 -245
rect 7924 -276 7956 -275
rect 7924 -325 7956 -324
rect 7924 -355 7925 -325
rect 7925 -355 7955 -325
rect 7955 -355 7956 -325
rect 7924 -356 7956 -355
rect 7924 -436 7956 -404
rect 7924 -485 7956 -484
rect 7924 -515 7925 -485
rect 7925 -515 7955 -485
rect 7955 -515 7956 -485
rect 7924 -516 7956 -515
rect 7924 -596 7956 -564
rect 7924 -645 7956 -644
rect 7924 -675 7925 -645
rect 7925 -675 7955 -645
rect 7955 -675 7956 -645
rect 7924 -676 7956 -675
rect 7924 -756 7956 -724
rect 7924 -805 7956 -804
rect 7924 -835 7925 -805
rect 7925 -835 7955 -805
rect 7955 -835 7956 -805
rect 7924 -836 7956 -835
rect 7924 -885 7956 -884
rect 7924 -915 7925 -885
rect 7925 -915 7955 -885
rect 7955 -915 7956 -885
rect 7924 -916 7956 -915
rect 7924 -996 7956 -964
rect 7924 -1076 7956 -1044
rect 7924 -1125 7956 -1124
rect 7924 -1155 7925 -1125
rect 7925 -1155 7955 -1125
rect 7955 -1155 7956 -1125
rect 7924 -1156 7956 -1155
rect 7924 -1205 7956 -1204
rect 7924 -1235 7925 -1205
rect 7925 -1235 7955 -1205
rect 7955 -1235 7956 -1205
rect 7924 -1236 7956 -1235
rect 7924 -1285 7956 -1284
rect 7924 -1315 7925 -1285
rect 7925 -1315 7955 -1285
rect 7955 -1315 7956 -1285
rect 7924 -1316 7956 -1315
rect 7924 -1365 7956 -1364
rect 7924 -1395 7925 -1365
rect 7925 -1395 7955 -1365
rect 7955 -1395 7956 -1365
rect 7924 -1396 7956 -1395
rect 7924 -1445 7956 -1444
rect 7924 -1475 7925 -1445
rect 7925 -1475 7955 -1445
rect 7955 -1475 7956 -1445
rect 7924 -1476 7956 -1475
rect 7924 -1525 7956 -1524
rect 7924 -1555 7925 -1525
rect 7925 -1555 7955 -1525
rect 7955 -1555 7956 -1525
rect 7924 -1556 7956 -1555
rect 7924 -1636 7956 -1604
rect 7924 -1716 7956 -1684
rect 7924 -1765 7956 -1764
rect 7924 -1795 7925 -1765
rect 7925 -1795 7955 -1765
rect 7955 -1795 7956 -1765
rect 7924 -1796 7956 -1795
rect 7924 -1845 7956 -1844
rect 7924 -1875 7925 -1845
rect 7925 -1875 7955 -1845
rect 7955 -1875 7956 -1845
rect 7924 -1876 7956 -1875
rect 7924 -1956 7956 -1924
rect 7924 -2005 7956 -2004
rect 7924 -2035 7925 -2005
rect 7925 -2035 7955 -2005
rect 7955 -2035 7956 -2005
rect 7924 -2036 7956 -2035
rect 7924 -2116 7956 -2084
rect 7924 -2165 7956 -2164
rect 7924 -2195 7925 -2165
rect 7925 -2195 7955 -2165
rect 7955 -2195 7956 -2165
rect 7924 -2196 7956 -2195
rect 7924 -2276 7956 -2244
rect 7924 -2325 7956 -2324
rect 7924 -2355 7925 -2325
rect 7925 -2355 7955 -2325
rect 7955 -2355 7956 -2325
rect 7924 -2356 7956 -2355
rect 7924 -2405 7956 -2404
rect 7924 -2435 7925 -2405
rect 7925 -2435 7955 -2405
rect 7955 -2435 7956 -2405
rect 7924 -2436 7956 -2435
rect 7924 -2485 7956 -2484
rect 7924 -2515 7925 -2485
rect 7925 -2515 7955 -2485
rect 7955 -2515 7956 -2485
rect 7924 -2516 7956 -2515
rect 7924 -2565 7956 -2564
rect 7924 -2595 7925 -2565
rect 7925 -2595 7955 -2565
rect 7955 -2595 7956 -2565
rect 7924 -2596 7956 -2595
rect 7924 -2645 7956 -2644
rect 7924 -2675 7925 -2645
rect 7925 -2675 7955 -2645
rect 7955 -2675 7956 -2645
rect 7924 -2676 7956 -2675
rect 7924 -2725 7956 -2724
rect 7924 -2755 7925 -2725
rect 7925 -2755 7955 -2725
rect 7955 -2755 7956 -2725
rect 7924 -2756 7956 -2755
rect 7924 -2836 7956 -2804
rect 7924 -2885 7956 -2884
rect 7924 -2915 7925 -2885
rect 7925 -2915 7955 -2885
rect 7955 -2915 7956 -2885
rect 7924 -2916 7956 -2915
rect 7924 -2996 7956 -2964
rect 7924 -3045 7956 -3044
rect 7924 -3075 7925 -3045
rect 7925 -3075 7955 -3045
rect 7955 -3075 7956 -3045
rect 7924 -3076 7956 -3075
rect 7924 -3156 7956 -3124
rect 7924 -3205 7956 -3204
rect 7924 -3235 7925 -3205
rect 7925 -3235 7955 -3205
rect 7955 -3235 7956 -3205
rect 7924 -3236 7956 -3235
rect 7924 -3285 7956 -3284
rect 7924 -3315 7925 -3285
rect 7925 -3315 7955 -3285
rect 7955 -3315 7956 -3285
rect 7924 -3316 7956 -3315
rect 7924 -3396 7956 -3364
rect 7924 -3476 7956 -3444
rect 7924 -3525 7956 -3524
rect 7924 -3555 7925 -3525
rect 7925 -3555 7955 -3525
rect 7955 -3555 7956 -3525
rect 7924 -3556 7956 -3555
rect 7924 -3605 7956 -3604
rect 7924 -3635 7925 -3605
rect 7925 -3635 7955 -3605
rect 7955 -3635 7956 -3605
rect 7924 -3636 7956 -3635
rect 7924 -3685 7956 -3684
rect 7924 -3715 7925 -3685
rect 7925 -3715 7955 -3685
rect 7955 -3715 7956 -3685
rect 7924 -3716 7956 -3715
rect 8004 1035 8036 1036
rect 8004 1005 8005 1035
rect 8005 1005 8035 1035
rect 8035 1005 8036 1035
rect 8004 1004 8036 1005
rect 8004 955 8036 956
rect 8004 925 8005 955
rect 8005 925 8035 955
rect 8035 925 8036 955
rect 8004 924 8036 925
rect 8004 875 8036 876
rect 8004 845 8005 875
rect 8005 845 8035 875
rect 8035 845 8036 875
rect 8004 844 8036 845
rect 8004 764 8036 796
rect 8004 684 8036 716
rect 8004 635 8036 636
rect 8004 605 8005 635
rect 8005 605 8035 635
rect 8035 605 8036 635
rect 8004 604 8036 605
rect 8004 555 8036 556
rect 8004 525 8005 555
rect 8005 525 8035 555
rect 8035 525 8036 555
rect 8004 524 8036 525
rect 8004 444 8036 476
rect 8004 395 8036 396
rect 8004 365 8005 395
rect 8005 365 8035 395
rect 8035 365 8036 395
rect 8004 364 8036 365
rect 8004 284 8036 316
rect 8004 235 8036 236
rect 8004 205 8005 235
rect 8005 205 8035 235
rect 8035 205 8036 235
rect 8004 204 8036 205
rect 8004 124 8036 156
rect 8004 75 8036 76
rect 8004 45 8005 75
rect 8005 45 8035 75
rect 8035 45 8036 75
rect 8004 44 8036 45
rect 8004 -5 8036 -4
rect 8004 -35 8005 -5
rect 8005 -35 8035 -5
rect 8035 -35 8036 -5
rect 8004 -36 8036 -35
rect 8004 -85 8036 -84
rect 8004 -115 8005 -85
rect 8005 -115 8035 -85
rect 8035 -115 8036 -85
rect 8004 -116 8036 -115
rect 8004 -165 8036 -164
rect 8004 -195 8005 -165
rect 8005 -195 8035 -165
rect 8035 -195 8036 -165
rect 8004 -196 8036 -195
rect 8004 -245 8036 -244
rect 8004 -275 8005 -245
rect 8005 -275 8035 -245
rect 8035 -275 8036 -245
rect 8004 -276 8036 -275
rect 8004 -325 8036 -324
rect 8004 -355 8005 -325
rect 8005 -355 8035 -325
rect 8035 -355 8036 -325
rect 8004 -356 8036 -355
rect 8004 -436 8036 -404
rect 8004 -485 8036 -484
rect 8004 -515 8005 -485
rect 8005 -515 8035 -485
rect 8035 -515 8036 -485
rect 8004 -516 8036 -515
rect 8004 -596 8036 -564
rect 8004 -645 8036 -644
rect 8004 -675 8005 -645
rect 8005 -675 8035 -645
rect 8035 -675 8036 -645
rect 8004 -676 8036 -675
rect 8004 -756 8036 -724
rect 8004 -805 8036 -804
rect 8004 -835 8005 -805
rect 8005 -835 8035 -805
rect 8035 -835 8036 -805
rect 8004 -836 8036 -835
rect 8004 -885 8036 -884
rect 8004 -915 8005 -885
rect 8005 -915 8035 -885
rect 8035 -915 8036 -885
rect 8004 -916 8036 -915
rect 8004 -996 8036 -964
rect 8004 -1076 8036 -1044
rect 8004 -1125 8036 -1124
rect 8004 -1155 8005 -1125
rect 8005 -1155 8035 -1125
rect 8035 -1155 8036 -1125
rect 8004 -1156 8036 -1155
rect 8004 -1205 8036 -1204
rect 8004 -1235 8005 -1205
rect 8005 -1235 8035 -1205
rect 8035 -1235 8036 -1205
rect 8004 -1236 8036 -1235
rect 8004 -1285 8036 -1284
rect 8004 -1315 8005 -1285
rect 8005 -1315 8035 -1285
rect 8035 -1315 8036 -1285
rect 8004 -1316 8036 -1315
rect 8004 -1365 8036 -1364
rect 8004 -1395 8005 -1365
rect 8005 -1395 8035 -1365
rect 8035 -1395 8036 -1365
rect 8004 -1396 8036 -1395
rect 8004 -1445 8036 -1444
rect 8004 -1475 8005 -1445
rect 8005 -1475 8035 -1445
rect 8035 -1475 8036 -1445
rect 8004 -1476 8036 -1475
rect 8004 -1525 8036 -1524
rect 8004 -1555 8005 -1525
rect 8005 -1555 8035 -1525
rect 8035 -1555 8036 -1525
rect 8004 -1556 8036 -1555
rect 8004 -1636 8036 -1604
rect 8004 -1716 8036 -1684
rect 8004 -1765 8036 -1764
rect 8004 -1795 8005 -1765
rect 8005 -1795 8035 -1765
rect 8035 -1795 8036 -1765
rect 8004 -1796 8036 -1795
rect 8004 -1845 8036 -1844
rect 8004 -1875 8005 -1845
rect 8005 -1875 8035 -1845
rect 8035 -1875 8036 -1845
rect 8004 -1876 8036 -1875
rect 8004 -1956 8036 -1924
rect 8004 -2005 8036 -2004
rect 8004 -2035 8005 -2005
rect 8005 -2035 8035 -2005
rect 8035 -2035 8036 -2005
rect 8004 -2036 8036 -2035
rect 8004 -2116 8036 -2084
rect 8004 -2165 8036 -2164
rect 8004 -2195 8005 -2165
rect 8005 -2195 8035 -2165
rect 8035 -2195 8036 -2165
rect 8004 -2196 8036 -2195
rect 8004 -2276 8036 -2244
rect 8004 -2325 8036 -2324
rect 8004 -2355 8005 -2325
rect 8005 -2355 8035 -2325
rect 8035 -2355 8036 -2325
rect 8004 -2356 8036 -2355
rect 8004 -2405 8036 -2404
rect 8004 -2435 8005 -2405
rect 8005 -2435 8035 -2405
rect 8035 -2435 8036 -2405
rect 8004 -2436 8036 -2435
rect 8004 -2485 8036 -2484
rect 8004 -2515 8005 -2485
rect 8005 -2515 8035 -2485
rect 8035 -2515 8036 -2485
rect 8004 -2516 8036 -2515
rect 8004 -2565 8036 -2564
rect 8004 -2595 8005 -2565
rect 8005 -2595 8035 -2565
rect 8035 -2595 8036 -2565
rect 8004 -2596 8036 -2595
rect 8004 -2645 8036 -2644
rect 8004 -2675 8005 -2645
rect 8005 -2675 8035 -2645
rect 8035 -2675 8036 -2645
rect 8004 -2676 8036 -2675
rect 8004 -2725 8036 -2724
rect 8004 -2755 8005 -2725
rect 8005 -2755 8035 -2725
rect 8035 -2755 8036 -2725
rect 8004 -2756 8036 -2755
rect 8004 -2836 8036 -2804
rect 8004 -2885 8036 -2884
rect 8004 -2915 8005 -2885
rect 8005 -2915 8035 -2885
rect 8035 -2915 8036 -2885
rect 8004 -2916 8036 -2915
rect 8004 -2996 8036 -2964
rect 8004 -3045 8036 -3044
rect 8004 -3075 8005 -3045
rect 8005 -3075 8035 -3045
rect 8035 -3075 8036 -3045
rect 8004 -3076 8036 -3075
rect 8004 -3156 8036 -3124
rect 8004 -3205 8036 -3204
rect 8004 -3235 8005 -3205
rect 8005 -3235 8035 -3205
rect 8035 -3235 8036 -3205
rect 8004 -3236 8036 -3235
rect 8004 -3285 8036 -3284
rect 8004 -3315 8005 -3285
rect 8005 -3315 8035 -3285
rect 8035 -3315 8036 -3285
rect 8004 -3316 8036 -3315
rect 8004 -3396 8036 -3364
rect 8004 -3476 8036 -3444
rect 8004 -3525 8036 -3524
rect 8004 -3555 8005 -3525
rect 8005 -3555 8035 -3525
rect 8035 -3555 8036 -3525
rect 8004 -3556 8036 -3555
rect 8004 -3605 8036 -3604
rect 8004 -3635 8005 -3605
rect 8005 -3635 8035 -3605
rect 8035 -3635 8036 -3605
rect 8004 -3636 8036 -3635
rect 8004 -3685 8036 -3684
rect 8004 -3715 8005 -3685
rect 8005 -3715 8035 -3685
rect 8035 -3715 8036 -3685
rect 8004 -3716 8036 -3715
rect 8084 1035 8116 1036
rect 8084 1005 8085 1035
rect 8085 1005 8115 1035
rect 8115 1005 8116 1035
rect 8084 1004 8116 1005
rect 8084 955 8116 956
rect 8084 925 8085 955
rect 8085 925 8115 955
rect 8115 925 8116 955
rect 8084 924 8116 925
rect 8084 875 8116 876
rect 8084 845 8085 875
rect 8085 845 8115 875
rect 8115 845 8116 875
rect 8084 844 8116 845
rect 8084 764 8116 796
rect 8084 684 8116 716
rect 8084 635 8116 636
rect 8084 605 8085 635
rect 8085 605 8115 635
rect 8115 605 8116 635
rect 8084 604 8116 605
rect 8084 555 8116 556
rect 8084 525 8085 555
rect 8085 525 8115 555
rect 8115 525 8116 555
rect 8084 524 8116 525
rect 8084 444 8116 476
rect 8084 395 8116 396
rect 8084 365 8085 395
rect 8085 365 8115 395
rect 8115 365 8116 395
rect 8084 364 8116 365
rect 8084 284 8116 316
rect 8084 235 8116 236
rect 8084 205 8085 235
rect 8085 205 8115 235
rect 8115 205 8116 235
rect 8084 204 8116 205
rect 8084 124 8116 156
rect 8084 75 8116 76
rect 8084 45 8085 75
rect 8085 45 8115 75
rect 8115 45 8116 75
rect 8084 44 8116 45
rect 8084 -5 8116 -4
rect 8084 -35 8085 -5
rect 8085 -35 8115 -5
rect 8115 -35 8116 -5
rect 8084 -36 8116 -35
rect 8084 -85 8116 -84
rect 8084 -115 8085 -85
rect 8085 -115 8115 -85
rect 8115 -115 8116 -85
rect 8084 -116 8116 -115
rect 8084 -165 8116 -164
rect 8084 -195 8085 -165
rect 8085 -195 8115 -165
rect 8115 -195 8116 -165
rect 8084 -196 8116 -195
rect 8084 -245 8116 -244
rect 8084 -275 8085 -245
rect 8085 -275 8115 -245
rect 8115 -275 8116 -245
rect 8084 -276 8116 -275
rect 8084 -325 8116 -324
rect 8084 -355 8085 -325
rect 8085 -355 8115 -325
rect 8115 -355 8116 -325
rect 8084 -356 8116 -355
rect 8084 -436 8116 -404
rect 8084 -485 8116 -484
rect 8084 -515 8085 -485
rect 8085 -515 8115 -485
rect 8115 -515 8116 -485
rect 8084 -516 8116 -515
rect 8084 -596 8116 -564
rect 8084 -645 8116 -644
rect 8084 -675 8085 -645
rect 8085 -675 8115 -645
rect 8115 -675 8116 -645
rect 8084 -676 8116 -675
rect 8084 -756 8116 -724
rect 8084 -805 8116 -804
rect 8084 -835 8085 -805
rect 8085 -835 8115 -805
rect 8115 -835 8116 -805
rect 8084 -836 8116 -835
rect 8084 -885 8116 -884
rect 8084 -915 8085 -885
rect 8085 -915 8115 -885
rect 8115 -915 8116 -885
rect 8084 -916 8116 -915
rect 8084 -996 8116 -964
rect 8084 -1076 8116 -1044
rect 8084 -1125 8116 -1124
rect 8084 -1155 8085 -1125
rect 8085 -1155 8115 -1125
rect 8115 -1155 8116 -1125
rect 8084 -1156 8116 -1155
rect 8084 -1205 8116 -1204
rect 8084 -1235 8085 -1205
rect 8085 -1235 8115 -1205
rect 8115 -1235 8116 -1205
rect 8084 -1236 8116 -1235
rect 8084 -1285 8116 -1284
rect 8084 -1315 8085 -1285
rect 8085 -1315 8115 -1285
rect 8115 -1315 8116 -1285
rect 8084 -1316 8116 -1315
rect 8084 -1365 8116 -1364
rect 8084 -1395 8085 -1365
rect 8085 -1395 8115 -1365
rect 8115 -1395 8116 -1365
rect 8084 -1396 8116 -1395
rect 8084 -1445 8116 -1444
rect 8084 -1475 8085 -1445
rect 8085 -1475 8115 -1445
rect 8115 -1475 8116 -1445
rect 8084 -1476 8116 -1475
rect 8084 -1525 8116 -1524
rect 8084 -1555 8085 -1525
rect 8085 -1555 8115 -1525
rect 8115 -1555 8116 -1525
rect 8084 -1556 8116 -1555
rect 8084 -1636 8116 -1604
rect 8084 -1716 8116 -1684
rect 8084 -1765 8116 -1764
rect 8084 -1795 8085 -1765
rect 8085 -1795 8115 -1765
rect 8115 -1795 8116 -1765
rect 8084 -1796 8116 -1795
rect 8084 -1845 8116 -1844
rect 8084 -1875 8085 -1845
rect 8085 -1875 8115 -1845
rect 8115 -1875 8116 -1845
rect 8084 -1876 8116 -1875
rect 8084 -1956 8116 -1924
rect 8084 -2005 8116 -2004
rect 8084 -2035 8085 -2005
rect 8085 -2035 8115 -2005
rect 8115 -2035 8116 -2005
rect 8084 -2036 8116 -2035
rect 8084 -2116 8116 -2084
rect 8084 -2165 8116 -2164
rect 8084 -2195 8085 -2165
rect 8085 -2195 8115 -2165
rect 8115 -2195 8116 -2165
rect 8084 -2196 8116 -2195
rect 8084 -2276 8116 -2244
rect 8084 -2325 8116 -2324
rect 8084 -2355 8085 -2325
rect 8085 -2355 8115 -2325
rect 8115 -2355 8116 -2325
rect 8084 -2356 8116 -2355
rect 8084 -2405 8116 -2404
rect 8084 -2435 8085 -2405
rect 8085 -2435 8115 -2405
rect 8115 -2435 8116 -2405
rect 8084 -2436 8116 -2435
rect 8084 -2485 8116 -2484
rect 8084 -2515 8085 -2485
rect 8085 -2515 8115 -2485
rect 8115 -2515 8116 -2485
rect 8084 -2516 8116 -2515
rect 8084 -2565 8116 -2564
rect 8084 -2595 8085 -2565
rect 8085 -2595 8115 -2565
rect 8115 -2595 8116 -2565
rect 8084 -2596 8116 -2595
rect 8084 -2645 8116 -2644
rect 8084 -2675 8085 -2645
rect 8085 -2675 8115 -2645
rect 8115 -2675 8116 -2645
rect 8084 -2676 8116 -2675
rect 8084 -2725 8116 -2724
rect 8084 -2755 8085 -2725
rect 8085 -2755 8115 -2725
rect 8115 -2755 8116 -2725
rect 8084 -2756 8116 -2755
rect 8084 -2836 8116 -2804
rect 8084 -2885 8116 -2884
rect 8084 -2915 8085 -2885
rect 8085 -2915 8115 -2885
rect 8115 -2915 8116 -2885
rect 8084 -2916 8116 -2915
rect 8084 -2996 8116 -2964
rect 8084 -3045 8116 -3044
rect 8084 -3075 8085 -3045
rect 8085 -3075 8115 -3045
rect 8115 -3075 8116 -3045
rect 8084 -3076 8116 -3075
rect 8084 -3156 8116 -3124
rect 8084 -3205 8116 -3204
rect 8084 -3235 8085 -3205
rect 8085 -3235 8115 -3205
rect 8115 -3235 8116 -3205
rect 8084 -3236 8116 -3235
rect 8084 -3285 8116 -3284
rect 8084 -3315 8085 -3285
rect 8085 -3315 8115 -3285
rect 8115 -3315 8116 -3285
rect 8084 -3316 8116 -3315
rect 8084 -3396 8116 -3364
rect 8084 -3476 8116 -3444
rect 8084 -3525 8116 -3524
rect 8084 -3555 8085 -3525
rect 8085 -3555 8115 -3525
rect 8115 -3555 8116 -3525
rect 8084 -3556 8116 -3555
rect 8084 -3605 8116 -3604
rect 8084 -3635 8085 -3605
rect 8085 -3635 8115 -3605
rect 8115 -3635 8116 -3605
rect 8084 -3636 8116 -3635
rect 8084 -3685 8116 -3684
rect 8084 -3715 8085 -3685
rect 8085 -3715 8115 -3685
rect 8115 -3715 8116 -3685
rect 8084 -3716 8116 -3715
rect 8164 1035 8196 1036
rect 8164 1005 8165 1035
rect 8165 1005 8195 1035
rect 8195 1005 8196 1035
rect 8164 1004 8196 1005
rect 8164 955 8196 956
rect 8164 925 8165 955
rect 8165 925 8195 955
rect 8195 925 8196 955
rect 8164 924 8196 925
rect 8164 875 8196 876
rect 8164 845 8165 875
rect 8165 845 8195 875
rect 8195 845 8196 875
rect 8164 844 8196 845
rect 8164 764 8196 796
rect 8164 684 8196 716
rect 8164 635 8196 636
rect 8164 605 8165 635
rect 8165 605 8195 635
rect 8195 605 8196 635
rect 8164 604 8196 605
rect 8164 555 8196 556
rect 8164 525 8165 555
rect 8165 525 8195 555
rect 8195 525 8196 555
rect 8164 524 8196 525
rect 8164 444 8196 476
rect 8164 395 8196 396
rect 8164 365 8165 395
rect 8165 365 8195 395
rect 8195 365 8196 395
rect 8164 364 8196 365
rect 8164 284 8196 316
rect 8164 235 8196 236
rect 8164 205 8165 235
rect 8165 205 8195 235
rect 8195 205 8196 235
rect 8164 204 8196 205
rect 8164 124 8196 156
rect 8164 75 8196 76
rect 8164 45 8165 75
rect 8165 45 8195 75
rect 8195 45 8196 75
rect 8164 44 8196 45
rect 8164 -5 8196 -4
rect 8164 -35 8165 -5
rect 8165 -35 8195 -5
rect 8195 -35 8196 -5
rect 8164 -36 8196 -35
rect 8164 -85 8196 -84
rect 8164 -115 8165 -85
rect 8165 -115 8195 -85
rect 8195 -115 8196 -85
rect 8164 -116 8196 -115
rect 8164 -165 8196 -164
rect 8164 -195 8165 -165
rect 8165 -195 8195 -165
rect 8195 -195 8196 -165
rect 8164 -196 8196 -195
rect 8164 -245 8196 -244
rect 8164 -275 8165 -245
rect 8165 -275 8195 -245
rect 8195 -275 8196 -245
rect 8164 -276 8196 -275
rect 8164 -325 8196 -324
rect 8164 -355 8165 -325
rect 8165 -355 8195 -325
rect 8195 -355 8196 -325
rect 8164 -356 8196 -355
rect 8164 -436 8196 -404
rect 8164 -485 8196 -484
rect 8164 -515 8165 -485
rect 8165 -515 8195 -485
rect 8195 -515 8196 -485
rect 8164 -516 8196 -515
rect 8164 -596 8196 -564
rect 8164 -645 8196 -644
rect 8164 -675 8165 -645
rect 8165 -675 8195 -645
rect 8195 -675 8196 -645
rect 8164 -676 8196 -675
rect 8164 -756 8196 -724
rect 8164 -805 8196 -804
rect 8164 -835 8165 -805
rect 8165 -835 8195 -805
rect 8195 -835 8196 -805
rect 8164 -836 8196 -835
rect 8164 -885 8196 -884
rect 8164 -915 8165 -885
rect 8165 -915 8195 -885
rect 8195 -915 8196 -885
rect 8164 -916 8196 -915
rect 8164 -996 8196 -964
rect 8164 -1076 8196 -1044
rect 8164 -1125 8196 -1124
rect 8164 -1155 8165 -1125
rect 8165 -1155 8195 -1125
rect 8195 -1155 8196 -1125
rect 8164 -1156 8196 -1155
rect 8164 -1205 8196 -1204
rect 8164 -1235 8165 -1205
rect 8165 -1235 8195 -1205
rect 8195 -1235 8196 -1205
rect 8164 -1236 8196 -1235
rect 8164 -1285 8196 -1284
rect 8164 -1315 8165 -1285
rect 8165 -1315 8195 -1285
rect 8195 -1315 8196 -1285
rect 8164 -1316 8196 -1315
rect 8164 -1365 8196 -1364
rect 8164 -1395 8165 -1365
rect 8165 -1395 8195 -1365
rect 8195 -1395 8196 -1365
rect 8164 -1396 8196 -1395
rect 8164 -1445 8196 -1444
rect 8164 -1475 8165 -1445
rect 8165 -1475 8195 -1445
rect 8195 -1475 8196 -1445
rect 8164 -1476 8196 -1475
rect 8164 -1525 8196 -1524
rect 8164 -1555 8165 -1525
rect 8165 -1555 8195 -1525
rect 8195 -1555 8196 -1525
rect 8164 -1556 8196 -1555
rect 8164 -1636 8196 -1604
rect 8164 -1716 8196 -1684
rect 8164 -1765 8196 -1764
rect 8164 -1795 8165 -1765
rect 8165 -1795 8195 -1765
rect 8195 -1795 8196 -1765
rect 8164 -1796 8196 -1795
rect 8164 -1845 8196 -1844
rect 8164 -1875 8165 -1845
rect 8165 -1875 8195 -1845
rect 8195 -1875 8196 -1845
rect 8164 -1876 8196 -1875
rect 8164 -1956 8196 -1924
rect 8164 -2005 8196 -2004
rect 8164 -2035 8165 -2005
rect 8165 -2035 8195 -2005
rect 8195 -2035 8196 -2005
rect 8164 -2036 8196 -2035
rect 8164 -2116 8196 -2084
rect 8164 -2165 8196 -2164
rect 8164 -2195 8165 -2165
rect 8165 -2195 8195 -2165
rect 8195 -2195 8196 -2165
rect 8164 -2196 8196 -2195
rect 8164 -2276 8196 -2244
rect 8164 -2325 8196 -2324
rect 8164 -2355 8165 -2325
rect 8165 -2355 8195 -2325
rect 8195 -2355 8196 -2325
rect 8164 -2356 8196 -2355
rect 8164 -2405 8196 -2404
rect 8164 -2435 8165 -2405
rect 8165 -2435 8195 -2405
rect 8195 -2435 8196 -2405
rect 8164 -2436 8196 -2435
rect 8164 -2485 8196 -2484
rect 8164 -2515 8165 -2485
rect 8165 -2515 8195 -2485
rect 8195 -2515 8196 -2485
rect 8164 -2516 8196 -2515
rect 8164 -2565 8196 -2564
rect 8164 -2595 8165 -2565
rect 8165 -2595 8195 -2565
rect 8195 -2595 8196 -2565
rect 8164 -2596 8196 -2595
rect 8164 -2645 8196 -2644
rect 8164 -2675 8165 -2645
rect 8165 -2675 8195 -2645
rect 8195 -2675 8196 -2645
rect 8164 -2676 8196 -2675
rect 8164 -2725 8196 -2724
rect 8164 -2755 8165 -2725
rect 8165 -2755 8195 -2725
rect 8195 -2755 8196 -2725
rect 8164 -2756 8196 -2755
rect 8164 -2836 8196 -2804
rect 8164 -2885 8196 -2884
rect 8164 -2915 8165 -2885
rect 8165 -2915 8195 -2885
rect 8195 -2915 8196 -2885
rect 8164 -2916 8196 -2915
rect 8164 -2996 8196 -2964
rect 8164 -3045 8196 -3044
rect 8164 -3075 8165 -3045
rect 8165 -3075 8195 -3045
rect 8195 -3075 8196 -3045
rect 8164 -3076 8196 -3075
rect 8164 -3156 8196 -3124
rect 8164 -3205 8196 -3204
rect 8164 -3235 8165 -3205
rect 8165 -3235 8195 -3205
rect 8195 -3235 8196 -3205
rect 8164 -3236 8196 -3235
rect 8164 -3285 8196 -3284
rect 8164 -3315 8165 -3285
rect 8165 -3315 8195 -3285
rect 8195 -3315 8196 -3285
rect 8164 -3316 8196 -3315
rect 8164 -3396 8196 -3364
rect 8164 -3476 8196 -3444
rect 8164 -3525 8196 -3524
rect 8164 -3555 8165 -3525
rect 8165 -3555 8195 -3525
rect 8195 -3555 8196 -3525
rect 8164 -3556 8196 -3555
rect 8164 -3605 8196 -3604
rect 8164 -3635 8165 -3605
rect 8165 -3635 8195 -3605
rect 8195 -3635 8196 -3605
rect 8164 -3636 8196 -3635
rect 8164 -3685 8196 -3684
rect 8164 -3715 8165 -3685
rect 8165 -3715 8195 -3685
rect 8195 -3715 8196 -3685
rect 8164 -3716 8196 -3715
rect 8244 1035 8276 1036
rect 8244 1005 8245 1035
rect 8245 1005 8275 1035
rect 8275 1005 8276 1035
rect 8244 1004 8276 1005
rect 8244 955 8276 956
rect 8244 925 8245 955
rect 8245 925 8275 955
rect 8275 925 8276 955
rect 8244 924 8276 925
rect 8244 875 8276 876
rect 8244 845 8245 875
rect 8245 845 8275 875
rect 8275 845 8276 875
rect 8244 844 8276 845
rect 8244 764 8276 796
rect 8244 684 8276 716
rect 8244 635 8276 636
rect 8244 605 8245 635
rect 8245 605 8275 635
rect 8275 605 8276 635
rect 8244 604 8276 605
rect 8244 555 8276 556
rect 8244 525 8245 555
rect 8245 525 8275 555
rect 8275 525 8276 555
rect 8244 524 8276 525
rect 8244 444 8276 476
rect 8244 395 8276 396
rect 8244 365 8245 395
rect 8245 365 8275 395
rect 8275 365 8276 395
rect 8244 364 8276 365
rect 8244 284 8276 316
rect 8244 235 8276 236
rect 8244 205 8245 235
rect 8245 205 8275 235
rect 8275 205 8276 235
rect 8244 204 8276 205
rect 8244 124 8276 156
rect 8244 75 8276 76
rect 8244 45 8245 75
rect 8245 45 8275 75
rect 8275 45 8276 75
rect 8244 44 8276 45
rect 8244 -5 8276 -4
rect 8244 -35 8245 -5
rect 8245 -35 8275 -5
rect 8275 -35 8276 -5
rect 8244 -36 8276 -35
rect 8244 -85 8276 -84
rect 8244 -115 8245 -85
rect 8245 -115 8275 -85
rect 8275 -115 8276 -85
rect 8244 -116 8276 -115
rect 8244 -165 8276 -164
rect 8244 -195 8245 -165
rect 8245 -195 8275 -165
rect 8275 -195 8276 -165
rect 8244 -196 8276 -195
rect 8244 -245 8276 -244
rect 8244 -275 8245 -245
rect 8245 -275 8275 -245
rect 8275 -275 8276 -245
rect 8244 -276 8276 -275
rect 8244 -325 8276 -324
rect 8244 -355 8245 -325
rect 8245 -355 8275 -325
rect 8275 -355 8276 -325
rect 8244 -356 8276 -355
rect 8244 -436 8276 -404
rect 8244 -485 8276 -484
rect 8244 -515 8245 -485
rect 8245 -515 8275 -485
rect 8275 -515 8276 -485
rect 8244 -516 8276 -515
rect 8244 -596 8276 -564
rect 8244 -645 8276 -644
rect 8244 -675 8245 -645
rect 8245 -675 8275 -645
rect 8275 -675 8276 -645
rect 8244 -676 8276 -675
rect 8244 -756 8276 -724
rect 8244 -805 8276 -804
rect 8244 -835 8245 -805
rect 8245 -835 8275 -805
rect 8275 -835 8276 -805
rect 8244 -836 8276 -835
rect 8244 -885 8276 -884
rect 8244 -915 8245 -885
rect 8245 -915 8275 -885
rect 8275 -915 8276 -885
rect 8244 -916 8276 -915
rect 8244 -996 8276 -964
rect 8244 -1076 8276 -1044
rect 8244 -1125 8276 -1124
rect 8244 -1155 8245 -1125
rect 8245 -1155 8275 -1125
rect 8275 -1155 8276 -1125
rect 8244 -1156 8276 -1155
rect 8244 -1205 8276 -1204
rect 8244 -1235 8245 -1205
rect 8245 -1235 8275 -1205
rect 8275 -1235 8276 -1205
rect 8244 -1236 8276 -1235
rect 8244 -1285 8276 -1284
rect 8244 -1315 8245 -1285
rect 8245 -1315 8275 -1285
rect 8275 -1315 8276 -1285
rect 8244 -1316 8276 -1315
rect 8244 -1365 8276 -1364
rect 8244 -1395 8245 -1365
rect 8245 -1395 8275 -1365
rect 8275 -1395 8276 -1365
rect 8244 -1396 8276 -1395
rect 8244 -1445 8276 -1444
rect 8244 -1475 8245 -1445
rect 8245 -1475 8275 -1445
rect 8275 -1475 8276 -1445
rect 8244 -1476 8276 -1475
rect 8244 -1525 8276 -1524
rect 8244 -1555 8245 -1525
rect 8245 -1555 8275 -1525
rect 8275 -1555 8276 -1525
rect 8244 -1556 8276 -1555
rect 8244 -1636 8276 -1604
rect 8244 -1716 8276 -1684
rect 8244 -1765 8276 -1764
rect 8244 -1795 8245 -1765
rect 8245 -1795 8275 -1765
rect 8275 -1795 8276 -1765
rect 8244 -1796 8276 -1795
rect 8244 -1845 8276 -1844
rect 8244 -1875 8245 -1845
rect 8245 -1875 8275 -1845
rect 8275 -1875 8276 -1845
rect 8244 -1876 8276 -1875
rect 8244 -1956 8276 -1924
rect 8244 -2005 8276 -2004
rect 8244 -2035 8245 -2005
rect 8245 -2035 8275 -2005
rect 8275 -2035 8276 -2005
rect 8244 -2036 8276 -2035
rect 8244 -2116 8276 -2084
rect 8244 -2165 8276 -2164
rect 8244 -2195 8245 -2165
rect 8245 -2195 8275 -2165
rect 8275 -2195 8276 -2165
rect 8244 -2196 8276 -2195
rect 8244 -2276 8276 -2244
rect 8244 -2325 8276 -2324
rect 8244 -2355 8245 -2325
rect 8245 -2355 8275 -2325
rect 8275 -2355 8276 -2325
rect 8244 -2356 8276 -2355
rect 8244 -2405 8276 -2404
rect 8244 -2435 8245 -2405
rect 8245 -2435 8275 -2405
rect 8275 -2435 8276 -2405
rect 8244 -2436 8276 -2435
rect 8244 -2485 8276 -2484
rect 8244 -2515 8245 -2485
rect 8245 -2515 8275 -2485
rect 8275 -2515 8276 -2485
rect 8244 -2516 8276 -2515
rect 8244 -2565 8276 -2564
rect 8244 -2595 8245 -2565
rect 8245 -2595 8275 -2565
rect 8275 -2595 8276 -2565
rect 8244 -2596 8276 -2595
rect 8244 -2645 8276 -2644
rect 8244 -2675 8245 -2645
rect 8245 -2675 8275 -2645
rect 8275 -2675 8276 -2645
rect 8244 -2676 8276 -2675
rect 8244 -2725 8276 -2724
rect 8244 -2755 8245 -2725
rect 8245 -2755 8275 -2725
rect 8275 -2755 8276 -2725
rect 8244 -2756 8276 -2755
rect 8244 -2836 8276 -2804
rect 8244 -2885 8276 -2884
rect 8244 -2915 8245 -2885
rect 8245 -2915 8275 -2885
rect 8275 -2915 8276 -2885
rect 8244 -2916 8276 -2915
rect 8244 -2996 8276 -2964
rect 8244 -3045 8276 -3044
rect 8244 -3075 8245 -3045
rect 8245 -3075 8275 -3045
rect 8275 -3075 8276 -3045
rect 8244 -3076 8276 -3075
rect 8244 -3156 8276 -3124
rect 8244 -3205 8276 -3204
rect 8244 -3235 8245 -3205
rect 8245 -3235 8275 -3205
rect 8275 -3235 8276 -3205
rect 8244 -3236 8276 -3235
rect 8244 -3285 8276 -3284
rect 8244 -3315 8245 -3285
rect 8245 -3315 8275 -3285
rect 8275 -3315 8276 -3285
rect 8244 -3316 8276 -3315
rect 8244 -3396 8276 -3364
rect 8244 -3476 8276 -3444
rect 8244 -3525 8276 -3524
rect 8244 -3555 8245 -3525
rect 8245 -3555 8275 -3525
rect 8275 -3555 8276 -3525
rect 8244 -3556 8276 -3555
rect 8244 -3605 8276 -3604
rect 8244 -3635 8245 -3605
rect 8245 -3635 8275 -3605
rect 8275 -3635 8276 -3605
rect 8244 -3636 8276 -3635
rect 8244 -3685 8276 -3684
rect 8244 -3715 8245 -3685
rect 8245 -3715 8275 -3685
rect 8275 -3715 8276 -3685
rect 8244 -3716 8276 -3715
rect 8324 1035 8356 1036
rect 8324 1005 8325 1035
rect 8325 1005 8355 1035
rect 8355 1005 8356 1035
rect 8324 1004 8356 1005
rect 8324 955 8356 956
rect 8324 925 8325 955
rect 8325 925 8355 955
rect 8355 925 8356 955
rect 8324 924 8356 925
rect 8324 875 8356 876
rect 8324 845 8325 875
rect 8325 845 8355 875
rect 8355 845 8356 875
rect 8324 844 8356 845
rect 8324 764 8356 796
rect 8324 684 8356 716
rect 8324 635 8356 636
rect 8324 605 8325 635
rect 8325 605 8355 635
rect 8355 605 8356 635
rect 8324 604 8356 605
rect 8324 555 8356 556
rect 8324 525 8325 555
rect 8325 525 8355 555
rect 8355 525 8356 555
rect 8324 524 8356 525
rect 8324 444 8356 476
rect 8324 395 8356 396
rect 8324 365 8325 395
rect 8325 365 8355 395
rect 8355 365 8356 395
rect 8324 364 8356 365
rect 8324 284 8356 316
rect 8324 235 8356 236
rect 8324 205 8325 235
rect 8325 205 8355 235
rect 8355 205 8356 235
rect 8324 204 8356 205
rect 8324 124 8356 156
rect 8324 75 8356 76
rect 8324 45 8325 75
rect 8325 45 8355 75
rect 8355 45 8356 75
rect 8324 44 8356 45
rect 8324 -5 8356 -4
rect 8324 -35 8325 -5
rect 8325 -35 8355 -5
rect 8355 -35 8356 -5
rect 8324 -36 8356 -35
rect 8324 -85 8356 -84
rect 8324 -115 8325 -85
rect 8325 -115 8355 -85
rect 8355 -115 8356 -85
rect 8324 -116 8356 -115
rect 8324 -165 8356 -164
rect 8324 -195 8325 -165
rect 8325 -195 8355 -165
rect 8355 -195 8356 -165
rect 8324 -196 8356 -195
rect 8324 -245 8356 -244
rect 8324 -275 8325 -245
rect 8325 -275 8355 -245
rect 8355 -275 8356 -245
rect 8324 -276 8356 -275
rect 8324 -325 8356 -324
rect 8324 -355 8325 -325
rect 8325 -355 8355 -325
rect 8355 -355 8356 -325
rect 8324 -356 8356 -355
rect 8324 -436 8356 -404
rect 8324 -485 8356 -484
rect 8324 -515 8325 -485
rect 8325 -515 8355 -485
rect 8355 -515 8356 -485
rect 8324 -516 8356 -515
rect 8324 -596 8356 -564
rect 8324 -645 8356 -644
rect 8324 -675 8325 -645
rect 8325 -675 8355 -645
rect 8355 -675 8356 -645
rect 8324 -676 8356 -675
rect 8324 -756 8356 -724
rect 8324 -805 8356 -804
rect 8324 -835 8325 -805
rect 8325 -835 8355 -805
rect 8355 -835 8356 -805
rect 8324 -836 8356 -835
rect 8324 -885 8356 -884
rect 8324 -915 8325 -885
rect 8325 -915 8355 -885
rect 8355 -915 8356 -885
rect 8324 -916 8356 -915
rect 8324 -996 8356 -964
rect 8324 -1076 8356 -1044
rect 8324 -1125 8356 -1124
rect 8324 -1155 8325 -1125
rect 8325 -1155 8355 -1125
rect 8355 -1155 8356 -1125
rect 8324 -1156 8356 -1155
rect 8324 -1205 8356 -1204
rect 8324 -1235 8325 -1205
rect 8325 -1235 8355 -1205
rect 8355 -1235 8356 -1205
rect 8324 -1236 8356 -1235
rect 8324 -1285 8356 -1284
rect 8324 -1315 8325 -1285
rect 8325 -1315 8355 -1285
rect 8355 -1315 8356 -1285
rect 8324 -1316 8356 -1315
rect 8324 -1365 8356 -1364
rect 8324 -1395 8325 -1365
rect 8325 -1395 8355 -1365
rect 8355 -1395 8356 -1365
rect 8324 -1396 8356 -1395
rect 8324 -1445 8356 -1444
rect 8324 -1475 8325 -1445
rect 8325 -1475 8355 -1445
rect 8355 -1475 8356 -1445
rect 8324 -1476 8356 -1475
rect 8324 -1525 8356 -1524
rect 8324 -1555 8325 -1525
rect 8325 -1555 8355 -1525
rect 8355 -1555 8356 -1525
rect 8324 -1556 8356 -1555
rect 8324 -1636 8356 -1604
rect 8324 -1716 8356 -1684
rect 8324 -1765 8356 -1764
rect 8324 -1795 8325 -1765
rect 8325 -1795 8355 -1765
rect 8355 -1795 8356 -1765
rect 8324 -1796 8356 -1795
rect 8324 -1845 8356 -1844
rect 8324 -1875 8325 -1845
rect 8325 -1875 8355 -1845
rect 8355 -1875 8356 -1845
rect 8324 -1876 8356 -1875
rect 8324 -1956 8356 -1924
rect 8324 -2005 8356 -2004
rect 8324 -2035 8325 -2005
rect 8325 -2035 8355 -2005
rect 8355 -2035 8356 -2005
rect 8324 -2036 8356 -2035
rect 8324 -2116 8356 -2084
rect 8324 -2165 8356 -2164
rect 8324 -2195 8325 -2165
rect 8325 -2195 8355 -2165
rect 8355 -2195 8356 -2165
rect 8324 -2196 8356 -2195
rect 8324 -2276 8356 -2244
rect 8324 -2325 8356 -2324
rect 8324 -2355 8325 -2325
rect 8325 -2355 8355 -2325
rect 8355 -2355 8356 -2325
rect 8324 -2356 8356 -2355
rect 8324 -2405 8356 -2404
rect 8324 -2435 8325 -2405
rect 8325 -2435 8355 -2405
rect 8355 -2435 8356 -2405
rect 8324 -2436 8356 -2435
rect 8324 -2485 8356 -2484
rect 8324 -2515 8325 -2485
rect 8325 -2515 8355 -2485
rect 8355 -2515 8356 -2485
rect 8324 -2516 8356 -2515
rect 8324 -2565 8356 -2564
rect 8324 -2595 8325 -2565
rect 8325 -2595 8355 -2565
rect 8355 -2595 8356 -2565
rect 8324 -2596 8356 -2595
rect 8324 -2645 8356 -2644
rect 8324 -2675 8325 -2645
rect 8325 -2675 8355 -2645
rect 8355 -2675 8356 -2645
rect 8324 -2676 8356 -2675
rect 8324 -2725 8356 -2724
rect 8324 -2755 8325 -2725
rect 8325 -2755 8355 -2725
rect 8355 -2755 8356 -2725
rect 8324 -2756 8356 -2755
rect 8324 -2836 8356 -2804
rect 8324 -2885 8356 -2884
rect 8324 -2915 8325 -2885
rect 8325 -2915 8355 -2885
rect 8355 -2915 8356 -2885
rect 8324 -2916 8356 -2915
rect 8324 -2996 8356 -2964
rect 8324 -3045 8356 -3044
rect 8324 -3075 8325 -3045
rect 8325 -3075 8355 -3045
rect 8355 -3075 8356 -3045
rect 8324 -3076 8356 -3075
rect 8324 -3156 8356 -3124
rect 8324 -3205 8356 -3204
rect 8324 -3235 8325 -3205
rect 8325 -3235 8355 -3205
rect 8355 -3235 8356 -3205
rect 8324 -3236 8356 -3235
rect 8324 -3285 8356 -3284
rect 8324 -3315 8325 -3285
rect 8325 -3315 8355 -3285
rect 8355 -3315 8356 -3285
rect 8324 -3316 8356 -3315
rect 8324 -3396 8356 -3364
rect 8324 -3476 8356 -3444
rect 8324 -3525 8356 -3524
rect 8324 -3555 8325 -3525
rect 8325 -3555 8355 -3525
rect 8355 -3555 8356 -3525
rect 8324 -3556 8356 -3555
rect 8324 -3605 8356 -3604
rect 8324 -3635 8325 -3605
rect 8325 -3635 8355 -3605
rect 8355 -3635 8356 -3605
rect 8324 -3636 8356 -3635
rect 8324 -3685 8356 -3684
rect 8324 -3715 8325 -3685
rect 8325 -3715 8355 -3685
rect 8355 -3715 8356 -3685
rect 8324 -3716 8356 -3715
rect 8404 1035 8436 1036
rect 8404 1005 8405 1035
rect 8405 1005 8435 1035
rect 8435 1005 8436 1035
rect 8404 1004 8436 1005
rect 8404 955 8436 956
rect 8404 925 8405 955
rect 8405 925 8435 955
rect 8435 925 8436 955
rect 8404 924 8436 925
rect 8404 875 8436 876
rect 8404 845 8405 875
rect 8405 845 8435 875
rect 8435 845 8436 875
rect 8404 844 8436 845
rect 8404 764 8436 796
rect 8404 684 8436 716
rect 8404 635 8436 636
rect 8404 605 8405 635
rect 8405 605 8435 635
rect 8435 605 8436 635
rect 8404 604 8436 605
rect 8404 555 8436 556
rect 8404 525 8405 555
rect 8405 525 8435 555
rect 8435 525 8436 555
rect 8404 524 8436 525
rect 8404 444 8436 476
rect 8404 395 8436 396
rect 8404 365 8405 395
rect 8405 365 8435 395
rect 8435 365 8436 395
rect 8404 364 8436 365
rect 8404 284 8436 316
rect 8404 235 8436 236
rect 8404 205 8405 235
rect 8405 205 8435 235
rect 8435 205 8436 235
rect 8404 204 8436 205
rect 8404 124 8436 156
rect 8404 75 8436 76
rect 8404 45 8405 75
rect 8405 45 8435 75
rect 8435 45 8436 75
rect 8404 44 8436 45
rect 8404 -5 8436 -4
rect 8404 -35 8405 -5
rect 8405 -35 8435 -5
rect 8435 -35 8436 -5
rect 8404 -36 8436 -35
rect 8404 -85 8436 -84
rect 8404 -115 8405 -85
rect 8405 -115 8435 -85
rect 8435 -115 8436 -85
rect 8404 -116 8436 -115
rect 8404 -165 8436 -164
rect 8404 -195 8405 -165
rect 8405 -195 8435 -165
rect 8435 -195 8436 -165
rect 8404 -196 8436 -195
rect 8404 -245 8436 -244
rect 8404 -275 8405 -245
rect 8405 -275 8435 -245
rect 8435 -275 8436 -245
rect 8404 -276 8436 -275
rect 8404 -325 8436 -324
rect 8404 -355 8405 -325
rect 8405 -355 8435 -325
rect 8435 -355 8436 -325
rect 8404 -356 8436 -355
rect 8404 -436 8436 -404
rect 8404 -485 8436 -484
rect 8404 -515 8405 -485
rect 8405 -515 8435 -485
rect 8435 -515 8436 -485
rect 8404 -516 8436 -515
rect 8404 -596 8436 -564
rect 8404 -645 8436 -644
rect 8404 -675 8405 -645
rect 8405 -675 8435 -645
rect 8435 -675 8436 -645
rect 8404 -676 8436 -675
rect 8404 -756 8436 -724
rect 8404 -805 8436 -804
rect 8404 -835 8405 -805
rect 8405 -835 8435 -805
rect 8435 -835 8436 -805
rect 8404 -836 8436 -835
rect 8404 -885 8436 -884
rect 8404 -915 8405 -885
rect 8405 -915 8435 -885
rect 8435 -915 8436 -885
rect 8404 -916 8436 -915
rect 8404 -996 8436 -964
rect 8404 -1076 8436 -1044
rect 8404 -1125 8436 -1124
rect 8404 -1155 8405 -1125
rect 8405 -1155 8435 -1125
rect 8435 -1155 8436 -1125
rect 8404 -1156 8436 -1155
rect 8404 -1205 8436 -1204
rect 8404 -1235 8405 -1205
rect 8405 -1235 8435 -1205
rect 8435 -1235 8436 -1205
rect 8404 -1236 8436 -1235
rect 8404 -1285 8436 -1284
rect 8404 -1315 8405 -1285
rect 8405 -1315 8435 -1285
rect 8435 -1315 8436 -1285
rect 8404 -1316 8436 -1315
rect 8404 -1365 8436 -1364
rect 8404 -1395 8405 -1365
rect 8405 -1395 8435 -1365
rect 8435 -1395 8436 -1365
rect 8404 -1396 8436 -1395
rect 8404 -1445 8436 -1444
rect 8404 -1475 8405 -1445
rect 8405 -1475 8435 -1445
rect 8435 -1475 8436 -1445
rect 8404 -1476 8436 -1475
rect 8404 -1525 8436 -1524
rect 8404 -1555 8405 -1525
rect 8405 -1555 8435 -1525
rect 8435 -1555 8436 -1525
rect 8404 -1556 8436 -1555
rect 8404 -1636 8436 -1604
rect 8404 -1716 8436 -1684
rect 8404 -1765 8436 -1764
rect 8404 -1795 8405 -1765
rect 8405 -1795 8435 -1765
rect 8435 -1795 8436 -1765
rect 8404 -1796 8436 -1795
rect 8404 -1845 8436 -1844
rect 8404 -1875 8405 -1845
rect 8405 -1875 8435 -1845
rect 8435 -1875 8436 -1845
rect 8404 -1876 8436 -1875
rect 8404 -1956 8436 -1924
rect 8404 -2005 8436 -2004
rect 8404 -2035 8405 -2005
rect 8405 -2035 8435 -2005
rect 8435 -2035 8436 -2005
rect 8404 -2036 8436 -2035
rect 8404 -2116 8436 -2084
rect 8404 -2165 8436 -2164
rect 8404 -2195 8405 -2165
rect 8405 -2195 8435 -2165
rect 8435 -2195 8436 -2165
rect 8404 -2196 8436 -2195
rect 8404 -2276 8436 -2244
rect 8404 -2325 8436 -2324
rect 8404 -2355 8405 -2325
rect 8405 -2355 8435 -2325
rect 8435 -2355 8436 -2325
rect 8404 -2356 8436 -2355
rect 8404 -2405 8436 -2404
rect 8404 -2435 8405 -2405
rect 8405 -2435 8435 -2405
rect 8435 -2435 8436 -2405
rect 8404 -2436 8436 -2435
rect 8404 -2485 8436 -2484
rect 8404 -2515 8405 -2485
rect 8405 -2515 8435 -2485
rect 8435 -2515 8436 -2485
rect 8404 -2516 8436 -2515
rect 8404 -2565 8436 -2564
rect 8404 -2595 8405 -2565
rect 8405 -2595 8435 -2565
rect 8435 -2595 8436 -2565
rect 8404 -2596 8436 -2595
rect 8404 -2645 8436 -2644
rect 8404 -2675 8405 -2645
rect 8405 -2675 8435 -2645
rect 8435 -2675 8436 -2645
rect 8404 -2676 8436 -2675
rect 8404 -2725 8436 -2724
rect 8404 -2755 8405 -2725
rect 8405 -2755 8435 -2725
rect 8435 -2755 8436 -2725
rect 8404 -2756 8436 -2755
rect 8404 -2836 8436 -2804
rect 8404 -2885 8436 -2884
rect 8404 -2915 8405 -2885
rect 8405 -2915 8435 -2885
rect 8435 -2915 8436 -2885
rect 8404 -2916 8436 -2915
rect 8404 -2996 8436 -2964
rect 8404 -3045 8436 -3044
rect 8404 -3075 8405 -3045
rect 8405 -3075 8435 -3045
rect 8435 -3075 8436 -3045
rect 8404 -3076 8436 -3075
rect 8404 -3156 8436 -3124
rect 8404 -3205 8436 -3204
rect 8404 -3235 8405 -3205
rect 8405 -3235 8435 -3205
rect 8435 -3235 8436 -3205
rect 8404 -3236 8436 -3235
rect 8404 -3285 8436 -3284
rect 8404 -3315 8405 -3285
rect 8405 -3315 8435 -3285
rect 8435 -3315 8436 -3285
rect 8404 -3316 8436 -3315
rect 8404 -3396 8436 -3364
rect 8404 -3476 8436 -3444
rect 8404 -3525 8436 -3524
rect 8404 -3555 8405 -3525
rect 8405 -3555 8435 -3525
rect 8435 -3555 8436 -3525
rect 8404 -3556 8436 -3555
rect 8404 -3605 8436 -3604
rect 8404 -3635 8405 -3605
rect 8405 -3635 8435 -3605
rect 8435 -3635 8436 -3605
rect 8404 -3636 8436 -3635
rect 8404 -3685 8436 -3684
rect 8404 -3715 8405 -3685
rect 8405 -3715 8435 -3685
rect 8435 -3715 8436 -3685
rect 8404 -3716 8436 -3715
rect 8484 1035 8516 1036
rect 8484 1005 8485 1035
rect 8485 1005 8515 1035
rect 8515 1005 8516 1035
rect 8484 1004 8516 1005
rect 8484 955 8516 956
rect 8484 925 8485 955
rect 8485 925 8515 955
rect 8515 925 8516 955
rect 8484 924 8516 925
rect 8484 875 8516 876
rect 8484 845 8485 875
rect 8485 845 8515 875
rect 8515 845 8516 875
rect 8484 844 8516 845
rect 8484 764 8516 796
rect 8484 684 8516 716
rect 8484 635 8516 636
rect 8484 605 8485 635
rect 8485 605 8515 635
rect 8515 605 8516 635
rect 8484 604 8516 605
rect 8484 555 8516 556
rect 8484 525 8485 555
rect 8485 525 8515 555
rect 8515 525 8516 555
rect 8484 524 8516 525
rect 8484 444 8516 476
rect 8484 395 8516 396
rect 8484 365 8485 395
rect 8485 365 8515 395
rect 8515 365 8516 395
rect 8484 364 8516 365
rect 8484 284 8516 316
rect 8484 235 8516 236
rect 8484 205 8485 235
rect 8485 205 8515 235
rect 8515 205 8516 235
rect 8484 204 8516 205
rect 8484 124 8516 156
rect 8484 75 8516 76
rect 8484 45 8485 75
rect 8485 45 8515 75
rect 8515 45 8516 75
rect 8484 44 8516 45
rect 8484 -5 8516 -4
rect 8484 -35 8485 -5
rect 8485 -35 8515 -5
rect 8515 -35 8516 -5
rect 8484 -36 8516 -35
rect 8484 -85 8516 -84
rect 8484 -115 8485 -85
rect 8485 -115 8515 -85
rect 8515 -115 8516 -85
rect 8484 -116 8516 -115
rect 8484 -165 8516 -164
rect 8484 -195 8485 -165
rect 8485 -195 8515 -165
rect 8515 -195 8516 -165
rect 8484 -196 8516 -195
rect 8484 -245 8516 -244
rect 8484 -275 8485 -245
rect 8485 -275 8515 -245
rect 8515 -275 8516 -245
rect 8484 -276 8516 -275
rect 8484 -325 8516 -324
rect 8484 -355 8485 -325
rect 8485 -355 8515 -325
rect 8515 -355 8516 -325
rect 8484 -356 8516 -355
rect 8484 -436 8516 -404
rect 8484 -485 8516 -484
rect 8484 -515 8485 -485
rect 8485 -515 8515 -485
rect 8515 -515 8516 -485
rect 8484 -516 8516 -515
rect 8484 -596 8516 -564
rect 8484 -645 8516 -644
rect 8484 -675 8485 -645
rect 8485 -675 8515 -645
rect 8515 -675 8516 -645
rect 8484 -676 8516 -675
rect 8484 -756 8516 -724
rect 8484 -805 8516 -804
rect 8484 -835 8485 -805
rect 8485 -835 8515 -805
rect 8515 -835 8516 -805
rect 8484 -836 8516 -835
rect 8484 -885 8516 -884
rect 8484 -915 8485 -885
rect 8485 -915 8515 -885
rect 8515 -915 8516 -885
rect 8484 -916 8516 -915
rect 8484 -996 8516 -964
rect 8484 -1076 8516 -1044
rect 8484 -1125 8516 -1124
rect 8484 -1155 8485 -1125
rect 8485 -1155 8515 -1125
rect 8515 -1155 8516 -1125
rect 8484 -1156 8516 -1155
rect 8484 -1205 8516 -1204
rect 8484 -1235 8485 -1205
rect 8485 -1235 8515 -1205
rect 8515 -1235 8516 -1205
rect 8484 -1236 8516 -1235
rect 8484 -1285 8516 -1284
rect 8484 -1315 8485 -1285
rect 8485 -1315 8515 -1285
rect 8515 -1315 8516 -1285
rect 8484 -1316 8516 -1315
rect 8484 -1365 8516 -1364
rect 8484 -1395 8485 -1365
rect 8485 -1395 8515 -1365
rect 8515 -1395 8516 -1365
rect 8484 -1396 8516 -1395
rect 8484 -1445 8516 -1444
rect 8484 -1475 8485 -1445
rect 8485 -1475 8515 -1445
rect 8515 -1475 8516 -1445
rect 8484 -1476 8516 -1475
rect 8484 -1525 8516 -1524
rect 8484 -1555 8485 -1525
rect 8485 -1555 8515 -1525
rect 8515 -1555 8516 -1525
rect 8484 -1556 8516 -1555
rect 8484 -1636 8516 -1604
rect 8484 -1716 8516 -1684
rect 8484 -1765 8516 -1764
rect 8484 -1795 8485 -1765
rect 8485 -1795 8515 -1765
rect 8515 -1795 8516 -1765
rect 8484 -1796 8516 -1795
rect 8484 -1845 8516 -1844
rect 8484 -1875 8485 -1845
rect 8485 -1875 8515 -1845
rect 8515 -1875 8516 -1845
rect 8484 -1876 8516 -1875
rect 8484 -1956 8516 -1924
rect 8484 -2005 8516 -2004
rect 8484 -2035 8485 -2005
rect 8485 -2035 8515 -2005
rect 8515 -2035 8516 -2005
rect 8484 -2036 8516 -2035
rect 8484 -2116 8516 -2084
rect 8484 -2165 8516 -2164
rect 8484 -2195 8485 -2165
rect 8485 -2195 8515 -2165
rect 8515 -2195 8516 -2165
rect 8484 -2196 8516 -2195
rect 8484 -2276 8516 -2244
rect 8484 -2325 8516 -2324
rect 8484 -2355 8485 -2325
rect 8485 -2355 8515 -2325
rect 8515 -2355 8516 -2325
rect 8484 -2356 8516 -2355
rect 8484 -2405 8516 -2404
rect 8484 -2435 8485 -2405
rect 8485 -2435 8515 -2405
rect 8515 -2435 8516 -2405
rect 8484 -2436 8516 -2435
rect 8484 -2485 8516 -2484
rect 8484 -2515 8485 -2485
rect 8485 -2515 8515 -2485
rect 8515 -2515 8516 -2485
rect 8484 -2516 8516 -2515
rect 8484 -2565 8516 -2564
rect 8484 -2595 8485 -2565
rect 8485 -2595 8515 -2565
rect 8515 -2595 8516 -2565
rect 8484 -2596 8516 -2595
rect 8484 -2645 8516 -2644
rect 8484 -2675 8485 -2645
rect 8485 -2675 8515 -2645
rect 8515 -2675 8516 -2645
rect 8484 -2676 8516 -2675
rect 8484 -2725 8516 -2724
rect 8484 -2755 8485 -2725
rect 8485 -2755 8515 -2725
rect 8515 -2755 8516 -2725
rect 8484 -2756 8516 -2755
rect 8484 -2836 8516 -2804
rect 8484 -2885 8516 -2884
rect 8484 -2915 8485 -2885
rect 8485 -2915 8515 -2885
rect 8515 -2915 8516 -2885
rect 8484 -2916 8516 -2915
rect 8484 -2996 8516 -2964
rect 8484 -3045 8516 -3044
rect 8484 -3075 8485 -3045
rect 8485 -3075 8515 -3045
rect 8515 -3075 8516 -3045
rect 8484 -3076 8516 -3075
rect 8484 -3156 8516 -3124
rect 8484 -3205 8516 -3204
rect 8484 -3235 8485 -3205
rect 8485 -3235 8515 -3205
rect 8515 -3235 8516 -3205
rect 8484 -3236 8516 -3235
rect 8484 -3285 8516 -3284
rect 8484 -3315 8485 -3285
rect 8485 -3315 8515 -3285
rect 8515 -3315 8516 -3285
rect 8484 -3316 8516 -3315
rect 8484 -3396 8516 -3364
rect 8484 -3476 8516 -3444
rect 8484 -3525 8516 -3524
rect 8484 -3555 8485 -3525
rect 8485 -3555 8515 -3525
rect 8515 -3555 8516 -3525
rect 8484 -3556 8516 -3555
rect 8484 -3605 8516 -3604
rect 8484 -3635 8485 -3605
rect 8485 -3635 8515 -3605
rect 8515 -3635 8516 -3605
rect 8484 -3636 8516 -3635
rect 8484 -3685 8516 -3684
rect 8484 -3715 8485 -3685
rect 8485 -3715 8515 -3685
rect 8515 -3715 8516 -3685
rect 8484 -3716 8516 -3715
rect 8564 1035 8596 1036
rect 8564 1005 8565 1035
rect 8565 1005 8595 1035
rect 8595 1005 8596 1035
rect 8564 1004 8596 1005
rect 8564 955 8596 956
rect 8564 925 8565 955
rect 8565 925 8595 955
rect 8595 925 8596 955
rect 8564 924 8596 925
rect 8564 875 8596 876
rect 8564 845 8565 875
rect 8565 845 8595 875
rect 8595 845 8596 875
rect 8564 844 8596 845
rect 8564 764 8596 796
rect 8564 684 8596 716
rect 8564 635 8596 636
rect 8564 605 8565 635
rect 8565 605 8595 635
rect 8595 605 8596 635
rect 8564 604 8596 605
rect 8564 555 8596 556
rect 8564 525 8565 555
rect 8565 525 8595 555
rect 8595 525 8596 555
rect 8564 524 8596 525
rect 8564 444 8596 476
rect 8564 395 8596 396
rect 8564 365 8565 395
rect 8565 365 8595 395
rect 8595 365 8596 395
rect 8564 364 8596 365
rect 8564 284 8596 316
rect 8564 235 8596 236
rect 8564 205 8565 235
rect 8565 205 8595 235
rect 8595 205 8596 235
rect 8564 204 8596 205
rect 8564 124 8596 156
rect 8564 75 8596 76
rect 8564 45 8565 75
rect 8565 45 8595 75
rect 8595 45 8596 75
rect 8564 44 8596 45
rect 8564 -5 8596 -4
rect 8564 -35 8565 -5
rect 8565 -35 8595 -5
rect 8595 -35 8596 -5
rect 8564 -36 8596 -35
rect 8564 -85 8596 -84
rect 8564 -115 8565 -85
rect 8565 -115 8595 -85
rect 8595 -115 8596 -85
rect 8564 -116 8596 -115
rect 8564 -165 8596 -164
rect 8564 -195 8565 -165
rect 8565 -195 8595 -165
rect 8595 -195 8596 -165
rect 8564 -196 8596 -195
rect 8564 -245 8596 -244
rect 8564 -275 8565 -245
rect 8565 -275 8595 -245
rect 8595 -275 8596 -245
rect 8564 -276 8596 -275
rect 8564 -325 8596 -324
rect 8564 -355 8565 -325
rect 8565 -355 8595 -325
rect 8595 -355 8596 -325
rect 8564 -356 8596 -355
rect 8564 -436 8596 -404
rect 8564 -485 8596 -484
rect 8564 -515 8565 -485
rect 8565 -515 8595 -485
rect 8595 -515 8596 -485
rect 8564 -516 8596 -515
rect 8564 -596 8596 -564
rect 8564 -645 8596 -644
rect 8564 -675 8565 -645
rect 8565 -675 8595 -645
rect 8595 -675 8596 -645
rect 8564 -676 8596 -675
rect 8564 -756 8596 -724
rect 8564 -805 8596 -804
rect 8564 -835 8565 -805
rect 8565 -835 8595 -805
rect 8595 -835 8596 -805
rect 8564 -836 8596 -835
rect 8564 -885 8596 -884
rect 8564 -915 8565 -885
rect 8565 -915 8595 -885
rect 8595 -915 8596 -885
rect 8564 -916 8596 -915
rect 8564 -996 8596 -964
rect 8564 -1076 8596 -1044
rect 8564 -1125 8596 -1124
rect 8564 -1155 8565 -1125
rect 8565 -1155 8595 -1125
rect 8595 -1155 8596 -1125
rect 8564 -1156 8596 -1155
rect 8564 -1205 8596 -1204
rect 8564 -1235 8565 -1205
rect 8565 -1235 8595 -1205
rect 8595 -1235 8596 -1205
rect 8564 -1236 8596 -1235
rect 8564 -1285 8596 -1284
rect 8564 -1315 8565 -1285
rect 8565 -1315 8595 -1285
rect 8595 -1315 8596 -1285
rect 8564 -1316 8596 -1315
rect 8564 -1365 8596 -1364
rect 8564 -1395 8565 -1365
rect 8565 -1395 8595 -1365
rect 8595 -1395 8596 -1365
rect 8564 -1396 8596 -1395
rect 8564 -1445 8596 -1444
rect 8564 -1475 8565 -1445
rect 8565 -1475 8595 -1445
rect 8595 -1475 8596 -1445
rect 8564 -1476 8596 -1475
rect 8564 -1525 8596 -1524
rect 8564 -1555 8565 -1525
rect 8565 -1555 8595 -1525
rect 8595 -1555 8596 -1525
rect 8564 -1556 8596 -1555
rect 8564 -1636 8596 -1604
rect 8564 -1716 8596 -1684
rect 8564 -1765 8596 -1764
rect 8564 -1795 8565 -1765
rect 8565 -1795 8595 -1765
rect 8595 -1795 8596 -1765
rect 8564 -1796 8596 -1795
rect 8564 -1845 8596 -1844
rect 8564 -1875 8565 -1845
rect 8565 -1875 8595 -1845
rect 8595 -1875 8596 -1845
rect 8564 -1876 8596 -1875
rect 8564 -1956 8596 -1924
rect 8564 -2005 8596 -2004
rect 8564 -2035 8565 -2005
rect 8565 -2035 8595 -2005
rect 8595 -2035 8596 -2005
rect 8564 -2036 8596 -2035
rect 8564 -2116 8596 -2084
rect 8564 -2165 8596 -2164
rect 8564 -2195 8565 -2165
rect 8565 -2195 8595 -2165
rect 8595 -2195 8596 -2165
rect 8564 -2196 8596 -2195
rect 8564 -2276 8596 -2244
rect 8564 -2325 8596 -2324
rect 8564 -2355 8565 -2325
rect 8565 -2355 8595 -2325
rect 8595 -2355 8596 -2325
rect 8564 -2356 8596 -2355
rect 8564 -2405 8596 -2404
rect 8564 -2435 8565 -2405
rect 8565 -2435 8595 -2405
rect 8595 -2435 8596 -2405
rect 8564 -2436 8596 -2435
rect 8564 -2485 8596 -2484
rect 8564 -2515 8565 -2485
rect 8565 -2515 8595 -2485
rect 8595 -2515 8596 -2485
rect 8564 -2516 8596 -2515
rect 8564 -2565 8596 -2564
rect 8564 -2595 8565 -2565
rect 8565 -2595 8595 -2565
rect 8595 -2595 8596 -2565
rect 8564 -2596 8596 -2595
rect 8564 -2645 8596 -2644
rect 8564 -2675 8565 -2645
rect 8565 -2675 8595 -2645
rect 8595 -2675 8596 -2645
rect 8564 -2676 8596 -2675
rect 8564 -2725 8596 -2724
rect 8564 -2755 8565 -2725
rect 8565 -2755 8595 -2725
rect 8595 -2755 8596 -2725
rect 8564 -2756 8596 -2755
rect 8564 -2836 8596 -2804
rect 8564 -2885 8596 -2884
rect 8564 -2915 8565 -2885
rect 8565 -2915 8595 -2885
rect 8595 -2915 8596 -2885
rect 8564 -2916 8596 -2915
rect 8564 -2996 8596 -2964
rect 8564 -3045 8596 -3044
rect 8564 -3075 8565 -3045
rect 8565 -3075 8595 -3045
rect 8595 -3075 8596 -3045
rect 8564 -3076 8596 -3075
rect 8564 -3156 8596 -3124
rect 8564 -3205 8596 -3204
rect 8564 -3235 8565 -3205
rect 8565 -3235 8595 -3205
rect 8595 -3235 8596 -3205
rect 8564 -3236 8596 -3235
rect 8564 -3285 8596 -3284
rect 8564 -3315 8565 -3285
rect 8565 -3315 8595 -3285
rect 8595 -3315 8596 -3285
rect 8564 -3316 8596 -3315
rect 8564 -3396 8596 -3364
rect 8564 -3476 8596 -3444
rect 8564 -3525 8596 -3524
rect 8564 -3555 8565 -3525
rect 8565 -3555 8595 -3525
rect 8595 -3555 8596 -3525
rect 8564 -3556 8596 -3555
rect 8564 -3605 8596 -3604
rect 8564 -3635 8565 -3605
rect 8565 -3635 8595 -3605
rect 8595 -3635 8596 -3605
rect 8564 -3636 8596 -3635
rect 8564 -3685 8596 -3684
rect 8564 -3715 8565 -3685
rect 8565 -3715 8595 -3685
rect 8595 -3715 8596 -3685
rect 8564 -3716 8596 -3715
rect 8644 1035 8676 1036
rect 8644 1005 8645 1035
rect 8645 1005 8675 1035
rect 8675 1005 8676 1035
rect 8644 1004 8676 1005
rect 8644 955 8676 956
rect 8644 925 8645 955
rect 8645 925 8675 955
rect 8675 925 8676 955
rect 8644 924 8676 925
rect 8644 875 8676 876
rect 8644 845 8645 875
rect 8645 845 8675 875
rect 8675 845 8676 875
rect 8644 844 8676 845
rect 8644 764 8676 796
rect 8644 684 8676 716
rect 8644 635 8676 636
rect 8644 605 8645 635
rect 8645 605 8675 635
rect 8675 605 8676 635
rect 8644 604 8676 605
rect 8644 555 8676 556
rect 8644 525 8645 555
rect 8645 525 8675 555
rect 8675 525 8676 555
rect 8644 524 8676 525
rect 8644 444 8676 476
rect 8644 395 8676 396
rect 8644 365 8645 395
rect 8645 365 8675 395
rect 8675 365 8676 395
rect 8644 364 8676 365
rect 8644 284 8676 316
rect 8644 235 8676 236
rect 8644 205 8645 235
rect 8645 205 8675 235
rect 8675 205 8676 235
rect 8644 204 8676 205
rect 8644 124 8676 156
rect 8644 75 8676 76
rect 8644 45 8645 75
rect 8645 45 8675 75
rect 8675 45 8676 75
rect 8644 44 8676 45
rect 8644 -5 8676 -4
rect 8644 -35 8645 -5
rect 8645 -35 8675 -5
rect 8675 -35 8676 -5
rect 8644 -36 8676 -35
rect 8644 -85 8676 -84
rect 8644 -115 8645 -85
rect 8645 -115 8675 -85
rect 8675 -115 8676 -85
rect 8644 -116 8676 -115
rect 8644 -165 8676 -164
rect 8644 -195 8645 -165
rect 8645 -195 8675 -165
rect 8675 -195 8676 -165
rect 8644 -196 8676 -195
rect 8644 -245 8676 -244
rect 8644 -275 8645 -245
rect 8645 -275 8675 -245
rect 8675 -275 8676 -245
rect 8644 -276 8676 -275
rect 8644 -325 8676 -324
rect 8644 -355 8645 -325
rect 8645 -355 8675 -325
rect 8675 -355 8676 -325
rect 8644 -356 8676 -355
rect 8644 -436 8676 -404
rect 8644 -485 8676 -484
rect 8644 -515 8645 -485
rect 8645 -515 8675 -485
rect 8675 -515 8676 -485
rect 8644 -516 8676 -515
rect 8644 -596 8676 -564
rect 8644 -645 8676 -644
rect 8644 -675 8645 -645
rect 8645 -675 8675 -645
rect 8675 -675 8676 -645
rect 8644 -676 8676 -675
rect 8644 -756 8676 -724
rect 8644 -805 8676 -804
rect 8644 -835 8645 -805
rect 8645 -835 8675 -805
rect 8675 -835 8676 -805
rect 8644 -836 8676 -835
rect 8644 -885 8676 -884
rect 8644 -915 8645 -885
rect 8645 -915 8675 -885
rect 8675 -915 8676 -885
rect 8644 -916 8676 -915
rect 8644 -996 8676 -964
rect 8644 -1076 8676 -1044
rect 8644 -1125 8676 -1124
rect 8644 -1155 8645 -1125
rect 8645 -1155 8675 -1125
rect 8675 -1155 8676 -1125
rect 8644 -1156 8676 -1155
rect 8644 -1205 8676 -1204
rect 8644 -1235 8645 -1205
rect 8645 -1235 8675 -1205
rect 8675 -1235 8676 -1205
rect 8644 -1236 8676 -1235
rect 8644 -1285 8676 -1284
rect 8644 -1315 8645 -1285
rect 8645 -1315 8675 -1285
rect 8675 -1315 8676 -1285
rect 8644 -1316 8676 -1315
rect 8644 -1365 8676 -1364
rect 8644 -1395 8645 -1365
rect 8645 -1395 8675 -1365
rect 8675 -1395 8676 -1365
rect 8644 -1396 8676 -1395
rect 8644 -1445 8676 -1444
rect 8644 -1475 8645 -1445
rect 8645 -1475 8675 -1445
rect 8675 -1475 8676 -1445
rect 8644 -1476 8676 -1475
rect 8644 -1525 8676 -1524
rect 8644 -1555 8645 -1525
rect 8645 -1555 8675 -1525
rect 8675 -1555 8676 -1525
rect 8644 -1556 8676 -1555
rect 8644 -1636 8676 -1604
rect 8644 -1716 8676 -1684
rect 8644 -1765 8676 -1764
rect 8644 -1795 8645 -1765
rect 8645 -1795 8675 -1765
rect 8675 -1795 8676 -1765
rect 8644 -1796 8676 -1795
rect 8644 -1845 8676 -1844
rect 8644 -1875 8645 -1845
rect 8645 -1875 8675 -1845
rect 8675 -1875 8676 -1845
rect 8644 -1876 8676 -1875
rect 8644 -1956 8676 -1924
rect 8644 -2005 8676 -2004
rect 8644 -2035 8645 -2005
rect 8645 -2035 8675 -2005
rect 8675 -2035 8676 -2005
rect 8644 -2036 8676 -2035
rect 8644 -2116 8676 -2084
rect 8644 -2165 8676 -2164
rect 8644 -2195 8645 -2165
rect 8645 -2195 8675 -2165
rect 8675 -2195 8676 -2165
rect 8644 -2196 8676 -2195
rect 8644 -2276 8676 -2244
rect 8644 -2325 8676 -2324
rect 8644 -2355 8645 -2325
rect 8645 -2355 8675 -2325
rect 8675 -2355 8676 -2325
rect 8644 -2356 8676 -2355
rect 8644 -2405 8676 -2404
rect 8644 -2435 8645 -2405
rect 8645 -2435 8675 -2405
rect 8675 -2435 8676 -2405
rect 8644 -2436 8676 -2435
rect 8644 -2485 8676 -2484
rect 8644 -2515 8645 -2485
rect 8645 -2515 8675 -2485
rect 8675 -2515 8676 -2485
rect 8644 -2516 8676 -2515
rect 8644 -2565 8676 -2564
rect 8644 -2595 8645 -2565
rect 8645 -2595 8675 -2565
rect 8675 -2595 8676 -2565
rect 8644 -2596 8676 -2595
rect 8644 -2645 8676 -2644
rect 8644 -2675 8645 -2645
rect 8645 -2675 8675 -2645
rect 8675 -2675 8676 -2645
rect 8644 -2676 8676 -2675
rect 8644 -2725 8676 -2724
rect 8644 -2755 8645 -2725
rect 8645 -2755 8675 -2725
rect 8675 -2755 8676 -2725
rect 8644 -2756 8676 -2755
rect 8644 -2836 8676 -2804
rect 8644 -2885 8676 -2884
rect 8644 -2915 8645 -2885
rect 8645 -2915 8675 -2885
rect 8675 -2915 8676 -2885
rect 8644 -2916 8676 -2915
rect 8644 -2996 8676 -2964
rect 8644 -3045 8676 -3044
rect 8644 -3075 8645 -3045
rect 8645 -3075 8675 -3045
rect 8675 -3075 8676 -3045
rect 8644 -3076 8676 -3075
rect 8644 -3156 8676 -3124
rect 8644 -3205 8676 -3204
rect 8644 -3235 8645 -3205
rect 8645 -3235 8675 -3205
rect 8675 -3235 8676 -3205
rect 8644 -3236 8676 -3235
rect 8644 -3285 8676 -3284
rect 8644 -3315 8645 -3285
rect 8645 -3315 8675 -3285
rect 8675 -3315 8676 -3285
rect 8644 -3316 8676 -3315
rect 8644 -3396 8676 -3364
rect 8644 -3476 8676 -3444
rect 8644 -3525 8676 -3524
rect 8644 -3555 8645 -3525
rect 8645 -3555 8675 -3525
rect 8675 -3555 8676 -3525
rect 8644 -3556 8676 -3555
rect 8644 -3605 8676 -3604
rect 8644 -3635 8645 -3605
rect 8645 -3635 8675 -3605
rect 8675 -3635 8676 -3605
rect 8644 -3636 8676 -3635
rect 8644 -3685 8676 -3684
rect 8644 -3715 8645 -3685
rect 8645 -3715 8675 -3685
rect 8675 -3715 8676 -3685
rect 8644 -3716 8676 -3715
rect 8724 1035 8756 1036
rect 8724 1005 8725 1035
rect 8725 1005 8755 1035
rect 8755 1005 8756 1035
rect 8724 1004 8756 1005
rect 8724 955 8756 956
rect 8724 925 8725 955
rect 8725 925 8755 955
rect 8755 925 8756 955
rect 8724 924 8756 925
rect 8724 875 8756 876
rect 8724 845 8725 875
rect 8725 845 8755 875
rect 8755 845 8756 875
rect 8724 844 8756 845
rect 8724 764 8756 796
rect 8724 684 8756 716
rect 8724 635 8756 636
rect 8724 605 8725 635
rect 8725 605 8755 635
rect 8755 605 8756 635
rect 8724 604 8756 605
rect 8724 555 8756 556
rect 8724 525 8725 555
rect 8725 525 8755 555
rect 8755 525 8756 555
rect 8724 524 8756 525
rect 8724 444 8756 476
rect 8724 395 8756 396
rect 8724 365 8725 395
rect 8725 365 8755 395
rect 8755 365 8756 395
rect 8724 364 8756 365
rect 8724 284 8756 316
rect 8724 235 8756 236
rect 8724 205 8725 235
rect 8725 205 8755 235
rect 8755 205 8756 235
rect 8724 204 8756 205
rect 8724 124 8756 156
rect 8724 75 8756 76
rect 8724 45 8725 75
rect 8725 45 8755 75
rect 8755 45 8756 75
rect 8724 44 8756 45
rect 8724 -5 8756 -4
rect 8724 -35 8725 -5
rect 8725 -35 8755 -5
rect 8755 -35 8756 -5
rect 8724 -36 8756 -35
rect 8724 -85 8756 -84
rect 8724 -115 8725 -85
rect 8725 -115 8755 -85
rect 8755 -115 8756 -85
rect 8724 -116 8756 -115
rect 8724 -165 8756 -164
rect 8724 -195 8725 -165
rect 8725 -195 8755 -165
rect 8755 -195 8756 -165
rect 8724 -196 8756 -195
rect 8724 -245 8756 -244
rect 8724 -275 8725 -245
rect 8725 -275 8755 -245
rect 8755 -275 8756 -245
rect 8724 -276 8756 -275
rect 8724 -325 8756 -324
rect 8724 -355 8725 -325
rect 8725 -355 8755 -325
rect 8755 -355 8756 -325
rect 8724 -356 8756 -355
rect 8724 -436 8756 -404
rect 8724 -485 8756 -484
rect 8724 -515 8725 -485
rect 8725 -515 8755 -485
rect 8755 -515 8756 -485
rect 8724 -516 8756 -515
rect 8724 -596 8756 -564
rect 8724 -645 8756 -644
rect 8724 -675 8725 -645
rect 8725 -675 8755 -645
rect 8755 -675 8756 -645
rect 8724 -676 8756 -675
rect 8724 -756 8756 -724
rect 8724 -805 8756 -804
rect 8724 -835 8725 -805
rect 8725 -835 8755 -805
rect 8755 -835 8756 -805
rect 8724 -836 8756 -835
rect 8724 -885 8756 -884
rect 8724 -915 8725 -885
rect 8725 -915 8755 -885
rect 8755 -915 8756 -885
rect 8724 -916 8756 -915
rect 8724 -996 8756 -964
rect 8724 -1076 8756 -1044
rect 8724 -1125 8756 -1124
rect 8724 -1155 8725 -1125
rect 8725 -1155 8755 -1125
rect 8755 -1155 8756 -1125
rect 8724 -1156 8756 -1155
rect 8724 -1205 8756 -1204
rect 8724 -1235 8725 -1205
rect 8725 -1235 8755 -1205
rect 8755 -1235 8756 -1205
rect 8724 -1236 8756 -1235
rect 8724 -1285 8756 -1284
rect 8724 -1315 8725 -1285
rect 8725 -1315 8755 -1285
rect 8755 -1315 8756 -1285
rect 8724 -1316 8756 -1315
rect 8724 -1365 8756 -1364
rect 8724 -1395 8725 -1365
rect 8725 -1395 8755 -1365
rect 8755 -1395 8756 -1365
rect 8724 -1396 8756 -1395
rect 8724 -1445 8756 -1444
rect 8724 -1475 8725 -1445
rect 8725 -1475 8755 -1445
rect 8755 -1475 8756 -1445
rect 8724 -1476 8756 -1475
rect 8724 -1525 8756 -1524
rect 8724 -1555 8725 -1525
rect 8725 -1555 8755 -1525
rect 8755 -1555 8756 -1525
rect 8724 -1556 8756 -1555
rect 8724 -1636 8756 -1604
rect 8724 -1716 8756 -1684
rect 8724 -1765 8756 -1764
rect 8724 -1795 8725 -1765
rect 8725 -1795 8755 -1765
rect 8755 -1795 8756 -1765
rect 8724 -1796 8756 -1795
rect 8724 -1845 8756 -1844
rect 8724 -1875 8725 -1845
rect 8725 -1875 8755 -1845
rect 8755 -1875 8756 -1845
rect 8724 -1876 8756 -1875
rect 8724 -1956 8756 -1924
rect 8724 -2005 8756 -2004
rect 8724 -2035 8725 -2005
rect 8725 -2035 8755 -2005
rect 8755 -2035 8756 -2005
rect 8724 -2036 8756 -2035
rect 8724 -2116 8756 -2084
rect 8724 -2165 8756 -2164
rect 8724 -2195 8725 -2165
rect 8725 -2195 8755 -2165
rect 8755 -2195 8756 -2165
rect 8724 -2196 8756 -2195
rect 8724 -2276 8756 -2244
rect 8724 -2325 8756 -2324
rect 8724 -2355 8725 -2325
rect 8725 -2355 8755 -2325
rect 8755 -2355 8756 -2325
rect 8724 -2356 8756 -2355
rect 8724 -2405 8756 -2404
rect 8724 -2435 8725 -2405
rect 8725 -2435 8755 -2405
rect 8755 -2435 8756 -2405
rect 8724 -2436 8756 -2435
rect 8724 -2485 8756 -2484
rect 8724 -2515 8725 -2485
rect 8725 -2515 8755 -2485
rect 8755 -2515 8756 -2485
rect 8724 -2516 8756 -2515
rect 8724 -2565 8756 -2564
rect 8724 -2595 8725 -2565
rect 8725 -2595 8755 -2565
rect 8755 -2595 8756 -2565
rect 8724 -2596 8756 -2595
rect 8724 -2645 8756 -2644
rect 8724 -2675 8725 -2645
rect 8725 -2675 8755 -2645
rect 8755 -2675 8756 -2645
rect 8724 -2676 8756 -2675
rect 8724 -2725 8756 -2724
rect 8724 -2755 8725 -2725
rect 8725 -2755 8755 -2725
rect 8755 -2755 8756 -2725
rect 8724 -2756 8756 -2755
rect 8724 -2836 8756 -2804
rect 8724 -2885 8756 -2884
rect 8724 -2915 8725 -2885
rect 8725 -2915 8755 -2885
rect 8755 -2915 8756 -2885
rect 8724 -2916 8756 -2915
rect 8724 -2996 8756 -2964
rect 8724 -3045 8756 -3044
rect 8724 -3075 8725 -3045
rect 8725 -3075 8755 -3045
rect 8755 -3075 8756 -3045
rect 8724 -3076 8756 -3075
rect 8724 -3156 8756 -3124
rect 8724 -3205 8756 -3204
rect 8724 -3235 8725 -3205
rect 8725 -3235 8755 -3205
rect 8755 -3235 8756 -3205
rect 8724 -3236 8756 -3235
rect 8724 -3285 8756 -3284
rect 8724 -3315 8725 -3285
rect 8725 -3315 8755 -3285
rect 8755 -3315 8756 -3285
rect 8724 -3316 8756 -3315
rect 8724 -3396 8756 -3364
rect 8724 -3476 8756 -3444
rect 8724 -3525 8756 -3524
rect 8724 -3555 8725 -3525
rect 8725 -3555 8755 -3525
rect 8755 -3555 8756 -3525
rect 8724 -3556 8756 -3555
rect 8724 -3605 8756 -3604
rect 8724 -3635 8725 -3605
rect 8725 -3635 8755 -3605
rect 8755 -3635 8756 -3605
rect 8724 -3636 8756 -3635
rect 8724 -3685 8756 -3684
rect 8724 -3715 8725 -3685
rect 8725 -3715 8755 -3685
rect 8755 -3715 8756 -3685
rect 8724 -3716 8756 -3715
rect 8804 1035 8836 1036
rect 8804 1005 8805 1035
rect 8805 1005 8835 1035
rect 8835 1005 8836 1035
rect 8804 1004 8836 1005
rect 8804 955 8836 956
rect 8804 925 8805 955
rect 8805 925 8835 955
rect 8835 925 8836 955
rect 8804 924 8836 925
rect 8804 875 8836 876
rect 8804 845 8805 875
rect 8805 845 8835 875
rect 8835 845 8836 875
rect 8804 844 8836 845
rect 8804 764 8836 796
rect 8804 684 8836 716
rect 8804 635 8836 636
rect 8804 605 8805 635
rect 8805 605 8835 635
rect 8835 605 8836 635
rect 8804 604 8836 605
rect 8804 555 8836 556
rect 8804 525 8805 555
rect 8805 525 8835 555
rect 8835 525 8836 555
rect 8804 524 8836 525
rect 8804 444 8836 476
rect 8804 395 8836 396
rect 8804 365 8805 395
rect 8805 365 8835 395
rect 8835 365 8836 395
rect 8804 364 8836 365
rect 8804 284 8836 316
rect 8804 235 8836 236
rect 8804 205 8805 235
rect 8805 205 8835 235
rect 8835 205 8836 235
rect 8804 204 8836 205
rect 8804 124 8836 156
rect 8804 75 8836 76
rect 8804 45 8805 75
rect 8805 45 8835 75
rect 8835 45 8836 75
rect 8804 44 8836 45
rect 8804 -5 8836 -4
rect 8804 -35 8805 -5
rect 8805 -35 8835 -5
rect 8835 -35 8836 -5
rect 8804 -36 8836 -35
rect 8804 -85 8836 -84
rect 8804 -115 8805 -85
rect 8805 -115 8835 -85
rect 8835 -115 8836 -85
rect 8804 -116 8836 -115
rect 8804 -165 8836 -164
rect 8804 -195 8805 -165
rect 8805 -195 8835 -165
rect 8835 -195 8836 -165
rect 8804 -196 8836 -195
rect 8804 -245 8836 -244
rect 8804 -275 8805 -245
rect 8805 -275 8835 -245
rect 8835 -275 8836 -245
rect 8804 -276 8836 -275
rect 8804 -325 8836 -324
rect 8804 -355 8805 -325
rect 8805 -355 8835 -325
rect 8835 -355 8836 -325
rect 8804 -356 8836 -355
rect 8804 -436 8836 -404
rect 8804 -485 8836 -484
rect 8804 -515 8805 -485
rect 8805 -515 8835 -485
rect 8835 -515 8836 -485
rect 8804 -516 8836 -515
rect 8804 -596 8836 -564
rect 8804 -645 8836 -644
rect 8804 -675 8805 -645
rect 8805 -675 8835 -645
rect 8835 -675 8836 -645
rect 8804 -676 8836 -675
rect 8804 -756 8836 -724
rect 8804 -805 8836 -804
rect 8804 -835 8805 -805
rect 8805 -835 8835 -805
rect 8835 -835 8836 -805
rect 8804 -836 8836 -835
rect 8804 -885 8836 -884
rect 8804 -915 8805 -885
rect 8805 -915 8835 -885
rect 8835 -915 8836 -885
rect 8804 -916 8836 -915
rect 8804 -996 8836 -964
rect 8804 -1076 8836 -1044
rect 8804 -1125 8836 -1124
rect 8804 -1155 8805 -1125
rect 8805 -1155 8835 -1125
rect 8835 -1155 8836 -1125
rect 8804 -1156 8836 -1155
rect 8804 -1205 8836 -1204
rect 8804 -1235 8805 -1205
rect 8805 -1235 8835 -1205
rect 8835 -1235 8836 -1205
rect 8804 -1236 8836 -1235
rect 8804 -1285 8836 -1284
rect 8804 -1315 8805 -1285
rect 8805 -1315 8835 -1285
rect 8835 -1315 8836 -1285
rect 8804 -1316 8836 -1315
rect 8804 -1365 8836 -1364
rect 8804 -1395 8805 -1365
rect 8805 -1395 8835 -1365
rect 8835 -1395 8836 -1365
rect 8804 -1396 8836 -1395
rect 8804 -1445 8836 -1444
rect 8804 -1475 8805 -1445
rect 8805 -1475 8835 -1445
rect 8835 -1475 8836 -1445
rect 8804 -1476 8836 -1475
rect 8804 -1525 8836 -1524
rect 8804 -1555 8805 -1525
rect 8805 -1555 8835 -1525
rect 8835 -1555 8836 -1525
rect 8804 -1556 8836 -1555
rect 8804 -1636 8836 -1604
rect 8804 -1716 8836 -1684
rect 8804 -1765 8836 -1764
rect 8804 -1795 8805 -1765
rect 8805 -1795 8835 -1765
rect 8835 -1795 8836 -1765
rect 8804 -1796 8836 -1795
rect 8804 -1845 8836 -1844
rect 8804 -1875 8805 -1845
rect 8805 -1875 8835 -1845
rect 8835 -1875 8836 -1845
rect 8804 -1876 8836 -1875
rect 8804 -1956 8836 -1924
rect 8804 -2005 8836 -2004
rect 8804 -2035 8805 -2005
rect 8805 -2035 8835 -2005
rect 8835 -2035 8836 -2005
rect 8804 -2036 8836 -2035
rect 8804 -2116 8836 -2084
rect 8804 -2165 8836 -2164
rect 8804 -2195 8805 -2165
rect 8805 -2195 8835 -2165
rect 8835 -2195 8836 -2165
rect 8804 -2196 8836 -2195
rect 8804 -2276 8836 -2244
rect 8804 -2325 8836 -2324
rect 8804 -2355 8805 -2325
rect 8805 -2355 8835 -2325
rect 8835 -2355 8836 -2325
rect 8804 -2356 8836 -2355
rect 8804 -2405 8836 -2404
rect 8804 -2435 8805 -2405
rect 8805 -2435 8835 -2405
rect 8835 -2435 8836 -2405
rect 8804 -2436 8836 -2435
rect 8804 -2485 8836 -2484
rect 8804 -2515 8805 -2485
rect 8805 -2515 8835 -2485
rect 8835 -2515 8836 -2485
rect 8804 -2516 8836 -2515
rect 8804 -2565 8836 -2564
rect 8804 -2595 8805 -2565
rect 8805 -2595 8835 -2565
rect 8835 -2595 8836 -2565
rect 8804 -2596 8836 -2595
rect 8804 -2645 8836 -2644
rect 8804 -2675 8805 -2645
rect 8805 -2675 8835 -2645
rect 8835 -2675 8836 -2645
rect 8804 -2676 8836 -2675
rect 8804 -2725 8836 -2724
rect 8804 -2755 8805 -2725
rect 8805 -2755 8835 -2725
rect 8835 -2755 8836 -2725
rect 8804 -2756 8836 -2755
rect 8804 -2836 8836 -2804
rect 8804 -2885 8836 -2884
rect 8804 -2915 8805 -2885
rect 8805 -2915 8835 -2885
rect 8835 -2915 8836 -2885
rect 8804 -2916 8836 -2915
rect 8804 -2996 8836 -2964
rect 8804 -3045 8836 -3044
rect 8804 -3075 8805 -3045
rect 8805 -3075 8835 -3045
rect 8835 -3075 8836 -3045
rect 8804 -3076 8836 -3075
rect 8804 -3156 8836 -3124
rect 8804 -3205 8836 -3204
rect 8804 -3235 8805 -3205
rect 8805 -3235 8835 -3205
rect 8835 -3235 8836 -3205
rect 8804 -3236 8836 -3235
rect 8804 -3285 8836 -3284
rect 8804 -3315 8805 -3285
rect 8805 -3315 8835 -3285
rect 8835 -3315 8836 -3285
rect 8804 -3316 8836 -3315
rect 8804 -3396 8836 -3364
rect 8804 -3476 8836 -3444
rect 8804 -3525 8836 -3524
rect 8804 -3555 8805 -3525
rect 8805 -3555 8835 -3525
rect 8835 -3555 8836 -3525
rect 8804 -3556 8836 -3555
rect 8804 -3605 8836 -3604
rect 8804 -3635 8805 -3605
rect 8805 -3635 8835 -3605
rect 8835 -3635 8836 -3605
rect 8804 -3636 8836 -3635
rect 8804 -3685 8836 -3684
rect 8804 -3715 8805 -3685
rect 8805 -3715 8835 -3685
rect 8835 -3715 8836 -3685
rect 8804 -3716 8836 -3715
rect 8884 1035 8916 1036
rect 8884 1005 8885 1035
rect 8885 1005 8915 1035
rect 8915 1005 8916 1035
rect 8884 1004 8916 1005
rect 8884 955 8916 956
rect 8884 925 8885 955
rect 8885 925 8915 955
rect 8915 925 8916 955
rect 8884 924 8916 925
rect 8884 875 8916 876
rect 8884 845 8885 875
rect 8885 845 8915 875
rect 8915 845 8916 875
rect 8884 844 8916 845
rect 8884 764 8916 796
rect 8884 684 8916 716
rect 8884 635 8916 636
rect 8884 605 8885 635
rect 8885 605 8915 635
rect 8915 605 8916 635
rect 8884 604 8916 605
rect 8884 555 8916 556
rect 8884 525 8885 555
rect 8885 525 8915 555
rect 8915 525 8916 555
rect 8884 524 8916 525
rect 8884 444 8916 476
rect 8884 395 8916 396
rect 8884 365 8885 395
rect 8885 365 8915 395
rect 8915 365 8916 395
rect 8884 364 8916 365
rect 8884 284 8916 316
rect 8884 235 8916 236
rect 8884 205 8885 235
rect 8885 205 8915 235
rect 8915 205 8916 235
rect 8884 204 8916 205
rect 8884 124 8916 156
rect 8884 75 8916 76
rect 8884 45 8885 75
rect 8885 45 8915 75
rect 8915 45 8916 75
rect 8884 44 8916 45
rect 8884 -5 8916 -4
rect 8884 -35 8885 -5
rect 8885 -35 8915 -5
rect 8915 -35 8916 -5
rect 8884 -36 8916 -35
rect 8884 -85 8916 -84
rect 8884 -115 8885 -85
rect 8885 -115 8915 -85
rect 8915 -115 8916 -85
rect 8884 -116 8916 -115
rect 8884 -165 8916 -164
rect 8884 -195 8885 -165
rect 8885 -195 8915 -165
rect 8915 -195 8916 -165
rect 8884 -196 8916 -195
rect 8884 -245 8916 -244
rect 8884 -275 8885 -245
rect 8885 -275 8915 -245
rect 8915 -275 8916 -245
rect 8884 -276 8916 -275
rect 8884 -325 8916 -324
rect 8884 -355 8885 -325
rect 8885 -355 8915 -325
rect 8915 -355 8916 -325
rect 8884 -356 8916 -355
rect 8884 -436 8916 -404
rect 8884 -485 8916 -484
rect 8884 -515 8885 -485
rect 8885 -515 8915 -485
rect 8915 -515 8916 -485
rect 8884 -516 8916 -515
rect 8884 -596 8916 -564
rect 8884 -645 8916 -644
rect 8884 -675 8885 -645
rect 8885 -675 8915 -645
rect 8915 -675 8916 -645
rect 8884 -676 8916 -675
rect 8884 -756 8916 -724
rect 8884 -805 8916 -804
rect 8884 -835 8885 -805
rect 8885 -835 8915 -805
rect 8915 -835 8916 -805
rect 8884 -836 8916 -835
rect 8884 -885 8916 -884
rect 8884 -915 8885 -885
rect 8885 -915 8915 -885
rect 8915 -915 8916 -885
rect 8884 -916 8916 -915
rect 8884 -996 8916 -964
rect 8884 -1076 8916 -1044
rect 8884 -1125 8916 -1124
rect 8884 -1155 8885 -1125
rect 8885 -1155 8915 -1125
rect 8915 -1155 8916 -1125
rect 8884 -1156 8916 -1155
rect 8884 -1205 8916 -1204
rect 8884 -1235 8885 -1205
rect 8885 -1235 8915 -1205
rect 8915 -1235 8916 -1205
rect 8884 -1236 8916 -1235
rect 8884 -1285 8916 -1284
rect 8884 -1315 8885 -1285
rect 8885 -1315 8915 -1285
rect 8915 -1315 8916 -1285
rect 8884 -1316 8916 -1315
rect 8884 -1365 8916 -1364
rect 8884 -1395 8885 -1365
rect 8885 -1395 8915 -1365
rect 8915 -1395 8916 -1365
rect 8884 -1396 8916 -1395
rect 8884 -1445 8916 -1444
rect 8884 -1475 8885 -1445
rect 8885 -1475 8915 -1445
rect 8915 -1475 8916 -1445
rect 8884 -1476 8916 -1475
rect 8884 -1525 8916 -1524
rect 8884 -1555 8885 -1525
rect 8885 -1555 8915 -1525
rect 8915 -1555 8916 -1525
rect 8884 -1556 8916 -1555
rect 8884 -1636 8916 -1604
rect 8884 -1716 8916 -1684
rect 8884 -1765 8916 -1764
rect 8884 -1795 8885 -1765
rect 8885 -1795 8915 -1765
rect 8915 -1795 8916 -1765
rect 8884 -1796 8916 -1795
rect 8884 -1845 8916 -1844
rect 8884 -1875 8885 -1845
rect 8885 -1875 8915 -1845
rect 8915 -1875 8916 -1845
rect 8884 -1876 8916 -1875
rect 8884 -1956 8916 -1924
rect 8884 -2005 8916 -2004
rect 8884 -2035 8885 -2005
rect 8885 -2035 8915 -2005
rect 8915 -2035 8916 -2005
rect 8884 -2036 8916 -2035
rect 8884 -2116 8916 -2084
rect 8884 -2165 8916 -2164
rect 8884 -2195 8885 -2165
rect 8885 -2195 8915 -2165
rect 8915 -2195 8916 -2165
rect 8884 -2196 8916 -2195
rect 8884 -2276 8916 -2244
rect 8884 -2325 8916 -2324
rect 8884 -2355 8885 -2325
rect 8885 -2355 8915 -2325
rect 8915 -2355 8916 -2325
rect 8884 -2356 8916 -2355
rect 8884 -2405 8916 -2404
rect 8884 -2435 8885 -2405
rect 8885 -2435 8915 -2405
rect 8915 -2435 8916 -2405
rect 8884 -2436 8916 -2435
rect 8884 -2485 8916 -2484
rect 8884 -2515 8885 -2485
rect 8885 -2515 8915 -2485
rect 8915 -2515 8916 -2485
rect 8884 -2516 8916 -2515
rect 8884 -2565 8916 -2564
rect 8884 -2595 8885 -2565
rect 8885 -2595 8915 -2565
rect 8915 -2595 8916 -2565
rect 8884 -2596 8916 -2595
rect 8884 -2645 8916 -2644
rect 8884 -2675 8885 -2645
rect 8885 -2675 8915 -2645
rect 8915 -2675 8916 -2645
rect 8884 -2676 8916 -2675
rect 8884 -2725 8916 -2724
rect 8884 -2755 8885 -2725
rect 8885 -2755 8915 -2725
rect 8915 -2755 8916 -2725
rect 8884 -2756 8916 -2755
rect 8884 -2836 8916 -2804
rect 8884 -2885 8916 -2884
rect 8884 -2915 8885 -2885
rect 8885 -2915 8915 -2885
rect 8915 -2915 8916 -2885
rect 8884 -2916 8916 -2915
rect 8884 -2996 8916 -2964
rect 8884 -3045 8916 -3044
rect 8884 -3075 8885 -3045
rect 8885 -3075 8915 -3045
rect 8915 -3075 8916 -3045
rect 8884 -3076 8916 -3075
rect 8884 -3156 8916 -3124
rect 8884 -3205 8916 -3204
rect 8884 -3235 8885 -3205
rect 8885 -3235 8915 -3205
rect 8915 -3235 8916 -3205
rect 8884 -3236 8916 -3235
rect 8884 -3285 8916 -3284
rect 8884 -3315 8885 -3285
rect 8885 -3315 8915 -3285
rect 8915 -3315 8916 -3285
rect 8884 -3316 8916 -3315
rect 8884 -3396 8916 -3364
rect 8884 -3476 8916 -3444
rect 8884 -3525 8916 -3524
rect 8884 -3555 8885 -3525
rect 8885 -3555 8915 -3525
rect 8915 -3555 8916 -3525
rect 8884 -3556 8916 -3555
rect 8884 -3605 8916 -3604
rect 8884 -3635 8885 -3605
rect 8885 -3635 8915 -3605
rect 8915 -3635 8916 -3605
rect 8884 -3636 8916 -3635
rect 8884 -3685 8916 -3684
rect 8884 -3715 8885 -3685
rect 8885 -3715 8915 -3685
rect 8915 -3715 8916 -3685
rect 8884 -3716 8916 -3715
rect 8964 1035 8996 1036
rect 8964 1005 8965 1035
rect 8965 1005 8995 1035
rect 8995 1005 8996 1035
rect 8964 1004 8996 1005
rect 8964 955 8996 956
rect 8964 925 8965 955
rect 8965 925 8995 955
rect 8995 925 8996 955
rect 8964 924 8996 925
rect 8964 875 8996 876
rect 8964 845 8965 875
rect 8965 845 8995 875
rect 8995 845 8996 875
rect 8964 844 8996 845
rect 8964 764 8996 796
rect 8964 684 8996 716
rect 8964 635 8996 636
rect 8964 605 8965 635
rect 8965 605 8995 635
rect 8995 605 8996 635
rect 8964 604 8996 605
rect 8964 555 8996 556
rect 8964 525 8965 555
rect 8965 525 8995 555
rect 8995 525 8996 555
rect 8964 524 8996 525
rect 8964 444 8996 476
rect 8964 395 8996 396
rect 8964 365 8965 395
rect 8965 365 8995 395
rect 8995 365 8996 395
rect 8964 364 8996 365
rect 8964 284 8996 316
rect 8964 235 8996 236
rect 8964 205 8965 235
rect 8965 205 8995 235
rect 8995 205 8996 235
rect 8964 204 8996 205
rect 8964 124 8996 156
rect 8964 75 8996 76
rect 8964 45 8965 75
rect 8965 45 8995 75
rect 8995 45 8996 75
rect 8964 44 8996 45
rect 8964 -5 8996 -4
rect 8964 -35 8965 -5
rect 8965 -35 8995 -5
rect 8995 -35 8996 -5
rect 8964 -36 8996 -35
rect 8964 -85 8996 -84
rect 8964 -115 8965 -85
rect 8965 -115 8995 -85
rect 8995 -115 8996 -85
rect 8964 -116 8996 -115
rect 8964 -165 8996 -164
rect 8964 -195 8965 -165
rect 8965 -195 8995 -165
rect 8995 -195 8996 -165
rect 8964 -196 8996 -195
rect 8964 -245 8996 -244
rect 8964 -275 8965 -245
rect 8965 -275 8995 -245
rect 8995 -275 8996 -245
rect 8964 -276 8996 -275
rect 8964 -325 8996 -324
rect 8964 -355 8965 -325
rect 8965 -355 8995 -325
rect 8995 -355 8996 -325
rect 8964 -356 8996 -355
rect 8964 -436 8996 -404
rect 8964 -485 8996 -484
rect 8964 -515 8965 -485
rect 8965 -515 8995 -485
rect 8995 -515 8996 -485
rect 8964 -516 8996 -515
rect 8964 -596 8996 -564
rect 8964 -645 8996 -644
rect 8964 -675 8965 -645
rect 8965 -675 8995 -645
rect 8995 -675 8996 -645
rect 8964 -676 8996 -675
rect 8964 -756 8996 -724
rect 8964 -805 8996 -804
rect 8964 -835 8965 -805
rect 8965 -835 8995 -805
rect 8995 -835 8996 -805
rect 8964 -836 8996 -835
rect 8964 -885 8996 -884
rect 8964 -915 8965 -885
rect 8965 -915 8995 -885
rect 8995 -915 8996 -885
rect 8964 -916 8996 -915
rect 8964 -996 8996 -964
rect 8964 -1076 8996 -1044
rect 8964 -1125 8996 -1124
rect 8964 -1155 8965 -1125
rect 8965 -1155 8995 -1125
rect 8995 -1155 8996 -1125
rect 8964 -1156 8996 -1155
rect 8964 -1205 8996 -1204
rect 8964 -1235 8965 -1205
rect 8965 -1235 8995 -1205
rect 8995 -1235 8996 -1205
rect 8964 -1236 8996 -1235
rect 8964 -1285 8996 -1284
rect 8964 -1315 8965 -1285
rect 8965 -1315 8995 -1285
rect 8995 -1315 8996 -1285
rect 8964 -1316 8996 -1315
rect 8964 -1365 8996 -1364
rect 8964 -1395 8965 -1365
rect 8965 -1395 8995 -1365
rect 8995 -1395 8996 -1365
rect 8964 -1396 8996 -1395
rect 8964 -1445 8996 -1444
rect 8964 -1475 8965 -1445
rect 8965 -1475 8995 -1445
rect 8995 -1475 8996 -1445
rect 8964 -1476 8996 -1475
rect 8964 -1525 8996 -1524
rect 8964 -1555 8965 -1525
rect 8965 -1555 8995 -1525
rect 8995 -1555 8996 -1525
rect 8964 -1556 8996 -1555
rect 8964 -1636 8996 -1604
rect 8964 -1716 8996 -1684
rect 8964 -1765 8996 -1764
rect 8964 -1795 8965 -1765
rect 8965 -1795 8995 -1765
rect 8995 -1795 8996 -1765
rect 8964 -1796 8996 -1795
rect 8964 -1845 8996 -1844
rect 8964 -1875 8965 -1845
rect 8965 -1875 8995 -1845
rect 8995 -1875 8996 -1845
rect 8964 -1876 8996 -1875
rect 8964 -1956 8996 -1924
rect 8964 -2005 8996 -2004
rect 8964 -2035 8965 -2005
rect 8965 -2035 8995 -2005
rect 8995 -2035 8996 -2005
rect 8964 -2036 8996 -2035
rect 8964 -2116 8996 -2084
rect 8964 -2165 8996 -2164
rect 8964 -2195 8965 -2165
rect 8965 -2195 8995 -2165
rect 8995 -2195 8996 -2165
rect 8964 -2196 8996 -2195
rect 8964 -2276 8996 -2244
rect 8964 -2325 8996 -2324
rect 8964 -2355 8965 -2325
rect 8965 -2355 8995 -2325
rect 8995 -2355 8996 -2325
rect 8964 -2356 8996 -2355
rect 8964 -2405 8996 -2404
rect 8964 -2435 8965 -2405
rect 8965 -2435 8995 -2405
rect 8995 -2435 8996 -2405
rect 8964 -2436 8996 -2435
rect 8964 -2485 8996 -2484
rect 8964 -2515 8965 -2485
rect 8965 -2515 8995 -2485
rect 8995 -2515 8996 -2485
rect 8964 -2516 8996 -2515
rect 8964 -2565 8996 -2564
rect 8964 -2595 8965 -2565
rect 8965 -2595 8995 -2565
rect 8995 -2595 8996 -2565
rect 8964 -2596 8996 -2595
rect 8964 -2645 8996 -2644
rect 8964 -2675 8965 -2645
rect 8965 -2675 8995 -2645
rect 8995 -2675 8996 -2645
rect 8964 -2676 8996 -2675
rect 8964 -2725 8996 -2724
rect 8964 -2755 8965 -2725
rect 8965 -2755 8995 -2725
rect 8995 -2755 8996 -2725
rect 8964 -2756 8996 -2755
rect 8964 -2836 8996 -2804
rect 8964 -2885 8996 -2884
rect 8964 -2915 8965 -2885
rect 8965 -2915 8995 -2885
rect 8995 -2915 8996 -2885
rect 8964 -2916 8996 -2915
rect 8964 -2996 8996 -2964
rect 8964 -3045 8996 -3044
rect 8964 -3075 8965 -3045
rect 8965 -3075 8995 -3045
rect 8995 -3075 8996 -3045
rect 8964 -3076 8996 -3075
rect 8964 -3156 8996 -3124
rect 8964 -3205 8996 -3204
rect 8964 -3235 8965 -3205
rect 8965 -3235 8995 -3205
rect 8995 -3235 8996 -3205
rect 8964 -3236 8996 -3235
rect 8964 -3285 8996 -3284
rect 8964 -3315 8965 -3285
rect 8965 -3315 8995 -3285
rect 8995 -3315 8996 -3285
rect 8964 -3316 8996 -3315
rect 8964 -3396 8996 -3364
rect 8964 -3476 8996 -3444
rect 8964 -3525 8996 -3524
rect 8964 -3555 8965 -3525
rect 8965 -3555 8995 -3525
rect 8995 -3555 8996 -3525
rect 8964 -3556 8996 -3555
rect 8964 -3605 8996 -3604
rect 8964 -3635 8965 -3605
rect 8965 -3635 8995 -3605
rect 8995 -3635 8996 -3605
rect 8964 -3636 8996 -3635
rect 8964 -3685 8996 -3684
rect 8964 -3715 8965 -3685
rect 8965 -3715 8995 -3685
rect 8995 -3715 8996 -3685
rect 8964 -3716 8996 -3715
rect 9044 1035 9076 1036
rect 9044 1005 9045 1035
rect 9045 1005 9075 1035
rect 9075 1005 9076 1035
rect 9044 1004 9076 1005
rect 9044 955 9076 956
rect 9044 925 9045 955
rect 9045 925 9075 955
rect 9075 925 9076 955
rect 9044 924 9076 925
rect 9044 875 9076 876
rect 9044 845 9045 875
rect 9045 845 9075 875
rect 9075 845 9076 875
rect 9044 844 9076 845
rect 9044 764 9076 796
rect 9044 684 9076 716
rect 9044 635 9076 636
rect 9044 605 9045 635
rect 9045 605 9075 635
rect 9075 605 9076 635
rect 9044 604 9076 605
rect 9044 555 9076 556
rect 9044 525 9045 555
rect 9045 525 9075 555
rect 9075 525 9076 555
rect 9044 524 9076 525
rect 9044 444 9076 476
rect 9044 395 9076 396
rect 9044 365 9045 395
rect 9045 365 9075 395
rect 9075 365 9076 395
rect 9044 364 9076 365
rect 9044 284 9076 316
rect 9044 235 9076 236
rect 9044 205 9045 235
rect 9045 205 9075 235
rect 9075 205 9076 235
rect 9044 204 9076 205
rect 9044 124 9076 156
rect 9044 75 9076 76
rect 9044 45 9045 75
rect 9045 45 9075 75
rect 9075 45 9076 75
rect 9044 44 9076 45
rect 9044 -5 9076 -4
rect 9044 -35 9045 -5
rect 9045 -35 9075 -5
rect 9075 -35 9076 -5
rect 9044 -36 9076 -35
rect 9044 -85 9076 -84
rect 9044 -115 9045 -85
rect 9045 -115 9075 -85
rect 9075 -115 9076 -85
rect 9044 -116 9076 -115
rect 9044 -165 9076 -164
rect 9044 -195 9045 -165
rect 9045 -195 9075 -165
rect 9075 -195 9076 -165
rect 9044 -196 9076 -195
rect 9044 -245 9076 -244
rect 9044 -275 9045 -245
rect 9045 -275 9075 -245
rect 9075 -275 9076 -245
rect 9044 -276 9076 -275
rect 9044 -325 9076 -324
rect 9044 -355 9045 -325
rect 9045 -355 9075 -325
rect 9075 -355 9076 -325
rect 9044 -356 9076 -355
rect 9044 -436 9076 -404
rect 9044 -485 9076 -484
rect 9044 -515 9045 -485
rect 9045 -515 9075 -485
rect 9075 -515 9076 -485
rect 9044 -516 9076 -515
rect 9044 -596 9076 -564
rect 9044 -645 9076 -644
rect 9044 -675 9045 -645
rect 9045 -675 9075 -645
rect 9075 -675 9076 -645
rect 9044 -676 9076 -675
rect 9044 -756 9076 -724
rect 9044 -805 9076 -804
rect 9044 -835 9045 -805
rect 9045 -835 9075 -805
rect 9075 -835 9076 -805
rect 9044 -836 9076 -835
rect 9044 -885 9076 -884
rect 9044 -915 9045 -885
rect 9045 -915 9075 -885
rect 9075 -915 9076 -885
rect 9044 -916 9076 -915
rect 9044 -996 9076 -964
rect 9044 -1076 9076 -1044
rect 9044 -1125 9076 -1124
rect 9044 -1155 9045 -1125
rect 9045 -1155 9075 -1125
rect 9075 -1155 9076 -1125
rect 9044 -1156 9076 -1155
rect 9044 -1205 9076 -1204
rect 9044 -1235 9045 -1205
rect 9045 -1235 9075 -1205
rect 9075 -1235 9076 -1205
rect 9044 -1236 9076 -1235
rect 9044 -1285 9076 -1284
rect 9044 -1315 9045 -1285
rect 9045 -1315 9075 -1285
rect 9075 -1315 9076 -1285
rect 9044 -1316 9076 -1315
rect 9044 -1365 9076 -1364
rect 9044 -1395 9045 -1365
rect 9045 -1395 9075 -1365
rect 9075 -1395 9076 -1365
rect 9044 -1396 9076 -1395
rect 9044 -1445 9076 -1444
rect 9044 -1475 9045 -1445
rect 9045 -1475 9075 -1445
rect 9075 -1475 9076 -1445
rect 9044 -1476 9076 -1475
rect 9044 -1525 9076 -1524
rect 9044 -1555 9045 -1525
rect 9045 -1555 9075 -1525
rect 9075 -1555 9076 -1525
rect 9044 -1556 9076 -1555
rect 9044 -1636 9076 -1604
rect 9044 -1716 9076 -1684
rect 9044 -1765 9076 -1764
rect 9044 -1795 9045 -1765
rect 9045 -1795 9075 -1765
rect 9075 -1795 9076 -1765
rect 9044 -1796 9076 -1795
rect 9044 -1845 9076 -1844
rect 9044 -1875 9045 -1845
rect 9045 -1875 9075 -1845
rect 9075 -1875 9076 -1845
rect 9044 -1876 9076 -1875
rect 9044 -1956 9076 -1924
rect 9044 -2005 9076 -2004
rect 9044 -2035 9045 -2005
rect 9045 -2035 9075 -2005
rect 9075 -2035 9076 -2005
rect 9044 -2036 9076 -2035
rect 9044 -2116 9076 -2084
rect 9044 -2165 9076 -2164
rect 9044 -2195 9045 -2165
rect 9045 -2195 9075 -2165
rect 9075 -2195 9076 -2165
rect 9044 -2196 9076 -2195
rect 9044 -2276 9076 -2244
rect 9044 -2325 9076 -2324
rect 9044 -2355 9045 -2325
rect 9045 -2355 9075 -2325
rect 9075 -2355 9076 -2325
rect 9044 -2356 9076 -2355
rect 9044 -2405 9076 -2404
rect 9044 -2435 9045 -2405
rect 9045 -2435 9075 -2405
rect 9075 -2435 9076 -2405
rect 9044 -2436 9076 -2435
rect 9044 -2485 9076 -2484
rect 9044 -2515 9045 -2485
rect 9045 -2515 9075 -2485
rect 9075 -2515 9076 -2485
rect 9044 -2516 9076 -2515
rect 9044 -2565 9076 -2564
rect 9044 -2595 9045 -2565
rect 9045 -2595 9075 -2565
rect 9075 -2595 9076 -2565
rect 9044 -2596 9076 -2595
rect 9044 -2645 9076 -2644
rect 9044 -2675 9045 -2645
rect 9045 -2675 9075 -2645
rect 9075 -2675 9076 -2645
rect 9044 -2676 9076 -2675
rect 9044 -2725 9076 -2724
rect 9044 -2755 9045 -2725
rect 9045 -2755 9075 -2725
rect 9075 -2755 9076 -2725
rect 9044 -2756 9076 -2755
rect 9044 -2836 9076 -2804
rect 9044 -2885 9076 -2884
rect 9044 -2915 9045 -2885
rect 9045 -2915 9075 -2885
rect 9075 -2915 9076 -2885
rect 9044 -2916 9076 -2915
rect 9044 -2996 9076 -2964
rect 9044 -3045 9076 -3044
rect 9044 -3075 9045 -3045
rect 9045 -3075 9075 -3045
rect 9075 -3075 9076 -3045
rect 9044 -3076 9076 -3075
rect 9044 -3156 9076 -3124
rect 9044 -3205 9076 -3204
rect 9044 -3235 9045 -3205
rect 9045 -3235 9075 -3205
rect 9075 -3235 9076 -3205
rect 9044 -3236 9076 -3235
rect 9044 -3285 9076 -3284
rect 9044 -3315 9045 -3285
rect 9045 -3315 9075 -3285
rect 9075 -3315 9076 -3285
rect 9044 -3316 9076 -3315
rect 9044 -3396 9076 -3364
rect 9044 -3476 9076 -3444
rect 9044 -3525 9076 -3524
rect 9044 -3555 9045 -3525
rect 9045 -3555 9075 -3525
rect 9075 -3555 9076 -3525
rect 9044 -3556 9076 -3555
rect 9044 -3605 9076 -3604
rect 9044 -3635 9045 -3605
rect 9045 -3635 9075 -3605
rect 9075 -3635 9076 -3605
rect 9044 -3636 9076 -3635
rect 9044 -3685 9076 -3684
rect 9044 -3715 9045 -3685
rect 9045 -3715 9075 -3685
rect 9075 -3715 9076 -3685
rect 9044 -3716 9076 -3715
rect 9124 1035 9156 1036
rect 9124 1005 9125 1035
rect 9125 1005 9155 1035
rect 9155 1005 9156 1035
rect 9124 1004 9156 1005
rect 9124 955 9156 956
rect 9124 925 9125 955
rect 9125 925 9155 955
rect 9155 925 9156 955
rect 9124 924 9156 925
rect 9124 875 9156 876
rect 9124 845 9125 875
rect 9125 845 9155 875
rect 9155 845 9156 875
rect 9124 844 9156 845
rect 9124 764 9156 796
rect 9124 684 9156 716
rect 9124 635 9156 636
rect 9124 605 9125 635
rect 9125 605 9155 635
rect 9155 605 9156 635
rect 9124 604 9156 605
rect 9124 555 9156 556
rect 9124 525 9125 555
rect 9125 525 9155 555
rect 9155 525 9156 555
rect 9124 524 9156 525
rect 9124 444 9156 476
rect 9124 395 9156 396
rect 9124 365 9125 395
rect 9125 365 9155 395
rect 9155 365 9156 395
rect 9124 364 9156 365
rect 9124 284 9156 316
rect 9124 235 9156 236
rect 9124 205 9125 235
rect 9125 205 9155 235
rect 9155 205 9156 235
rect 9124 204 9156 205
rect 9124 124 9156 156
rect 9124 75 9156 76
rect 9124 45 9125 75
rect 9125 45 9155 75
rect 9155 45 9156 75
rect 9124 44 9156 45
rect 9124 -5 9156 -4
rect 9124 -35 9125 -5
rect 9125 -35 9155 -5
rect 9155 -35 9156 -5
rect 9124 -36 9156 -35
rect 9124 -85 9156 -84
rect 9124 -115 9125 -85
rect 9125 -115 9155 -85
rect 9155 -115 9156 -85
rect 9124 -116 9156 -115
rect 9124 -165 9156 -164
rect 9124 -195 9125 -165
rect 9125 -195 9155 -165
rect 9155 -195 9156 -165
rect 9124 -196 9156 -195
rect 9124 -245 9156 -244
rect 9124 -275 9125 -245
rect 9125 -275 9155 -245
rect 9155 -275 9156 -245
rect 9124 -276 9156 -275
rect 9124 -325 9156 -324
rect 9124 -355 9125 -325
rect 9125 -355 9155 -325
rect 9155 -355 9156 -325
rect 9124 -356 9156 -355
rect 9124 -436 9156 -404
rect 9124 -485 9156 -484
rect 9124 -515 9125 -485
rect 9125 -515 9155 -485
rect 9155 -515 9156 -485
rect 9124 -516 9156 -515
rect 9124 -596 9156 -564
rect 9124 -645 9156 -644
rect 9124 -675 9125 -645
rect 9125 -675 9155 -645
rect 9155 -675 9156 -645
rect 9124 -676 9156 -675
rect 9124 -756 9156 -724
rect 9124 -805 9156 -804
rect 9124 -835 9125 -805
rect 9125 -835 9155 -805
rect 9155 -835 9156 -805
rect 9124 -836 9156 -835
rect 9124 -885 9156 -884
rect 9124 -915 9125 -885
rect 9125 -915 9155 -885
rect 9155 -915 9156 -885
rect 9124 -916 9156 -915
rect 9124 -996 9156 -964
rect 9124 -1076 9156 -1044
rect 9124 -1125 9156 -1124
rect 9124 -1155 9125 -1125
rect 9125 -1155 9155 -1125
rect 9155 -1155 9156 -1125
rect 9124 -1156 9156 -1155
rect 9124 -1205 9156 -1204
rect 9124 -1235 9125 -1205
rect 9125 -1235 9155 -1205
rect 9155 -1235 9156 -1205
rect 9124 -1236 9156 -1235
rect 9124 -1285 9156 -1284
rect 9124 -1315 9125 -1285
rect 9125 -1315 9155 -1285
rect 9155 -1315 9156 -1285
rect 9124 -1316 9156 -1315
rect 9124 -1365 9156 -1364
rect 9124 -1395 9125 -1365
rect 9125 -1395 9155 -1365
rect 9155 -1395 9156 -1365
rect 9124 -1396 9156 -1395
rect 9124 -1445 9156 -1444
rect 9124 -1475 9125 -1445
rect 9125 -1475 9155 -1445
rect 9155 -1475 9156 -1445
rect 9124 -1476 9156 -1475
rect 9124 -1525 9156 -1524
rect 9124 -1555 9125 -1525
rect 9125 -1555 9155 -1525
rect 9155 -1555 9156 -1525
rect 9124 -1556 9156 -1555
rect 9124 -1636 9156 -1604
rect 9124 -1716 9156 -1684
rect 9124 -1765 9156 -1764
rect 9124 -1795 9125 -1765
rect 9125 -1795 9155 -1765
rect 9155 -1795 9156 -1765
rect 9124 -1796 9156 -1795
rect 9124 -1845 9156 -1844
rect 9124 -1875 9125 -1845
rect 9125 -1875 9155 -1845
rect 9155 -1875 9156 -1845
rect 9124 -1876 9156 -1875
rect 9124 -1956 9156 -1924
rect 9124 -2005 9156 -2004
rect 9124 -2035 9125 -2005
rect 9125 -2035 9155 -2005
rect 9155 -2035 9156 -2005
rect 9124 -2036 9156 -2035
rect 9124 -2116 9156 -2084
rect 9124 -2165 9156 -2164
rect 9124 -2195 9125 -2165
rect 9125 -2195 9155 -2165
rect 9155 -2195 9156 -2165
rect 9124 -2196 9156 -2195
rect 9124 -2276 9156 -2244
rect 9124 -2325 9156 -2324
rect 9124 -2355 9125 -2325
rect 9125 -2355 9155 -2325
rect 9155 -2355 9156 -2325
rect 9124 -2356 9156 -2355
rect 9124 -2405 9156 -2404
rect 9124 -2435 9125 -2405
rect 9125 -2435 9155 -2405
rect 9155 -2435 9156 -2405
rect 9124 -2436 9156 -2435
rect 9124 -2485 9156 -2484
rect 9124 -2515 9125 -2485
rect 9125 -2515 9155 -2485
rect 9155 -2515 9156 -2485
rect 9124 -2516 9156 -2515
rect 9124 -2565 9156 -2564
rect 9124 -2595 9125 -2565
rect 9125 -2595 9155 -2565
rect 9155 -2595 9156 -2565
rect 9124 -2596 9156 -2595
rect 9124 -2645 9156 -2644
rect 9124 -2675 9125 -2645
rect 9125 -2675 9155 -2645
rect 9155 -2675 9156 -2645
rect 9124 -2676 9156 -2675
rect 9124 -2725 9156 -2724
rect 9124 -2755 9125 -2725
rect 9125 -2755 9155 -2725
rect 9155 -2755 9156 -2725
rect 9124 -2756 9156 -2755
rect 9124 -2836 9156 -2804
rect 9124 -2885 9156 -2884
rect 9124 -2915 9125 -2885
rect 9125 -2915 9155 -2885
rect 9155 -2915 9156 -2885
rect 9124 -2916 9156 -2915
rect 9124 -2996 9156 -2964
rect 9124 -3045 9156 -3044
rect 9124 -3075 9125 -3045
rect 9125 -3075 9155 -3045
rect 9155 -3075 9156 -3045
rect 9124 -3076 9156 -3075
rect 9124 -3156 9156 -3124
rect 9124 -3205 9156 -3204
rect 9124 -3235 9125 -3205
rect 9125 -3235 9155 -3205
rect 9155 -3235 9156 -3205
rect 9124 -3236 9156 -3235
rect 9124 -3285 9156 -3284
rect 9124 -3315 9125 -3285
rect 9125 -3315 9155 -3285
rect 9155 -3315 9156 -3285
rect 9124 -3316 9156 -3315
rect 9124 -3396 9156 -3364
rect 9124 -3476 9156 -3444
rect 9124 -3525 9156 -3524
rect 9124 -3555 9125 -3525
rect 9125 -3555 9155 -3525
rect 9155 -3555 9156 -3525
rect 9124 -3556 9156 -3555
rect 9124 -3605 9156 -3604
rect 9124 -3635 9125 -3605
rect 9125 -3635 9155 -3605
rect 9155 -3635 9156 -3605
rect 9124 -3636 9156 -3635
rect 9124 -3685 9156 -3684
rect 9124 -3715 9125 -3685
rect 9125 -3715 9155 -3685
rect 9155 -3715 9156 -3685
rect 9124 -3716 9156 -3715
rect 9204 1035 9236 1036
rect 9204 1005 9205 1035
rect 9205 1005 9235 1035
rect 9235 1005 9236 1035
rect 9204 1004 9236 1005
rect 9204 955 9236 956
rect 9204 925 9205 955
rect 9205 925 9235 955
rect 9235 925 9236 955
rect 9204 924 9236 925
rect 9204 875 9236 876
rect 9204 845 9205 875
rect 9205 845 9235 875
rect 9235 845 9236 875
rect 9204 844 9236 845
rect 9204 764 9236 796
rect 9204 684 9236 716
rect 9204 635 9236 636
rect 9204 605 9205 635
rect 9205 605 9235 635
rect 9235 605 9236 635
rect 9204 604 9236 605
rect 9204 555 9236 556
rect 9204 525 9205 555
rect 9205 525 9235 555
rect 9235 525 9236 555
rect 9204 524 9236 525
rect 9204 444 9236 476
rect 9204 395 9236 396
rect 9204 365 9205 395
rect 9205 365 9235 395
rect 9235 365 9236 395
rect 9204 364 9236 365
rect 9204 284 9236 316
rect 9204 235 9236 236
rect 9204 205 9205 235
rect 9205 205 9235 235
rect 9235 205 9236 235
rect 9204 204 9236 205
rect 9204 124 9236 156
rect 9204 75 9236 76
rect 9204 45 9205 75
rect 9205 45 9235 75
rect 9235 45 9236 75
rect 9204 44 9236 45
rect 9204 -5 9236 -4
rect 9204 -35 9205 -5
rect 9205 -35 9235 -5
rect 9235 -35 9236 -5
rect 9204 -36 9236 -35
rect 9204 -85 9236 -84
rect 9204 -115 9205 -85
rect 9205 -115 9235 -85
rect 9235 -115 9236 -85
rect 9204 -116 9236 -115
rect 9204 -165 9236 -164
rect 9204 -195 9205 -165
rect 9205 -195 9235 -165
rect 9235 -195 9236 -165
rect 9204 -196 9236 -195
rect 9204 -245 9236 -244
rect 9204 -275 9205 -245
rect 9205 -275 9235 -245
rect 9235 -275 9236 -245
rect 9204 -276 9236 -275
rect 9204 -325 9236 -324
rect 9204 -355 9205 -325
rect 9205 -355 9235 -325
rect 9235 -355 9236 -325
rect 9204 -356 9236 -355
rect 9204 -436 9236 -404
rect 9204 -485 9236 -484
rect 9204 -515 9205 -485
rect 9205 -515 9235 -485
rect 9235 -515 9236 -485
rect 9204 -516 9236 -515
rect 9204 -596 9236 -564
rect 9204 -645 9236 -644
rect 9204 -675 9205 -645
rect 9205 -675 9235 -645
rect 9235 -675 9236 -645
rect 9204 -676 9236 -675
rect 9204 -756 9236 -724
rect 9204 -805 9236 -804
rect 9204 -835 9205 -805
rect 9205 -835 9235 -805
rect 9235 -835 9236 -805
rect 9204 -836 9236 -835
rect 9204 -885 9236 -884
rect 9204 -915 9205 -885
rect 9205 -915 9235 -885
rect 9235 -915 9236 -885
rect 9204 -916 9236 -915
rect 9204 -996 9236 -964
rect 9204 -1076 9236 -1044
rect 9204 -1125 9236 -1124
rect 9204 -1155 9205 -1125
rect 9205 -1155 9235 -1125
rect 9235 -1155 9236 -1125
rect 9204 -1156 9236 -1155
rect 9204 -1205 9236 -1204
rect 9204 -1235 9205 -1205
rect 9205 -1235 9235 -1205
rect 9235 -1235 9236 -1205
rect 9204 -1236 9236 -1235
rect 9204 -1285 9236 -1284
rect 9204 -1315 9205 -1285
rect 9205 -1315 9235 -1285
rect 9235 -1315 9236 -1285
rect 9204 -1316 9236 -1315
rect 9204 -1365 9236 -1364
rect 9204 -1395 9205 -1365
rect 9205 -1395 9235 -1365
rect 9235 -1395 9236 -1365
rect 9204 -1396 9236 -1395
rect 9204 -1445 9236 -1444
rect 9204 -1475 9205 -1445
rect 9205 -1475 9235 -1445
rect 9235 -1475 9236 -1445
rect 9204 -1476 9236 -1475
rect 9204 -1525 9236 -1524
rect 9204 -1555 9205 -1525
rect 9205 -1555 9235 -1525
rect 9235 -1555 9236 -1525
rect 9204 -1556 9236 -1555
rect 9204 -1636 9236 -1604
rect 9204 -1716 9236 -1684
rect 9204 -1765 9236 -1764
rect 9204 -1795 9205 -1765
rect 9205 -1795 9235 -1765
rect 9235 -1795 9236 -1765
rect 9204 -1796 9236 -1795
rect 9204 -1845 9236 -1844
rect 9204 -1875 9205 -1845
rect 9205 -1875 9235 -1845
rect 9235 -1875 9236 -1845
rect 9204 -1876 9236 -1875
rect 9204 -1956 9236 -1924
rect 9204 -2005 9236 -2004
rect 9204 -2035 9205 -2005
rect 9205 -2035 9235 -2005
rect 9235 -2035 9236 -2005
rect 9204 -2036 9236 -2035
rect 9204 -2116 9236 -2084
rect 9204 -2165 9236 -2164
rect 9204 -2195 9205 -2165
rect 9205 -2195 9235 -2165
rect 9235 -2195 9236 -2165
rect 9204 -2196 9236 -2195
rect 9204 -2276 9236 -2244
rect 9204 -2325 9236 -2324
rect 9204 -2355 9205 -2325
rect 9205 -2355 9235 -2325
rect 9235 -2355 9236 -2325
rect 9204 -2356 9236 -2355
rect 9204 -2405 9236 -2404
rect 9204 -2435 9205 -2405
rect 9205 -2435 9235 -2405
rect 9235 -2435 9236 -2405
rect 9204 -2436 9236 -2435
rect 9204 -2485 9236 -2484
rect 9204 -2515 9205 -2485
rect 9205 -2515 9235 -2485
rect 9235 -2515 9236 -2485
rect 9204 -2516 9236 -2515
rect 9204 -2565 9236 -2564
rect 9204 -2595 9205 -2565
rect 9205 -2595 9235 -2565
rect 9235 -2595 9236 -2565
rect 9204 -2596 9236 -2595
rect 9204 -2645 9236 -2644
rect 9204 -2675 9205 -2645
rect 9205 -2675 9235 -2645
rect 9235 -2675 9236 -2645
rect 9204 -2676 9236 -2675
rect 9204 -2725 9236 -2724
rect 9204 -2755 9205 -2725
rect 9205 -2755 9235 -2725
rect 9235 -2755 9236 -2725
rect 9204 -2756 9236 -2755
rect 9204 -2836 9236 -2804
rect 9204 -2885 9236 -2884
rect 9204 -2915 9205 -2885
rect 9205 -2915 9235 -2885
rect 9235 -2915 9236 -2885
rect 9204 -2916 9236 -2915
rect 9204 -2996 9236 -2964
rect 9204 -3045 9236 -3044
rect 9204 -3075 9205 -3045
rect 9205 -3075 9235 -3045
rect 9235 -3075 9236 -3045
rect 9204 -3076 9236 -3075
rect 9204 -3156 9236 -3124
rect 9204 -3205 9236 -3204
rect 9204 -3235 9205 -3205
rect 9205 -3235 9235 -3205
rect 9235 -3235 9236 -3205
rect 9204 -3236 9236 -3235
rect 9204 -3285 9236 -3284
rect 9204 -3315 9205 -3285
rect 9205 -3315 9235 -3285
rect 9235 -3315 9236 -3285
rect 9204 -3316 9236 -3315
rect 9204 -3396 9236 -3364
rect 9204 -3476 9236 -3444
rect 9204 -3525 9236 -3524
rect 9204 -3555 9205 -3525
rect 9205 -3555 9235 -3525
rect 9235 -3555 9236 -3525
rect 9204 -3556 9236 -3555
rect 9204 -3605 9236 -3604
rect 9204 -3635 9205 -3605
rect 9205 -3635 9235 -3605
rect 9235 -3635 9236 -3605
rect 9204 -3636 9236 -3635
rect 9204 -3685 9236 -3684
rect 9204 -3715 9205 -3685
rect 9205 -3715 9235 -3685
rect 9235 -3715 9236 -3685
rect 9204 -3716 9236 -3715
rect 9284 1035 9316 1036
rect 9284 1005 9285 1035
rect 9285 1005 9315 1035
rect 9315 1005 9316 1035
rect 9284 1004 9316 1005
rect 9284 955 9316 956
rect 9284 925 9285 955
rect 9285 925 9315 955
rect 9315 925 9316 955
rect 9284 924 9316 925
rect 9284 875 9316 876
rect 9284 845 9285 875
rect 9285 845 9315 875
rect 9315 845 9316 875
rect 9284 844 9316 845
rect 9284 764 9316 796
rect 9284 684 9316 716
rect 9284 635 9316 636
rect 9284 605 9285 635
rect 9285 605 9315 635
rect 9315 605 9316 635
rect 9284 604 9316 605
rect 9284 555 9316 556
rect 9284 525 9285 555
rect 9285 525 9315 555
rect 9315 525 9316 555
rect 9284 524 9316 525
rect 9284 444 9316 476
rect 9284 395 9316 396
rect 9284 365 9285 395
rect 9285 365 9315 395
rect 9315 365 9316 395
rect 9284 364 9316 365
rect 9284 284 9316 316
rect 9284 235 9316 236
rect 9284 205 9285 235
rect 9285 205 9315 235
rect 9315 205 9316 235
rect 9284 204 9316 205
rect 9284 124 9316 156
rect 9284 75 9316 76
rect 9284 45 9285 75
rect 9285 45 9315 75
rect 9315 45 9316 75
rect 9284 44 9316 45
rect 9284 -5 9316 -4
rect 9284 -35 9285 -5
rect 9285 -35 9315 -5
rect 9315 -35 9316 -5
rect 9284 -36 9316 -35
rect 9284 -85 9316 -84
rect 9284 -115 9285 -85
rect 9285 -115 9315 -85
rect 9315 -115 9316 -85
rect 9284 -116 9316 -115
rect 9284 -165 9316 -164
rect 9284 -195 9285 -165
rect 9285 -195 9315 -165
rect 9315 -195 9316 -165
rect 9284 -196 9316 -195
rect 9284 -245 9316 -244
rect 9284 -275 9285 -245
rect 9285 -275 9315 -245
rect 9315 -275 9316 -245
rect 9284 -276 9316 -275
rect 9284 -325 9316 -324
rect 9284 -355 9285 -325
rect 9285 -355 9315 -325
rect 9315 -355 9316 -325
rect 9284 -356 9316 -355
rect 9284 -436 9316 -404
rect 9284 -485 9316 -484
rect 9284 -515 9285 -485
rect 9285 -515 9315 -485
rect 9315 -515 9316 -485
rect 9284 -516 9316 -515
rect 9284 -596 9316 -564
rect 9284 -645 9316 -644
rect 9284 -675 9285 -645
rect 9285 -675 9315 -645
rect 9315 -675 9316 -645
rect 9284 -676 9316 -675
rect 9284 -756 9316 -724
rect 9284 -805 9316 -804
rect 9284 -835 9285 -805
rect 9285 -835 9315 -805
rect 9315 -835 9316 -805
rect 9284 -836 9316 -835
rect 9284 -885 9316 -884
rect 9284 -915 9285 -885
rect 9285 -915 9315 -885
rect 9315 -915 9316 -885
rect 9284 -916 9316 -915
rect 9284 -996 9316 -964
rect 9284 -1076 9316 -1044
rect 9284 -1125 9316 -1124
rect 9284 -1155 9285 -1125
rect 9285 -1155 9315 -1125
rect 9315 -1155 9316 -1125
rect 9284 -1156 9316 -1155
rect 9284 -1205 9316 -1204
rect 9284 -1235 9285 -1205
rect 9285 -1235 9315 -1205
rect 9315 -1235 9316 -1205
rect 9284 -1236 9316 -1235
rect 9284 -1285 9316 -1284
rect 9284 -1315 9285 -1285
rect 9285 -1315 9315 -1285
rect 9315 -1315 9316 -1285
rect 9284 -1316 9316 -1315
rect 9284 -1365 9316 -1364
rect 9284 -1395 9285 -1365
rect 9285 -1395 9315 -1365
rect 9315 -1395 9316 -1365
rect 9284 -1396 9316 -1395
rect 9284 -1445 9316 -1444
rect 9284 -1475 9285 -1445
rect 9285 -1475 9315 -1445
rect 9315 -1475 9316 -1445
rect 9284 -1476 9316 -1475
rect 9284 -1525 9316 -1524
rect 9284 -1555 9285 -1525
rect 9285 -1555 9315 -1525
rect 9315 -1555 9316 -1525
rect 9284 -1556 9316 -1555
rect 9284 -1636 9316 -1604
rect 9284 -1716 9316 -1684
rect 9284 -1765 9316 -1764
rect 9284 -1795 9285 -1765
rect 9285 -1795 9315 -1765
rect 9315 -1795 9316 -1765
rect 9284 -1796 9316 -1795
rect 9284 -1845 9316 -1844
rect 9284 -1875 9285 -1845
rect 9285 -1875 9315 -1845
rect 9315 -1875 9316 -1845
rect 9284 -1876 9316 -1875
rect 9284 -1956 9316 -1924
rect 9284 -2005 9316 -2004
rect 9284 -2035 9285 -2005
rect 9285 -2035 9315 -2005
rect 9315 -2035 9316 -2005
rect 9284 -2036 9316 -2035
rect 9284 -2116 9316 -2084
rect 9284 -2165 9316 -2164
rect 9284 -2195 9285 -2165
rect 9285 -2195 9315 -2165
rect 9315 -2195 9316 -2165
rect 9284 -2196 9316 -2195
rect 9284 -2276 9316 -2244
rect 9284 -2325 9316 -2324
rect 9284 -2355 9285 -2325
rect 9285 -2355 9315 -2325
rect 9315 -2355 9316 -2325
rect 9284 -2356 9316 -2355
rect 9284 -2405 9316 -2404
rect 9284 -2435 9285 -2405
rect 9285 -2435 9315 -2405
rect 9315 -2435 9316 -2405
rect 9284 -2436 9316 -2435
rect 9284 -2485 9316 -2484
rect 9284 -2515 9285 -2485
rect 9285 -2515 9315 -2485
rect 9315 -2515 9316 -2485
rect 9284 -2516 9316 -2515
rect 9284 -2565 9316 -2564
rect 9284 -2595 9285 -2565
rect 9285 -2595 9315 -2565
rect 9315 -2595 9316 -2565
rect 9284 -2596 9316 -2595
rect 9284 -2645 9316 -2644
rect 9284 -2675 9285 -2645
rect 9285 -2675 9315 -2645
rect 9315 -2675 9316 -2645
rect 9284 -2676 9316 -2675
rect 9284 -2725 9316 -2724
rect 9284 -2755 9285 -2725
rect 9285 -2755 9315 -2725
rect 9315 -2755 9316 -2725
rect 9284 -2756 9316 -2755
rect 9284 -2836 9316 -2804
rect 9284 -2885 9316 -2884
rect 9284 -2915 9285 -2885
rect 9285 -2915 9315 -2885
rect 9315 -2915 9316 -2885
rect 9284 -2916 9316 -2915
rect 9284 -2996 9316 -2964
rect 9284 -3045 9316 -3044
rect 9284 -3075 9285 -3045
rect 9285 -3075 9315 -3045
rect 9315 -3075 9316 -3045
rect 9284 -3076 9316 -3075
rect 9284 -3156 9316 -3124
rect 9284 -3205 9316 -3204
rect 9284 -3235 9285 -3205
rect 9285 -3235 9315 -3205
rect 9315 -3235 9316 -3205
rect 9284 -3236 9316 -3235
rect 9284 -3285 9316 -3284
rect 9284 -3315 9285 -3285
rect 9285 -3315 9315 -3285
rect 9315 -3315 9316 -3285
rect 9284 -3316 9316 -3315
rect 9284 -3396 9316 -3364
rect 9284 -3476 9316 -3444
rect 9284 -3525 9316 -3524
rect 9284 -3555 9285 -3525
rect 9285 -3555 9315 -3525
rect 9315 -3555 9316 -3525
rect 9284 -3556 9316 -3555
rect 9284 -3605 9316 -3604
rect 9284 -3635 9285 -3605
rect 9285 -3635 9315 -3605
rect 9315 -3635 9316 -3605
rect 9284 -3636 9316 -3635
rect 9284 -3685 9316 -3684
rect 9284 -3715 9285 -3685
rect 9285 -3715 9315 -3685
rect 9315 -3715 9316 -3685
rect 9284 -3716 9316 -3715
rect 9364 1035 9396 1036
rect 9364 1005 9365 1035
rect 9365 1005 9395 1035
rect 9395 1005 9396 1035
rect 9364 1004 9396 1005
rect 9364 955 9396 956
rect 9364 925 9365 955
rect 9365 925 9395 955
rect 9395 925 9396 955
rect 9364 924 9396 925
rect 9364 875 9396 876
rect 9364 845 9365 875
rect 9365 845 9395 875
rect 9395 845 9396 875
rect 9364 844 9396 845
rect 9364 764 9396 796
rect 9364 684 9396 716
rect 9364 635 9396 636
rect 9364 605 9365 635
rect 9365 605 9395 635
rect 9395 605 9396 635
rect 9364 604 9396 605
rect 9364 555 9396 556
rect 9364 525 9365 555
rect 9365 525 9395 555
rect 9395 525 9396 555
rect 9364 524 9396 525
rect 9364 444 9396 476
rect 9364 395 9396 396
rect 9364 365 9365 395
rect 9365 365 9395 395
rect 9395 365 9396 395
rect 9364 364 9396 365
rect 9364 284 9396 316
rect 9364 235 9396 236
rect 9364 205 9365 235
rect 9365 205 9395 235
rect 9395 205 9396 235
rect 9364 204 9396 205
rect 9364 124 9396 156
rect 9364 75 9396 76
rect 9364 45 9365 75
rect 9365 45 9395 75
rect 9395 45 9396 75
rect 9364 44 9396 45
rect 9364 -5 9396 -4
rect 9364 -35 9365 -5
rect 9365 -35 9395 -5
rect 9395 -35 9396 -5
rect 9364 -36 9396 -35
rect 9364 -85 9396 -84
rect 9364 -115 9365 -85
rect 9365 -115 9395 -85
rect 9395 -115 9396 -85
rect 9364 -116 9396 -115
rect 9364 -165 9396 -164
rect 9364 -195 9365 -165
rect 9365 -195 9395 -165
rect 9395 -195 9396 -165
rect 9364 -196 9396 -195
rect 9364 -245 9396 -244
rect 9364 -275 9365 -245
rect 9365 -275 9395 -245
rect 9395 -275 9396 -245
rect 9364 -276 9396 -275
rect 9364 -325 9396 -324
rect 9364 -355 9365 -325
rect 9365 -355 9395 -325
rect 9395 -355 9396 -325
rect 9364 -356 9396 -355
rect 9364 -436 9396 -404
rect 9364 -485 9396 -484
rect 9364 -515 9365 -485
rect 9365 -515 9395 -485
rect 9395 -515 9396 -485
rect 9364 -516 9396 -515
rect 9364 -596 9396 -564
rect 9364 -645 9396 -644
rect 9364 -675 9365 -645
rect 9365 -675 9395 -645
rect 9395 -675 9396 -645
rect 9364 -676 9396 -675
rect 9364 -756 9396 -724
rect 9364 -805 9396 -804
rect 9364 -835 9365 -805
rect 9365 -835 9395 -805
rect 9395 -835 9396 -805
rect 9364 -836 9396 -835
rect 9364 -885 9396 -884
rect 9364 -915 9365 -885
rect 9365 -915 9395 -885
rect 9395 -915 9396 -885
rect 9364 -916 9396 -915
rect 9364 -996 9396 -964
rect 9364 -1076 9396 -1044
rect 9364 -1125 9396 -1124
rect 9364 -1155 9365 -1125
rect 9365 -1155 9395 -1125
rect 9395 -1155 9396 -1125
rect 9364 -1156 9396 -1155
rect 9364 -1205 9396 -1204
rect 9364 -1235 9365 -1205
rect 9365 -1235 9395 -1205
rect 9395 -1235 9396 -1205
rect 9364 -1236 9396 -1235
rect 9364 -1285 9396 -1284
rect 9364 -1315 9365 -1285
rect 9365 -1315 9395 -1285
rect 9395 -1315 9396 -1285
rect 9364 -1316 9396 -1315
rect 9364 -1365 9396 -1364
rect 9364 -1395 9365 -1365
rect 9365 -1395 9395 -1365
rect 9395 -1395 9396 -1365
rect 9364 -1396 9396 -1395
rect 9364 -1445 9396 -1444
rect 9364 -1475 9365 -1445
rect 9365 -1475 9395 -1445
rect 9395 -1475 9396 -1445
rect 9364 -1476 9396 -1475
rect 9364 -1525 9396 -1524
rect 9364 -1555 9365 -1525
rect 9365 -1555 9395 -1525
rect 9395 -1555 9396 -1525
rect 9364 -1556 9396 -1555
rect 9364 -1636 9396 -1604
rect 9364 -1716 9396 -1684
rect 9364 -1765 9396 -1764
rect 9364 -1795 9365 -1765
rect 9365 -1795 9395 -1765
rect 9395 -1795 9396 -1765
rect 9364 -1796 9396 -1795
rect 9364 -1845 9396 -1844
rect 9364 -1875 9365 -1845
rect 9365 -1875 9395 -1845
rect 9395 -1875 9396 -1845
rect 9364 -1876 9396 -1875
rect 9364 -1956 9396 -1924
rect 9364 -2005 9396 -2004
rect 9364 -2035 9365 -2005
rect 9365 -2035 9395 -2005
rect 9395 -2035 9396 -2005
rect 9364 -2036 9396 -2035
rect 9364 -2116 9396 -2084
rect 9364 -2165 9396 -2164
rect 9364 -2195 9365 -2165
rect 9365 -2195 9395 -2165
rect 9395 -2195 9396 -2165
rect 9364 -2196 9396 -2195
rect 9364 -2276 9396 -2244
rect 9364 -2325 9396 -2324
rect 9364 -2355 9365 -2325
rect 9365 -2355 9395 -2325
rect 9395 -2355 9396 -2325
rect 9364 -2356 9396 -2355
rect 9364 -2405 9396 -2404
rect 9364 -2435 9365 -2405
rect 9365 -2435 9395 -2405
rect 9395 -2435 9396 -2405
rect 9364 -2436 9396 -2435
rect 9364 -2485 9396 -2484
rect 9364 -2515 9365 -2485
rect 9365 -2515 9395 -2485
rect 9395 -2515 9396 -2485
rect 9364 -2516 9396 -2515
rect 9364 -2565 9396 -2564
rect 9364 -2595 9365 -2565
rect 9365 -2595 9395 -2565
rect 9395 -2595 9396 -2565
rect 9364 -2596 9396 -2595
rect 9364 -2645 9396 -2644
rect 9364 -2675 9365 -2645
rect 9365 -2675 9395 -2645
rect 9395 -2675 9396 -2645
rect 9364 -2676 9396 -2675
rect 9364 -2725 9396 -2724
rect 9364 -2755 9365 -2725
rect 9365 -2755 9395 -2725
rect 9395 -2755 9396 -2725
rect 9364 -2756 9396 -2755
rect 9364 -2836 9396 -2804
rect 9364 -2885 9396 -2884
rect 9364 -2915 9365 -2885
rect 9365 -2915 9395 -2885
rect 9395 -2915 9396 -2885
rect 9364 -2916 9396 -2915
rect 9364 -2996 9396 -2964
rect 9364 -3045 9396 -3044
rect 9364 -3075 9365 -3045
rect 9365 -3075 9395 -3045
rect 9395 -3075 9396 -3045
rect 9364 -3076 9396 -3075
rect 9364 -3156 9396 -3124
rect 9364 -3205 9396 -3204
rect 9364 -3235 9365 -3205
rect 9365 -3235 9395 -3205
rect 9395 -3235 9396 -3205
rect 9364 -3236 9396 -3235
rect 9364 -3285 9396 -3284
rect 9364 -3315 9365 -3285
rect 9365 -3315 9395 -3285
rect 9395 -3315 9396 -3285
rect 9364 -3316 9396 -3315
rect 9364 -3396 9396 -3364
rect 9364 -3476 9396 -3444
rect 9364 -3525 9396 -3524
rect 9364 -3555 9365 -3525
rect 9365 -3555 9395 -3525
rect 9395 -3555 9396 -3525
rect 9364 -3556 9396 -3555
rect 9364 -3605 9396 -3604
rect 9364 -3635 9365 -3605
rect 9365 -3635 9395 -3605
rect 9395 -3635 9396 -3605
rect 9364 -3636 9396 -3635
rect 9364 -3685 9396 -3684
rect 9364 -3715 9365 -3685
rect 9365 -3715 9395 -3685
rect 9395 -3715 9396 -3685
rect 9364 -3716 9396 -3715
rect 9444 1035 9476 1036
rect 9444 1005 9445 1035
rect 9445 1005 9475 1035
rect 9475 1005 9476 1035
rect 9444 1004 9476 1005
rect 9444 955 9476 956
rect 9444 925 9445 955
rect 9445 925 9475 955
rect 9475 925 9476 955
rect 9444 924 9476 925
rect 9444 875 9476 876
rect 9444 845 9445 875
rect 9445 845 9475 875
rect 9475 845 9476 875
rect 9444 844 9476 845
rect 9444 764 9476 796
rect 9444 684 9476 716
rect 9444 635 9476 636
rect 9444 605 9445 635
rect 9445 605 9475 635
rect 9475 605 9476 635
rect 9444 604 9476 605
rect 9444 555 9476 556
rect 9444 525 9445 555
rect 9445 525 9475 555
rect 9475 525 9476 555
rect 9444 524 9476 525
rect 9444 444 9476 476
rect 9444 395 9476 396
rect 9444 365 9445 395
rect 9445 365 9475 395
rect 9475 365 9476 395
rect 9444 364 9476 365
rect 9444 284 9476 316
rect 9444 235 9476 236
rect 9444 205 9445 235
rect 9445 205 9475 235
rect 9475 205 9476 235
rect 9444 204 9476 205
rect 9444 124 9476 156
rect 9444 75 9476 76
rect 9444 45 9445 75
rect 9445 45 9475 75
rect 9475 45 9476 75
rect 9444 44 9476 45
rect 9444 -5 9476 -4
rect 9444 -35 9445 -5
rect 9445 -35 9475 -5
rect 9475 -35 9476 -5
rect 9444 -36 9476 -35
rect 9444 -85 9476 -84
rect 9444 -115 9445 -85
rect 9445 -115 9475 -85
rect 9475 -115 9476 -85
rect 9444 -116 9476 -115
rect 9444 -165 9476 -164
rect 9444 -195 9445 -165
rect 9445 -195 9475 -165
rect 9475 -195 9476 -165
rect 9444 -196 9476 -195
rect 9444 -245 9476 -244
rect 9444 -275 9445 -245
rect 9445 -275 9475 -245
rect 9475 -275 9476 -245
rect 9444 -276 9476 -275
rect 9444 -325 9476 -324
rect 9444 -355 9445 -325
rect 9445 -355 9475 -325
rect 9475 -355 9476 -325
rect 9444 -356 9476 -355
rect 9444 -436 9476 -404
rect 9444 -485 9476 -484
rect 9444 -515 9445 -485
rect 9445 -515 9475 -485
rect 9475 -515 9476 -485
rect 9444 -516 9476 -515
rect 9444 -596 9476 -564
rect 9444 -645 9476 -644
rect 9444 -675 9445 -645
rect 9445 -675 9475 -645
rect 9475 -675 9476 -645
rect 9444 -676 9476 -675
rect 9444 -756 9476 -724
rect 9444 -805 9476 -804
rect 9444 -835 9445 -805
rect 9445 -835 9475 -805
rect 9475 -835 9476 -805
rect 9444 -836 9476 -835
rect 9444 -885 9476 -884
rect 9444 -915 9445 -885
rect 9445 -915 9475 -885
rect 9475 -915 9476 -885
rect 9444 -916 9476 -915
rect 9444 -996 9476 -964
rect 9444 -1076 9476 -1044
rect 9444 -1125 9476 -1124
rect 9444 -1155 9445 -1125
rect 9445 -1155 9475 -1125
rect 9475 -1155 9476 -1125
rect 9444 -1156 9476 -1155
rect 9444 -1205 9476 -1204
rect 9444 -1235 9445 -1205
rect 9445 -1235 9475 -1205
rect 9475 -1235 9476 -1205
rect 9444 -1236 9476 -1235
rect 9444 -1285 9476 -1284
rect 9444 -1315 9445 -1285
rect 9445 -1315 9475 -1285
rect 9475 -1315 9476 -1285
rect 9444 -1316 9476 -1315
rect 9444 -1365 9476 -1364
rect 9444 -1395 9445 -1365
rect 9445 -1395 9475 -1365
rect 9475 -1395 9476 -1365
rect 9444 -1396 9476 -1395
rect 9444 -1445 9476 -1444
rect 9444 -1475 9445 -1445
rect 9445 -1475 9475 -1445
rect 9475 -1475 9476 -1445
rect 9444 -1476 9476 -1475
rect 9444 -1525 9476 -1524
rect 9444 -1555 9445 -1525
rect 9445 -1555 9475 -1525
rect 9475 -1555 9476 -1525
rect 9444 -1556 9476 -1555
rect 9444 -1636 9476 -1604
rect 9444 -1716 9476 -1684
rect 9444 -1765 9476 -1764
rect 9444 -1795 9445 -1765
rect 9445 -1795 9475 -1765
rect 9475 -1795 9476 -1765
rect 9444 -1796 9476 -1795
rect 9444 -1845 9476 -1844
rect 9444 -1875 9445 -1845
rect 9445 -1875 9475 -1845
rect 9475 -1875 9476 -1845
rect 9444 -1876 9476 -1875
rect 9444 -1956 9476 -1924
rect 9444 -2005 9476 -2004
rect 9444 -2035 9445 -2005
rect 9445 -2035 9475 -2005
rect 9475 -2035 9476 -2005
rect 9444 -2036 9476 -2035
rect 9444 -2116 9476 -2084
rect 9444 -2165 9476 -2164
rect 9444 -2195 9445 -2165
rect 9445 -2195 9475 -2165
rect 9475 -2195 9476 -2165
rect 9444 -2196 9476 -2195
rect 9444 -2276 9476 -2244
rect 9444 -2325 9476 -2324
rect 9444 -2355 9445 -2325
rect 9445 -2355 9475 -2325
rect 9475 -2355 9476 -2325
rect 9444 -2356 9476 -2355
rect 9444 -2405 9476 -2404
rect 9444 -2435 9445 -2405
rect 9445 -2435 9475 -2405
rect 9475 -2435 9476 -2405
rect 9444 -2436 9476 -2435
rect 9444 -2485 9476 -2484
rect 9444 -2515 9445 -2485
rect 9445 -2515 9475 -2485
rect 9475 -2515 9476 -2485
rect 9444 -2516 9476 -2515
rect 9444 -2565 9476 -2564
rect 9444 -2595 9445 -2565
rect 9445 -2595 9475 -2565
rect 9475 -2595 9476 -2565
rect 9444 -2596 9476 -2595
rect 9444 -2645 9476 -2644
rect 9444 -2675 9445 -2645
rect 9445 -2675 9475 -2645
rect 9475 -2675 9476 -2645
rect 9444 -2676 9476 -2675
rect 9444 -2725 9476 -2724
rect 9444 -2755 9445 -2725
rect 9445 -2755 9475 -2725
rect 9475 -2755 9476 -2725
rect 9444 -2756 9476 -2755
rect 9444 -2836 9476 -2804
rect 9444 -2885 9476 -2884
rect 9444 -2915 9445 -2885
rect 9445 -2915 9475 -2885
rect 9475 -2915 9476 -2885
rect 9444 -2916 9476 -2915
rect 9444 -2996 9476 -2964
rect 9444 -3045 9476 -3044
rect 9444 -3075 9445 -3045
rect 9445 -3075 9475 -3045
rect 9475 -3075 9476 -3045
rect 9444 -3076 9476 -3075
rect 9444 -3156 9476 -3124
rect 9444 -3205 9476 -3204
rect 9444 -3235 9445 -3205
rect 9445 -3235 9475 -3205
rect 9475 -3235 9476 -3205
rect 9444 -3236 9476 -3235
rect 9444 -3285 9476 -3284
rect 9444 -3315 9445 -3285
rect 9445 -3315 9475 -3285
rect 9475 -3315 9476 -3285
rect 9444 -3316 9476 -3315
rect 9444 -3396 9476 -3364
rect 9444 -3476 9476 -3444
rect 9444 -3525 9476 -3524
rect 9444 -3555 9445 -3525
rect 9445 -3555 9475 -3525
rect 9475 -3555 9476 -3525
rect 9444 -3556 9476 -3555
rect 9444 -3605 9476 -3604
rect 9444 -3635 9445 -3605
rect 9445 -3635 9475 -3605
rect 9475 -3635 9476 -3605
rect 9444 -3636 9476 -3635
rect 9444 -3685 9476 -3684
rect 9444 -3715 9445 -3685
rect 9445 -3715 9475 -3685
rect 9475 -3715 9476 -3685
rect 9444 -3716 9476 -3715
rect 9524 1035 9556 1036
rect 9524 1005 9525 1035
rect 9525 1005 9555 1035
rect 9555 1005 9556 1035
rect 9524 1004 9556 1005
rect 9524 955 9556 956
rect 9524 925 9525 955
rect 9525 925 9555 955
rect 9555 925 9556 955
rect 9524 924 9556 925
rect 9524 875 9556 876
rect 9524 845 9525 875
rect 9525 845 9555 875
rect 9555 845 9556 875
rect 9524 844 9556 845
rect 9524 764 9556 796
rect 9524 684 9556 716
rect 9524 635 9556 636
rect 9524 605 9525 635
rect 9525 605 9555 635
rect 9555 605 9556 635
rect 9524 604 9556 605
rect 9524 555 9556 556
rect 9524 525 9525 555
rect 9525 525 9555 555
rect 9555 525 9556 555
rect 9524 524 9556 525
rect 9524 444 9556 476
rect 9524 395 9556 396
rect 9524 365 9525 395
rect 9525 365 9555 395
rect 9555 365 9556 395
rect 9524 364 9556 365
rect 9524 284 9556 316
rect 9524 235 9556 236
rect 9524 205 9525 235
rect 9525 205 9555 235
rect 9555 205 9556 235
rect 9524 204 9556 205
rect 9524 124 9556 156
rect 9524 75 9556 76
rect 9524 45 9525 75
rect 9525 45 9555 75
rect 9555 45 9556 75
rect 9524 44 9556 45
rect 9524 -5 9556 -4
rect 9524 -35 9525 -5
rect 9525 -35 9555 -5
rect 9555 -35 9556 -5
rect 9524 -36 9556 -35
rect 9524 -85 9556 -84
rect 9524 -115 9525 -85
rect 9525 -115 9555 -85
rect 9555 -115 9556 -85
rect 9524 -116 9556 -115
rect 9524 -165 9556 -164
rect 9524 -195 9525 -165
rect 9525 -195 9555 -165
rect 9555 -195 9556 -165
rect 9524 -196 9556 -195
rect 9524 -245 9556 -244
rect 9524 -275 9525 -245
rect 9525 -275 9555 -245
rect 9555 -275 9556 -245
rect 9524 -276 9556 -275
rect 9524 -325 9556 -324
rect 9524 -355 9525 -325
rect 9525 -355 9555 -325
rect 9555 -355 9556 -325
rect 9524 -356 9556 -355
rect 9524 -436 9556 -404
rect 9524 -485 9556 -484
rect 9524 -515 9525 -485
rect 9525 -515 9555 -485
rect 9555 -515 9556 -485
rect 9524 -516 9556 -515
rect 9524 -596 9556 -564
rect 9524 -645 9556 -644
rect 9524 -675 9525 -645
rect 9525 -675 9555 -645
rect 9555 -675 9556 -645
rect 9524 -676 9556 -675
rect 9524 -756 9556 -724
rect 9524 -805 9556 -804
rect 9524 -835 9525 -805
rect 9525 -835 9555 -805
rect 9555 -835 9556 -805
rect 9524 -836 9556 -835
rect 9524 -885 9556 -884
rect 9524 -915 9525 -885
rect 9525 -915 9555 -885
rect 9555 -915 9556 -885
rect 9524 -916 9556 -915
rect 9524 -996 9556 -964
rect 9524 -1076 9556 -1044
rect 9524 -1125 9556 -1124
rect 9524 -1155 9525 -1125
rect 9525 -1155 9555 -1125
rect 9555 -1155 9556 -1125
rect 9524 -1156 9556 -1155
rect 9524 -1205 9556 -1204
rect 9524 -1235 9525 -1205
rect 9525 -1235 9555 -1205
rect 9555 -1235 9556 -1205
rect 9524 -1236 9556 -1235
rect 9524 -1285 9556 -1284
rect 9524 -1315 9525 -1285
rect 9525 -1315 9555 -1285
rect 9555 -1315 9556 -1285
rect 9524 -1316 9556 -1315
rect 9524 -1365 9556 -1364
rect 9524 -1395 9525 -1365
rect 9525 -1395 9555 -1365
rect 9555 -1395 9556 -1365
rect 9524 -1396 9556 -1395
rect 9524 -1445 9556 -1444
rect 9524 -1475 9525 -1445
rect 9525 -1475 9555 -1445
rect 9555 -1475 9556 -1445
rect 9524 -1476 9556 -1475
rect 9524 -1525 9556 -1524
rect 9524 -1555 9525 -1525
rect 9525 -1555 9555 -1525
rect 9555 -1555 9556 -1525
rect 9524 -1556 9556 -1555
rect 9524 -1636 9556 -1604
rect 9524 -1716 9556 -1684
rect 9524 -1765 9556 -1764
rect 9524 -1795 9525 -1765
rect 9525 -1795 9555 -1765
rect 9555 -1795 9556 -1765
rect 9524 -1796 9556 -1795
rect 9524 -1845 9556 -1844
rect 9524 -1875 9525 -1845
rect 9525 -1875 9555 -1845
rect 9555 -1875 9556 -1845
rect 9524 -1876 9556 -1875
rect 9524 -1956 9556 -1924
rect 9524 -2005 9556 -2004
rect 9524 -2035 9525 -2005
rect 9525 -2035 9555 -2005
rect 9555 -2035 9556 -2005
rect 9524 -2036 9556 -2035
rect 9524 -2116 9556 -2084
rect 9524 -2165 9556 -2164
rect 9524 -2195 9525 -2165
rect 9525 -2195 9555 -2165
rect 9555 -2195 9556 -2165
rect 9524 -2196 9556 -2195
rect 9524 -2276 9556 -2244
rect 9524 -2325 9556 -2324
rect 9524 -2355 9525 -2325
rect 9525 -2355 9555 -2325
rect 9555 -2355 9556 -2325
rect 9524 -2356 9556 -2355
rect 9524 -2405 9556 -2404
rect 9524 -2435 9525 -2405
rect 9525 -2435 9555 -2405
rect 9555 -2435 9556 -2405
rect 9524 -2436 9556 -2435
rect 9524 -2485 9556 -2484
rect 9524 -2515 9525 -2485
rect 9525 -2515 9555 -2485
rect 9555 -2515 9556 -2485
rect 9524 -2516 9556 -2515
rect 9524 -2565 9556 -2564
rect 9524 -2595 9525 -2565
rect 9525 -2595 9555 -2565
rect 9555 -2595 9556 -2565
rect 9524 -2596 9556 -2595
rect 9524 -2645 9556 -2644
rect 9524 -2675 9525 -2645
rect 9525 -2675 9555 -2645
rect 9555 -2675 9556 -2645
rect 9524 -2676 9556 -2675
rect 9524 -2725 9556 -2724
rect 9524 -2755 9525 -2725
rect 9525 -2755 9555 -2725
rect 9555 -2755 9556 -2725
rect 9524 -2756 9556 -2755
rect 9524 -2836 9556 -2804
rect 9524 -2885 9556 -2884
rect 9524 -2915 9525 -2885
rect 9525 -2915 9555 -2885
rect 9555 -2915 9556 -2885
rect 9524 -2916 9556 -2915
rect 9524 -2996 9556 -2964
rect 9524 -3045 9556 -3044
rect 9524 -3075 9525 -3045
rect 9525 -3075 9555 -3045
rect 9555 -3075 9556 -3045
rect 9524 -3076 9556 -3075
rect 9524 -3156 9556 -3124
rect 9524 -3205 9556 -3204
rect 9524 -3235 9525 -3205
rect 9525 -3235 9555 -3205
rect 9555 -3235 9556 -3205
rect 9524 -3236 9556 -3235
rect 9524 -3285 9556 -3284
rect 9524 -3315 9525 -3285
rect 9525 -3315 9555 -3285
rect 9555 -3315 9556 -3285
rect 9524 -3316 9556 -3315
rect 9524 -3396 9556 -3364
rect 9524 -3476 9556 -3444
rect 9524 -3525 9556 -3524
rect 9524 -3555 9525 -3525
rect 9525 -3555 9555 -3525
rect 9555 -3555 9556 -3525
rect 9524 -3556 9556 -3555
rect 9524 -3605 9556 -3604
rect 9524 -3635 9525 -3605
rect 9525 -3635 9555 -3605
rect 9555 -3635 9556 -3605
rect 9524 -3636 9556 -3635
rect 9524 -3685 9556 -3684
rect 9524 -3715 9525 -3685
rect 9525 -3715 9555 -3685
rect 9555 -3715 9556 -3685
rect 9524 -3716 9556 -3715
rect 9604 1035 9636 1036
rect 9604 1005 9605 1035
rect 9605 1005 9635 1035
rect 9635 1005 9636 1035
rect 9604 1004 9636 1005
rect 9604 955 9636 956
rect 9604 925 9605 955
rect 9605 925 9635 955
rect 9635 925 9636 955
rect 9604 924 9636 925
rect 9604 875 9636 876
rect 9604 845 9605 875
rect 9605 845 9635 875
rect 9635 845 9636 875
rect 9604 844 9636 845
rect 9604 764 9636 796
rect 9604 684 9636 716
rect 9604 635 9636 636
rect 9604 605 9605 635
rect 9605 605 9635 635
rect 9635 605 9636 635
rect 9604 604 9636 605
rect 9604 555 9636 556
rect 9604 525 9605 555
rect 9605 525 9635 555
rect 9635 525 9636 555
rect 9604 524 9636 525
rect 9604 444 9636 476
rect 9604 395 9636 396
rect 9604 365 9605 395
rect 9605 365 9635 395
rect 9635 365 9636 395
rect 9604 364 9636 365
rect 9604 284 9636 316
rect 9604 235 9636 236
rect 9604 205 9605 235
rect 9605 205 9635 235
rect 9635 205 9636 235
rect 9604 204 9636 205
rect 9604 124 9636 156
rect 9604 75 9636 76
rect 9604 45 9605 75
rect 9605 45 9635 75
rect 9635 45 9636 75
rect 9604 44 9636 45
rect 9604 -5 9636 -4
rect 9604 -35 9605 -5
rect 9605 -35 9635 -5
rect 9635 -35 9636 -5
rect 9604 -36 9636 -35
rect 9604 -85 9636 -84
rect 9604 -115 9605 -85
rect 9605 -115 9635 -85
rect 9635 -115 9636 -85
rect 9604 -116 9636 -115
rect 9604 -165 9636 -164
rect 9604 -195 9605 -165
rect 9605 -195 9635 -165
rect 9635 -195 9636 -165
rect 9604 -196 9636 -195
rect 9604 -245 9636 -244
rect 9604 -275 9605 -245
rect 9605 -275 9635 -245
rect 9635 -275 9636 -245
rect 9604 -276 9636 -275
rect 9604 -325 9636 -324
rect 9604 -355 9605 -325
rect 9605 -355 9635 -325
rect 9635 -355 9636 -325
rect 9604 -356 9636 -355
rect 9604 -436 9636 -404
rect 9604 -485 9636 -484
rect 9604 -515 9605 -485
rect 9605 -515 9635 -485
rect 9635 -515 9636 -485
rect 9604 -516 9636 -515
rect 9604 -596 9636 -564
rect 9604 -645 9636 -644
rect 9604 -675 9605 -645
rect 9605 -675 9635 -645
rect 9635 -675 9636 -645
rect 9604 -676 9636 -675
rect 9604 -756 9636 -724
rect 9604 -805 9636 -804
rect 9604 -835 9605 -805
rect 9605 -835 9635 -805
rect 9635 -835 9636 -805
rect 9604 -836 9636 -835
rect 9604 -885 9636 -884
rect 9604 -915 9605 -885
rect 9605 -915 9635 -885
rect 9635 -915 9636 -885
rect 9604 -916 9636 -915
rect 9604 -996 9636 -964
rect 9604 -1076 9636 -1044
rect 9604 -1125 9636 -1124
rect 9604 -1155 9605 -1125
rect 9605 -1155 9635 -1125
rect 9635 -1155 9636 -1125
rect 9604 -1156 9636 -1155
rect 9604 -1205 9636 -1204
rect 9604 -1235 9605 -1205
rect 9605 -1235 9635 -1205
rect 9635 -1235 9636 -1205
rect 9604 -1236 9636 -1235
rect 9604 -1285 9636 -1284
rect 9604 -1315 9605 -1285
rect 9605 -1315 9635 -1285
rect 9635 -1315 9636 -1285
rect 9604 -1316 9636 -1315
rect 9604 -1365 9636 -1364
rect 9604 -1395 9605 -1365
rect 9605 -1395 9635 -1365
rect 9635 -1395 9636 -1365
rect 9604 -1396 9636 -1395
rect 9604 -1445 9636 -1444
rect 9604 -1475 9605 -1445
rect 9605 -1475 9635 -1445
rect 9635 -1475 9636 -1445
rect 9604 -1476 9636 -1475
rect 9604 -1525 9636 -1524
rect 9604 -1555 9605 -1525
rect 9605 -1555 9635 -1525
rect 9635 -1555 9636 -1525
rect 9604 -1556 9636 -1555
rect 9604 -1636 9636 -1604
rect 9604 -1716 9636 -1684
rect 9604 -1765 9636 -1764
rect 9604 -1795 9605 -1765
rect 9605 -1795 9635 -1765
rect 9635 -1795 9636 -1765
rect 9604 -1796 9636 -1795
rect 9604 -1845 9636 -1844
rect 9604 -1875 9605 -1845
rect 9605 -1875 9635 -1845
rect 9635 -1875 9636 -1845
rect 9604 -1876 9636 -1875
rect 9604 -1956 9636 -1924
rect 9604 -2005 9636 -2004
rect 9604 -2035 9605 -2005
rect 9605 -2035 9635 -2005
rect 9635 -2035 9636 -2005
rect 9604 -2036 9636 -2035
rect 9604 -2116 9636 -2084
rect 9604 -2165 9636 -2164
rect 9604 -2195 9605 -2165
rect 9605 -2195 9635 -2165
rect 9635 -2195 9636 -2165
rect 9604 -2196 9636 -2195
rect 9604 -2276 9636 -2244
rect 9604 -2325 9636 -2324
rect 9604 -2355 9605 -2325
rect 9605 -2355 9635 -2325
rect 9635 -2355 9636 -2325
rect 9604 -2356 9636 -2355
rect 9604 -2405 9636 -2404
rect 9604 -2435 9605 -2405
rect 9605 -2435 9635 -2405
rect 9635 -2435 9636 -2405
rect 9604 -2436 9636 -2435
rect 9604 -2485 9636 -2484
rect 9604 -2515 9605 -2485
rect 9605 -2515 9635 -2485
rect 9635 -2515 9636 -2485
rect 9604 -2516 9636 -2515
rect 9604 -2565 9636 -2564
rect 9604 -2595 9605 -2565
rect 9605 -2595 9635 -2565
rect 9635 -2595 9636 -2565
rect 9604 -2596 9636 -2595
rect 9604 -2645 9636 -2644
rect 9604 -2675 9605 -2645
rect 9605 -2675 9635 -2645
rect 9635 -2675 9636 -2645
rect 9604 -2676 9636 -2675
rect 9604 -2725 9636 -2724
rect 9604 -2755 9605 -2725
rect 9605 -2755 9635 -2725
rect 9635 -2755 9636 -2725
rect 9604 -2756 9636 -2755
rect 9604 -2836 9636 -2804
rect 9604 -2885 9636 -2884
rect 9604 -2915 9605 -2885
rect 9605 -2915 9635 -2885
rect 9635 -2915 9636 -2885
rect 9604 -2916 9636 -2915
rect 9604 -2996 9636 -2964
rect 9604 -3045 9636 -3044
rect 9604 -3075 9605 -3045
rect 9605 -3075 9635 -3045
rect 9635 -3075 9636 -3045
rect 9604 -3076 9636 -3075
rect 9604 -3156 9636 -3124
rect 9604 -3205 9636 -3204
rect 9604 -3235 9605 -3205
rect 9605 -3235 9635 -3205
rect 9635 -3235 9636 -3205
rect 9604 -3236 9636 -3235
rect 9604 -3285 9636 -3284
rect 9604 -3315 9605 -3285
rect 9605 -3315 9635 -3285
rect 9635 -3315 9636 -3285
rect 9604 -3316 9636 -3315
rect 9604 -3396 9636 -3364
rect 9604 -3476 9636 -3444
rect 9604 -3525 9636 -3524
rect 9604 -3555 9605 -3525
rect 9605 -3555 9635 -3525
rect 9635 -3555 9636 -3525
rect 9604 -3556 9636 -3555
rect 9604 -3605 9636 -3604
rect 9604 -3635 9605 -3605
rect 9605 -3635 9635 -3605
rect 9635 -3635 9636 -3605
rect 9604 -3636 9636 -3635
rect 9604 -3685 9636 -3684
rect 9604 -3715 9605 -3685
rect 9605 -3715 9635 -3685
rect 9635 -3715 9636 -3685
rect 9604 -3716 9636 -3715
rect 9684 1035 9716 1036
rect 9684 1005 9685 1035
rect 9685 1005 9715 1035
rect 9715 1005 9716 1035
rect 9684 1004 9716 1005
rect 9684 955 9716 956
rect 9684 925 9685 955
rect 9685 925 9715 955
rect 9715 925 9716 955
rect 9684 924 9716 925
rect 9684 875 9716 876
rect 9684 845 9685 875
rect 9685 845 9715 875
rect 9715 845 9716 875
rect 9684 844 9716 845
rect 9684 764 9716 796
rect 9684 684 9716 716
rect 9684 635 9716 636
rect 9684 605 9685 635
rect 9685 605 9715 635
rect 9715 605 9716 635
rect 9684 604 9716 605
rect 9684 555 9716 556
rect 9684 525 9685 555
rect 9685 525 9715 555
rect 9715 525 9716 555
rect 9684 524 9716 525
rect 9684 444 9716 476
rect 9684 395 9716 396
rect 9684 365 9685 395
rect 9685 365 9715 395
rect 9715 365 9716 395
rect 9684 364 9716 365
rect 9684 284 9716 316
rect 9684 235 9716 236
rect 9684 205 9685 235
rect 9685 205 9715 235
rect 9715 205 9716 235
rect 9684 204 9716 205
rect 9684 124 9716 156
rect 9684 75 9716 76
rect 9684 45 9685 75
rect 9685 45 9715 75
rect 9715 45 9716 75
rect 9684 44 9716 45
rect 9684 -5 9716 -4
rect 9684 -35 9685 -5
rect 9685 -35 9715 -5
rect 9715 -35 9716 -5
rect 9684 -36 9716 -35
rect 9684 -85 9716 -84
rect 9684 -115 9685 -85
rect 9685 -115 9715 -85
rect 9715 -115 9716 -85
rect 9684 -116 9716 -115
rect 9684 -165 9716 -164
rect 9684 -195 9685 -165
rect 9685 -195 9715 -165
rect 9715 -195 9716 -165
rect 9684 -196 9716 -195
rect 9684 -245 9716 -244
rect 9684 -275 9685 -245
rect 9685 -275 9715 -245
rect 9715 -275 9716 -245
rect 9684 -276 9716 -275
rect 9684 -325 9716 -324
rect 9684 -355 9685 -325
rect 9685 -355 9715 -325
rect 9715 -355 9716 -325
rect 9684 -356 9716 -355
rect 9684 -436 9716 -404
rect 9684 -485 9716 -484
rect 9684 -515 9685 -485
rect 9685 -515 9715 -485
rect 9715 -515 9716 -485
rect 9684 -516 9716 -515
rect 9684 -596 9716 -564
rect 9684 -645 9716 -644
rect 9684 -675 9685 -645
rect 9685 -675 9715 -645
rect 9715 -675 9716 -645
rect 9684 -676 9716 -675
rect 9684 -756 9716 -724
rect 9684 -805 9716 -804
rect 9684 -835 9685 -805
rect 9685 -835 9715 -805
rect 9715 -835 9716 -805
rect 9684 -836 9716 -835
rect 9684 -885 9716 -884
rect 9684 -915 9685 -885
rect 9685 -915 9715 -885
rect 9715 -915 9716 -885
rect 9684 -916 9716 -915
rect 9684 -996 9716 -964
rect 9684 -1076 9716 -1044
rect 9684 -1125 9716 -1124
rect 9684 -1155 9685 -1125
rect 9685 -1155 9715 -1125
rect 9715 -1155 9716 -1125
rect 9684 -1156 9716 -1155
rect 9684 -1205 9716 -1204
rect 9684 -1235 9685 -1205
rect 9685 -1235 9715 -1205
rect 9715 -1235 9716 -1205
rect 9684 -1236 9716 -1235
rect 9684 -1285 9716 -1284
rect 9684 -1315 9685 -1285
rect 9685 -1315 9715 -1285
rect 9715 -1315 9716 -1285
rect 9684 -1316 9716 -1315
rect 9684 -1365 9716 -1364
rect 9684 -1395 9685 -1365
rect 9685 -1395 9715 -1365
rect 9715 -1395 9716 -1365
rect 9684 -1396 9716 -1395
rect 9684 -1445 9716 -1444
rect 9684 -1475 9685 -1445
rect 9685 -1475 9715 -1445
rect 9715 -1475 9716 -1445
rect 9684 -1476 9716 -1475
rect 9684 -1525 9716 -1524
rect 9684 -1555 9685 -1525
rect 9685 -1555 9715 -1525
rect 9715 -1555 9716 -1525
rect 9684 -1556 9716 -1555
rect 9684 -1636 9716 -1604
rect 9684 -1716 9716 -1684
rect 9684 -1765 9716 -1764
rect 9684 -1795 9685 -1765
rect 9685 -1795 9715 -1765
rect 9715 -1795 9716 -1765
rect 9684 -1796 9716 -1795
rect 9684 -1845 9716 -1844
rect 9684 -1875 9685 -1845
rect 9685 -1875 9715 -1845
rect 9715 -1875 9716 -1845
rect 9684 -1876 9716 -1875
rect 9684 -1956 9716 -1924
rect 9684 -2005 9716 -2004
rect 9684 -2035 9685 -2005
rect 9685 -2035 9715 -2005
rect 9715 -2035 9716 -2005
rect 9684 -2036 9716 -2035
rect 9684 -2116 9716 -2084
rect 9684 -2165 9716 -2164
rect 9684 -2195 9685 -2165
rect 9685 -2195 9715 -2165
rect 9715 -2195 9716 -2165
rect 9684 -2196 9716 -2195
rect 9684 -2276 9716 -2244
rect 9684 -2325 9716 -2324
rect 9684 -2355 9685 -2325
rect 9685 -2355 9715 -2325
rect 9715 -2355 9716 -2325
rect 9684 -2356 9716 -2355
rect 9684 -2405 9716 -2404
rect 9684 -2435 9685 -2405
rect 9685 -2435 9715 -2405
rect 9715 -2435 9716 -2405
rect 9684 -2436 9716 -2435
rect 9684 -2485 9716 -2484
rect 9684 -2515 9685 -2485
rect 9685 -2515 9715 -2485
rect 9715 -2515 9716 -2485
rect 9684 -2516 9716 -2515
rect 9684 -2565 9716 -2564
rect 9684 -2595 9685 -2565
rect 9685 -2595 9715 -2565
rect 9715 -2595 9716 -2565
rect 9684 -2596 9716 -2595
rect 9684 -2645 9716 -2644
rect 9684 -2675 9685 -2645
rect 9685 -2675 9715 -2645
rect 9715 -2675 9716 -2645
rect 9684 -2676 9716 -2675
rect 9684 -2725 9716 -2724
rect 9684 -2755 9685 -2725
rect 9685 -2755 9715 -2725
rect 9715 -2755 9716 -2725
rect 9684 -2756 9716 -2755
rect 9684 -2836 9716 -2804
rect 9684 -2885 9716 -2884
rect 9684 -2915 9685 -2885
rect 9685 -2915 9715 -2885
rect 9715 -2915 9716 -2885
rect 9684 -2916 9716 -2915
rect 9684 -2996 9716 -2964
rect 9684 -3045 9716 -3044
rect 9684 -3075 9685 -3045
rect 9685 -3075 9715 -3045
rect 9715 -3075 9716 -3045
rect 9684 -3076 9716 -3075
rect 9684 -3156 9716 -3124
rect 9684 -3205 9716 -3204
rect 9684 -3235 9685 -3205
rect 9685 -3235 9715 -3205
rect 9715 -3235 9716 -3205
rect 9684 -3236 9716 -3235
rect 9684 -3285 9716 -3284
rect 9684 -3315 9685 -3285
rect 9685 -3315 9715 -3285
rect 9715 -3315 9716 -3285
rect 9684 -3316 9716 -3315
rect 9684 -3396 9716 -3364
rect 9684 -3476 9716 -3444
rect 9684 -3525 9716 -3524
rect 9684 -3555 9685 -3525
rect 9685 -3555 9715 -3525
rect 9715 -3555 9716 -3525
rect 9684 -3556 9716 -3555
rect 9684 -3605 9716 -3604
rect 9684 -3635 9685 -3605
rect 9685 -3635 9715 -3605
rect 9715 -3635 9716 -3605
rect 9684 -3636 9716 -3635
rect 9684 -3685 9716 -3684
rect 9684 -3715 9685 -3685
rect 9685 -3715 9715 -3685
rect 9715 -3715 9716 -3685
rect 9684 -3716 9716 -3715
rect 9764 1035 9796 1036
rect 9764 1005 9765 1035
rect 9765 1005 9795 1035
rect 9795 1005 9796 1035
rect 9764 1004 9796 1005
rect 9764 955 9796 956
rect 9764 925 9765 955
rect 9765 925 9795 955
rect 9795 925 9796 955
rect 9764 924 9796 925
rect 9764 875 9796 876
rect 9764 845 9765 875
rect 9765 845 9795 875
rect 9795 845 9796 875
rect 9764 844 9796 845
rect 9764 764 9796 796
rect 9764 684 9796 716
rect 9764 635 9796 636
rect 9764 605 9765 635
rect 9765 605 9795 635
rect 9795 605 9796 635
rect 9764 604 9796 605
rect 9764 555 9796 556
rect 9764 525 9765 555
rect 9765 525 9795 555
rect 9795 525 9796 555
rect 9764 524 9796 525
rect 9764 444 9796 476
rect 9764 395 9796 396
rect 9764 365 9765 395
rect 9765 365 9795 395
rect 9795 365 9796 395
rect 9764 364 9796 365
rect 9764 284 9796 316
rect 9764 235 9796 236
rect 9764 205 9765 235
rect 9765 205 9795 235
rect 9795 205 9796 235
rect 9764 204 9796 205
rect 9764 124 9796 156
rect 9764 75 9796 76
rect 9764 45 9765 75
rect 9765 45 9795 75
rect 9795 45 9796 75
rect 9764 44 9796 45
rect 9764 -5 9796 -4
rect 9764 -35 9765 -5
rect 9765 -35 9795 -5
rect 9795 -35 9796 -5
rect 9764 -36 9796 -35
rect 9764 -85 9796 -84
rect 9764 -115 9765 -85
rect 9765 -115 9795 -85
rect 9795 -115 9796 -85
rect 9764 -116 9796 -115
rect 9764 -165 9796 -164
rect 9764 -195 9765 -165
rect 9765 -195 9795 -165
rect 9795 -195 9796 -165
rect 9764 -196 9796 -195
rect 9764 -245 9796 -244
rect 9764 -275 9765 -245
rect 9765 -275 9795 -245
rect 9795 -275 9796 -245
rect 9764 -276 9796 -275
rect 9764 -325 9796 -324
rect 9764 -355 9765 -325
rect 9765 -355 9795 -325
rect 9795 -355 9796 -325
rect 9764 -356 9796 -355
rect 9764 -436 9796 -404
rect 9764 -485 9796 -484
rect 9764 -515 9765 -485
rect 9765 -515 9795 -485
rect 9795 -515 9796 -485
rect 9764 -516 9796 -515
rect 9764 -596 9796 -564
rect 9764 -645 9796 -644
rect 9764 -675 9765 -645
rect 9765 -675 9795 -645
rect 9795 -675 9796 -645
rect 9764 -676 9796 -675
rect 9764 -756 9796 -724
rect 9764 -805 9796 -804
rect 9764 -835 9765 -805
rect 9765 -835 9795 -805
rect 9795 -835 9796 -805
rect 9764 -836 9796 -835
rect 9764 -885 9796 -884
rect 9764 -915 9765 -885
rect 9765 -915 9795 -885
rect 9795 -915 9796 -885
rect 9764 -916 9796 -915
rect 9764 -996 9796 -964
rect 9764 -1076 9796 -1044
rect 9764 -1125 9796 -1124
rect 9764 -1155 9765 -1125
rect 9765 -1155 9795 -1125
rect 9795 -1155 9796 -1125
rect 9764 -1156 9796 -1155
rect 9764 -1205 9796 -1204
rect 9764 -1235 9765 -1205
rect 9765 -1235 9795 -1205
rect 9795 -1235 9796 -1205
rect 9764 -1236 9796 -1235
rect 9764 -1285 9796 -1284
rect 9764 -1315 9765 -1285
rect 9765 -1315 9795 -1285
rect 9795 -1315 9796 -1285
rect 9764 -1316 9796 -1315
rect 9764 -1365 9796 -1364
rect 9764 -1395 9765 -1365
rect 9765 -1395 9795 -1365
rect 9795 -1395 9796 -1365
rect 9764 -1396 9796 -1395
rect 9764 -1445 9796 -1444
rect 9764 -1475 9765 -1445
rect 9765 -1475 9795 -1445
rect 9795 -1475 9796 -1445
rect 9764 -1476 9796 -1475
rect 9764 -1525 9796 -1524
rect 9764 -1555 9765 -1525
rect 9765 -1555 9795 -1525
rect 9795 -1555 9796 -1525
rect 9764 -1556 9796 -1555
rect 9764 -1636 9796 -1604
rect 9764 -1716 9796 -1684
rect 9764 -1765 9796 -1764
rect 9764 -1795 9765 -1765
rect 9765 -1795 9795 -1765
rect 9795 -1795 9796 -1765
rect 9764 -1796 9796 -1795
rect 9764 -1845 9796 -1844
rect 9764 -1875 9765 -1845
rect 9765 -1875 9795 -1845
rect 9795 -1875 9796 -1845
rect 9764 -1876 9796 -1875
rect 9764 -1956 9796 -1924
rect 9764 -2005 9796 -2004
rect 9764 -2035 9765 -2005
rect 9765 -2035 9795 -2005
rect 9795 -2035 9796 -2005
rect 9764 -2036 9796 -2035
rect 9764 -2116 9796 -2084
rect 9764 -2165 9796 -2164
rect 9764 -2195 9765 -2165
rect 9765 -2195 9795 -2165
rect 9795 -2195 9796 -2165
rect 9764 -2196 9796 -2195
rect 9764 -2276 9796 -2244
rect 9764 -2325 9796 -2324
rect 9764 -2355 9765 -2325
rect 9765 -2355 9795 -2325
rect 9795 -2355 9796 -2325
rect 9764 -2356 9796 -2355
rect 9764 -2405 9796 -2404
rect 9764 -2435 9765 -2405
rect 9765 -2435 9795 -2405
rect 9795 -2435 9796 -2405
rect 9764 -2436 9796 -2435
rect 9764 -2485 9796 -2484
rect 9764 -2515 9765 -2485
rect 9765 -2515 9795 -2485
rect 9795 -2515 9796 -2485
rect 9764 -2516 9796 -2515
rect 9764 -2565 9796 -2564
rect 9764 -2595 9765 -2565
rect 9765 -2595 9795 -2565
rect 9795 -2595 9796 -2565
rect 9764 -2596 9796 -2595
rect 9764 -2645 9796 -2644
rect 9764 -2675 9765 -2645
rect 9765 -2675 9795 -2645
rect 9795 -2675 9796 -2645
rect 9764 -2676 9796 -2675
rect 9764 -2725 9796 -2724
rect 9764 -2755 9765 -2725
rect 9765 -2755 9795 -2725
rect 9795 -2755 9796 -2725
rect 9764 -2756 9796 -2755
rect 9764 -2836 9796 -2804
rect 9764 -2885 9796 -2884
rect 9764 -2915 9765 -2885
rect 9765 -2915 9795 -2885
rect 9795 -2915 9796 -2885
rect 9764 -2916 9796 -2915
rect 9764 -2996 9796 -2964
rect 9764 -3045 9796 -3044
rect 9764 -3075 9765 -3045
rect 9765 -3075 9795 -3045
rect 9795 -3075 9796 -3045
rect 9764 -3076 9796 -3075
rect 9764 -3156 9796 -3124
rect 9764 -3205 9796 -3204
rect 9764 -3235 9765 -3205
rect 9765 -3235 9795 -3205
rect 9795 -3235 9796 -3205
rect 9764 -3236 9796 -3235
rect 9764 -3285 9796 -3284
rect 9764 -3315 9765 -3285
rect 9765 -3315 9795 -3285
rect 9795 -3315 9796 -3285
rect 9764 -3316 9796 -3315
rect 9764 -3396 9796 -3364
rect 9764 -3476 9796 -3444
rect 9764 -3525 9796 -3524
rect 9764 -3555 9765 -3525
rect 9765 -3555 9795 -3525
rect 9795 -3555 9796 -3525
rect 9764 -3556 9796 -3555
rect 9764 -3605 9796 -3604
rect 9764 -3635 9765 -3605
rect 9765 -3635 9795 -3605
rect 9795 -3635 9796 -3605
rect 9764 -3636 9796 -3635
rect 9764 -3685 9796 -3684
rect 9764 -3715 9765 -3685
rect 9765 -3715 9795 -3685
rect 9795 -3715 9796 -3685
rect 9764 -3716 9796 -3715
rect 9844 1035 9876 1036
rect 9844 1005 9845 1035
rect 9845 1005 9875 1035
rect 9875 1005 9876 1035
rect 9844 1004 9876 1005
rect 9844 955 9876 956
rect 9844 925 9845 955
rect 9845 925 9875 955
rect 9875 925 9876 955
rect 9844 924 9876 925
rect 9844 875 9876 876
rect 9844 845 9845 875
rect 9845 845 9875 875
rect 9875 845 9876 875
rect 9844 844 9876 845
rect 9844 764 9876 796
rect 9844 684 9876 716
rect 9844 635 9876 636
rect 9844 605 9845 635
rect 9845 605 9875 635
rect 9875 605 9876 635
rect 9844 604 9876 605
rect 9844 555 9876 556
rect 9844 525 9845 555
rect 9845 525 9875 555
rect 9875 525 9876 555
rect 9844 524 9876 525
rect 9844 444 9876 476
rect 9844 395 9876 396
rect 9844 365 9845 395
rect 9845 365 9875 395
rect 9875 365 9876 395
rect 9844 364 9876 365
rect 9844 284 9876 316
rect 9844 235 9876 236
rect 9844 205 9845 235
rect 9845 205 9875 235
rect 9875 205 9876 235
rect 9844 204 9876 205
rect 9844 124 9876 156
rect 9844 75 9876 76
rect 9844 45 9845 75
rect 9845 45 9875 75
rect 9875 45 9876 75
rect 9844 44 9876 45
rect 9844 -5 9876 -4
rect 9844 -35 9845 -5
rect 9845 -35 9875 -5
rect 9875 -35 9876 -5
rect 9844 -36 9876 -35
rect 9844 -85 9876 -84
rect 9844 -115 9845 -85
rect 9845 -115 9875 -85
rect 9875 -115 9876 -85
rect 9844 -116 9876 -115
rect 9844 -165 9876 -164
rect 9844 -195 9845 -165
rect 9845 -195 9875 -165
rect 9875 -195 9876 -165
rect 9844 -196 9876 -195
rect 9844 -245 9876 -244
rect 9844 -275 9845 -245
rect 9845 -275 9875 -245
rect 9875 -275 9876 -245
rect 9844 -276 9876 -275
rect 9844 -325 9876 -324
rect 9844 -355 9845 -325
rect 9845 -355 9875 -325
rect 9875 -355 9876 -325
rect 9844 -356 9876 -355
rect 9844 -436 9876 -404
rect 9844 -485 9876 -484
rect 9844 -515 9845 -485
rect 9845 -515 9875 -485
rect 9875 -515 9876 -485
rect 9844 -516 9876 -515
rect 9844 -596 9876 -564
rect 9844 -645 9876 -644
rect 9844 -675 9845 -645
rect 9845 -675 9875 -645
rect 9875 -675 9876 -645
rect 9844 -676 9876 -675
rect 9844 -756 9876 -724
rect 9844 -805 9876 -804
rect 9844 -835 9845 -805
rect 9845 -835 9875 -805
rect 9875 -835 9876 -805
rect 9844 -836 9876 -835
rect 9844 -885 9876 -884
rect 9844 -915 9845 -885
rect 9845 -915 9875 -885
rect 9875 -915 9876 -885
rect 9844 -916 9876 -915
rect 9844 -996 9876 -964
rect 9844 -1076 9876 -1044
rect 9844 -1125 9876 -1124
rect 9844 -1155 9845 -1125
rect 9845 -1155 9875 -1125
rect 9875 -1155 9876 -1125
rect 9844 -1156 9876 -1155
rect 9844 -1205 9876 -1204
rect 9844 -1235 9845 -1205
rect 9845 -1235 9875 -1205
rect 9875 -1235 9876 -1205
rect 9844 -1236 9876 -1235
rect 9844 -1285 9876 -1284
rect 9844 -1315 9845 -1285
rect 9845 -1315 9875 -1285
rect 9875 -1315 9876 -1285
rect 9844 -1316 9876 -1315
rect 9844 -1365 9876 -1364
rect 9844 -1395 9845 -1365
rect 9845 -1395 9875 -1365
rect 9875 -1395 9876 -1365
rect 9844 -1396 9876 -1395
rect 9844 -1445 9876 -1444
rect 9844 -1475 9845 -1445
rect 9845 -1475 9875 -1445
rect 9875 -1475 9876 -1445
rect 9844 -1476 9876 -1475
rect 9844 -1525 9876 -1524
rect 9844 -1555 9845 -1525
rect 9845 -1555 9875 -1525
rect 9875 -1555 9876 -1525
rect 9844 -1556 9876 -1555
rect 9844 -1636 9876 -1604
rect 9844 -1716 9876 -1684
rect 9844 -1765 9876 -1764
rect 9844 -1795 9845 -1765
rect 9845 -1795 9875 -1765
rect 9875 -1795 9876 -1765
rect 9844 -1796 9876 -1795
rect 9844 -1845 9876 -1844
rect 9844 -1875 9845 -1845
rect 9845 -1875 9875 -1845
rect 9875 -1875 9876 -1845
rect 9844 -1876 9876 -1875
rect 9844 -1956 9876 -1924
rect 9844 -2005 9876 -2004
rect 9844 -2035 9845 -2005
rect 9845 -2035 9875 -2005
rect 9875 -2035 9876 -2005
rect 9844 -2036 9876 -2035
rect 9844 -2116 9876 -2084
rect 9844 -2165 9876 -2164
rect 9844 -2195 9845 -2165
rect 9845 -2195 9875 -2165
rect 9875 -2195 9876 -2165
rect 9844 -2196 9876 -2195
rect 9844 -2276 9876 -2244
rect 9844 -2325 9876 -2324
rect 9844 -2355 9845 -2325
rect 9845 -2355 9875 -2325
rect 9875 -2355 9876 -2325
rect 9844 -2356 9876 -2355
rect 9844 -2405 9876 -2404
rect 9844 -2435 9845 -2405
rect 9845 -2435 9875 -2405
rect 9875 -2435 9876 -2405
rect 9844 -2436 9876 -2435
rect 9844 -2485 9876 -2484
rect 9844 -2515 9845 -2485
rect 9845 -2515 9875 -2485
rect 9875 -2515 9876 -2485
rect 9844 -2516 9876 -2515
rect 9844 -2565 9876 -2564
rect 9844 -2595 9845 -2565
rect 9845 -2595 9875 -2565
rect 9875 -2595 9876 -2565
rect 9844 -2596 9876 -2595
rect 9844 -2645 9876 -2644
rect 9844 -2675 9845 -2645
rect 9845 -2675 9875 -2645
rect 9875 -2675 9876 -2645
rect 9844 -2676 9876 -2675
rect 9844 -2725 9876 -2724
rect 9844 -2755 9845 -2725
rect 9845 -2755 9875 -2725
rect 9875 -2755 9876 -2725
rect 9844 -2756 9876 -2755
rect 9844 -2836 9876 -2804
rect 9844 -2885 9876 -2884
rect 9844 -2915 9845 -2885
rect 9845 -2915 9875 -2885
rect 9875 -2915 9876 -2885
rect 9844 -2916 9876 -2915
rect 9844 -2996 9876 -2964
rect 9844 -3045 9876 -3044
rect 9844 -3075 9845 -3045
rect 9845 -3075 9875 -3045
rect 9875 -3075 9876 -3045
rect 9844 -3076 9876 -3075
rect 9844 -3156 9876 -3124
rect 9844 -3205 9876 -3204
rect 9844 -3235 9845 -3205
rect 9845 -3235 9875 -3205
rect 9875 -3235 9876 -3205
rect 9844 -3236 9876 -3235
rect 9844 -3285 9876 -3284
rect 9844 -3315 9845 -3285
rect 9845 -3315 9875 -3285
rect 9875 -3315 9876 -3285
rect 9844 -3316 9876 -3315
rect 9844 -3396 9876 -3364
rect 9844 -3476 9876 -3444
rect 9844 -3525 9876 -3524
rect 9844 -3555 9845 -3525
rect 9845 -3555 9875 -3525
rect 9875 -3555 9876 -3525
rect 9844 -3556 9876 -3555
rect 9844 -3605 9876 -3604
rect 9844 -3635 9845 -3605
rect 9845 -3635 9875 -3605
rect 9875 -3635 9876 -3605
rect 9844 -3636 9876 -3635
rect 9844 -3685 9876 -3684
rect 9844 -3715 9845 -3685
rect 9845 -3715 9875 -3685
rect 9875 -3715 9876 -3685
rect 9844 -3716 9876 -3715
rect 9924 1035 9956 1036
rect 9924 1005 9925 1035
rect 9925 1005 9955 1035
rect 9955 1005 9956 1035
rect 9924 1004 9956 1005
rect 9924 955 9956 956
rect 9924 925 9925 955
rect 9925 925 9955 955
rect 9955 925 9956 955
rect 9924 924 9956 925
rect 9924 875 9956 876
rect 9924 845 9925 875
rect 9925 845 9955 875
rect 9955 845 9956 875
rect 9924 844 9956 845
rect 9924 764 9956 796
rect 9924 684 9956 716
rect 9924 635 9956 636
rect 9924 605 9925 635
rect 9925 605 9955 635
rect 9955 605 9956 635
rect 9924 604 9956 605
rect 9924 555 9956 556
rect 9924 525 9925 555
rect 9925 525 9955 555
rect 9955 525 9956 555
rect 9924 524 9956 525
rect 9924 444 9956 476
rect 9924 395 9956 396
rect 9924 365 9925 395
rect 9925 365 9955 395
rect 9955 365 9956 395
rect 9924 364 9956 365
rect 9924 284 9956 316
rect 9924 235 9956 236
rect 9924 205 9925 235
rect 9925 205 9955 235
rect 9955 205 9956 235
rect 9924 204 9956 205
rect 9924 124 9956 156
rect 9924 75 9956 76
rect 9924 45 9925 75
rect 9925 45 9955 75
rect 9955 45 9956 75
rect 9924 44 9956 45
rect 9924 -5 9956 -4
rect 9924 -35 9925 -5
rect 9925 -35 9955 -5
rect 9955 -35 9956 -5
rect 9924 -36 9956 -35
rect 9924 -85 9956 -84
rect 9924 -115 9925 -85
rect 9925 -115 9955 -85
rect 9955 -115 9956 -85
rect 9924 -116 9956 -115
rect 9924 -165 9956 -164
rect 9924 -195 9925 -165
rect 9925 -195 9955 -165
rect 9955 -195 9956 -165
rect 9924 -196 9956 -195
rect 9924 -245 9956 -244
rect 9924 -275 9925 -245
rect 9925 -275 9955 -245
rect 9955 -275 9956 -245
rect 9924 -276 9956 -275
rect 9924 -325 9956 -324
rect 9924 -355 9925 -325
rect 9925 -355 9955 -325
rect 9955 -355 9956 -325
rect 9924 -356 9956 -355
rect 9924 -436 9956 -404
rect 9924 -485 9956 -484
rect 9924 -515 9925 -485
rect 9925 -515 9955 -485
rect 9955 -515 9956 -485
rect 9924 -516 9956 -515
rect 9924 -596 9956 -564
rect 9924 -645 9956 -644
rect 9924 -675 9925 -645
rect 9925 -675 9955 -645
rect 9955 -675 9956 -645
rect 9924 -676 9956 -675
rect 9924 -756 9956 -724
rect 9924 -805 9956 -804
rect 9924 -835 9925 -805
rect 9925 -835 9955 -805
rect 9955 -835 9956 -805
rect 9924 -836 9956 -835
rect 9924 -885 9956 -884
rect 9924 -915 9925 -885
rect 9925 -915 9955 -885
rect 9955 -915 9956 -885
rect 9924 -916 9956 -915
rect 9924 -996 9956 -964
rect 9924 -1076 9956 -1044
rect 9924 -1125 9956 -1124
rect 9924 -1155 9925 -1125
rect 9925 -1155 9955 -1125
rect 9955 -1155 9956 -1125
rect 9924 -1156 9956 -1155
rect 9924 -1205 9956 -1204
rect 9924 -1235 9925 -1205
rect 9925 -1235 9955 -1205
rect 9955 -1235 9956 -1205
rect 9924 -1236 9956 -1235
rect 9924 -1285 9956 -1284
rect 9924 -1315 9925 -1285
rect 9925 -1315 9955 -1285
rect 9955 -1315 9956 -1285
rect 9924 -1316 9956 -1315
rect 9924 -1365 9956 -1364
rect 9924 -1395 9925 -1365
rect 9925 -1395 9955 -1365
rect 9955 -1395 9956 -1365
rect 9924 -1396 9956 -1395
rect 9924 -1445 9956 -1444
rect 9924 -1475 9925 -1445
rect 9925 -1475 9955 -1445
rect 9955 -1475 9956 -1445
rect 9924 -1476 9956 -1475
rect 9924 -1525 9956 -1524
rect 9924 -1555 9925 -1525
rect 9925 -1555 9955 -1525
rect 9955 -1555 9956 -1525
rect 9924 -1556 9956 -1555
rect 9924 -1636 9956 -1604
rect 9924 -1716 9956 -1684
rect 9924 -1765 9956 -1764
rect 9924 -1795 9925 -1765
rect 9925 -1795 9955 -1765
rect 9955 -1795 9956 -1765
rect 9924 -1796 9956 -1795
rect 9924 -1845 9956 -1844
rect 9924 -1875 9925 -1845
rect 9925 -1875 9955 -1845
rect 9955 -1875 9956 -1845
rect 9924 -1876 9956 -1875
rect 9924 -1956 9956 -1924
rect 9924 -2005 9956 -2004
rect 9924 -2035 9925 -2005
rect 9925 -2035 9955 -2005
rect 9955 -2035 9956 -2005
rect 9924 -2036 9956 -2035
rect 9924 -2116 9956 -2084
rect 9924 -2165 9956 -2164
rect 9924 -2195 9925 -2165
rect 9925 -2195 9955 -2165
rect 9955 -2195 9956 -2165
rect 9924 -2196 9956 -2195
rect 9924 -2276 9956 -2244
rect 9924 -2325 9956 -2324
rect 9924 -2355 9925 -2325
rect 9925 -2355 9955 -2325
rect 9955 -2355 9956 -2325
rect 9924 -2356 9956 -2355
rect 9924 -2405 9956 -2404
rect 9924 -2435 9925 -2405
rect 9925 -2435 9955 -2405
rect 9955 -2435 9956 -2405
rect 9924 -2436 9956 -2435
rect 9924 -2485 9956 -2484
rect 9924 -2515 9925 -2485
rect 9925 -2515 9955 -2485
rect 9955 -2515 9956 -2485
rect 9924 -2516 9956 -2515
rect 9924 -2565 9956 -2564
rect 9924 -2595 9925 -2565
rect 9925 -2595 9955 -2565
rect 9955 -2595 9956 -2565
rect 9924 -2596 9956 -2595
rect 9924 -2645 9956 -2644
rect 9924 -2675 9925 -2645
rect 9925 -2675 9955 -2645
rect 9955 -2675 9956 -2645
rect 9924 -2676 9956 -2675
rect 9924 -2725 9956 -2724
rect 9924 -2755 9925 -2725
rect 9925 -2755 9955 -2725
rect 9955 -2755 9956 -2725
rect 9924 -2756 9956 -2755
rect 9924 -2836 9956 -2804
rect 9924 -2885 9956 -2884
rect 9924 -2915 9925 -2885
rect 9925 -2915 9955 -2885
rect 9955 -2915 9956 -2885
rect 9924 -2916 9956 -2915
rect 9924 -2996 9956 -2964
rect 9924 -3045 9956 -3044
rect 9924 -3075 9925 -3045
rect 9925 -3075 9955 -3045
rect 9955 -3075 9956 -3045
rect 9924 -3076 9956 -3075
rect 9924 -3156 9956 -3124
rect 9924 -3205 9956 -3204
rect 9924 -3235 9925 -3205
rect 9925 -3235 9955 -3205
rect 9955 -3235 9956 -3205
rect 9924 -3236 9956 -3235
rect 9924 -3285 9956 -3284
rect 9924 -3315 9925 -3285
rect 9925 -3315 9955 -3285
rect 9955 -3315 9956 -3285
rect 9924 -3316 9956 -3315
rect 9924 -3396 9956 -3364
rect 9924 -3476 9956 -3444
rect 9924 -3525 9956 -3524
rect 9924 -3555 9925 -3525
rect 9925 -3555 9955 -3525
rect 9955 -3555 9956 -3525
rect 9924 -3556 9956 -3555
rect 9924 -3605 9956 -3604
rect 9924 -3635 9925 -3605
rect 9925 -3635 9955 -3605
rect 9955 -3635 9956 -3605
rect 9924 -3636 9956 -3635
rect 9924 -3685 9956 -3684
rect 9924 -3715 9925 -3685
rect 9925 -3715 9955 -3685
rect 9955 -3715 9956 -3685
rect 9924 -3716 9956 -3715
rect 10004 1035 10036 1036
rect 10004 1005 10005 1035
rect 10005 1005 10035 1035
rect 10035 1005 10036 1035
rect 10004 1004 10036 1005
rect 10004 955 10036 956
rect 10004 925 10005 955
rect 10005 925 10035 955
rect 10035 925 10036 955
rect 10004 924 10036 925
rect 10004 875 10036 876
rect 10004 845 10005 875
rect 10005 845 10035 875
rect 10035 845 10036 875
rect 10004 844 10036 845
rect 10004 764 10036 796
rect 10004 684 10036 716
rect 10004 635 10036 636
rect 10004 605 10005 635
rect 10005 605 10035 635
rect 10035 605 10036 635
rect 10004 604 10036 605
rect 10004 555 10036 556
rect 10004 525 10005 555
rect 10005 525 10035 555
rect 10035 525 10036 555
rect 10004 524 10036 525
rect 10004 444 10036 476
rect 10004 395 10036 396
rect 10004 365 10005 395
rect 10005 365 10035 395
rect 10035 365 10036 395
rect 10004 364 10036 365
rect 10004 284 10036 316
rect 10004 235 10036 236
rect 10004 205 10005 235
rect 10005 205 10035 235
rect 10035 205 10036 235
rect 10004 204 10036 205
rect 10004 124 10036 156
rect 10004 75 10036 76
rect 10004 45 10005 75
rect 10005 45 10035 75
rect 10035 45 10036 75
rect 10004 44 10036 45
rect 10004 -5 10036 -4
rect 10004 -35 10005 -5
rect 10005 -35 10035 -5
rect 10035 -35 10036 -5
rect 10004 -36 10036 -35
rect 10004 -85 10036 -84
rect 10004 -115 10005 -85
rect 10005 -115 10035 -85
rect 10035 -115 10036 -85
rect 10004 -116 10036 -115
rect 10004 -165 10036 -164
rect 10004 -195 10005 -165
rect 10005 -195 10035 -165
rect 10035 -195 10036 -165
rect 10004 -196 10036 -195
rect 10004 -245 10036 -244
rect 10004 -275 10005 -245
rect 10005 -275 10035 -245
rect 10035 -275 10036 -245
rect 10004 -276 10036 -275
rect 10004 -325 10036 -324
rect 10004 -355 10005 -325
rect 10005 -355 10035 -325
rect 10035 -355 10036 -325
rect 10004 -356 10036 -355
rect 10004 -436 10036 -404
rect 10004 -485 10036 -484
rect 10004 -515 10005 -485
rect 10005 -515 10035 -485
rect 10035 -515 10036 -485
rect 10004 -516 10036 -515
rect 10004 -596 10036 -564
rect 10004 -645 10036 -644
rect 10004 -675 10005 -645
rect 10005 -675 10035 -645
rect 10035 -675 10036 -645
rect 10004 -676 10036 -675
rect 10004 -756 10036 -724
rect 10004 -805 10036 -804
rect 10004 -835 10005 -805
rect 10005 -835 10035 -805
rect 10035 -835 10036 -805
rect 10004 -836 10036 -835
rect 10004 -885 10036 -884
rect 10004 -915 10005 -885
rect 10005 -915 10035 -885
rect 10035 -915 10036 -885
rect 10004 -916 10036 -915
rect 10004 -996 10036 -964
rect 10004 -1076 10036 -1044
rect 10004 -1125 10036 -1124
rect 10004 -1155 10005 -1125
rect 10005 -1155 10035 -1125
rect 10035 -1155 10036 -1125
rect 10004 -1156 10036 -1155
rect 10004 -1205 10036 -1204
rect 10004 -1235 10005 -1205
rect 10005 -1235 10035 -1205
rect 10035 -1235 10036 -1205
rect 10004 -1236 10036 -1235
rect 10004 -1285 10036 -1284
rect 10004 -1315 10005 -1285
rect 10005 -1315 10035 -1285
rect 10035 -1315 10036 -1285
rect 10004 -1316 10036 -1315
rect 10004 -1365 10036 -1364
rect 10004 -1395 10005 -1365
rect 10005 -1395 10035 -1365
rect 10035 -1395 10036 -1365
rect 10004 -1396 10036 -1395
rect 10004 -1445 10036 -1444
rect 10004 -1475 10005 -1445
rect 10005 -1475 10035 -1445
rect 10035 -1475 10036 -1445
rect 10004 -1476 10036 -1475
rect 10004 -1525 10036 -1524
rect 10004 -1555 10005 -1525
rect 10005 -1555 10035 -1525
rect 10035 -1555 10036 -1525
rect 10004 -1556 10036 -1555
rect 10004 -1636 10036 -1604
rect 10004 -1716 10036 -1684
rect 10004 -1765 10036 -1764
rect 10004 -1795 10005 -1765
rect 10005 -1795 10035 -1765
rect 10035 -1795 10036 -1765
rect 10004 -1796 10036 -1795
rect 10004 -1845 10036 -1844
rect 10004 -1875 10005 -1845
rect 10005 -1875 10035 -1845
rect 10035 -1875 10036 -1845
rect 10004 -1876 10036 -1875
rect 10004 -1956 10036 -1924
rect 10004 -2005 10036 -2004
rect 10004 -2035 10005 -2005
rect 10005 -2035 10035 -2005
rect 10035 -2035 10036 -2005
rect 10004 -2036 10036 -2035
rect 10004 -2116 10036 -2084
rect 10004 -2165 10036 -2164
rect 10004 -2195 10005 -2165
rect 10005 -2195 10035 -2165
rect 10035 -2195 10036 -2165
rect 10004 -2196 10036 -2195
rect 10004 -2276 10036 -2244
rect 10004 -2325 10036 -2324
rect 10004 -2355 10005 -2325
rect 10005 -2355 10035 -2325
rect 10035 -2355 10036 -2325
rect 10004 -2356 10036 -2355
rect 10004 -2405 10036 -2404
rect 10004 -2435 10005 -2405
rect 10005 -2435 10035 -2405
rect 10035 -2435 10036 -2405
rect 10004 -2436 10036 -2435
rect 10004 -2485 10036 -2484
rect 10004 -2515 10005 -2485
rect 10005 -2515 10035 -2485
rect 10035 -2515 10036 -2485
rect 10004 -2516 10036 -2515
rect 10004 -2565 10036 -2564
rect 10004 -2595 10005 -2565
rect 10005 -2595 10035 -2565
rect 10035 -2595 10036 -2565
rect 10004 -2596 10036 -2595
rect 10004 -2645 10036 -2644
rect 10004 -2675 10005 -2645
rect 10005 -2675 10035 -2645
rect 10035 -2675 10036 -2645
rect 10004 -2676 10036 -2675
rect 10004 -2725 10036 -2724
rect 10004 -2755 10005 -2725
rect 10005 -2755 10035 -2725
rect 10035 -2755 10036 -2725
rect 10004 -2756 10036 -2755
rect 10004 -2836 10036 -2804
rect 10004 -2885 10036 -2884
rect 10004 -2915 10005 -2885
rect 10005 -2915 10035 -2885
rect 10035 -2915 10036 -2885
rect 10004 -2916 10036 -2915
rect 10004 -2996 10036 -2964
rect 10004 -3045 10036 -3044
rect 10004 -3075 10005 -3045
rect 10005 -3075 10035 -3045
rect 10035 -3075 10036 -3045
rect 10004 -3076 10036 -3075
rect 10004 -3156 10036 -3124
rect 10004 -3205 10036 -3204
rect 10004 -3235 10005 -3205
rect 10005 -3235 10035 -3205
rect 10035 -3235 10036 -3205
rect 10004 -3236 10036 -3235
rect 10004 -3285 10036 -3284
rect 10004 -3315 10005 -3285
rect 10005 -3315 10035 -3285
rect 10035 -3315 10036 -3285
rect 10004 -3316 10036 -3315
rect 10004 -3396 10036 -3364
rect 10004 -3476 10036 -3444
rect 10004 -3525 10036 -3524
rect 10004 -3555 10005 -3525
rect 10005 -3555 10035 -3525
rect 10035 -3555 10036 -3525
rect 10004 -3556 10036 -3555
rect 10004 -3605 10036 -3604
rect 10004 -3635 10005 -3605
rect 10005 -3635 10035 -3605
rect 10035 -3635 10036 -3605
rect 10004 -3636 10036 -3635
rect 10004 -3685 10036 -3684
rect 10004 -3715 10005 -3685
rect 10005 -3715 10035 -3685
rect 10035 -3715 10036 -3685
rect 10004 -3716 10036 -3715
rect 10084 1035 10116 1036
rect 10084 1005 10085 1035
rect 10085 1005 10115 1035
rect 10115 1005 10116 1035
rect 10084 1004 10116 1005
rect 10084 955 10116 956
rect 10084 925 10085 955
rect 10085 925 10115 955
rect 10115 925 10116 955
rect 10084 924 10116 925
rect 10084 875 10116 876
rect 10084 845 10085 875
rect 10085 845 10115 875
rect 10115 845 10116 875
rect 10084 844 10116 845
rect 10084 764 10116 796
rect 10084 684 10116 716
rect 10084 635 10116 636
rect 10084 605 10085 635
rect 10085 605 10115 635
rect 10115 605 10116 635
rect 10084 604 10116 605
rect 10084 555 10116 556
rect 10084 525 10085 555
rect 10085 525 10115 555
rect 10115 525 10116 555
rect 10084 524 10116 525
rect 10084 444 10116 476
rect 10084 395 10116 396
rect 10084 365 10085 395
rect 10085 365 10115 395
rect 10115 365 10116 395
rect 10084 364 10116 365
rect 10084 284 10116 316
rect 10084 235 10116 236
rect 10084 205 10085 235
rect 10085 205 10115 235
rect 10115 205 10116 235
rect 10084 204 10116 205
rect 10084 124 10116 156
rect 10084 75 10116 76
rect 10084 45 10085 75
rect 10085 45 10115 75
rect 10115 45 10116 75
rect 10084 44 10116 45
rect 10084 -5 10116 -4
rect 10084 -35 10085 -5
rect 10085 -35 10115 -5
rect 10115 -35 10116 -5
rect 10084 -36 10116 -35
rect 10084 -85 10116 -84
rect 10084 -115 10085 -85
rect 10085 -115 10115 -85
rect 10115 -115 10116 -85
rect 10084 -116 10116 -115
rect 10084 -165 10116 -164
rect 10084 -195 10085 -165
rect 10085 -195 10115 -165
rect 10115 -195 10116 -165
rect 10084 -196 10116 -195
rect 10084 -245 10116 -244
rect 10084 -275 10085 -245
rect 10085 -275 10115 -245
rect 10115 -275 10116 -245
rect 10084 -276 10116 -275
rect 10084 -325 10116 -324
rect 10084 -355 10085 -325
rect 10085 -355 10115 -325
rect 10115 -355 10116 -325
rect 10084 -356 10116 -355
rect 10084 -436 10116 -404
rect 10084 -485 10116 -484
rect 10084 -515 10085 -485
rect 10085 -515 10115 -485
rect 10115 -515 10116 -485
rect 10084 -516 10116 -515
rect 10084 -596 10116 -564
rect 10084 -645 10116 -644
rect 10084 -675 10085 -645
rect 10085 -675 10115 -645
rect 10115 -675 10116 -645
rect 10084 -676 10116 -675
rect 10084 -756 10116 -724
rect 10084 -805 10116 -804
rect 10084 -835 10085 -805
rect 10085 -835 10115 -805
rect 10115 -835 10116 -805
rect 10084 -836 10116 -835
rect 10084 -885 10116 -884
rect 10084 -915 10085 -885
rect 10085 -915 10115 -885
rect 10115 -915 10116 -885
rect 10084 -916 10116 -915
rect 10084 -996 10116 -964
rect 10084 -1076 10116 -1044
rect 10084 -1125 10116 -1124
rect 10084 -1155 10085 -1125
rect 10085 -1155 10115 -1125
rect 10115 -1155 10116 -1125
rect 10084 -1156 10116 -1155
rect 10084 -1205 10116 -1204
rect 10084 -1235 10085 -1205
rect 10085 -1235 10115 -1205
rect 10115 -1235 10116 -1205
rect 10084 -1236 10116 -1235
rect 10084 -1285 10116 -1284
rect 10084 -1315 10085 -1285
rect 10085 -1315 10115 -1285
rect 10115 -1315 10116 -1285
rect 10084 -1316 10116 -1315
rect 10084 -1365 10116 -1364
rect 10084 -1395 10085 -1365
rect 10085 -1395 10115 -1365
rect 10115 -1395 10116 -1365
rect 10084 -1396 10116 -1395
rect 10084 -1445 10116 -1444
rect 10084 -1475 10085 -1445
rect 10085 -1475 10115 -1445
rect 10115 -1475 10116 -1445
rect 10084 -1476 10116 -1475
rect 10084 -1525 10116 -1524
rect 10084 -1555 10085 -1525
rect 10085 -1555 10115 -1525
rect 10115 -1555 10116 -1525
rect 10084 -1556 10116 -1555
rect 10084 -1636 10116 -1604
rect 10084 -1716 10116 -1684
rect 10084 -1765 10116 -1764
rect 10084 -1795 10085 -1765
rect 10085 -1795 10115 -1765
rect 10115 -1795 10116 -1765
rect 10084 -1796 10116 -1795
rect 10084 -1845 10116 -1844
rect 10084 -1875 10085 -1845
rect 10085 -1875 10115 -1845
rect 10115 -1875 10116 -1845
rect 10084 -1876 10116 -1875
rect 10084 -1956 10116 -1924
rect 10084 -2005 10116 -2004
rect 10084 -2035 10085 -2005
rect 10085 -2035 10115 -2005
rect 10115 -2035 10116 -2005
rect 10084 -2036 10116 -2035
rect 10084 -2116 10116 -2084
rect 10084 -2165 10116 -2164
rect 10084 -2195 10085 -2165
rect 10085 -2195 10115 -2165
rect 10115 -2195 10116 -2165
rect 10084 -2196 10116 -2195
rect 10084 -2276 10116 -2244
rect 10084 -2325 10116 -2324
rect 10084 -2355 10085 -2325
rect 10085 -2355 10115 -2325
rect 10115 -2355 10116 -2325
rect 10084 -2356 10116 -2355
rect 10084 -2405 10116 -2404
rect 10084 -2435 10085 -2405
rect 10085 -2435 10115 -2405
rect 10115 -2435 10116 -2405
rect 10084 -2436 10116 -2435
rect 10084 -2485 10116 -2484
rect 10084 -2515 10085 -2485
rect 10085 -2515 10115 -2485
rect 10115 -2515 10116 -2485
rect 10084 -2516 10116 -2515
rect 10084 -2565 10116 -2564
rect 10084 -2595 10085 -2565
rect 10085 -2595 10115 -2565
rect 10115 -2595 10116 -2565
rect 10084 -2596 10116 -2595
rect 10084 -2645 10116 -2644
rect 10084 -2675 10085 -2645
rect 10085 -2675 10115 -2645
rect 10115 -2675 10116 -2645
rect 10084 -2676 10116 -2675
rect 10084 -2725 10116 -2724
rect 10084 -2755 10085 -2725
rect 10085 -2755 10115 -2725
rect 10115 -2755 10116 -2725
rect 10084 -2756 10116 -2755
rect 10084 -2836 10116 -2804
rect 10084 -2885 10116 -2884
rect 10084 -2915 10085 -2885
rect 10085 -2915 10115 -2885
rect 10115 -2915 10116 -2885
rect 10084 -2916 10116 -2915
rect 10084 -2996 10116 -2964
rect 10084 -3045 10116 -3044
rect 10084 -3075 10085 -3045
rect 10085 -3075 10115 -3045
rect 10115 -3075 10116 -3045
rect 10084 -3076 10116 -3075
rect 10084 -3156 10116 -3124
rect 10084 -3205 10116 -3204
rect 10084 -3235 10085 -3205
rect 10085 -3235 10115 -3205
rect 10115 -3235 10116 -3205
rect 10084 -3236 10116 -3235
rect 10084 -3285 10116 -3284
rect 10084 -3315 10085 -3285
rect 10085 -3315 10115 -3285
rect 10115 -3315 10116 -3285
rect 10084 -3316 10116 -3315
rect 10084 -3396 10116 -3364
rect 10084 -3476 10116 -3444
rect 10084 -3525 10116 -3524
rect 10084 -3555 10085 -3525
rect 10085 -3555 10115 -3525
rect 10115 -3555 10116 -3525
rect 10084 -3556 10116 -3555
rect 10084 -3605 10116 -3604
rect 10084 -3635 10085 -3605
rect 10085 -3635 10115 -3605
rect 10115 -3635 10116 -3605
rect 10084 -3636 10116 -3635
rect 10084 -3685 10116 -3684
rect 10084 -3715 10085 -3685
rect 10085 -3715 10115 -3685
rect 10115 -3715 10116 -3685
rect 10084 -3716 10116 -3715
rect 10164 1035 10196 1036
rect 10164 1005 10165 1035
rect 10165 1005 10195 1035
rect 10195 1005 10196 1035
rect 10164 1004 10196 1005
rect 10164 955 10196 956
rect 10164 925 10165 955
rect 10165 925 10195 955
rect 10195 925 10196 955
rect 10164 924 10196 925
rect 10164 875 10196 876
rect 10164 845 10165 875
rect 10165 845 10195 875
rect 10195 845 10196 875
rect 10164 844 10196 845
rect 10164 764 10196 796
rect 10164 684 10196 716
rect 10164 635 10196 636
rect 10164 605 10165 635
rect 10165 605 10195 635
rect 10195 605 10196 635
rect 10164 604 10196 605
rect 10164 555 10196 556
rect 10164 525 10165 555
rect 10165 525 10195 555
rect 10195 525 10196 555
rect 10164 524 10196 525
rect 10164 444 10196 476
rect 10164 395 10196 396
rect 10164 365 10165 395
rect 10165 365 10195 395
rect 10195 365 10196 395
rect 10164 364 10196 365
rect 10164 284 10196 316
rect 10164 235 10196 236
rect 10164 205 10165 235
rect 10165 205 10195 235
rect 10195 205 10196 235
rect 10164 204 10196 205
rect 10164 124 10196 156
rect 10164 75 10196 76
rect 10164 45 10165 75
rect 10165 45 10195 75
rect 10195 45 10196 75
rect 10164 44 10196 45
rect 10164 -5 10196 -4
rect 10164 -35 10165 -5
rect 10165 -35 10195 -5
rect 10195 -35 10196 -5
rect 10164 -36 10196 -35
rect 10164 -85 10196 -84
rect 10164 -115 10165 -85
rect 10165 -115 10195 -85
rect 10195 -115 10196 -85
rect 10164 -116 10196 -115
rect 10164 -165 10196 -164
rect 10164 -195 10165 -165
rect 10165 -195 10195 -165
rect 10195 -195 10196 -165
rect 10164 -196 10196 -195
rect 10164 -245 10196 -244
rect 10164 -275 10165 -245
rect 10165 -275 10195 -245
rect 10195 -275 10196 -245
rect 10164 -276 10196 -275
rect 10164 -325 10196 -324
rect 10164 -355 10165 -325
rect 10165 -355 10195 -325
rect 10195 -355 10196 -325
rect 10164 -356 10196 -355
rect 10164 -436 10196 -404
rect 10164 -485 10196 -484
rect 10164 -515 10165 -485
rect 10165 -515 10195 -485
rect 10195 -515 10196 -485
rect 10164 -516 10196 -515
rect 10164 -596 10196 -564
rect 10164 -645 10196 -644
rect 10164 -675 10165 -645
rect 10165 -675 10195 -645
rect 10195 -675 10196 -645
rect 10164 -676 10196 -675
rect 10164 -756 10196 -724
rect 10164 -805 10196 -804
rect 10164 -835 10165 -805
rect 10165 -835 10195 -805
rect 10195 -835 10196 -805
rect 10164 -836 10196 -835
rect 10164 -885 10196 -884
rect 10164 -915 10165 -885
rect 10165 -915 10195 -885
rect 10195 -915 10196 -885
rect 10164 -916 10196 -915
rect 10164 -996 10196 -964
rect 10164 -1076 10196 -1044
rect 10164 -1125 10196 -1124
rect 10164 -1155 10165 -1125
rect 10165 -1155 10195 -1125
rect 10195 -1155 10196 -1125
rect 10164 -1156 10196 -1155
rect 10164 -1205 10196 -1204
rect 10164 -1235 10165 -1205
rect 10165 -1235 10195 -1205
rect 10195 -1235 10196 -1205
rect 10164 -1236 10196 -1235
rect 10164 -1285 10196 -1284
rect 10164 -1315 10165 -1285
rect 10165 -1315 10195 -1285
rect 10195 -1315 10196 -1285
rect 10164 -1316 10196 -1315
rect 10164 -1365 10196 -1364
rect 10164 -1395 10165 -1365
rect 10165 -1395 10195 -1365
rect 10195 -1395 10196 -1365
rect 10164 -1396 10196 -1395
rect 10164 -1445 10196 -1444
rect 10164 -1475 10165 -1445
rect 10165 -1475 10195 -1445
rect 10195 -1475 10196 -1445
rect 10164 -1476 10196 -1475
rect 10164 -1525 10196 -1524
rect 10164 -1555 10165 -1525
rect 10165 -1555 10195 -1525
rect 10195 -1555 10196 -1525
rect 10164 -1556 10196 -1555
rect 10164 -1636 10196 -1604
rect 10164 -1716 10196 -1684
rect 10164 -1765 10196 -1764
rect 10164 -1795 10165 -1765
rect 10165 -1795 10195 -1765
rect 10195 -1795 10196 -1765
rect 10164 -1796 10196 -1795
rect 10164 -1845 10196 -1844
rect 10164 -1875 10165 -1845
rect 10165 -1875 10195 -1845
rect 10195 -1875 10196 -1845
rect 10164 -1876 10196 -1875
rect 10164 -1956 10196 -1924
rect 10164 -2005 10196 -2004
rect 10164 -2035 10165 -2005
rect 10165 -2035 10195 -2005
rect 10195 -2035 10196 -2005
rect 10164 -2036 10196 -2035
rect 10164 -2116 10196 -2084
rect 10164 -2165 10196 -2164
rect 10164 -2195 10165 -2165
rect 10165 -2195 10195 -2165
rect 10195 -2195 10196 -2165
rect 10164 -2196 10196 -2195
rect 10164 -2276 10196 -2244
rect 10164 -2325 10196 -2324
rect 10164 -2355 10165 -2325
rect 10165 -2355 10195 -2325
rect 10195 -2355 10196 -2325
rect 10164 -2356 10196 -2355
rect 10164 -2405 10196 -2404
rect 10164 -2435 10165 -2405
rect 10165 -2435 10195 -2405
rect 10195 -2435 10196 -2405
rect 10164 -2436 10196 -2435
rect 10164 -2485 10196 -2484
rect 10164 -2515 10165 -2485
rect 10165 -2515 10195 -2485
rect 10195 -2515 10196 -2485
rect 10164 -2516 10196 -2515
rect 10164 -2565 10196 -2564
rect 10164 -2595 10165 -2565
rect 10165 -2595 10195 -2565
rect 10195 -2595 10196 -2565
rect 10164 -2596 10196 -2595
rect 10164 -2645 10196 -2644
rect 10164 -2675 10165 -2645
rect 10165 -2675 10195 -2645
rect 10195 -2675 10196 -2645
rect 10164 -2676 10196 -2675
rect 10164 -2725 10196 -2724
rect 10164 -2755 10165 -2725
rect 10165 -2755 10195 -2725
rect 10195 -2755 10196 -2725
rect 10164 -2756 10196 -2755
rect 10164 -2836 10196 -2804
rect 10164 -2885 10196 -2884
rect 10164 -2915 10165 -2885
rect 10165 -2915 10195 -2885
rect 10195 -2915 10196 -2885
rect 10164 -2916 10196 -2915
rect 10164 -2996 10196 -2964
rect 10164 -3045 10196 -3044
rect 10164 -3075 10165 -3045
rect 10165 -3075 10195 -3045
rect 10195 -3075 10196 -3045
rect 10164 -3076 10196 -3075
rect 10164 -3156 10196 -3124
rect 10164 -3205 10196 -3204
rect 10164 -3235 10165 -3205
rect 10165 -3235 10195 -3205
rect 10195 -3235 10196 -3205
rect 10164 -3236 10196 -3235
rect 10164 -3285 10196 -3284
rect 10164 -3315 10165 -3285
rect 10165 -3315 10195 -3285
rect 10195 -3315 10196 -3285
rect 10164 -3316 10196 -3315
rect 10164 -3396 10196 -3364
rect 10164 -3476 10196 -3444
rect 10164 -3525 10196 -3524
rect 10164 -3555 10165 -3525
rect 10165 -3555 10195 -3525
rect 10195 -3555 10196 -3525
rect 10164 -3556 10196 -3555
rect 10164 -3605 10196 -3604
rect 10164 -3635 10165 -3605
rect 10165 -3635 10195 -3605
rect 10195 -3635 10196 -3605
rect 10164 -3636 10196 -3635
rect 10164 -3685 10196 -3684
rect 10164 -3715 10165 -3685
rect 10165 -3715 10195 -3685
rect 10195 -3715 10196 -3685
rect 10164 -3716 10196 -3715
rect 10244 1035 10276 1036
rect 10244 1005 10245 1035
rect 10245 1005 10275 1035
rect 10275 1005 10276 1035
rect 10244 1004 10276 1005
rect 10244 955 10276 956
rect 10244 925 10245 955
rect 10245 925 10275 955
rect 10275 925 10276 955
rect 10244 924 10276 925
rect 10244 875 10276 876
rect 10244 845 10245 875
rect 10245 845 10275 875
rect 10275 845 10276 875
rect 10244 844 10276 845
rect 10244 764 10276 796
rect 10244 684 10276 716
rect 10244 635 10276 636
rect 10244 605 10245 635
rect 10245 605 10275 635
rect 10275 605 10276 635
rect 10244 604 10276 605
rect 10244 555 10276 556
rect 10244 525 10245 555
rect 10245 525 10275 555
rect 10275 525 10276 555
rect 10244 524 10276 525
rect 10244 444 10276 476
rect 10244 395 10276 396
rect 10244 365 10245 395
rect 10245 365 10275 395
rect 10275 365 10276 395
rect 10244 364 10276 365
rect 10244 284 10276 316
rect 10244 235 10276 236
rect 10244 205 10245 235
rect 10245 205 10275 235
rect 10275 205 10276 235
rect 10244 204 10276 205
rect 10244 124 10276 156
rect 10244 75 10276 76
rect 10244 45 10245 75
rect 10245 45 10275 75
rect 10275 45 10276 75
rect 10244 44 10276 45
rect 10244 -5 10276 -4
rect 10244 -35 10245 -5
rect 10245 -35 10275 -5
rect 10275 -35 10276 -5
rect 10244 -36 10276 -35
rect 10244 -85 10276 -84
rect 10244 -115 10245 -85
rect 10245 -115 10275 -85
rect 10275 -115 10276 -85
rect 10244 -116 10276 -115
rect 10244 -165 10276 -164
rect 10244 -195 10245 -165
rect 10245 -195 10275 -165
rect 10275 -195 10276 -165
rect 10244 -196 10276 -195
rect 10244 -245 10276 -244
rect 10244 -275 10245 -245
rect 10245 -275 10275 -245
rect 10275 -275 10276 -245
rect 10244 -276 10276 -275
rect 10244 -325 10276 -324
rect 10244 -355 10245 -325
rect 10245 -355 10275 -325
rect 10275 -355 10276 -325
rect 10244 -356 10276 -355
rect 10244 -436 10276 -404
rect 10244 -485 10276 -484
rect 10244 -515 10245 -485
rect 10245 -515 10275 -485
rect 10275 -515 10276 -485
rect 10244 -516 10276 -515
rect 10244 -596 10276 -564
rect 10244 -645 10276 -644
rect 10244 -675 10245 -645
rect 10245 -675 10275 -645
rect 10275 -675 10276 -645
rect 10244 -676 10276 -675
rect 10244 -756 10276 -724
rect 10244 -805 10276 -804
rect 10244 -835 10245 -805
rect 10245 -835 10275 -805
rect 10275 -835 10276 -805
rect 10244 -836 10276 -835
rect 10244 -885 10276 -884
rect 10244 -915 10245 -885
rect 10245 -915 10275 -885
rect 10275 -915 10276 -885
rect 10244 -916 10276 -915
rect 10244 -996 10276 -964
rect 10244 -1076 10276 -1044
rect 10244 -1125 10276 -1124
rect 10244 -1155 10245 -1125
rect 10245 -1155 10275 -1125
rect 10275 -1155 10276 -1125
rect 10244 -1156 10276 -1155
rect 10244 -1205 10276 -1204
rect 10244 -1235 10245 -1205
rect 10245 -1235 10275 -1205
rect 10275 -1235 10276 -1205
rect 10244 -1236 10276 -1235
rect 10244 -1285 10276 -1284
rect 10244 -1315 10245 -1285
rect 10245 -1315 10275 -1285
rect 10275 -1315 10276 -1285
rect 10244 -1316 10276 -1315
rect 10244 -1365 10276 -1364
rect 10244 -1395 10245 -1365
rect 10245 -1395 10275 -1365
rect 10275 -1395 10276 -1365
rect 10244 -1396 10276 -1395
rect 10244 -1445 10276 -1444
rect 10244 -1475 10245 -1445
rect 10245 -1475 10275 -1445
rect 10275 -1475 10276 -1445
rect 10244 -1476 10276 -1475
rect 10244 -1525 10276 -1524
rect 10244 -1555 10245 -1525
rect 10245 -1555 10275 -1525
rect 10275 -1555 10276 -1525
rect 10244 -1556 10276 -1555
rect 10244 -1636 10276 -1604
rect 10244 -1716 10276 -1684
rect 10244 -1765 10276 -1764
rect 10244 -1795 10245 -1765
rect 10245 -1795 10275 -1765
rect 10275 -1795 10276 -1765
rect 10244 -1796 10276 -1795
rect 10244 -1845 10276 -1844
rect 10244 -1875 10245 -1845
rect 10245 -1875 10275 -1845
rect 10275 -1875 10276 -1845
rect 10244 -1876 10276 -1875
rect 10244 -1956 10276 -1924
rect 10244 -2005 10276 -2004
rect 10244 -2035 10245 -2005
rect 10245 -2035 10275 -2005
rect 10275 -2035 10276 -2005
rect 10244 -2036 10276 -2035
rect 10244 -2116 10276 -2084
rect 10244 -2165 10276 -2164
rect 10244 -2195 10245 -2165
rect 10245 -2195 10275 -2165
rect 10275 -2195 10276 -2165
rect 10244 -2196 10276 -2195
rect 10244 -2276 10276 -2244
rect 10244 -2325 10276 -2324
rect 10244 -2355 10245 -2325
rect 10245 -2355 10275 -2325
rect 10275 -2355 10276 -2325
rect 10244 -2356 10276 -2355
rect 10244 -2405 10276 -2404
rect 10244 -2435 10245 -2405
rect 10245 -2435 10275 -2405
rect 10275 -2435 10276 -2405
rect 10244 -2436 10276 -2435
rect 10244 -2485 10276 -2484
rect 10244 -2515 10245 -2485
rect 10245 -2515 10275 -2485
rect 10275 -2515 10276 -2485
rect 10244 -2516 10276 -2515
rect 10244 -2565 10276 -2564
rect 10244 -2595 10245 -2565
rect 10245 -2595 10275 -2565
rect 10275 -2595 10276 -2565
rect 10244 -2596 10276 -2595
rect 10244 -2645 10276 -2644
rect 10244 -2675 10245 -2645
rect 10245 -2675 10275 -2645
rect 10275 -2675 10276 -2645
rect 10244 -2676 10276 -2675
rect 10244 -2725 10276 -2724
rect 10244 -2755 10245 -2725
rect 10245 -2755 10275 -2725
rect 10275 -2755 10276 -2725
rect 10244 -2756 10276 -2755
rect 10244 -2836 10276 -2804
rect 10244 -2885 10276 -2884
rect 10244 -2915 10245 -2885
rect 10245 -2915 10275 -2885
rect 10275 -2915 10276 -2885
rect 10244 -2916 10276 -2915
rect 10244 -2996 10276 -2964
rect 10244 -3045 10276 -3044
rect 10244 -3075 10245 -3045
rect 10245 -3075 10275 -3045
rect 10275 -3075 10276 -3045
rect 10244 -3076 10276 -3075
rect 10244 -3156 10276 -3124
rect 10244 -3205 10276 -3204
rect 10244 -3235 10245 -3205
rect 10245 -3235 10275 -3205
rect 10275 -3235 10276 -3205
rect 10244 -3236 10276 -3235
rect 10244 -3285 10276 -3284
rect 10244 -3315 10245 -3285
rect 10245 -3315 10275 -3285
rect 10275 -3315 10276 -3285
rect 10244 -3316 10276 -3315
rect 10244 -3396 10276 -3364
rect 10244 -3476 10276 -3444
rect 10244 -3525 10276 -3524
rect 10244 -3555 10245 -3525
rect 10245 -3555 10275 -3525
rect 10275 -3555 10276 -3525
rect 10244 -3556 10276 -3555
rect 10244 -3605 10276 -3604
rect 10244 -3635 10245 -3605
rect 10245 -3635 10275 -3605
rect 10275 -3635 10276 -3605
rect 10244 -3636 10276 -3635
rect 10244 -3685 10276 -3684
rect 10244 -3715 10245 -3685
rect 10245 -3715 10275 -3685
rect 10275 -3715 10276 -3685
rect 10244 -3716 10276 -3715
rect 10324 1035 10356 1036
rect 10324 1005 10325 1035
rect 10325 1005 10355 1035
rect 10355 1005 10356 1035
rect 10324 1004 10356 1005
rect 10324 955 10356 956
rect 10324 925 10325 955
rect 10325 925 10355 955
rect 10355 925 10356 955
rect 10324 924 10356 925
rect 10324 875 10356 876
rect 10324 845 10325 875
rect 10325 845 10355 875
rect 10355 845 10356 875
rect 10324 844 10356 845
rect 10324 764 10356 796
rect 10324 684 10356 716
rect 10324 635 10356 636
rect 10324 605 10325 635
rect 10325 605 10355 635
rect 10355 605 10356 635
rect 10324 604 10356 605
rect 10324 555 10356 556
rect 10324 525 10325 555
rect 10325 525 10355 555
rect 10355 525 10356 555
rect 10324 524 10356 525
rect 10324 444 10356 476
rect 10324 395 10356 396
rect 10324 365 10325 395
rect 10325 365 10355 395
rect 10355 365 10356 395
rect 10324 364 10356 365
rect 10324 284 10356 316
rect 10324 235 10356 236
rect 10324 205 10325 235
rect 10325 205 10355 235
rect 10355 205 10356 235
rect 10324 204 10356 205
rect 10324 124 10356 156
rect 10324 75 10356 76
rect 10324 45 10325 75
rect 10325 45 10355 75
rect 10355 45 10356 75
rect 10324 44 10356 45
rect 10324 -5 10356 -4
rect 10324 -35 10325 -5
rect 10325 -35 10355 -5
rect 10355 -35 10356 -5
rect 10324 -36 10356 -35
rect 10324 -85 10356 -84
rect 10324 -115 10325 -85
rect 10325 -115 10355 -85
rect 10355 -115 10356 -85
rect 10324 -116 10356 -115
rect 10324 -165 10356 -164
rect 10324 -195 10325 -165
rect 10325 -195 10355 -165
rect 10355 -195 10356 -165
rect 10324 -196 10356 -195
rect 10324 -245 10356 -244
rect 10324 -275 10325 -245
rect 10325 -275 10355 -245
rect 10355 -275 10356 -245
rect 10324 -276 10356 -275
rect 10324 -325 10356 -324
rect 10324 -355 10325 -325
rect 10325 -355 10355 -325
rect 10355 -355 10356 -325
rect 10324 -356 10356 -355
rect 10324 -436 10356 -404
rect 10324 -485 10356 -484
rect 10324 -515 10325 -485
rect 10325 -515 10355 -485
rect 10355 -515 10356 -485
rect 10324 -516 10356 -515
rect 10324 -596 10356 -564
rect 10324 -645 10356 -644
rect 10324 -675 10325 -645
rect 10325 -675 10355 -645
rect 10355 -675 10356 -645
rect 10324 -676 10356 -675
rect 10324 -756 10356 -724
rect 10324 -805 10356 -804
rect 10324 -835 10325 -805
rect 10325 -835 10355 -805
rect 10355 -835 10356 -805
rect 10324 -836 10356 -835
rect 10324 -885 10356 -884
rect 10324 -915 10325 -885
rect 10325 -915 10355 -885
rect 10355 -915 10356 -885
rect 10324 -916 10356 -915
rect 10324 -996 10356 -964
rect 10324 -1076 10356 -1044
rect 10324 -1125 10356 -1124
rect 10324 -1155 10325 -1125
rect 10325 -1155 10355 -1125
rect 10355 -1155 10356 -1125
rect 10324 -1156 10356 -1155
rect 10324 -1205 10356 -1204
rect 10324 -1235 10325 -1205
rect 10325 -1235 10355 -1205
rect 10355 -1235 10356 -1205
rect 10324 -1236 10356 -1235
rect 10324 -1285 10356 -1284
rect 10324 -1315 10325 -1285
rect 10325 -1315 10355 -1285
rect 10355 -1315 10356 -1285
rect 10324 -1316 10356 -1315
rect 10324 -1365 10356 -1364
rect 10324 -1395 10325 -1365
rect 10325 -1395 10355 -1365
rect 10355 -1395 10356 -1365
rect 10324 -1396 10356 -1395
rect 10324 -1445 10356 -1444
rect 10324 -1475 10325 -1445
rect 10325 -1475 10355 -1445
rect 10355 -1475 10356 -1445
rect 10324 -1476 10356 -1475
rect 10324 -1525 10356 -1524
rect 10324 -1555 10325 -1525
rect 10325 -1555 10355 -1525
rect 10355 -1555 10356 -1525
rect 10324 -1556 10356 -1555
rect 10324 -1636 10356 -1604
rect 10324 -1716 10356 -1684
rect 10324 -1765 10356 -1764
rect 10324 -1795 10325 -1765
rect 10325 -1795 10355 -1765
rect 10355 -1795 10356 -1765
rect 10324 -1796 10356 -1795
rect 10324 -1845 10356 -1844
rect 10324 -1875 10325 -1845
rect 10325 -1875 10355 -1845
rect 10355 -1875 10356 -1845
rect 10324 -1876 10356 -1875
rect 10324 -1956 10356 -1924
rect 10324 -2005 10356 -2004
rect 10324 -2035 10325 -2005
rect 10325 -2035 10355 -2005
rect 10355 -2035 10356 -2005
rect 10324 -2036 10356 -2035
rect 10324 -2116 10356 -2084
rect 10324 -2165 10356 -2164
rect 10324 -2195 10325 -2165
rect 10325 -2195 10355 -2165
rect 10355 -2195 10356 -2165
rect 10324 -2196 10356 -2195
rect 10324 -2276 10356 -2244
rect 10324 -2325 10356 -2324
rect 10324 -2355 10325 -2325
rect 10325 -2355 10355 -2325
rect 10355 -2355 10356 -2325
rect 10324 -2356 10356 -2355
rect 10324 -2405 10356 -2404
rect 10324 -2435 10325 -2405
rect 10325 -2435 10355 -2405
rect 10355 -2435 10356 -2405
rect 10324 -2436 10356 -2435
rect 10324 -2485 10356 -2484
rect 10324 -2515 10325 -2485
rect 10325 -2515 10355 -2485
rect 10355 -2515 10356 -2485
rect 10324 -2516 10356 -2515
rect 10324 -2565 10356 -2564
rect 10324 -2595 10325 -2565
rect 10325 -2595 10355 -2565
rect 10355 -2595 10356 -2565
rect 10324 -2596 10356 -2595
rect 10324 -2645 10356 -2644
rect 10324 -2675 10325 -2645
rect 10325 -2675 10355 -2645
rect 10355 -2675 10356 -2645
rect 10324 -2676 10356 -2675
rect 10324 -2725 10356 -2724
rect 10324 -2755 10325 -2725
rect 10325 -2755 10355 -2725
rect 10355 -2755 10356 -2725
rect 10324 -2756 10356 -2755
rect 10324 -2836 10356 -2804
rect 10324 -2885 10356 -2884
rect 10324 -2915 10325 -2885
rect 10325 -2915 10355 -2885
rect 10355 -2915 10356 -2885
rect 10324 -2916 10356 -2915
rect 10324 -2996 10356 -2964
rect 10324 -3045 10356 -3044
rect 10324 -3075 10325 -3045
rect 10325 -3075 10355 -3045
rect 10355 -3075 10356 -3045
rect 10324 -3076 10356 -3075
rect 10324 -3156 10356 -3124
rect 10324 -3205 10356 -3204
rect 10324 -3235 10325 -3205
rect 10325 -3235 10355 -3205
rect 10355 -3235 10356 -3205
rect 10324 -3236 10356 -3235
rect 10324 -3285 10356 -3284
rect 10324 -3315 10325 -3285
rect 10325 -3315 10355 -3285
rect 10355 -3315 10356 -3285
rect 10324 -3316 10356 -3315
rect 10324 -3396 10356 -3364
rect 10324 -3476 10356 -3444
rect 10324 -3525 10356 -3524
rect 10324 -3555 10325 -3525
rect 10325 -3555 10355 -3525
rect 10355 -3555 10356 -3525
rect 10324 -3556 10356 -3555
rect 10324 -3605 10356 -3604
rect 10324 -3635 10325 -3605
rect 10325 -3635 10355 -3605
rect 10355 -3635 10356 -3605
rect 10324 -3636 10356 -3635
rect 10324 -3685 10356 -3684
rect 10324 -3715 10325 -3685
rect 10325 -3715 10355 -3685
rect 10355 -3715 10356 -3685
rect 10324 -3716 10356 -3715
rect 10404 1035 10436 1036
rect 10404 1005 10405 1035
rect 10405 1005 10435 1035
rect 10435 1005 10436 1035
rect 10404 1004 10436 1005
rect 10404 955 10436 956
rect 10404 925 10405 955
rect 10405 925 10435 955
rect 10435 925 10436 955
rect 10404 924 10436 925
rect 10404 875 10436 876
rect 10404 845 10405 875
rect 10405 845 10435 875
rect 10435 845 10436 875
rect 10404 844 10436 845
rect 10404 764 10436 796
rect 10404 684 10436 716
rect 10404 635 10436 636
rect 10404 605 10405 635
rect 10405 605 10435 635
rect 10435 605 10436 635
rect 10404 604 10436 605
rect 10404 555 10436 556
rect 10404 525 10405 555
rect 10405 525 10435 555
rect 10435 525 10436 555
rect 10404 524 10436 525
rect 10404 444 10436 476
rect 10404 395 10436 396
rect 10404 365 10405 395
rect 10405 365 10435 395
rect 10435 365 10436 395
rect 10404 364 10436 365
rect 10404 284 10436 316
rect 10404 235 10436 236
rect 10404 205 10405 235
rect 10405 205 10435 235
rect 10435 205 10436 235
rect 10404 204 10436 205
rect 10404 124 10436 156
rect 10404 75 10436 76
rect 10404 45 10405 75
rect 10405 45 10435 75
rect 10435 45 10436 75
rect 10404 44 10436 45
rect 10404 -5 10436 -4
rect 10404 -35 10405 -5
rect 10405 -35 10435 -5
rect 10435 -35 10436 -5
rect 10404 -36 10436 -35
rect 10404 -85 10436 -84
rect 10404 -115 10405 -85
rect 10405 -115 10435 -85
rect 10435 -115 10436 -85
rect 10404 -116 10436 -115
rect 10404 -165 10436 -164
rect 10404 -195 10405 -165
rect 10405 -195 10435 -165
rect 10435 -195 10436 -165
rect 10404 -196 10436 -195
rect 10404 -245 10436 -244
rect 10404 -275 10405 -245
rect 10405 -275 10435 -245
rect 10435 -275 10436 -245
rect 10404 -276 10436 -275
rect 10404 -325 10436 -324
rect 10404 -355 10405 -325
rect 10405 -355 10435 -325
rect 10435 -355 10436 -325
rect 10404 -356 10436 -355
rect 10404 -436 10436 -404
rect 10404 -485 10436 -484
rect 10404 -515 10405 -485
rect 10405 -515 10435 -485
rect 10435 -515 10436 -485
rect 10404 -516 10436 -515
rect 10404 -596 10436 -564
rect 10404 -645 10436 -644
rect 10404 -675 10405 -645
rect 10405 -675 10435 -645
rect 10435 -675 10436 -645
rect 10404 -676 10436 -675
rect 10404 -756 10436 -724
rect 10404 -805 10436 -804
rect 10404 -835 10405 -805
rect 10405 -835 10435 -805
rect 10435 -835 10436 -805
rect 10404 -836 10436 -835
rect 10404 -885 10436 -884
rect 10404 -915 10405 -885
rect 10405 -915 10435 -885
rect 10435 -915 10436 -885
rect 10404 -916 10436 -915
rect 10404 -996 10436 -964
rect 10404 -1076 10436 -1044
rect 10404 -1125 10436 -1124
rect 10404 -1155 10405 -1125
rect 10405 -1155 10435 -1125
rect 10435 -1155 10436 -1125
rect 10404 -1156 10436 -1155
rect 10404 -1205 10436 -1204
rect 10404 -1235 10405 -1205
rect 10405 -1235 10435 -1205
rect 10435 -1235 10436 -1205
rect 10404 -1236 10436 -1235
rect 10404 -1285 10436 -1284
rect 10404 -1315 10405 -1285
rect 10405 -1315 10435 -1285
rect 10435 -1315 10436 -1285
rect 10404 -1316 10436 -1315
rect 10404 -1365 10436 -1364
rect 10404 -1395 10405 -1365
rect 10405 -1395 10435 -1365
rect 10435 -1395 10436 -1365
rect 10404 -1396 10436 -1395
rect 10404 -1445 10436 -1444
rect 10404 -1475 10405 -1445
rect 10405 -1475 10435 -1445
rect 10435 -1475 10436 -1445
rect 10404 -1476 10436 -1475
rect 10404 -1525 10436 -1524
rect 10404 -1555 10405 -1525
rect 10405 -1555 10435 -1525
rect 10435 -1555 10436 -1525
rect 10404 -1556 10436 -1555
rect 10404 -1636 10436 -1604
rect 10404 -1716 10436 -1684
rect 10404 -1765 10436 -1764
rect 10404 -1795 10405 -1765
rect 10405 -1795 10435 -1765
rect 10435 -1795 10436 -1765
rect 10404 -1796 10436 -1795
rect 10404 -1845 10436 -1844
rect 10404 -1875 10405 -1845
rect 10405 -1875 10435 -1845
rect 10435 -1875 10436 -1845
rect 10404 -1876 10436 -1875
rect 10404 -1956 10436 -1924
rect 10404 -2005 10436 -2004
rect 10404 -2035 10405 -2005
rect 10405 -2035 10435 -2005
rect 10435 -2035 10436 -2005
rect 10404 -2036 10436 -2035
rect 10404 -2116 10436 -2084
rect 10404 -2165 10436 -2164
rect 10404 -2195 10405 -2165
rect 10405 -2195 10435 -2165
rect 10435 -2195 10436 -2165
rect 10404 -2196 10436 -2195
rect 10404 -2276 10436 -2244
rect 10404 -2325 10436 -2324
rect 10404 -2355 10405 -2325
rect 10405 -2355 10435 -2325
rect 10435 -2355 10436 -2325
rect 10404 -2356 10436 -2355
rect 10404 -2405 10436 -2404
rect 10404 -2435 10405 -2405
rect 10405 -2435 10435 -2405
rect 10435 -2435 10436 -2405
rect 10404 -2436 10436 -2435
rect 10404 -2485 10436 -2484
rect 10404 -2515 10405 -2485
rect 10405 -2515 10435 -2485
rect 10435 -2515 10436 -2485
rect 10404 -2516 10436 -2515
rect 10404 -2565 10436 -2564
rect 10404 -2595 10405 -2565
rect 10405 -2595 10435 -2565
rect 10435 -2595 10436 -2565
rect 10404 -2596 10436 -2595
rect 10404 -2645 10436 -2644
rect 10404 -2675 10405 -2645
rect 10405 -2675 10435 -2645
rect 10435 -2675 10436 -2645
rect 10404 -2676 10436 -2675
rect 10404 -2725 10436 -2724
rect 10404 -2755 10405 -2725
rect 10405 -2755 10435 -2725
rect 10435 -2755 10436 -2725
rect 10404 -2756 10436 -2755
rect 10404 -2836 10436 -2804
rect 10404 -2885 10436 -2884
rect 10404 -2915 10405 -2885
rect 10405 -2915 10435 -2885
rect 10435 -2915 10436 -2885
rect 10404 -2916 10436 -2915
rect 10404 -2996 10436 -2964
rect 10404 -3045 10436 -3044
rect 10404 -3075 10405 -3045
rect 10405 -3075 10435 -3045
rect 10435 -3075 10436 -3045
rect 10404 -3076 10436 -3075
rect 10404 -3156 10436 -3124
rect 10404 -3205 10436 -3204
rect 10404 -3235 10405 -3205
rect 10405 -3235 10435 -3205
rect 10435 -3235 10436 -3205
rect 10404 -3236 10436 -3235
rect 10404 -3285 10436 -3284
rect 10404 -3315 10405 -3285
rect 10405 -3315 10435 -3285
rect 10435 -3315 10436 -3285
rect 10404 -3316 10436 -3315
rect 10404 -3396 10436 -3364
rect 10404 -3476 10436 -3444
rect 10404 -3525 10436 -3524
rect 10404 -3555 10405 -3525
rect 10405 -3555 10435 -3525
rect 10435 -3555 10436 -3525
rect 10404 -3556 10436 -3555
rect 10404 -3605 10436 -3604
rect 10404 -3635 10405 -3605
rect 10405 -3635 10435 -3605
rect 10435 -3635 10436 -3605
rect 10404 -3636 10436 -3635
rect 10404 -3685 10436 -3684
rect 10404 -3715 10405 -3685
rect 10405 -3715 10435 -3685
rect 10435 -3715 10436 -3685
rect 10404 -3716 10436 -3715
rect 10484 1035 10516 1036
rect 10484 1005 10485 1035
rect 10485 1005 10515 1035
rect 10515 1005 10516 1035
rect 10484 1004 10516 1005
rect 10484 955 10516 956
rect 10484 925 10485 955
rect 10485 925 10515 955
rect 10515 925 10516 955
rect 10484 924 10516 925
rect 10484 875 10516 876
rect 10484 845 10485 875
rect 10485 845 10515 875
rect 10515 845 10516 875
rect 10484 844 10516 845
rect 10484 764 10516 796
rect 10484 684 10516 716
rect 10484 635 10516 636
rect 10484 605 10485 635
rect 10485 605 10515 635
rect 10515 605 10516 635
rect 10484 604 10516 605
rect 10484 555 10516 556
rect 10484 525 10485 555
rect 10485 525 10515 555
rect 10515 525 10516 555
rect 10484 524 10516 525
rect 10484 444 10516 476
rect 10484 395 10516 396
rect 10484 365 10485 395
rect 10485 365 10515 395
rect 10515 365 10516 395
rect 10484 364 10516 365
rect 10484 284 10516 316
rect 10484 235 10516 236
rect 10484 205 10485 235
rect 10485 205 10515 235
rect 10515 205 10516 235
rect 10484 204 10516 205
rect 10484 124 10516 156
rect 10484 75 10516 76
rect 10484 45 10485 75
rect 10485 45 10515 75
rect 10515 45 10516 75
rect 10484 44 10516 45
rect 10484 -5 10516 -4
rect 10484 -35 10485 -5
rect 10485 -35 10515 -5
rect 10515 -35 10516 -5
rect 10484 -36 10516 -35
rect 10484 -85 10516 -84
rect 10484 -115 10485 -85
rect 10485 -115 10515 -85
rect 10515 -115 10516 -85
rect 10484 -116 10516 -115
rect 10484 -165 10516 -164
rect 10484 -195 10485 -165
rect 10485 -195 10515 -165
rect 10515 -195 10516 -165
rect 10484 -196 10516 -195
rect 10484 -245 10516 -244
rect 10484 -275 10485 -245
rect 10485 -275 10515 -245
rect 10515 -275 10516 -245
rect 10484 -276 10516 -275
rect 10484 -325 10516 -324
rect 10484 -355 10485 -325
rect 10485 -355 10515 -325
rect 10515 -355 10516 -325
rect 10484 -356 10516 -355
rect 10484 -436 10516 -404
rect 10484 -485 10516 -484
rect 10484 -515 10485 -485
rect 10485 -515 10515 -485
rect 10515 -515 10516 -485
rect 10484 -516 10516 -515
rect 10484 -596 10516 -564
rect 10484 -645 10516 -644
rect 10484 -675 10485 -645
rect 10485 -675 10515 -645
rect 10515 -675 10516 -645
rect 10484 -676 10516 -675
rect 10484 -756 10516 -724
rect 10484 -805 10516 -804
rect 10484 -835 10485 -805
rect 10485 -835 10515 -805
rect 10515 -835 10516 -805
rect 10484 -836 10516 -835
rect 10484 -885 10516 -884
rect 10484 -915 10485 -885
rect 10485 -915 10515 -885
rect 10515 -915 10516 -885
rect 10484 -916 10516 -915
rect 10484 -996 10516 -964
rect 10484 -1076 10516 -1044
rect 10484 -1125 10516 -1124
rect 10484 -1155 10485 -1125
rect 10485 -1155 10515 -1125
rect 10515 -1155 10516 -1125
rect 10484 -1156 10516 -1155
rect 10484 -1205 10516 -1204
rect 10484 -1235 10485 -1205
rect 10485 -1235 10515 -1205
rect 10515 -1235 10516 -1205
rect 10484 -1236 10516 -1235
rect 10484 -1285 10516 -1284
rect 10484 -1315 10485 -1285
rect 10485 -1315 10515 -1285
rect 10515 -1315 10516 -1285
rect 10484 -1316 10516 -1315
rect 10484 -1365 10516 -1364
rect 10484 -1395 10485 -1365
rect 10485 -1395 10515 -1365
rect 10515 -1395 10516 -1365
rect 10484 -1396 10516 -1395
rect 10484 -1445 10516 -1444
rect 10484 -1475 10485 -1445
rect 10485 -1475 10515 -1445
rect 10515 -1475 10516 -1445
rect 10484 -1476 10516 -1475
rect 10484 -1525 10516 -1524
rect 10484 -1555 10485 -1525
rect 10485 -1555 10515 -1525
rect 10515 -1555 10516 -1525
rect 10484 -1556 10516 -1555
rect 10484 -1636 10516 -1604
rect 10484 -1716 10516 -1684
rect 10484 -1765 10516 -1764
rect 10484 -1795 10485 -1765
rect 10485 -1795 10515 -1765
rect 10515 -1795 10516 -1765
rect 10484 -1796 10516 -1795
rect 10484 -1845 10516 -1844
rect 10484 -1875 10485 -1845
rect 10485 -1875 10515 -1845
rect 10515 -1875 10516 -1845
rect 10484 -1876 10516 -1875
rect 10484 -1956 10516 -1924
rect 10484 -2005 10516 -2004
rect 10484 -2035 10485 -2005
rect 10485 -2035 10515 -2005
rect 10515 -2035 10516 -2005
rect 10484 -2036 10516 -2035
rect 10484 -2116 10516 -2084
rect 10484 -2165 10516 -2164
rect 10484 -2195 10485 -2165
rect 10485 -2195 10515 -2165
rect 10515 -2195 10516 -2165
rect 10484 -2196 10516 -2195
rect 10484 -2276 10516 -2244
rect 10484 -2325 10516 -2324
rect 10484 -2355 10485 -2325
rect 10485 -2355 10515 -2325
rect 10515 -2355 10516 -2325
rect 10484 -2356 10516 -2355
rect 10484 -2405 10516 -2404
rect 10484 -2435 10485 -2405
rect 10485 -2435 10515 -2405
rect 10515 -2435 10516 -2405
rect 10484 -2436 10516 -2435
rect 10484 -2485 10516 -2484
rect 10484 -2515 10485 -2485
rect 10485 -2515 10515 -2485
rect 10515 -2515 10516 -2485
rect 10484 -2516 10516 -2515
rect 10484 -2565 10516 -2564
rect 10484 -2595 10485 -2565
rect 10485 -2595 10515 -2565
rect 10515 -2595 10516 -2565
rect 10484 -2596 10516 -2595
rect 10484 -2645 10516 -2644
rect 10484 -2675 10485 -2645
rect 10485 -2675 10515 -2645
rect 10515 -2675 10516 -2645
rect 10484 -2676 10516 -2675
rect 10484 -2725 10516 -2724
rect 10484 -2755 10485 -2725
rect 10485 -2755 10515 -2725
rect 10515 -2755 10516 -2725
rect 10484 -2756 10516 -2755
rect 10484 -2836 10516 -2804
rect 10484 -2885 10516 -2884
rect 10484 -2915 10485 -2885
rect 10485 -2915 10515 -2885
rect 10515 -2915 10516 -2885
rect 10484 -2916 10516 -2915
rect 10484 -2996 10516 -2964
rect 10484 -3045 10516 -3044
rect 10484 -3075 10485 -3045
rect 10485 -3075 10515 -3045
rect 10515 -3075 10516 -3045
rect 10484 -3076 10516 -3075
rect 10484 -3156 10516 -3124
rect 10484 -3205 10516 -3204
rect 10484 -3235 10485 -3205
rect 10485 -3235 10515 -3205
rect 10515 -3235 10516 -3205
rect 10484 -3236 10516 -3235
rect 10484 -3285 10516 -3284
rect 10484 -3315 10485 -3285
rect 10485 -3315 10515 -3285
rect 10515 -3315 10516 -3285
rect 10484 -3316 10516 -3315
rect 10484 -3396 10516 -3364
rect 10484 -3476 10516 -3444
rect 10484 -3525 10516 -3524
rect 10484 -3555 10485 -3525
rect 10485 -3555 10515 -3525
rect 10515 -3555 10516 -3525
rect 10484 -3556 10516 -3555
rect 10484 -3605 10516 -3604
rect 10484 -3635 10485 -3605
rect 10485 -3635 10515 -3605
rect 10515 -3635 10516 -3605
rect 10484 -3636 10516 -3635
rect 10484 -3685 10516 -3684
rect 10484 -3715 10485 -3685
rect 10485 -3715 10515 -3685
rect 10515 -3715 10516 -3685
rect 10484 -3716 10516 -3715
rect 10564 -165 10596 -164
rect 10564 -195 10565 -165
rect 10565 -195 10595 -165
rect 10595 -195 10596 -165
rect 10564 -196 10596 -195
rect 10564 -245 10596 -244
rect 10564 -275 10565 -245
rect 10565 -275 10595 -245
rect 10595 -275 10596 -245
rect 10564 -276 10596 -275
rect 10564 -325 10596 -324
rect 10564 -355 10565 -325
rect 10565 -355 10595 -325
rect 10595 -355 10596 -325
rect 10564 -356 10596 -355
rect 10564 -436 10596 -404
rect 10564 -485 10596 -484
rect 10564 -515 10565 -485
rect 10565 -515 10595 -485
rect 10595 -515 10596 -485
rect 10564 -516 10596 -515
rect 10564 -596 10596 -564
rect 10564 -645 10596 -644
rect 10564 -675 10565 -645
rect 10565 -675 10595 -645
rect 10595 -675 10596 -645
rect 10564 -676 10596 -675
rect 10564 -756 10596 -724
rect 10564 -805 10596 -804
rect 10564 -835 10565 -805
rect 10565 -835 10595 -805
rect 10595 -835 10596 -805
rect 10564 -836 10596 -835
rect 10564 -885 10596 -884
rect 10564 -915 10565 -885
rect 10565 -915 10595 -885
rect 10595 -915 10596 -885
rect 10564 -916 10596 -915
rect 10564 -996 10596 -964
rect 10564 -1076 10596 -1044
rect 10564 -1125 10596 -1124
rect 10564 -1155 10565 -1125
rect 10565 -1155 10595 -1125
rect 10595 -1155 10596 -1125
rect 10564 -1156 10596 -1155
rect 10564 -1205 10596 -1204
rect 10564 -1235 10565 -1205
rect 10565 -1235 10595 -1205
rect 10595 -1235 10596 -1205
rect 10564 -1236 10596 -1235
rect 10564 -1285 10596 -1284
rect 10564 -1315 10565 -1285
rect 10565 -1315 10595 -1285
rect 10595 -1315 10596 -1285
rect 10564 -1316 10596 -1315
rect 10564 -1365 10596 -1364
rect 10564 -1395 10565 -1365
rect 10565 -1395 10595 -1365
rect 10595 -1395 10596 -1365
rect 10564 -1396 10596 -1395
rect 10564 -1445 10596 -1444
rect 10564 -1475 10565 -1445
rect 10565 -1475 10595 -1445
rect 10595 -1475 10596 -1445
rect 10564 -1476 10596 -1475
rect 10564 -1525 10596 -1524
rect 10564 -1555 10565 -1525
rect 10565 -1555 10595 -1525
rect 10595 -1555 10596 -1525
rect 10564 -1556 10596 -1555
rect 10564 -1636 10596 -1604
rect 10564 -1716 10596 -1684
rect 10564 -1765 10596 -1764
rect 10564 -1795 10565 -1765
rect 10565 -1795 10595 -1765
rect 10595 -1795 10596 -1765
rect 10564 -1796 10596 -1795
rect 10564 -1845 10596 -1844
rect 10564 -1875 10565 -1845
rect 10565 -1875 10595 -1845
rect 10595 -1875 10596 -1845
rect 10564 -1876 10596 -1875
rect 10564 -1956 10596 -1924
rect 10564 -2005 10596 -2004
rect 10564 -2035 10565 -2005
rect 10565 -2035 10595 -2005
rect 10595 -2035 10596 -2005
rect 10564 -2036 10596 -2035
rect 10564 -2116 10596 -2084
rect 10564 -2165 10596 -2164
rect 10564 -2195 10565 -2165
rect 10565 -2195 10595 -2165
rect 10595 -2195 10596 -2165
rect 10564 -2196 10596 -2195
rect 10564 -2276 10596 -2244
rect 10564 -2325 10596 -2324
rect 10564 -2355 10565 -2325
rect 10565 -2355 10595 -2325
rect 10595 -2355 10596 -2325
rect 10564 -2356 10596 -2355
rect 10564 -2405 10596 -2404
rect 10564 -2435 10565 -2405
rect 10565 -2435 10595 -2405
rect 10595 -2435 10596 -2405
rect 10564 -2436 10596 -2435
rect 10564 -2485 10596 -2484
rect 10564 -2515 10565 -2485
rect 10565 -2515 10595 -2485
rect 10595 -2515 10596 -2485
rect 10564 -2516 10596 -2515
rect 10644 1035 10676 1036
rect 10644 1005 10645 1035
rect 10645 1005 10675 1035
rect 10675 1005 10676 1035
rect 10644 1004 10676 1005
rect 10644 955 10676 956
rect 10644 925 10645 955
rect 10645 925 10675 955
rect 10675 925 10676 955
rect 10644 924 10676 925
rect 10644 875 10676 876
rect 10644 845 10645 875
rect 10645 845 10675 875
rect 10675 845 10676 875
rect 10644 844 10676 845
rect 10644 795 10676 796
rect 10644 765 10645 795
rect 10645 765 10675 795
rect 10675 765 10676 795
rect 10644 764 10676 765
rect 10644 715 10676 716
rect 10644 685 10645 715
rect 10645 685 10675 715
rect 10675 685 10676 715
rect 10644 684 10676 685
rect 10644 635 10676 636
rect 10644 605 10645 635
rect 10645 605 10675 635
rect 10675 605 10676 635
rect 10644 604 10676 605
rect 10644 555 10676 556
rect 10644 525 10645 555
rect 10645 525 10675 555
rect 10675 525 10676 555
rect 10644 524 10676 525
rect 10644 475 10676 476
rect 10644 445 10645 475
rect 10645 445 10675 475
rect 10675 445 10676 475
rect 10644 444 10676 445
rect 10644 395 10676 396
rect 10644 365 10645 395
rect 10645 365 10675 395
rect 10675 365 10676 395
rect 10644 364 10676 365
rect 10644 284 10676 316
rect 10644 235 10676 236
rect 10644 205 10645 235
rect 10645 205 10675 235
rect 10675 205 10676 235
rect 10644 204 10676 205
rect 10644 124 10676 156
rect 10644 75 10676 76
rect 10644 45 10645 75
rect 10645 45 10675 75
rect 10675 45 10676 75
rect 10644 44 10676 45
rect 10644 -5 10676 -4
rect 10644 -35 10645 -5
rect 10645 -35 10675 -5
rect 10675 -35 10676 -5
rect 10644 -36 10676 -35
rect 10644 -85 10676 -84
rect 10644 -115 10645 -85
rect 10645 -115 10675 -85
rect 10675 -115 10676 -85
rect 10644 -116 10676 -115
rect 10644 -165 10676 -164
rect 10644 -195 10645 -165
rect 10645 -195 10675 -165
rect 10675 -195 10676 -165
rect 10644 -196 10676 -195
rect 10644 -245 10676 -244
rect 10644 -275 10645 -245
rect 10645 -275 10675 -245
rect 10675 -275 10676 -245
rect 10644 -276 10676 -275
rect 10644 -325 10676 -324
rect 10644 -355 10645 -325
rect 10645 -355 10675 -325
rect 10675 -355 10676 -325
rect 10644 -356 10676 -355
rect 10644 -436 10676 -404
rect 10644 -485 10676 -484
rect 10644 -515 10645 -485
rect 10645 -515 10675 -485
rect 10675 -515 10676 -485
rect 10644 -516 10676 -515
rect 10644 -596 10676 -564
rect 10644 -645 10676 -644
rect 10644 -675 10645 -645
rect 10645 -675 10675 -645
rect 10675 -675 10676 -645
rect 10644 -676 10676 -675
rect 10644 -725 10676 -724
rect 10644 -755 10645 -725
rect 10645 -755 10675 -725
rect 10675 -755 10676 -725
rect 10644 -756 10676 -755
rect 10644 -805 10676 -804
rect 10644 -835 10645 -805
rect 10645 -835 10675 -805
rect 10675 -835 10676 -805
rect 10644 -836 10676 -835
rect 10644 -885 10676 -884
rect 10644 -915 10645 -885
rect 10645 -915 10675 -885
rect 10675 -915 10676 -885
rect 10644 -916 10676 -915
rect 10644 -965 10676 -964
rect 10644 -995 10645 -965
rect 10645 -995 10675 -965
rect 10675 -995 10676 -965
rect 10644 -996 10676 -995
rect 10644 -1045 10676 -1044
rect 10644 -1075 10645 -1045
rect 10645 -1075 10675 -1045
rect 10675 -1075 10676 -1045
rect 10644 -1076 10676 -1075
rect 10644 -1125 10676 -1124
rect 10644 -1155 10645 -1125
rect 10645 -1155 10675 -1125
rect 10675 -1155 10676 -1125
rect 10644 -1156 10676 -1155
rect 10644 -1205 10676 -1204
rect 10644 -1235 10645 -1205
rect 10645 -1235 10675 -1205
rect 10675 -1235 10676 -1205
rect 10644 -1236 10676 -1235
rect 10644 -1285 10676 -1284
rect 10644 -1315 10645 -1285
rect 10645 -1315 10675 -1285
rect 10675 -1315 10676 -1285
rect 10644 -1316 10676 -1315
rect 10644 -1365 10676 -1364
rect 10644 -1395 10645 -1365
rect 10645 -1395 10675 -1365
rect 10675 -1395 10676 -1365
rect 10644 -1396 10676 -1395
rect 10644 -1445 10676 -1444
rect 10644 -1475 10645 -1445
rect 10645 -1475 10675 -1445
rect 10675 -1475 10676 -1445
rect 10644 -1476 10676 -1475
rect 10644 -1525 10676 -1524
rect 10644 -1555 10645 -1525
rect 10645 -1555 10675 -1525
rect 10675 -1555 10676 -1525
rect 10644 -1556 10676 -1555
rect 10644 -1605 10676 -1604
rect 10644 -1635 10645 -1605
rect 10645 -1635 10675 -1605
rect 10675 -1635 10676 -1605
rect 10644 -1636 10676 -1635
rect 10644 -1685 10676 -1684
rect 10644 -1715 10645 -1685
rect 10645 -1715 10675 -1685
rect 10675 -1715 10676 -1685
rect 10644 -1716 10676 -1715
rect 10644 -1765 10676 -1764
rect 10644 -1795 10645 -1765
rect 10645 -1795 10675 -1765
rect 10675 -1795 10676 -1765
rect 10644 -1796 10676 -1795
rect 10644 -1845 10676 -1844
rect 10644 -1875 10645 -1845
rect 10645 -1875 10675 -1845
rect 10675 -1875 10676 -1845
rect 10644 -1876 10676 -1875
rect 10644 -1925 10676 -1924
rect 10644 -1955 10645 -1925
rect 10645 -1955 10675 -1925
rect 10675 -1955 10676 -1925
rect 10644 -1956 10676 -1955
rect 10644 -2005 10676 -2004
rect 10644 -2035 10645 -2005
rect 10645 -2035 10675 -2005
rect 10675 -2035 10676 -2005
rect 10644 -2036 10676 -2035
rect 10644 -2116 10676 -2084
rect 10644 -2165 10676 -2164
rect 10644 -2195 10645 -2165
rect 10645 -2195 10675 -2165
rect 10675 -2195 10676 -2165
rect 10644 -2196 10676 -2195
rect 10644 -2276 10676 -2244
rect 10644 -2325 10676 -2324
rect 10644 -2355 10645 -2325
rect 10645 -2355 10675 -2325
rect 10675 -2355 10676 -2325
rect 10644 -2356 10676 -2355
rect 10644 -2405 10676 -2404
rect 10644 -2435 10645 -2405
rect 10645 -2435 10675 -2405
rect 10675 -2435 10676 -2405
rect 10644 -2436 10676 -2435
rect 10644 -2485 10676 -2484
rect 10644 -2515 10645 -2485
rect 10645 -2515 10675 -2485
rect 10675 -2515 10676 -2485
rect 10644 -2516 10676 -2515
rect 10644 -2565 10676 -2564
rect 10644 -2595 10645 -2565
rect 10645 -2595 10675 -2565
rect 10675 -2595 10676 -2565
rect 10644 -2596 10676 -2595
rect 10644 -2645 10676 -2644
rect 10644 -2675 10645 -2645
rect 10645 -2675 10675 -2645
rect 10675 -2675 10676 -2645
rect 10644 -2676 10676 -2675
rect 10644 -2725 10676 -2724
rect 10644 -2755 10645 -2725
rect 10645 -2755 10675 -2725
rect 10675 -2755 10676 -2725
rect 10644 -2756 10676 -2755
rect 10644 -2836 10676 -2804
rect 10644 -2885 10676 -2884
rect 10644 -2915 10645 -2885
rect 10645 -2915 10675 -2885
rect 10675 -2915 10676 -2885
rect 10644 -2916 10676 -2915
rect 10644 -2996 10676 -2964
rect 10644 -3045 10676 -3044
rect 10644 -3075 10645 -3045
rect 10645 -3075 10675 -3045
rect 10675 -3075 10676 -3045
rect 10644 -3076 10676 -3075
rect 10644 -3125 10676 -3124
rect 10644 -3155 10645 -3125
rect 10645 -3155 10675 -3125
rect 10675 -3155 10676 -3125
rect 10644 -3156 10676 -3155
rect 10644 -3205 10676 -3204
rect 10644 -3235 10645 -3205
rect 10645 -3235 10675 -3205
rect 10675 -3235 10676 -3205
rect 10644 -3236 10676 -3235
rect 10644 -3285 10676 -3284
rect 10644 -3315 10645 -3285
rect 10645 -3315 10675 -3285
rect 10675 -3315 10676 -3285
rect 10644 -3316 10676 -3315
rect 10644 -3365 10676 -3364
rect 10644 -3395 10645 -3365
rect 10645 -3395 10675 -3365
rect 10675 -3395 10676 -3365
rect 10644 -3396 10676 -3395
rect 10644 -3445 10676 -3444
rect 10644 -3475 10645 -3445
rect 10645 -3475 10675 -3445
rect 10675 -3475 10676 -3445
rect 10644 -3476 10676 -3475
rect 10644 -3525 10676 -3524
rect 10644 -3555 10645 -3525
rect 10645 -3555 10675 -3525
rect 10675 -3555 10676 -3525
rect 10644 -3556 10676 -3555
rect 10644 -3605 10676 -3604
rect 10644 -3635 10645 -3605
rect 10645 -3635 10675 -3605
rect 10675 -3635 10676 -3605
rect 10644 -3636 10676 -3635
rect 10644 -3685 10676 -3684
rect 10644 -3715 10645 -3685
rect 10645 -3715 10675 -3685
rect 10675 -3715 10676 -3685
rect 10644 -3716 10676 -3715
rect 10804 1035 10836 1036
rect 10804 1005 10805 1035
rect 10805 1005 10835 1035
rect 10835 1005 10836 1035
rect 10804 1004 10836 1005
rect 10804 955 10836 956
rect 10804 925 10805 955
rect 10805 925 10835 955
rect 10835 925 10836 955
rect 10804 924 10836 925
rect 10804 875 10836 876
rect 10804 845 10805 875
rect 10805 845 10835 875
rect 10835 845 10836 875
rect 10804 844 10836 845
rect 10804 795 10836 796
rect 10804 765 10805 795
rect 10805 765 10835 795
rect 10835 765 10836 795
rect 10804 764 10836 765
rect 10804 715 10836 716
rect 10804 685 10805 715
rect 10805 685 10835 715
rect 10835 685 10836 715
rect 10804 684 10836 685
rect 10804 635 10836 636
rect 10804 605 10805 635
rect 10805 605 10835 635
rect 10835 605 10836 635
rect 10804 604 10836 605
rect 10804 555 10836 556
rect 10804 525 10805 555
rect 10805 525 10835 555
rect 10835 525 10836 555
rect 10804 524 10836 525
rect 10804 475 10836 476
rect 10804 445 10805 475
rect 10805 445 10835 475
rect 10835 445 10836 475
rect 10804 444 10836 445
rect 10804 395 10836 396
rect 10804 365 10805 395
rect 10805 365 10835 395
rect 10835 365 10836 395
rect 10804 364 10836 365
rect 10804 284 10836 316
rect 10804 235 10836 236
rect 10804 205 10805 235
rect 10805 205 10835 235
rect 10835 205 10836 235
rect 10804 204 10836 205
rect 10804 155 10836 156
rect 10804 125 10805 155
rect 10805 125 10835 155
rect 10835 125 10836 155
rect 10804 124 10836 125
rect 10804 75 10836 76
rect 10804 45 10805 75
rect 10805 45 10835 75
rect 10835 45 10836 75
rect 10804 44 10836 45
rect 10804 -5 10836 -4
rect 10804 -35 10805 -5
rect 10805 -35 10835 -5
rect 10835 -35 10836 -5
rect 10804 -36 10836 -35
rect 10804 -85 10836 -84
rect 10804 -115 10805 -85
rect 10805 -115 10835 -85
rect 10835 -115 10836 -85
rect 10804 -116 10836 -115
rect 10804 -165 10836 -164
rect 10804 -195 10805 -165
rect 10805 -195 10835 -165
rect 10835 -195 10836 -165
rect 10804 -196 10836 -195
rect 10804 -245 10836 -244
rect 10804 -275 10805 -245
rect 10805 -275 10835 -245
rect 10835 -275 10836 -245
rect 10804 -276 10836 -275
rect 10804 -325 10836 -324
rect 10804 -355 10805 -325
rect 10805 -355 10835 -325
rect 10835 -355 10836 -325
rect 10804 -356 10836 -355
rect 10804 -405 10836 -404
rect 10804 -435 10805 -405
rect 10805 -435 10835 -405
rect 10835 -435 10836 -405
rect 10804 -436 10836 -435
rect 10804 -485 10836 -484
rect 10804 -515 10805 -485
rect 10805 -515 10835 -485
rect 10835 -515 10836 -485
rect 10804 -516 10836 -515
rect 10804 -596 10836 -564
rect 10804 -645 10836 -644
rect 10804 -675 10805 -645
rect 10805 -675 10835 -645
rect 10835 -675 10836 -645
rect 10804 -676 10836 -675
rect 10804 -725 10836 -724
rect 10804 -755 10805 -725
rect 10805 -755 10835 -725
rect 10835 -755 10836 -725
rect 10804 -756 10836 -755
rect 10804 -805 10836 -804
rect 10804 -835 10805 -805
rect 10805 -835 10835 -805
rect 10835 -835 10836 -805
rect 10804 -836 10836 -835
rect 10804 -885 10836 -884
rect 10804 -915 10805 -885
rect 10805 -915 10835 -885
rect 10835 -915 10836 -885
rect 10804 -916 10836 -915
rect 10804 -965 10836 -964
rect 10804 -995 10805 -965
rect 10805 -995 10835 -965
rect 10835 -995 10836 -965
rect 10804 -996 10836 -995
rect 10804 -1045 10836 -1044
rect 10804 -1075 10805 -1045
rect 10805 -1075 10835 -1045
rect 10835 -1075 10836 -1045
rect 10804 -1076 10836 -1075
rect 10804 -1125 10836 -1124
rect 10804 -1155 10805 -1125
rect 10805 -1155 10835 -1125
rect 10835 -1155 10836 -1125
rect 10804 -1156 10836 -1155
rect 10804 -1205 10836 -1204
rect 10804 -1235 10805 -1205
rect 10805 -1235 10835 -1205
rect 10835 -1235 10836 -1205
rect 10804 -1236 10836 -1235
rect 10804 -1285 10836 -1284
rect 10804 -1315 10805 -1285
rect 10805 -1315 10835 -1285
rect 10835 -1315 10836 -1285
rect 10804 -1316 10836 -1315
rect 10804 -1365 10836 -1364
rect 10804 -1395 10805 -1365
rect 10805 -1395 10835 -1365
rect 10835 -1395 10836 -1365
rect 10804 -1396 10836 -1395
rect 10804 -1445 10836 -1444
rect 10804 -1475 10805 -1445
rect 10805 -1475 10835 -1445
rect 10835 -1475 10836 -1445
rect 10804 -1476 10836 -1475
rect 10804 -1525 10836 -1524
rect 10804 -1555 10805 -1525
rect 10805 -1555 10835 -1525
rect 10835 -1555 10836 -1525
rect 10804 -1556 10836 -1555
rect 10804 -1605 10836 -1604
rect 10804 -1635 10805 -1605
rect 10805 -1635 10835 -1605
rect 10835 -1635 10836 -1605
rect 10804 -1636 10836 -1635
rect 10804 -1685 10836 -1684
rect 10804 -1715 10805 -1685
rect 10805 -1715 10835 -1685
rect 10835 -1715 10836 -1685
rect 10804 -1716 10836 -1715
rect 10804 -1765 10836 -1764
rect 10804 -1795 10805 -1765
rect 10805 -1795 10835 -1765
rect 10835 -1795 10836 -1765
rect 10804 -1796 10836 -1795
rect 10804 -1845 10836 -1844
rect 10804 -1875 10805 -1845
rect 10805 -1875 10835 -1845
rect 10835 -1875 10836 -1845
rect 10804 -1876 10836 -1875
rect 10804 -1925 10836 -1924
rect 10804 -1955 10805 -1925
rect 10805 -1955 10835 -1925
rect 10835 -1955 10836 -1925
rect 10804 -1956 10836 -1955
rect 10804 -2005 10836 -2004
rect 10804 -2035 10805 -2005
rect 10805 -2035 10835 -2005
rect 10835 -2035 10836 -2005
rect 10804 -2036 10836 -2035
rect 10804 -2116 10836 -2084
rect 10804 -2165 10836 -2164
rect 10804 -2195 10805 -2165
rect 10805 -2195 10835 -2165
rect 10835 -2195 10836 -2165
rect 10804 -2196 10836 -2195
rect 10804 -2245 10836 -2244
rect 10804 -2275 10805 -2245
rect 10805 -2275 10835 -2245
rect 10835 -2275 10836 -2245
rect 10804 -2276 10836 -2275
rect 10804 -2325 10836 -2324
rect 10804 -2355 10805 -2325
rect 10805 -2355 10835 -2325
rect 10835 -2355 10836 -2325
rect 10804 -2356 10836 -2355
rect 10804 -2405 10836 -2404
rect 10804 -2435 10805 -2405
rect 10805 -2435 10835 -2405
rect 10835 -2435 10836 -2405
rect 10804 -2436 10836 -2435
rect 10804 -2485 10836 -2484
rect 10804 -2515 10805 -2485
rect 10805 -2515 10835 -2485
rect 10835 -2515 10836 -2485
rect 10804 -2516 10836 -2515
rect 10804 -2565 10836 -2564
rect 10804 -2595 10805 -2565
rect 10805 -2595 10835 -2565
rect 10835 -2595 10836 -2565
rect 10804 -2596 10836 -2595
rect 10804 -2645 10836 -2644
rect 10804 -2675 10805 -2645
rect 10805 -2675 10835 -2645
rect 10835 -2675 10836 -2645
rect 10804 -2676 10836 -2675
rect 10804 -2725 10836 -2724
rect 10804 -2755 10805 -2725
rect 10805 -2755 10835 -2725
rect 10835 -2755 10836 -2725
rect 10804 -2756 10836 -2755
rect 10804 -2805 10836 -2804
rect 10804 -2835 10805 -2805
rect 10805 -2835 10835 -2805
rect 10835 -2835 10836 -2805
rect 10804 -2836 10836 -2835
rect 10804 -2885 10836 -2884
rect 10804 -2915 10805 -2885
rect 10805 -2915 10835 -2885
rect 10835 -2915 10836 -2885
rect 10804 -2916 10836 -2915
rect 10804 -2996 10836 -2964
rect 10804 -3045 10836 -3044
rect 10804 -3075 10805 -3045
rect 10805 -3075 10835 -3045
rect 10835 -3075 10836 -3045
rect 10804 -3076 10836 -3075
rect 10804 -3125 10836 -3124
rect 10804 -3155 10805 -3125
rect 10805 -3155 10835 -3125
rect 10835 -3155 10836 -3125
rect 10804 -3156 10836 -3155
rect 10804 -3205 10836 -3204
rect 10804 -3235 10805 -3205
rect 10805 -3235 10835 -3205
rect 10835 -3235 10836 -3205
rect 10804 -3236 10836 -3235
rect 10804 -3285 10836 -3284
rect 10804 -3315 10805 -3285
rect 10805 -3315 10835 -3285
rect 10835 -3315 10836 -3285
rect 10804 -3316 10836 -3315
rect 10804 -3365 10836 -3364
rect 10804 -3395 10805 -3365
rect 10805 -3395 10835 -3365
rect 10835 -3395 10836 -3365
rect 10804 -3396 10836 -3395
rect 10804 -3445 10836 -3444
rect 10804 -3475 10805 -3445
rect 10805 -3475 10835 -3445
rect 10835 -3475 10836 -3445
rect 10804 -3476 10836 -3475
rect 10804 -3525 10836 -3524
rect 10804 -3555 10805 -3525
rect 10805 -3555 10835 -3525
rect 10835 -3555 10836 -3525
rect 10804 -3556 10836 -3555
rect 10804 -3605 10836 -3604
rect 10804 -3635 10805 -3605
rect 10805 -3635 10835 -3605
rect 10835 -3635 10836 -3605
rect 10804 -3636 10836 -3635
rect 10804 -3685 10836 -3684
rect 10804 -3715 10805 -3685
rect 10805 -3715 10835 -3685
rect 10835 -3715 10836 -3685
rect 10804 -3716 10836 -3715
rect 10964 1035 10996 1036
rect 10964 1005 10965 1035
rect 10965 1005 10995 1035
rect 10995 1005 10996 1035
rect 10964 1004 10996 1005
rect 10964 955 10996 956
rect 10964 925 10965 955
rect 10965 925 10995 955
rect 10995 925 10996 955
rect 10964 924 10996 925
rect 10964 875 10996 876
rect 10964 845 10965 875
rect 10965 845 10995 875
rect 10995 845 10996 875
rect 10964 844 10996 845
rect 10964 795 10996 796
rect 10964 765 10965 795
rect 10965 765 10995 795
rect 10995 765 10996 795
rect 10964 764 10996 765
rect 10964 715 10996 716
rect 10964 685 10965 715
rect 10965 685 10995 715
rect 10995 685 10996 715
rect 10964 684 10996 685
rect 10964 635 10996 636
rect 10964 605 10965 635
rect 10965 605 10995 635
rect 10995 605 10996 635
rect 10964 604 10996 605
rect 10964 555 10996 556
rect 10964 525 10965 555
rect 10965 525 10995 555
rect 10995 525 10996 555
rect 10964 524 10996 525
rect 10964 475 10996 476
rect 10964 445 10965 475
rect 10965 445 10995 475
rect 10995 445 10996 475
rect 10964 444 10996 445
rect 10964 395 10996 396
rect 10964 365 10965 395
rect 10965 365 10995 395
rect 10995 365 10996 395
rect 10964 364 10996 365
rect 10964 284 10996 316
rect 10964 235 10996 236
rect 10964 205 10965 235
rect 10965 205 10995 235
rect 10995 205 10996 235
rect 10964 204 10996 205
rect 10964 155 10996 156
rect 10964 125 10965 155
rect 10965 125 10995 155
rect 10995 125 10996 155
rect 10964 124 10996 125
rect 10964 75 10996 76
rect 10964 45 10965 75
rect 10965 45 10995 75
rect 10995 45 10996 75
rect 10964 44 10996 45
rect 10964 -5 10996 -4
rect 10964 -35 10965 -5
rect 10965 -35 10995 -5
rect 10995 -35 10996 -5
rect 10964 -36 10996 -35
rect 10964 -85 10996 -84
rect 10964 -115 10965 -85
rect 10965 -115 10995 -85
rect 10995 -115 10996 -85
rect 10964 -116 10996 -115
rect 10964 -165 10996 -164
rect 10964 -195 10965 -165
rect 10965 -195 10995 -165
rect 10995 -195 10996 -165
rect 10964 -196 10996 -195
rect 10964 -245 10996 -244
rect 10964 -275 10965 -245
rect 10965 -275 10995 -245
rect 10995 -275 10996 -245
rect 10964 -276 10996 -275
rect 10964 -325 10996 -324
rect 10964 -355 10965 -325
rect 10965 -355 10995 -325
rect 10995 -355 10996 -325
rect 10964 -356 10996 -355
rect 10964 -405 10996 -404
rect 10964 -435 10965 -405
rect 10965 -435 10995 -405
rect 10995 -435 10996 -405
rect 10964 -436 10996 -435
rect 10964 -485 10996 -484
rect 10964 -515 10965 -485
rect 10965 -515 10995 -485
rect 10995 -515 10996 -485
rect 10964 -516 10996 -515
rect 10964 -596 10996 -564
rect 10964 -645 10996 -644
rect 10964 -675 10965 -645
rect 10965 -675 10995 -645
rect 10995 -675 10996 -645
rect 10964 -676 10996 -675
rect 10964 -725 10996 -724
rect 10964 -755 10965 -725
rect 10965 -755 10995 -725
rect 10995 -755 10996 -725
rect 10964 -756 10996 -755
rect 10964 -805 10996 -804
rect 10964 -835 10965 -805
rect 10965 -835 10995 -805
rect 10995 -835 10996 -805
rect 10964 -836 10996 -835
rect 10964 -885 10996 -884
rect 10964 -915 10965 -885
rect 10965 -915 10995 -885
rect 10995 -915 10996 -885
rect 10964 -916 10996 -915
rect 10964 -965 10996 -964
rect 10964 -995 10965 -965
rect 10965 -995 10995 -965
rect 10995 -995 10996 -965
rect 10964 -996 10996 -995
rect 10964 -1045 10996 -1044
rect 10964 -1075 10965 -1045
rect 10965 -1075 10995 -1045
rect 10995 -1075 10996 -1045
rect 10964 -1076 10996 -1075
rect 10964 -1125 10996 -1124
rect 10964 -1155 10965 -1125
rect 10965 -1155 10995 -1125
rect 10995 -1155 10996 -1125
rect 10964 -1156 10996 -1155
rect 10964 -1205 10996 -1204
rect 10964 -1235 10965 -1205
rect 10965 -1235 10995 -1205
rect 10995 -1235 10996 -1205
rect 10964 -1236 10996 -1235
rect 10964 -1285 10996 -1284
rect 10964 -1315 10965 -1285
rect 10965 -1315 10995 -1285
rect 10995 -1315 10996 -1285
rect 10964 -1316 10996 -1315
rect 10964 -1365 10996 -1364
rect 10964 -1395 10965 -1365
rect 10965 -1395 10995 -1365
rect 10995 -1395 10996 -1365
rect 10964 -1396 10996 -1395
rect 10964 -1445 10996 -1444
rect 10964 -1475 10965 -1445
rect 10965 -1475 10995 -1445
rect 10995 -1475 10996 -1445
rect 10964 -1476 10996 -1475
rect 10964 -1525 10996 -1524
rect 10964 -1555 10965 -1525
rect 10965 -1555 10995 -1525
rect 10995 -1555 10996 -1525
rect 10964 -1556 10996 -1555
rect 10964 -1605 10996 -1604
rect 10964 -1635 10965 -1605
rect 10965 -1635 10995 -1605
rect 10995 -1635 10996 -1605
rect 10964 -1636 10996 -1635
rect 10964 -1685 10996 -1684
rect 10964 -1715 10965 -1685
rect 10965 -1715 10995 -1685
rect 10995 -1715 10996 -1685
rect 10964 -1716 10996 -1715
rect 10964 -1765 10996 -1764
rect 10964 -1795 10965 -1765
rect 10965 -1795 10995 -1765
rect 10995 -1795 10996 -1765
rect 10964 -1796 10996 -1795
rect 10964 -1845 10996 -1844
rect 10964 -1875 10965 -1845
rect 10965 -1875 10995 -1845
rect 10995 -1875 10996 -1845
rect 10964 -1876 10996 -1875
rect 10964 -1925 10996 -1924
rect 10964 -1955 10965 -1925
rect 10965 -1955 10995 -1925
rect 10995 -1955 10996 -1925
rect 10964 -1956 10996 -1955
rect 10964 -2005 10996 -2004
rect 10964 -2035 10965 -2005
rect 10965 -2035 10995 -2005
rect 10995 -2035 10996 -2005
rect 10964 -2036 10996 -2035
rect 10964 -2116 10996 -2084
rect 10964 -2165 10996 -2164
rect 10964 -2195 10965 -2165
rect 10965 -2195 10995 -2165
rect 10995 -2195 10996 -2165
rect 10964 -2196 10996 -2195
rect 10964 -2245 10996 -2244
rect 10964 -2275 10965 -2245
rect 10965 -2275 10995 -2245
rect 10995 -2275 10996 -2245
rect 10964 -2276 10996 -2275
rect 10964 -2325 10996 -2324
rect 10964 -2355 10965 -2325
rect 10965 -2355 10995 -2325
rect 10995 -2355 10996 -2325
rect 10964 -2356 10996 -2355
rect 10964 -2405 10996 -2404
rect 10964 -2435 10965 -2405
rect 10965 -2435 10995 -2405
rect 10995 -2435 10996 -2405
rect 10964 -2436 10996 -2435
rect 10964 -2485 10996 -2484
rect 10964 -2515 10965 -2485
rect 10965 -2515 10995 -2485
rect 10995 -2515 10996 -2485
rect 10964 -2516 10996 -2515
rect 10964 -2565 10996 -2564
rect 10964 -2595 10965 -2565
rect 10965 -2595 10995 -2565
rect 10995 -2595 10996 -2565
rect 10964 -2596 10996 -2595
rect 10964 -2645 10996 -2644
rect 10964 -2675 10965 -2645
rect 10965 -2675 10995 -2645
rect 10995 -2675 10996 -2645
rect 10964 -2676 10996 -2675
rect 10964 -2725 10996 -2724
rect 10964 -2755 10965 -2725
rect 10965 -2755 10995 -2725
rect 10995 -2755 10996 -2725
rect 10964 -2756 10996 -2755
rect 10964 -2805 10996 -2804
rect 10964 -2835 10965 -2805
rect 10965 -2835 10995 -2805
rect 10995 -2835 10996 -2805
rect 10964 -2836 10996 -2835
rect 10964 -2885 10996 -2884
rect 10964 -2915 10965 -2885
rect 10965 -2915 10995 -2885
rect 10995 -2915 10996 -2885
rect 10964 -2916 10996 -2915
rect 10964 -2996 10996 -2964
rect 10964 -3045 10996 -3044
rect 10964 -3075 10965 -3045
rect 10965 -3075 10995 -3045
rect 10995 -3075 10996 -3045
rect 10964 -3076 10996 -3075
rect 10964 -3125 10996 -3124
rect 10964 -3155 10965 -3125
rect 10965 -3155 10995 -3125
rect 10995 -3155 10996 -3125
rect 10964 -3156 10996 -3155
rect 10964 -3205 10996 -3204
rect 10964 -3235 10965 -3205
rect 10965 -3235 10995 -3205
rect 10995 -3235 10996 -3205
rect 10964 -3236 10996 -3235
rect 10964 -3285 10996 -3284
rect 10964 -3315 10965 -3285
rect 10965 -3315 10995 -3285
rect 10995 -3315 10996 -3285
rect 10964 -3316 10996 -3315
rect 10964 -3365 10996 -3364
rect 10964 -3395 10965 -3365
rect 10965 -3395 10995 -3365
rect 10995 -3395 10996 -3365
rect 10964 -3396 10996 -3395
rect 10964 -3445 10996 -3444
rect 10964 -3475 10965 -3445
rect 10965 -3475 10995 -3445
rect 10995 -3475 10996 -3445
rect 10964 -3476 10996 -3475
rect 10964 -3525 10996 -3524
rect 10964 -3555 10965 -3525
rect 10965 -3555 10995 -3525
rect 10995 -3555 10996 -3525
rect 10964 -3556 10996 -3555
rect 10964 -3605 10996 -3604
rect 10964 -3635 10965 -3605
rect 10965 -3635 10995 -3605
rect 10995 -3635 10996 -3605
rect 10964 -3636 10996 -3635
rect 10964 -3685 10996 -3684
rect 10964 -3715 10965 -3685
rect 10965 -3715 10995 -3685
rect 10995 -3715 10996 -3685
rect 10964 -3716 10996 -3715
<< metal4 >>
rect -720 1036 11000 1040
rect -720 1004 -716 1036
rect -684 1004 -556 1036
rect -524 1004 -396 1036
rect -364 1004 -316 1036
rect -284 1004 -236 1036
rect -204 1004 -156 1036
rect -124 1004 -76 1036
rect -44 1004 4 1036
rect 36 1004 84 1036
rect 116 1004 164 1036
rect 196 1004 244 1036
rect 276 1004 324 1036
rect 356 1004 404 1036
rect 436 1004 484 1036
rect 516 1004 564 1036
rect 596 1004 644 1036
rect 676 1004 724 1036
rect 756 1004 804 1036
rect 836 1004 884 1036
rect 916 1004 964 1036
rect 996 1004 1044 1036
rect 1076 1004 1124 1036
rect 1156 1004 1204 1036
rect 1236 1004 1284 1036
rect 1316 1004 1364 1036
rect 1396 1004 1444 1036
rect 1476 1004 1524 1036
rect 1556 1004 1604 1036
rect 1636 1004 1684 1036
rect 1716 1004 1764 1036
rect 1796 1004 1844 1036
rect 1876 1004 1924 1036
rect 1956 1004 2004 1036
rect 2036 1004 2084 1036
rect 2116 1004 2164 1036
rect 2196 1004 2244 1036
rect 2276 1004 2324 1036
rect 2356 1004 2404 1036
rect 2436 1004 2484 1036
rect 2516 1004 2564 1036
rect 2596 1004 2644 1036
rect 2676 1004 2724 1036
rect 2756 1004 2804 1036
rect 2836 1004 2884 1036
rect 2916 1004 2964 1036
rect 2996 1004 3044 1036
rect 3076 1004 3124 1036
rect 3156 1004 3204 1036
rect 3236 1004 3284 1036
rect 3316 1004 3364 1036
rect 3396 1004 3444 1036
rect 3476 1004 3524 1036
rect 3556 1004 3604 1036
rect 3636 1004 3684 1036
rect 3716 1004 3764 1036
rect 3796 1004 3844 1036
rect 3876 1004 3924 1036
rect 3956 1004 4004 1036
rect 4036 1004 4084 1036
rect 4116 1004 4164 1036
rect 4196 1004 4244 1036
rect 4276 1004 4324 1036
rect 4356 1004 4404 1036
rect 4436 1004 4484 1036
rect 4516 1004 4564 1036
rect 4596 1004 4644 1036
rect 4676 1004 4724 1036
rect 4756 1004 4804 1036
rect 4836 1004 4884 1036
rect 4916 1004 4964 1036
rect 4996 1004 5044 1036
rect 5076 1004 5124 1036
rect 5156 1004 5204 1036
rect 5236 1004 5284 1036
rect 5316 1004 5364 1036
rect 5396 1004 5444 1036
rect 5476 1004 5524 1036
rect 5556 1004 5604 1036
rect 5636 1004 5684 1036
rect 5716 1004 5764 1036
rect 5796 1004 5844 1036
rect 5876 1004 5924 1036
rect 5956 1004 6004 1036
rect 6036 1004 6084 1036
rect 6116 1004 6164 1036
rect 6196 1004 6244 1036
rect 6276 1004 6324 1036
rect 6356 1004 6404 1036
rect 6436 1004 6484 1036
rect 6516 1004 6564 1036
rect 6596 1004 6644 1036
rect 6676 1004 6724 1036
rect 6756 1004 6804 1036
rect 6836 1004 6884 1036
rect 6916 1004 6964 1036
rect 6996 1004 7044 1036
rect 7076 1004 7124 1036
rect 7156 1004 7204 1036
rect 7236 1004 7284 1036
rect 7316 1004 7364 1036
rect 7396 1004 7444 1036
rect 7476 1004 7524 1036
rect 7556 1004 7604 1036
rect 7636 1004 7684 1036
rect 7716 1004 7764 1036
rect 7796 1004 7844 1036
rect 7876 1004 7924 1036
rect 7956 1004 8004 1036
rect 8036 1004 8084 1036
rect 8116 1004 8164 1036
rect 8196 1004 8244 1036
rect 8276 1004 8324 1036
rect 8356 1004 8404 1036
rect 8436 1004 8484 1036
rect 8516 1004 8564 1036
rect 8596 1004 8644 1036
rect 8676 1004 8724 1036
rect 8756 1004 8804 1036
rect 8836 1004 8884 1036
rect 8916 1004 8964 1036
rect 8996 1004 9044 1036
rect 9076 1004 9124 1036
rect 9156 1004 9204 1036
rect 9236 1004 9284 1036
rect 9316 1004 9364 1036
rect 9396 1004 9444 1036
rect 9476 1004 9524 1036
rect 9556 1004 9604 1036
rect 9636 1004 9684 1036
rect 9716 1004 9764 1036
rect 9796 1004 9844 1036
rect 9876 1004 9924 1036
rect 9956 1004 10004 1036
rect 10036 1004 10084 1036
rect 10116 1004 10164 1036
rect 10196 1004 10244 1036
rect 10276 1004 10324 1036
rect 10356 1004 10404 1036
rect 10436 1004 10484 1036
rect 10516 1004 10644 1036
rect 10676 1004 10804 1036
rect 10836 1004 10964 1036
rect 10996 1004 11000 1036
rect -720 1000 11000 1004
rect -720 956 11000 960
rect -720 924 -716 956
rect -684 924 -556 956
rect -524 924 -396 956
rect -364 924 -316 956
rect -284 924 -236 956
rect -204 924 -156 956
rect -124 924 -76 956
rect -44 924 4 956
rect 36 924 84 956
rect 116 924 164 956
rect 196 924 244 956
rect 276 924 324 956
rect 356 924 404 956
rect 436 924 484 956
rect 516 924 564 956
rect 596 924 644 956
rect 676 924 724 956
rect 756 924 804 956
rect 836 924 884 956
rect 916 924 964 956
rect 996 924 1044 956
rect 1076 924 1124 956
rect 1156 924 1204 956
rect 1236 924 1284 956
rect 1316 924 1364 956
rect 1396 924 1444 956
rect 1476 924 1524 956
rect 1556 924 1604 956
rect 1636 924 1684 956
rect 1716 924 1764 956
rect 1796 924 1844 956
rect 1876 924 1924 956
rect 1956 924 2004 956
rect 2036 924 2084 956
rect 2116 924 2164 956
rect 2196 924 2244 956
rect 2276 924 2324 956
rect 2356 924 2404 956
rect 2436 924 2484 956
rect 2516 924 2564 956
rect 2596 924 2644 956
rect 2676 924 2724 956
rect 2756 924 2804 956
rect 2836 924 2884 956
rect 2916 924 2964 956
rect 2996 924 3044 956
rect 3076 924 3124 956
rect 3156 924 3204 956
rect 3236 924 3284 956
rect 3316 924 3364 956
rect 3396 924 3444 956
rect 3476 924 3524 956
rect 3556 924 3604 956
rect 3636 924 3684 956
rect 3716 924 3764 956
rect 3796 924 3844 956
rect 3876 924 3924 956
rect 3956 924 4004 956
rect 4036 924 4084 956
rect 4116 924 4164 956
rect 4196 924 4244 956
rect 4276 924 4324 956
rect 4356 924 4404 956
rect 4436 924 4484 956
rect 4516 924 4564 956
rect 4596 924 4644 956
rect 4676 924 4724 956
rect 4756 924 4804 956
rect 4836 924 4884 956
rect 4916 924 4964 956
rect 4996 924 5044 956
rect 5076 924 5124 956
rect 5156 924 5204 956
rect 5236 924 5284 956
rect 5316 924 5364 956
rect 5396 924 5444 956
rect 5476 924 5524 956
rect 5556 924 5604 956
rect 5636 924 5684 956
rect 5716 924 5764 956
rect 5796 924 5844 956
rect 5876 924 5924 956
rect 5956 924 6004 956
rect 6036 924 6084 956
rect 6116 924 6164 956
rect 6196 924 6244 956
rect 6276 924 6324 956
rect 6356 924 6404 956
rect 6436 924 6484 956
rect 6516 924 6564 956
rect 6596 924 6644 956
rect 6676 924 6724 956
rect 6756 924 6804 956
rect 6836 924 6884 956
rect 6916 924 6964 956
rect 6996 924 7044 956
rect 7076 924 7124 956
rect 7156 924 7204 956
rect 7236 924 7284 956
rect 7316 924 7364 956
rect 7396 924 7444 956
rect 7476 924 7524 956
rect 7556 924 7604 956
rect 7636 924 7684 956
rect 7716 924 7764 956
rect 7796 924 7844 956
rect 7876 924 7924 956
rect 7956 924 8004 956
rect 8036 924 8084 956
rect 8116 924 8164 956
rect 8196 924 8244 956
rect 8276 924 8324 956
rect 8356 924 8404 956
rect 8436 924 8484 956
rect 8516 924 8564 956
rect 8596 924 8644 956
rect 8676 924 8724 956
rect 8756 924 8804 956
rect 8836 924 8884 956
rect 8916 924 8964 956
rect 8996 924 9044 956
rect 9076 924 9124 956
rect 9156 924 9204 956
rect 9236 924 9284 956
rect 9316 924 9364 956
rect 9396 924 9444 956
rect 9476 924 9524 956
rect 9556 924 9604 956
rect 9636 924 9684 956
rect 9716 924 9764 956
rect 9796 924 9844 956
rect 9876 924 9924 956
rect 9956 924 10004 956
rect 10036 924 10084 956
rect 10116 924 10164 956
rect 10196 924 10244 956
rect 10276 924 10324 956
rect 10356 924 10404 956
rect 10436 924 10484 956
rect 10516 924 10644 956
rect 10676 924 10804 956
rect 10836 924 10964 956
rect 10996 924 11000 956
rect -720 920 11000 924
rect -720 876 11000 880
rect -720 844 -716 876
rect -684 844 -556 876
rect -524 844 -396 876
rect -364 844 -316 876
rect -284 844 -236 876
rect -204 844 -156 876
rect -124 844 -76 876
rect -44 844 4 876
rect 36 844 84 876
rect 116 844 164 876
rect 196 844 244 876
rect 276 844 324 876
rect 356 844 404 876
rect 436 844 484 876
rect 516 844 564 876
rect 596 844 644 876
rect 676 844 724 876
rect 756 844 804 876
rect 836 844 884 876
rect 916 844 964 876
rect 996 844 1044 876
rect 1076 844 1124 876
rect 1156 844 1204 876
rect 1236 844 1284 876
rect 1316 844 1364 876
rect 1396 844 1444 876
rect 1476 844 1524 876
rect 1556 844 1604 876
rect 1636 844 1684 876
rect 1716 844 1764 876
rect 1796 844 1844 876
rect 1876 844 1924 876
rect 1956 844 2004 876
rect 2036 844 2084 876
rect 2116 844 2164 876
rect 2196 844 2244 876
rect 2276 844 2324 876
rect 2356 844 2404 876
rect 2436 844 2484 876
rect 2516 844 2564 876
rect 2596 844 2644 876
rect 2676 844 2724 876
rect 2756 844 2804 876
rect 2836 844 2884 876
rect 2916 844 2964 876
rect 2996 844 3044 876
rect 3076 844 3124 876
rect 3156 844 3204 876
rect 3236 844 3284 876
rect 3316 844 3364 876
rect 3396 844 3444 876
rect 3476 844 3524 876
rect 3556 844 3604 876
rect 3636 844 3684 876
rect 3716 844 3764 876
rect 3796 844 3844 876
rect 3876 844 3924 876
rect 3956 844 4004 876
rect 4036 844 4084 876
rect 4116 844 4164 876
rect 4196 844 4244 876
rect 4276 844 4324 876
rect 4356 844 4404 876
rect 4436 844 4484 876
rect 4516 844 4564 876
rect 4596 844 4644 876
rect 4676 844 4724 876
rect 4756 844 4804 876
rect 4836 844 4884 876
rect 4916 844 4964 876
rect 4996 844 5044 876
rect 5076 844 5124 876
rect 5156 844 5204 876
rect 5236 844 5284 876
rect 5316 844 5364 876
rect 5396 844 5444 876
rect 5476 844 5524 876
rect 5556 844 5604 876
rect 5636 844 5684 876
rect 5716 844 5764 876
rect 5796 844 5844 876
rect 5876 844 5924 876
rect 5956 844 6004 876
rect 6036 844 6084 876
rect 6116 844 6164 876
rect 6196 844 6244 876
rect 6276 844 6324 876
rect 6356 844 6404 876
rect 6436 844 6484 876
rect 6516 844 6564 876
rect 6596 844 6644 876
rect 6676 844 6724 876
rect 6756 844 6804 876
rect 6836 844 6884 876
rect 6916 844 6964 876
rect 6996 844 7044 876
rect 7076 844 7124 876
rect 7156 844 7204 876
rect 7236 844 7284 876
rect 7316 844 7364 876
rect 7396 844 7444 876
rect 7476 844 7524 876
rect 7556 844 7604 876
rect 7636 844 7684 876
rect 7716 844 7764 876
rect 7796 844 7844 876
rect 7876 844 7924 876
rect 7956 844 8004 876
rect 8036 844 8084 876
rect 8116 844 8164 876
rect 8196 844 8244 876
rect 8276 844 8324 876
rect 8356 844 8404 876
rect 8436 844 8484 876
rect 8516 844 8564 876
rect 8596 844 8644 876
rect 8676 844 8724 876
rect 8756 844 8804 876
rect 8836 844 8884 876
rect 8916 844 8964 876
rect 8996 844 9044 876
rect 9076 844 9124 876
rect 9156 844 9204 876
rect 9236 844 9284 876
rect 9316 844 9364 876
rect 9396 844 9444 876
rect 9476 844 9524 876
rect 9556 844 9604 876
rect 9636 844 9684 876
rect 9716 844 9764 876
rect 9796 844 9844 876
rect 9876 844 9924 876
rect 9956 844 10004 876
rect 10036 844 10084 876
rect 10116 844 10164 876
rect 10196 844 10244 876
rect 10276 844 10324 876
rect 10356 844 10404 876
rect 10436 844 10484 876
rect 10516 844 10644 876
rect 10676 844 10804 876
rect 10836 844 10964 876
rect 10996 844 11000 876
rect -720 840 11000 844
rect -720 796 10600 800
rect -720 764 -716 796
rect -684 764 -556 796
rect -524 764 -396 796
rect -364 764 -316 796
rect -284 764 -236 796
rect -204 764 -156 796
rect -124 764 -76 796
rect -44 764 4 796
rect 36 764 84 796
rect 116 764 164 796
rect 196 764 244 796
rect 276 764 324 796
rect 356 764 404 796
rect 436 764 484 796
rect 516 764 564 796
rect 596 764 644 796
rect 676 764 724 796
rect 756 764 804 796
rect 836 764 884 796
rect 916 764 964 796
rect 996 764 1044 796
rect 1076 764 1124 796
rect 1156 764 1204 796
rect 1236 764 1284 796
rect 1316 764 1364 796
rect 1396 764 1444 796
rect 1476 764 1524 796
rect 1556 764 1604 796
rect 1636 764 1684 796
rect 1716 764 1764 796
rect 1796 764 1844 796
rect 1876 764 1924 796
rect 1956 764 2004 796
rect 2036 764 2084 796
rect 2116 764 2164 796
rect 2196 764 2244 796
rect 2276 764 2324 796
rect 2356 764 2404 796
rect 2436 764 2484 796
rect 2516 764 2564 796
rect 2596 764 2644 796
rect 2676 764 2724 796
rect 2756 764 2804 796
rect 2836 764 2884 796
rect 2916 764 2964 796
rect 2996 764 3044 796
rect 3076 764 3124 796
rect 3156 764 3204 796
rect 3236 764 3284 796
rect 3316 764 3364 796
rect 3396 764 3444 796
rect 3476 764 3524 796
rect 3556 764 3604 796
rect 3636 764 3684 796
rect 3716 764 3764 796
rect 3796 764 3844 796
rect 3876 764 3924 796
rect 3956 764 4004 796
rect 4036 764 4084 796
rect 4116 764 4164 796
rect 4196 764 4244 796
rect 4276 764 4324 796
rect 4356 764 4404 796
rect 4436 764 4484 796
rect 4516 764 4564 796
rect 4596 764 4644 796
rect 4676 764 4724 796
rect 4756 764 4804 796
rect 4836 764 4884 796
rect 4916 764 4964 796
rect 4996 764 5044 796
rect 5076 764 5124 796
rect 5156 764 5204 796
rect 5236 764 5284 796
rect 5316 764 5364 796
rect 5396 764 5444 796
rect 5476 764 5524 796
rect 5556 764 5604 796
rect 5636 764 5684 796
rect 5716 764 5764 796
rect 5796 764 5844 796
rect 5876 764 5924 796
rect 5956 764 6004 796
rect 6036 764 6084 796
rect 6116 764 6164 796
rect 6196 764 6244 796
rect 6276 764 6324 796
rect 6356 764 6404 796
rect 6436 764 6484 796
rect 6516 764 6564 796
rect 6596 764 6644 796
rect 6676 764 6724 796
rect 6756 764 6804 796
rect 6836 764 6884 796
rect 6916 764 6964 796
rect 6996 764 7044 796
rect 7076 764 7124 796
rect 7156 764 7204 796
rect 7236 764 7284 796
rect 7316 764 7364 796
rect 7396 764 7444 796
rect 7476 764 7524 796
rect 7556 764 7604 796
rect 7636 764 7684 796
rect 7716 764 7764 796
rect 7796 764 7844 796
rect 7876 764 7924 796
rect 7956 764 8004 796
rect 8036 764 8084 796
rect 8116 764 8164 796
rect 8196 764 8244 796
rect 8276 764 8324 796
rect 8356 764 8404 796
rect 8436 764 8484 796
rect 8516 764 8564 796
rect 8596 764 8644 796
rect 8676 764 8724 796
rect 8756 764 8804 796
rect 8836 764 8884 796
rect 8916 764 8964 796
rect 8996 764 9044 796
rect 9076 764 9124 796
rect 9156 764 9204 796
rect 9236 764 9284 796
rect 9316 764 9364 796
rect 9396 764 9444 796
rect 9476 764 9524 796
rect 9556 764 9604 796
rect 9636 764 9684 796
rect 9716 764 9764 796
rect 9796 764 9844 796
rect 9876 764 9924 796
rect 9956 764 10004 796
rect 10036 764 10084 796
rect 10116 764 10164 796
rect 10196 764 10244 796
rect 10276 764 10324 796
rect 10356 764 10404 796
rect 10436 764 10484 796
rect 10516 764 10600 796
rect -720 760 10600 764
rect 10640 796 11000 800
rect 10640 764 10644 796
rect 10676 764 10804 796
rect 10836 764 10964 796
rect 10996 764 11000 796
rect 10640 760 11000 764
rect -720 716 10600 720
rect -720 684 -716 716
rect -684 684 -556 716
rect -524 684 -396 716
rect -364 684 -316 716
rect -284 684 -236 716
rect -204 684 -156 716
rect -124 684 -76 716
rect -44 684 4 716
rect 36 684 84 716
rect 116 684 164 716
rect 196 684 244 716
rect 276 684 324 716
rect 356 684 404 716
rect 436 684 484 716
rect 516 684 564 716
rect 596 684 644 716
rect 676 684 724 716
rect 756 684 804 716
rect 836 684 884 716
rect 916 684 964 716
rect 996 684 1044 716
rect 1076 684 1124 716
rect 1156 684 1204 716
rect 1236 684 1284 716
rect 1316 684 1364 716
rect 1396 684 1444 716
rect 1476 684 1524 716
rect 1556 684 1604 716
rect 1636 684 1684 716
rect 1716 684 1764 716
rect 1796 684 1844 716
rect 1876 684 1924 716
rect 1956 684 2004 716
rect 2036 684 2084 716
rect 2116 684 2164 716
rect 2196 684 2244 716
rect 2276 684 2324 716
rect 2356 684 2404 716
rect 2436 684 2484 716
rect 2516 684 2564 716
rect 2596 684 2644 716
rect 2676 684 2724 716
rect 2756 684 2804 716
rect 2836 684 2884 716
rect 2916 684 2964 716
rect 2996 684 3044 716
rect 3076 684 3124 716
rect 3156 684 3204 716
rect 3236 684 3284 716
rect 3316 684 3364 716
rect 3396 684 3444 716
rect 3476 684 3524 716
rect 3556 684 3604 716
rect 3636 684 3684 716
rect 3716 684 3764 716
rect 3796 684 3844 716
rect 3876 684 3924 716
rect 3956 684 4004 716
rect 4036 684 4084 716
rect 4116 684 4164 716
rect 4196 684 4244 716
rect 4276 684 4324 716
rect 4356 684 4404 716
rect 4436 684 4484 716
rect 4516 684 4564 716
rect 4596 684 4644 716
rect 4676 684 4724 716
rect 4756 684 4804 716
rect 4836 684 4884 716
rect 4916 684 4964 716
rect 4996 684 5044 716
rect 5076 684 5124 716
rect 5156 684 5204 716
rect 5236 684 5284 716
rect 5316 684 5364 716
rect 5396 684 5444 716
rect 5476 684 5524 716
rect 5556 684 5604 716
rect 5636 684 5684 716
rect 5716 684 5764 716
rect 5796 684 5844 716
rect 5876 684 5924 716
rect 5956 684 6004 716
rect 6036 684 6084 716
rect 6116 684 6164 716
rect 6196 684 6244 716
rect 6276 684 6324 716
rect 6356 684 6404 716
rect 6436 684 6484 716
rect 6516 684 6564 716
rect 6596 684 6644 716
rect 6676 684 6724 716
rect 6756 684 6804 716
rect 6836 684 6884 716
rect 6916 684 6964 716
rect 6996 684 7044 716
rect 7076 684 7124 716
rect 7156 684 7204 716
rect 7236 684 7284 716
rect 7316 684 7364 716
rect 7396 684 7444 716
rect 7476 684 7524 716
rect 7556 684 7604 716
rect 7636 684 7684 716
rect 7716 684 7764 716
rect 7796 684 7844 716
rect 7876 684 7924 716
rect 7956 684 8004 716
rect 8036 684 8084 716
rect 8116 684 8164 716
rect 8196 684 8244 716
rect 8276 684 8324 716
rect 8356 684 8404 716
rect 8436 684 8484 716
rect 8516 684 8564 716
rect 8596 684 8644 716
rect 8676 684 8724 716
rect 8756 684 8804 716
rect 8836 684 8884 716
rect 8916 684 8964 716
rect 8996 684 9044 716
rect 9076 684 9124 716
rect 9156 684 9204 716
rect 9236 684 9284 716
rect 9316 684 9364 716
rect 9396 684 9444 716
rect 9476 684 9524 716
rect 9556 684 9604 716
rect 9636 684 9684 716
rect 9716 684 9764 716
rect 9796 684 9844 716
rect 9876 684 9924 716
rect 9956 684 10004 716
rect 10036 684 10084 716
rect 10116 684 10164 716
rect 10196 684 10244 716
rect 10276 684 10324 716
rect 10356 684 10404 716
rect 10436 684 10484 716
rect 10516 684 10600 716
rect -720 680 10600 684
rect 10640 716 11000 720
rect 10640 684 10644 716
rect 10676 684 10804 716
rect 10836 684 10964 716
rect 10996 684 11000 716
rect 10640 680 11000 684
rect -720 636 11000 640
rect -720 604 -716 636
rect -684 604 -556 636
rect -524 604 -396 636
rect -364 604 -316 636
rect -284 604 -236 636
rect -204 604 -156 636
rect -124 604 -76 636
rect -44 604 4 636
rect 36 604 84 636
rect 116 604 164 636
rect 196 604 244 636
rect 276 604 324 636
rect 356 604 404 636
rect 436 604 484 636
rect 516 604 564 636
rect 596 604 644 636
rect 676 604 724 636
rect 756 604 804 636
rect 836 604 884 636
rect 916 604 964 636
rect 996 604 1044 636
rect 1076 604 1124 636
rect 1156 604 1204 636
rect 1236 604 1284 636
rect 1316 604 1364 636
rect 1396 604 1444 636
rect 1476 604 1524 636
rect 1556 604 1604 636
rect 1636 604 1684 636
rect 1716 604 1764 636
rect 1796 604 1844 636
rect 1876 604 1924 636
rect 1956 604 2004 636
rect 2036 604 2084 636
rect 2116 604 2164 636
rect 2196 604 2244 636
rect 2276 604 2324 636
rect 2356 604 2404 636
rect 2436 604 2484 636
rect 2516 604 2564 636
rect 2596 604 2644 636
rect 2676 604 2724 636
rect 2756 604 2804 636
rect 2836 604 2884 636
rect 2916 604 2964 636
rect 2996 604 3044 636
rect 3076 604 3124 636
rect 3156 604 3204 636
rect 3236 604 3284 636
rect 3316 604 3364 636
rect 3396 604 3444 636
rect 3476 604 3524 636
rect 3556 604 3604 636
rect 3636 604 3684 636
rect 3716 604 3764 636
rect 3796 604 3844 636
rect 3876 604 3924 636
rect 3956 604 4004 636
rect 4036 604 4084 636
rect 4116 604 4164 636
rect 4196 604 4244 636
rect 4276 604 4324 636
rect 4356 604 4404 636
rect 4436 604 4484 636
rect 4516 604 4564 636
rect 4596 604 4644 636
rect 4676 604 4724 636
rect 4756 604 4804 636
rect 4836 604 4884 636
rect 4916 604 4964 636
rect 4996 604 5044 636
rect 5076 604 5124 636
rect 5156 604 5204 636
rect 5236 604 5284 636
rect 5316 604 5364 636
rect 5396 604 5444 636
rect 5476 604 5524 636
rect 5556 604 5604 636
rect 5636 604 5684 636
rect 5716 604 5764 636
rect 5796 604 5844 636
rect 5876 604 5924 636
rect 5956 604 6004 636
rect 6036 604 6084 636
rect 6116 604 6164 636
rect 6196 604 6244 636
rect 6276 604 6324 636
rect 6356 604 6404 636
rect 6436 604 6484 636
rect 6516 604 6564 636
rect 6596 604 6644 636
rect 6676 604 6724 636
rect 6756 604 6804 636
rect 6836 604 6884 636
rect 6916 604 6964 636
rect 6996 604 7044 636
rect 7076 604 7124 636
rect 7156 604 7204 636
rect 7236 604 7284 636
rect 7316 604 7364 636
rect 7396 604 7444 636
rect 7476 604 7524 636
rect 7556 604 7604 636
rect 7636 604 7684 636
rect 7716 604 7764 636
rect 7796 604 7844 636
rect 7876 604 7924 636
rect 7956 604 8004 636
rect 8036 604 8084 636
rect 8116 604 8164 636
rect 8196 604 8244 636
rect 8276 604 8324 636
rect 8356 604 8404 636
rect 8436 604 8484 636
rect 8516 604 8564 636
rect 8596 604 8644 636
rect 8676 604 8724 636
rect 8756 604 8804 636
rect 8836 604 8884 636
rect 8916 604 8964 636
rect 8996 604 9044 636
rect 9076 604 9124 636
rect 9156 604 9204 636
rect 9236 604 9284 636
rect 9316 604 9364 636
rect 9396 604 9444 636
rect 9476 604 9524 636
rect 9556 604 9604 636
rect 9636 604 9684 636
rect 9716 604 9764 636
rect 9796 604 9844 636
rect 9876 604 9924 636
rect 9956 604 10004 636
rect 10036 604 10084 636
rect 10116 604 10164 636
rect 10196 604 10244 636
rect 10276 604 10324 636
rect 10356 604 10404 636
rect 10436 604 10484 636
rect 10516 604 10644 636
rect 10676 604 10804 636
rect 10836 604 10964 636
rect 10996 604 11000 636
rect -720 600 11000 604
rect -720 556 11000 560
rect -720 524 -716 556
rect -684 524 -556 556
rect -524 524 -396 556
rect -364 524 -316 556
rect -284 524 -236 556
rect -204 524 -156 556
rect -124 524 -76 556
rect -44 524 4 556
rect 36 524 84 556
rect 116 524 164 556
rect 196 524 244 556
rect 276 524 324 556
rect 356 524 404 556
rect 436 524 484 556
rect 516 524 564 556
rect 596 524 644 556
rect 676 524 724 556
rect 756 524 804 556
rect 836 524 884 556
rect 916 524 964 556
rect 996 524 1044 556
rect 1076 524 1124 556
rect 1156 524 1204 556
rect 1236 524 1284 556
rect 1316 524 1364 556
rect 1396 524 1444 556
rect 1476 524 1524 556
rect 1556 524 1604 556
rect 1636 524 1684 556
rect 1716 524 1764 556
rect 1796 524 1844 556
rect 1876 524 1924 556
rect 1956 524 2004 556
rect 2036 524 2084 556
rect 2116 524 2164 556
rect 2196 524 2244 556
rect 2276 524 2324 556
rect 2356 524 2404 556
rect 2436 524 2484 556
rect 2516 524 2564 556
rect 2596 524 2644 556
rect 2676 524 2724 556
rect 2756 524 2804 556
rect 2836 524 2884 556
rect 2916 524 2964 556
rect 2996 524 3044 556
rect 3076 524 3124 556
rect 3156 524 3204 556
rect 3236 524 3284 556
rect 3316 524 3364 556
rect 3396 524 3444 556
rect 3476 524 3524 556
rect 3556 524 3604 556
rect 3636 524 3684 556
rect 3716 524 3764 556
rect 3796 524 3844 556
rect 3876 524 3924 556
rect 3956 524 4004 556
rect 4036 524 4084 556
rect 4116 524 4164 556
rect 4196 524 4244 556
rect 4276 524 4324 556
rect 4356 524 4404 556
rect 4436 524 4484 556
rect 4516 524 4564 556
rect 4596 524 4644 556
rect 4676 524 4724 556
rect 4756 524 4804 556
rect 4836 524 4884 556
rect 4916 524 4964 556
rect 4996 524 5044 556
rect 5076 524 5124 556
rect 5156 524 5204 556
rect 5236 524 5284 556
rect 5316 524 5364 556
rect 5396 524 5444 556
rect 5476 524 5524 556
rect 5556 524 5604 556
rect 5636 524 5684 556
rect 5716 524 5764 556
rect 5796 524 5844 556
rect 5876 524 5924 556
rect 5956 524 6004 556
rect 6036 524 6084 556
rect 6116 524 6164 556
rect 6196 524 6244 556
rect 6276 524 6324 556
rect 6356 524 6404 556
rect 6436 524 6484 556
rect 6516 524 6564 556
rect 6596 524 6644 556
rect 6676 524 6724 556
rect 6756 524 6804 556
rect 6836 524 6884 556
rect 6916 524 6964 556
rect 6996 524 7044 556
rect 7076 524 7124 556
rect 7156 524 7204 556
rect 7236 524 7284 556
rect 7316 524 7364 556
rect 7396 524 7444 556
rect 7476 524 7524 556
rect 7556 524 7604 556
rect 7636 524 7684 556
rect 7716 524 7764 556
rect 7796 524 7844 556
rect 7876 524 7924 556
rect 7956 524 8004 556
rect 8036 524 8084 556
rect 8116 524 8164 556
rect 8196 524 8244 556
rect 8276 524 8324 556
rect 8356 524 8404 556
rect 8436 524 8484 556
rect 8516 524 8564 556
rect 8596 524 8644 556
rect 8676 524 8724 556
rect 8756 524 8804 556
rect 8836 524 8884 556
rect 8916 524 8964 556
rect 8996 524 9044 556
rect 9076 524 9124 556
rect 9156 524 9204 556
rect 9236 524 9284 556
rect 9316 524 9364 556
rect 9396 524 9444 556
rect 9476 524 9524 556
rect 9556 524 9604 556
rect 9636 524 9684 556
rect 9716 524 9764 556
rect 9796 524 9844 556
rect 9876 524 9924 556
rect 9956 524 10004 556
rect 10036 524 10084 556
rect 10116 524 10164 556
rect 10196 524 10244 556
rect 10276 524 10324 556
rect 10356 524 10404 556
rect 10436 524 10484 556
rect 10516 524 10644 556
rect 10676 524 10804 556
rect 10836 524 10964 556
rect 10996 524 11000 556
rect -720 520 11000 524
rect -720 476 10600 480
rect -720 444 -716 476
rect -684 444 -556 476
rect -524 444 -396 476
rect -364 444 -316 476
rect -284 444 -236 476
rect -204 444 -156 476
rect -124 444 -76 476
rect -44 444 4 476
rect 36 444 84 476
rect 116 444 164 476
rect 196 444 244 476
rect 276 444 324 476
rect 356 444 404 476
rect 436 444 484 476
rect 516 444 564 476
rect 596 444 644 476
rect 676 444 724 476
rect 756 444 804 476
rect 836 444 884 476
rect 916 444 964 476
rect 996 444 1044 476
rect 1076 444 1124 476
rect 1156 444 1204 476
rect 1236 444 1284 476
rect 1316 444 1364 476
rect 1396 444 1444 476
rect 1476 444 1524 476
rect 1556 444 1604 476
rect 1636 444 1684 476
rect 1716 444 1764 476
rect 1796 444 1844 476
rect 1876 444 1924 476
rect 1956 444 2004 476
rect 2036 444 2084 476
rect 2116 444 2164 476
rect 2196 444 2244 476
rect 2276 444 2324 476
rect 2356 444 2404 476
rect 2436 444 2484 476
rect 2516 444 2564 476
rect 2596 444 2644 476
rect 2676 444 2724 476
rect 2756 444 2804 476
rect 2836 444 2884 476
rect 2916 444 2964 476
rect 2996 444 3044 476
rect 3076 444 3124 476
rect 3156 444 3204 476
rect 3236 444 3284 476
rect 3316 444 3364 476
rect 3396 444 3444 476
rect 3476 444 3524 476
rect 3556 444 3604 476
rect 3636 444 3684 476
rect 3716 444 3764 476
rect 3796 444 3844 476
rect 3876 444 3924 476
rect 3956 444 4004 476
rect 4036 444 4084 476
rect 4116 444 4164 476
rect 4196 444 4244 476
rect 4276 444 4324 476
rect 4356 444 4404 476
rect 4436 444 4484 476
rect 4516 444 4564 476
rect 4596 444 4644 476
rect 4676 444 4724 476
rect 4756 444 4804 476
rect 4836 444 4884 476
rect 4916 444 4964 476
rect 4996 444 5044 476
rect 5076 444 5124 476
rect 5156 444 5204 476
rect 5236 444 5284 476
rect 5316 444 5364 476
rect 5396 444 5444 476
rect 5476 444 5524 476
rect 5556 444 5604 476
rect 5636 444 5684 476
rect 5716 444 5764 476
rect 5796 444 5844 476
rect 5876 444 5924 476
rect 5956 444 6004 476
rect 6036 444 6084 476
rect 6116 444 6164 476
rect 6196 444 6244 476
rect 6276 444 6324 476
rect 6356 444 6404 476
rect 6436 444 6484 476
rect 6516 444 6564 476
rect 6596 444 6644 476
rect 6676 444 6724 476
rect 6756 444 6804 476
rect 6836 444 6884 476
rect 6916 444 6964 476
rect 6996 444 7044 476
rect 7076 444 7124 476
rect 7156 444 7204 476
rect 7236 444 7284 476
rect 7316 444 7364 476
rect 7396 444 7444 476
rect 7476 444 7524 476
rect 7556 444 7604 476
rect 7636 444 7684 476
rect 7716 444 7764 476
rect 7796 444 7844 476
rect 7876 444 7924 476
rect 7956 444 8004 476
rect 8036 444 8084 476
rect 8116 444 8164 476
rect 8196 444 8244 476
rect 8276 444 8324 476
rect 8356 444 8404 476
rect 8436 444 8484 476
rect 8516 444 8564 476
rect 8596 444 8644 476
rect 8676 444 8724 476
rect 8756 444 8804 476
rect 8836 444 8884 476
rect 8916 444 8964 476
rect 8996 444 9044 476
rect 9076 444 9124 476
rect 9156 444 9204 476
rect 9236 444 9284 476
rect 9316 444 9364 476
rect 9396 444 9444 476
rect 9476 444 9524 476
rect 9556 444 9604 476
rect 9636 444 9684 476
rect 9716 444 9764 476
rect 9796 444 9844 476
rect 9876 444 9924 476
rect 9956 444 10004 476
rect 10036 444 10084 476
rect 10116 444 10164 476
rect 10196 444 10244 476
rect 10276 444 10324 476
rect 10356 444 10404 476
rect 10436 444 10484 476
rect 10516 444 10600 476
rect -720 440 10600 444
rect 10640 476 11000 480
rect 10640 444 10644 476
rect 10676 444 10804 476
rect 10836 444 10964 476
rect 10996 444 11000 476
rect 10640 440 11000 444
rect -720 396 11000 400
rect -720 364 -716 396
rect -684 364 -556 396
rect -524 364 -396 396
rect -364 364 -316 396
rect -284 364 -236 396
rect -204 364 -156 396
rect -124 364 -76 396
rect -44 364 4 396
rect 36 364 84 396
rect 116 364 164 396
rect 196 364 244 396
rect 276 364 324 396
rect 356 364 404 396
rect 436 364 484 396
rect 516 364 564 396
rect 596 364 644 396
rect 676 364 724 396
rect 756 364 804 396
rect 836 364 884 396
rect 916 364 964 396
rect 996 364 1044 396
rect 1076 364 1124 396
rect 1156 364 1204 396
rect 1236 364 1284 396
rect 1316 364 1364 396
rect 1396 364 1444 396
rect 1476 364 1524 396
rect 1556 364 1604 396
rect 1636 364 1684 396
rect 1716 364 1764 396
rect 1796 364 1844 396
rect 1876 364 1924 396
rect 1956 364 2004 396
rect 2036 364 2084 396
rect 2116 364 2164 396
rect 2196 364 2244 396
rect 2276 364 2324 396
rect 2356 364 2404 396
rect 2436 364 2484 396
rect 2516 364 2564 396
rect 2596 364 2644 396
rect 2676 364 2724 396
rect 2756 364 2804 396
rect 2836 364 2884 396
rect 2916 364 2964 396
rect 2996 364 3044 396
rect 3076 364 3124 396
rect 3156 364 3204 396
rect 3236 364 3284 396
rect 3316 364 3364 396
rect 3396 364 3444 396
rect 3476 364 3524 396
rect 3556 364 3604 396
rect 3636 364 3684 396
rect 3716 364 3764 396
rect 3796 364 3844 396
rect 3876 364 3924 396
rect 3956 364 4004 396
rect 4036 364 4084 396
rect 4116 364 4164 396
rect 4196 364 4244 396
rect 4276 364 4324 396
rect 4356 364 4404 396
rect 4436 364 4484 396
rect 4516 364 4564 396
rect 4596 364 4644 396
rect 4676 364 4724 396
rect 4756 364 4804 396
rect 4836 364 4884 396
rect 4916 364 4964 396
rect 4996 364 5044 396
rect 5076 364 5124 396
rect 5156 364 5204 396
rect 5236 364 5284 396
rect 5316 364 5364 396
rect 5396 364 5444 396
rect 5476 364 5524 396
rect 5556 364 5604 396
rect 5636 364 5684 396
rect 5716 364 5764 396
rect 5796 364 5844 396
rect 5876 364 5924 396
rect 5956 364 6004 396
rect 6036 364 6084 396
rect 6116 364 6164 396
rect 6196 364 6244 396
rect 6276 364 6324 396
rect 6356 364 6404 396
rect 6436 364 6484 396
rect 6516 364 6564 396
rect 6596 364 6644 396
rect 6676 364 6724 396
rect 6756 364 6804 396
rect 6836 364 6884 396
rect 6916 364 6964 396
rect 6996 364 7044 396
rect 7076 364 7124 396
rect 7156 364 7204 396
rect 7236 364 7284 396
rect 7316 364 7364 396
rect 7396 364 7444 396
rect 7476 364 7524 396
rect 7556 364 7604 396
rect 7636 364 7684 396
rect 7716 364 7764 396
rect 7796 364 7844 396
rect 7876 364 7924 396
rect 7956 364 8004 396
rect 8036 364 8084 396
rect 8116 364 8164 396
rect 8196 364 8244 396
rect 8276 364 8324 396
rect 8356 364 8404 396
rect 8436 364 8484 396
rect 8516 364 8564 396
rect 8596 364 8644 396
rect 8676 364 8724 396
rect 8756 364 8804 396
rect 8836 364 8884 396
rect 8916 364 8964 396
rect 8996 364 9044 396
rect 9076 364 9124 396
rect 9156 364 9204 396
rect 9236 364 9284 396
rect 9316 364 9364 396
rect 9396 364 9444 396
rect 9476 364 9524 396
rect 9556 364 9604 396
rect 9636 364 9684 396
rect 9716 364 9764 396
rect 9796 364 9844 396
rect 9876 364 9924 396
rect 9956 364 10004 396
rect 10036 364 10084 396
rect 10116 364 10164 396
rect 10196 364 10244 396
rect 10276 364 10324 396
rect 10356 364 10404 396
rect 10436 364 10484 396
rect 10516 364 10644 396
rect 10676 364 10804 396
rect 10836 364 10964 396
rect 10996 364 11000 396
rect -720 360 11000 364
rect -720 316 -360 320
rect -720 284 -716 316
rect -684 284 -556 316
rect -524 284 -396 316
rect -364 284 -360 316
rect -720 280 -360 284
rect -320 316 11000 320
rect -320 284 -316 316
rect -284 284 -236 316
rect -204 284 -156 316
rect -124 284 -76 316
rect -44 284 4 316
rect 36 284 84 316
rect 116 284 164 316
rect 196 284 244 316
rect 276 284 324 316
rect 356 284 404 316
rect 436 284 484 316
rect 516 284 564 316
rect 596 284 644 316
rect 676 284 724 316
rect 756 284 804 316
rect 836 284 884 316
rect 916 284 964 316
rect 996 284 1044 316
rect 1076 284 1124 316
rect 1156 284 1204 316
rect 1236 284 1284 316
rect 1316 284 1364 316
rect 1396 284 1444 316
rect 1476 284 1524 316
rect 1556 284 1604 316
rect 1636 284 1684 316
rect 1716 284 1764 316
rect 1796 284 1844 316
rect 1876 284 1924 316
rect 1956 284 2004 316
rect 2036 284 2084 316
rect 2116 284 2164 316
rect 2196 284 2244 316
rect 2276 284 2324 316
rect 2356 284 2404 316
rect 2436 284 2484 316
rect 2516 284 2564 316
rect 2596 284 2644 316
rect 2676 284 2724 316
rect 2756 284 2804 316
rect 2836 284 2884 316
rect 2916 284 2964 316
rect 2996 284 3044 316
rect 3076 284 3124 316
rect 3156 284 3204 316
rect 3236 284 3284 316
rect 3316 284 3364 316
rect 3396 284 3444 316
rect 3476 284 3524 316
rect 3556 284 3604 316
rect 3636 284 3684 316
rect 3716 284 3764 316
rect 3796 284 3844 316
rect 3876 284 3924 316
rect 3956 284 4004 316
rect 4036 284 4084 316
rect 4116 284 4164 316
rect 4196 284 4244 316
rect 4276 284 4324 316
rect 4356 284 4404 316
rect 4436 284 4484 316
rect 4516 284 4564 316
rect 4596 284 4644 316
rect 4676 284 4724 316
rect 4756 284 4804 316
rect 4836 284 4884 316
rect 4916 284 4964 316
rect 4996 284 5044 316
rect 5076 284 5124 316
rect 5156 284 5204 316
rect 5236 284 5284 316
rect 5316 284 5364 316
rect 5396 284 5444 316
rect 5476 284 5524 316
rect 5556 284 5604 316
rect 5636 284 5684 316
rect 5716 284 5764 316
rect 5796 284 5844 316
rect 5876 284 5924 316
rect 5956 284 6004 316
rect 6036 284 6084 316
rect 6116 284 6164 316
rect 6196 284 6244 316
rect 6276 284 6324 316
rect 6356 284 6404 316
rect 6436 284 6484 316
rect 6516 284 6564 316
rect 6596 284 6644 316
rect 6676 284 6724 316
rect 6756 284 6804 316
rect 6836 284 6884 316
rect 6916 284 6964 316
rect 6996 284 7044 316
rect 7076 284 7124 316
rect 7156 284 7204 316
rect 7236 284 7284 316
rect 7316 284 7364 316
rect 7396 284 7444 316
rect 7476 284 7524 316
rect 7556 284 7604 316
rect 7636 284 7684 316
rect 7716 284 7764 316
rect 7796 284 7844 316
rect 7876 284 7924 316
rect 7956 284 8004 316
rect 8036 284 8084 316
rect 8116 284 8164 316
rect 8196 284 8244 316
rect 8276 284 8324 316
rect 8356 284 8404 316
rect 8436 284 8484 316
rect 8516 284 8564 316
rect 8596 284 8644 316
rect 8676 284 8724 316
rect 8756 284 8804 316
rect 8836 284 8884 316
rect 8916 284 8964 316
rect 8996 284 9044 316
rect 9076 284 9124 316
rect 9156 284 9204 316
rect 9236 284 9284 316
rect 9316 284 9364 316
rect 9396 284 9444 316
rect 9476 284 9524 316
rect 9556 284 9604 316
rect 9636 284 9684 316
rect 9716 284 9764 316
rect 9796 284 9844 316
rect 9876 284 9924 316
rect 9956 284 10004 316
rect 10036 284 10084 316
rect 10116 284 10164 316
rect 10196 284 10244 316
rect 10276 284 10324 316
rect 10356 284 10404 316
rect 10436 284 10484 316
rect 10516 284 10644 316
rect 10676 284 10804 316
rect 10836 284 10964 316
rect 10996 284 11000 316
rect -320 280 11000 284
rect -720 236 11000 240
rect -720 204 -716 236
rect -684 204 -556 236
rect -524 204 -396 236
rect -364 204 -316 236
rect -284 204 -236 236
rect -204 204 -156 236
rect -124 204 -76 236
rect -44 204 4 236
rect 36 204 84 236
rect 116 204 164 236
rect 196 204 244 236
rect 276 204 324 236
rect 356 204 404 236
rect 436 204 484 236
rect 516 204 564 236
rect 596 204 644 236
rect 676 204 724 236
rect 756 204 804 236
rect 836 204 884 236
rect 916 204 964 236
rect 996 204 1044 236
rect 1076 204 1124 236
rect 1156 204 1204 236
rect 1236 204 1284 236
rect 1316 204 1364 236
rect 1396 204 1444 236
rect 1476 204 1524 236
rect 1556 204 1604 236
rect 1636 204 1684 236
rect 1716 204 1764 236
rect 1796 204 1844 236
rect 1876 204 1924 236
rect 1956 204 2004 236
rect 2036 204 2084 236
rect 2116 204 2164 236
rect 2196 204 2244 236
rect 2276 204 2324 236
rect 2356 204 2404 236
rect 2436 204 2484 236
rect 2516 204 2564 236
rect 2596 204 2644 236
rect 2676 204 2724 236
rect 2756 204 2804 236
rect 2836 204 2884 236
rect 2916 204 2964 236
rect 2996 204 3044 236
rect 3076 204 3124 236
rect 3156 204 3204 236
rect 3236 204 3284 236
rect 3316 204 3364 236
rect 3396 204 3444 236
rect 3476 204 3524 236
rect 3556 204 3604 236
rect 3636 204 3684 236
rect 3716 204 3764 236
rect 3796 204 3844 236
rect 3876 204 3924 236
rect 3956 204 4004 236
rect 4036 204 4084 236
rect 4116 204 4164 236
rect 4196 204 4244 236
rect 4276 204 4324 236
rect 4356 204 4404 236
rect 4436 204 4484 236
rect 4516 204 4564 236
rect 4596 204 4644 236
rect 4676 204 4724 236
rect 4756 204 4804 236
rect 4836 204 4884 236
rect 4916 204 4964 236
rect 4996 204 5044 236
rect 5076 204 5124 236
rect 5156 204 5204 236
rect 5236 204 5284 236
rect 5316 204 5364 236
rect 5396 204 5444 236
rect 5476 204 5524 236
rect 5556 204 5604 236
rect 5636 204 5684 236
rect 5716 204 5764 236
rect 5796 204 5844 236
rect 5876 204 5924 236
rect 5956 204 6004 236
rect 6036 204 6084 236
rect 6116 204 6164 236
rect 6196 204 6244 236
rect 6276 204 6324 236
rect 6356 204 6404 236
rect 6436 204 6484 236
rect 6516 204 6564 236
rect 6596 204 6644 236
rect 6676 204 6724 236
rect 6756 204 6804 236
rect 6836 204 6884 236
rect 6916 204 6964 236
rect 6996 204 7044 236
rect 7076 204 7124 236
rect 7156 204 7204 236
rect 7236 204 7284 236
rect 7316 204 7364 236
rect 7396 204 7444 236
rect 7476 204 7524 236
rect 7556 204 7604 236
rect 7636 204 7684 236
rect 7716 204 7764 236
rect 7796 204 7844 236
rect 7876 204 7924 236
rect 7956 204 8004 236
rect 8036 204 8084 236
rect 8116 204 8164 236
rect 8196 204 8244 236
rect 8276 204 8324 236
rect 8356 204 8404 236
rect 8436 204 8484 236
rect 8516 204 8564 236
rect 8596 204 8644 236
rect 8676 204 8724 236
rect 8756 204 8804 236
rect 8836 204 8884 236
rect 8916 204 8964 236
rect 8996 204 9044 236
rect 9076 204 9124 236
rect 9156 204 9204 236
rect 9236 204 9284 236
rect 9316 204 9364 236
rect 9396 204 9444 236
rect 9476 204 9524 236
rect 9556 204 9604 236
rect 9636 204 9684 236
rect 9716 204 9764 236
rect 9796 204 9844 236
rect 9876 204 9924 236
rect 9956 204 10004 236
rect 10036 204 10084 236
rect 10116 204 10164 236
rect 10196 204 10244 236
rect 10276 204 10324 236
rect 10356 204 10404 236
rect 10436 204 10484 236
rect 10516 204 10644 236
rect 10676 204 10804 236
rect 10836 204 10964 236
rect 10996 204 11000 236
rect -720 200 11000 204
rect -720 156 -360 160
rect -720 124 -716 156
rect -684 124 -556 156
rect -524 124 -396 156
rect -364 124 -360 156
rect -720 120 -360 124
rect -320 156 11000 160
rect -320 124 -316 156
rect -284 124 -236 156
rect -204 124 -156 156
rect -124 124 -76 156
rect -44 124 4 156
rect 36 124 84 156
rect 116 124 164 156
rect 196 124 244 156
rect 276 124 324 156
rect 356 124 404 156
rect 436 124 484 156
rect 516 124 564 156
rect 596 124 644 156
rect 676 124 724 156
rect 756 124 804 156
rect 836 124 884 156
rect 916 124 964 156
rect 996 124 1044 156
rect 1076 124 1124 156
rect 1156 124 1204 156
rect 1236 124 1284 156
rect 1316 124 1364 156
rect 1396 124 1444 156
rect 1476 124 1524 156
rect 1556 124 1604 156
rect 1636 124 1684 156
rect 1716 124 1764 156
rect 1796 124 1844 156
rect 1876 124 1924 156
rect 1956 124 2004 156
rect 2036 124 2084 156
rect 2116 124 2164 156
rect 2196 124 2244 156
rect 2276 124 2324 156
rect 2356 124 2404 156
rect 2436 124 2484 156
rect 2516 124 2564 156
rect 2596 124 2644 156
rect 2676 124 2724 156
rect 2756 124 2804 156
rect 2836 124 2884 156
rect 2916 124 2964 156
rect 2996 124 3044 156
rect 3076 124 3124 156
rect 3156 124 3204 156
rect 3236 124 3284 156
rect 3316 124 3364 156
rect 3396 124 3444 156
rect 3476 124 3524 156
rect 3556 124 3604 156
rect 3636 124 3684 156
rect 3716 124 3764 156
rect 3796 124 3844 156
rect 3876 124 3924 156
rect 3956 124 4004 156
rect 4036 124 4084 156
rect 4116 124 4164 156
rect 4196 124 4244 156
rect 4276 124 4324 156
rect 4356 124 4404 156
rect 4436 124 4484 156
rect 4516 124 4564 156
rect 4596 124 4644 156
rect 4676 124 4724 156
rect 4756 124 4804 156
rect 4836 124 4884 156
rect 4916 124 4964 156
rect 4996 124 5044 156
rect 5076 124 5124 156
rect 5156 124 5204 156
rect 5236 124 5284 156
rect 5316 124 5364 156
rect 5396 124 5444 156
rect 5476 124 5524 156
rect 5556 124 5604 156
rect 5636 124 5684 156
rect 5716 124 5764 156
rect 5796 124 5844 156
rect 5876 124 5924 156
rect 5956 124 6004 156
rect 6036 124 6084 156
rect 6116 124 6164 156
rect 6196 124 6244 156
rect 6276 124 6324 156
rect 6356 124 6404 156
rect 6436 124 6484 156
rect 6516 124 6564 156
rect 6596 124 6644 156
rect 6676 124 6724 156
rect 6756 124 6804 156
rect 6836 124 6884 156
rect 6916 124 6964 156
rect 6996 124 7044 156
rect 7076 124 7124 156
rect 7156 124 7204 156
rect 7236 124 7284 156
rect 7316 124 7364 156
rect 7396 124 7444 156
rect 7476 124 7524 156
rect 7556 124 7604 156
rect 7636 124 7684 156
rect 7716 124 7764 156
rect 7796 124 7844 156
rect 7876 124 7924 156
rect 7956 124 8004 156
rect 8036 124 8084 156
rect 8116 124 8164 156
rect 8196 124 8244 156
rect 8276 124 8324 156
rect 8356 124 8404 156
rect 8436 124 8484 156
rect 8516 124 8564 156
rect 8596 124 8644 156
rect 8676 124 8724 156
rect 8756 124 8804 156
rect 8836 124 8884 156
rect 8916 124 8964 156
rect 8996 124 9044 156
rect 9076 124 9124 156
rect 9156 124 9204 156
rect 9236 124 9284 156
rect 9316 124 9364 156
rect 9396 124 9444 156
rect 9476 124 9524 156
rect 9556 124 9604 156
rect 9636 124 9684 156
rect 9716 124 9764 156
rect 9796 124 9844 156
rect 9876 124 9924 156
rect 9956 124 10004 156
rect 10036 124 10084 156
rect 10116 124 10164 156
rect 10196 124 10244 156
rect 10276 124 10324 156
rect 10356 124 10404 156
rect 10436 124 10484 156
rect 10516 124 10644 156
rect 10676 124 10804 156
rect 10836 124 10964 156
rect 10996 124 11000 156
rect -320 120 11000 124
rect -720 76 11000 80
rect -720 44 -716 76
rect -684 44 -556 76
rect -524 44 -396 76
rect -364 44 -316 76
rect -284 44 -236 76
rect -204 44 -156 76
rect -124 44 -76 76
rect -44 44 4 76
rect 36 44 84 76
rect 116 44 164 76
rect 196 44 244 76
rect 276 44 324 76
rect 356 44 404 76
rect 436 44 484 76
rect 516 44 564 76
rect 596 44 644 76
rect 676 44 724 76
rect 756 44 804 76
rect 836 44 884 76
rect 916 44 964 76
rect 996 44 1044 76
rect 1076 44 1124 76
rect 1156 44 1204 76
rect 1236 44 1284 76
rect 1316 44 1364 76
rect 1396 44 1444 76
rect 1476 44 1524 76
rect 1556 44 1604 76
rect 1636 44 1684 76
rect 1716 44 1764 76
rect 1796 44 1844 76
rect 1876 44 1924 76
rect 1956 44 2004 76
rect 2036 44 2084 76
rect 2116 44 2164 76
rect 2196 44 2244 76
rect 2276 44 2324 76
rect 2356 44 2404 76
rect 2436 44 2484 76
rect 2516 44 2564 76
rect 2596 44 2644 76
rect 2676 44 2724 76
rect 2756 44 2804 76
rect 2836 44 2884 76
rect 2916 44 2964 76
rect 2996 44 3044 76
rect 3076 44 3124 76
rect 3156 44 3204 76
rect 3236 44 3284 76
rect 3316 44 3364 76
rect 3396 44 3444 76
rect 3476 44 3524 76
rect 3556 44 3604 76
rect 3636 44 3684 76
rect 3716 44 3764 76
rect 3796 44 3844 76
rect 3876 44 3924 76
rect 3956 44 4004 76
rect 4036 44 4084 76
rect 4116 44 4164 76
rect 4196 44 4244 76
rect 4276 44 4324 76
rect 4356 44 4404 76
rect 4436 44 4484 76
rect 4516 44 4564 76
rect 4596 44 4644 76
rect 4676 44 4724 76
rect 4756 44 4804 76
rect 4836 44 4884 76
rect 4916 44 4964 76
rect 4996 44 5044 76
rect 5076 44 5124 76
rect 5156 44 5204 76
rect 5236 44 5284 76
rect 5316 44 5364 76
rect 5396 44 5444 76
rect 5476 44 5524 76
rect 5556 44 5604 76
rect 5636 44 5684 76
rect 5716 44 5764 76
rect 5796 44 5844 76
rect 5876 44 5924 76
rect 5956 44 6004 76
rect 6036 44 6084 76
rect 6116 44 6164 76
rect 6196 44 6244 76
rect 6276 44 6324 76
rect 6356 44 6404 76
rect 6436 44 6484 76
rect 6516 44 6564 76
rect 6596 44 6644 76
rect 6676 44 6724 76
rect 6756 44 6804 76
rect 6836 44 6884 76
rect 6916 44 6964 76
rect 6996 44 7044 76
rect 7076 44 7124 76
rect 7156 44 7204 76
rect 7236 44 7284 76
rect 7316 44 7364 76
rect 7396 44 7444 76
rect 7476 44 7524 76
rect 7556 44 7604 76
rect 7636 44 7684 76
rect 7716 44 7764 76
rect 7796 44 7844 76
rect 7876 44 7924 76
rect 7956 44 8004 76
rect 8036 44 8084 76
rect 8116 44 8164 76
rect 8196 44 8244 76
rect 8276 44 8324 76
rect 8356 44 8404 76
rect 8436 44 8484 76
rect 8516 44 8564 76
rect 8596 44 8644 76
rect 8676 44 8724 76
rect 8756 44 8804 76
rect 8836 44 8884 76
rect 8916 44 8964 76
rect 8996 44 9044 76
rect 9076 44 9124 76
rect 9156 44 9204 76
rect 9236 44 9284 76
rect 9316 44 9364 76
rect 9396 44 9444 76
rect 9476 44 9524 76
rect 9556 44 9604 76
rect 9636 44 9684 76
rect 9716 44 9764 76
rect 9796 44 9844 76
rect 9876 44 9924 76
rect 9956 44 10004 76
rect 10036 44 10084 76
rect 10116 44 10164 76
rect 10196 44 10244 76
rect 10276 44 10324 76
rect 10356 44 10404 76
rect 10436 44 10484 76
rect 10516 44 10644 76
rect 10676 44 10804 76
rect 10836 44 10964 76
rect 10996 44 11000 76
rect -720 40 11000 44
rect -720 -4 11000 0
rect -720 -36 -716 -4
rect -684 -36 -556 -4
rect -524 -36 -396 -4
rect -364 -36 -316 -4
rect -284 -36 -236 -4
rect -204 -36 -156 -4
rect -124 -36 -76 -4
rect -44 -36 4 -4
rect 36 -36 84 -4
rect 116 -36 164 -4
rect 196 -36 244 -4
rect 276 -36 324 -4
rect 356 -36 404 -4
rect 436 -36 484 -4
rect 516 -36 564 -4
rect 596 -36 644 -4
rect 676 -36 724 -4
rect 756 -36 804 -4
rect 836 -36 884 -4
rect 916 -36 964 -4
rect 996 -36 1044 -4
rect 1076 -36 1124 -4
rect 1156 -36 1204 -4
rect 1236 -36 1284 -4
rect 1316 -36 1364 -4
rect 1396 -36 1444 -4
rect 1476 -36 1524 -4
rect 1556 -36 1604 -4
rect 1636 -36 1684 -4
rect 1716 -36 1764 -4
rect 1796 -36 1844 -4
rect 1876 -36 1924 -4
rect 1956 -36 2004 -4
rect 2036 -36 2084 -4
rect 2116 -36 2164 -4
rect 2196 -36 2244 -4
rect 2276 -36 2324 -4
rect 2356 -36 2404 -4
rect 2436 -36 2484 -4
rect 2516 -36 2564 -4
rect 2596 -36 2644 -4
rect 2676 -36 2724 -4
rect 2756 -36 2804 -4
rect 2836 -36 2884 -4
rect 2916 -36 2964 -4
rect 2996 -36 3044 -4
rect 3076 -36 3124 -4
rect 3156 -36 3204 -4
rect 3236 -36 3284 -4
rect 3316 -36 3364 -4
rect 3396 -36 3444 -4
rect 3476 -36 3524 -4
rect 3556 -36 3604 -4
rect 3636 -36 3684 -4
rect 3716 -36 3764 -4
rect 3796 -36 3844 -4
rect 3876 -36 3924 -4
rect 3956 -36 4004 -4
rect 4036 -36 4084 -4
rect 4116 -36 4164 -4
rect 4196 -36 4244 -4
rect 4276 -36 4324 -4
rect 4356 -36 4404 -4
rect 4436 -36 4484 -4
rect 4516 -36 4564 -4
rect 4596 -36 4644 -4
rect 4676 -36 4724 -4
rect 4756 -36 4804 -4
rect 4836 -36 4884 -4
rect 4916 -36 4964 -4
rect 4996 -36 5044 -4
rect 5076 -36 5124 -4
rect 5156 -36 5204 -4
rect 5236 -36 5284 -4
rect 5316 -36 5364 -4
rect 5396 -36 5444 -4
rect 5476 -36 5524 -4
rect 5556 -36 5604 -4
rect 5636 -36 5684 -4
rect 5716 -36 5764 -4
rect 5796 -36 5844 -4
rect 5876 -36 5924 -4
rect 5956 -36 6004 -4
rect 6036 -36 6084 -4
rect 6116 -36 6164 -4
rect 6196 -36 6244 -4
rect 6276 -36 6324 -4
rect 6356 -36 6404 -4
rect 6436 -36 6484 -4
rect 6516 -36 6564 -4
rect 6596 -36 6644 -4
rect 6676 -36 6724 -4
rect 6756 -36 6804 -4
rect 6836 -36 6884 -4
rect 6916 -36 6964 -4
rect 6996 -36 7044 -4
rect 7076 -36 7124 -4
rect 7156 -36 7204 -4
rect 7236 -36 7284 -4
rect 7316 -36 7364 -4
rect 7396 -36 7444 -4
rect 7476 -36 7524 -4
rect 7556 -36 7604 -4
rect 7636 -36 7684 -4
rect 7716 -36 7764 -4
rect 7796 -36 7844 -4
rect 7876 -36 7924 -4
rect 7956 -36 8004 -4
rect 8036 -36 8084 -4
rect 8116 -36 8164 -4
rect 8196 -36 8244 -4
rect 8276 -36 8324 -4
rect 8356 -36 8404 -4
rect 8436 -36 8484 -4
rect 8516 -36 8564 -4
rect 8596 -36 8644 -4
rect 8676 -36 8724 -4
rect 8756 -36 8804 -4
rect 8836 -36 8884 -4
rect 8916 -36 8964 -4
rect 8996 -36 9044 -4
rect 9076 -36 9124 -4
rect 9156 -36 9204 -4
rect 9236 -36 9284 -4
rect 9316 -36 9364 -4
rect 9396 -36 9444 -4
rect 9476 -36 9524 -4
rect 9556 -36 9604 -4
rect 9636 -36 9684 -4
rect 9716 -36 9764 -4
rect 9796 -36 9844 -4
rect 9876 -36 9924 -4
rect 9956 -36 10004 -4
rect 10036 -36 10084 -4
rect 10116 -36 10164 -4
rect 10196 -36 10244 -4
rect 10276 -36 10324 -4
rect 10356 -36 10404 -4
rect 10436 -36 10484 -4
rect 10516 -36 10644 -4
rect 10676 -36 10804 -4
rect 10836 -36 10964 -4
rect 10996 -36 11000 -4
rect -720 -40 11000 -36
rect -720 -84 11000 -80
rect -720 -116 -716 -84
rect -684 -116 -556 -84
rect -524 -116 -396 -84
rect -364 -116 -316 -84
rect -284 -116 -236 -84
rect -204 -116 -156 -84
rect -124 -116 -76 -84
rect -44 -116 4 -84
rect 36 -116 84 -84
rect 116 -116 164 -84
rect 196 -116 244 -84
rect 276 -116 324 -84
rect 356 -116 404 -84
rect 436 -116 484 -84
rect 516 -116 564 -84
rect 596 -116 644 -84
rect 676 -116 724 -84
rect 756 -116 804 -84
rect 836 -116 884 -84
rect 916 -116 964 -84
rect 996 -116 1044 -84
rect 1076 -116 1124 -84
rect 1156 -116 1204 -84
rect 1236 -116 1284 -84
rect 1316 -116 1364 -84
rect 1396 -116 1444 -84
rect 1476 -116 1524 -84
rect 1556 -116 1604 -84
rect 1636 -116 1684 -84
rect 1716 -116 1764 -84
rect 1796 -116 1844 -84
rect 1876 -116 1924 -84
rect 1956 -116 2004 -84
rect 2036 -116 2084 -84
rect 2116 -116 2164 -84
rect 2196 -116 2244 -84
rect 2276 -116 2324 -84
rect 2356 -116 2404 -84
rect 2436 -116 2484 -84
rect 2516 -116 2564 -84
rect 2596 -116 2644 -84
rect 2676 -116 2724 -84
rect 2756 -116 2804 -84
rect 2836 -116 2884 -84
rect 2916 -116 2964 -84
rect 2996 -116 3044 -84
rect 3076 -116 3124 -84
rect 3156 -116 3204 -84
rect 3236 -116 3284 -84
rect 3316 -116 3364 -84
rect 3396 -116 3444 -84
rect 3476 -116 3524 -84
rect 3556 -116 3604 -84
rect 3636 -116 3684 -84
rect 3716 -116 3764 -84
rect 3796 -116 3844 -84
rect 3876 -116 3924 -84
rect 3956 -116 4004 -84
rect 4036 -116 4084 -84
rect 4116 -116 4164 -84
rect 4196 -116 4244 -84
rect 4276 -116 4324 -84
rect 4356 -116 4404 -84
rect 4436 -116 4484 -84
rect 4516 -116 4564 -84
rect 4596 -116 4644 -84
rect 4676 -116 4724 -84
rect 4756 -116 4804 -84
rect 4836 -116 4884 -84
rect 4916 -116 4964 -84
rect 4996 -116 5044 -84
rect 5076 -116 5124 -84
rect 5156 -116 5204 -84
rect 5236 -116 5284 -84
rect 5316 -116 5364 -84
rect 5396 -116 5444 -84
rect 5476 -116 5524 -84
rect 5556 -116 5604 -84
rect 5636 -116 5684 -84
rect 5716 -116 5764 -84
rect 5796 -116 5844 -84
rect 5876 -116 5924 -84
rect 5956 -116 6004 -84
rect 6036 -116 6084 -84
rect 6116 -116 6164 -84
rect 6196 -116 6244 -84
rect 6276 -116 6324 -84
rect 6356 -116 6404 -84
rect 6436 -116 6484 -84
rect 6516 -116 6564 -84
rect 6596 -116 6644 -84
rect 6676 -116 6724 -84
rect 6756 -116 6804 -84
rect 6836 -116 6884 -84
rect 6916 -116 6964 -84
rect 6996 -116 7044 -84
rect 7076 -116 7124 -84
rect 7156 -116 7204 -84
rect 7236 -116 7284 -84
rect 7316 -116 7364 -84
rect 7396 -116 7444 -84
rect 7476 -116 7524 -84
rect 7556 -116 7604 -84
rect 7636 -116 7684 -84
rect 7716 -116 7764 -84
rect 7796 -116 7844 -84
rect 7876 -116 7924 -84
rect 7956 -116 8004 -84
rect 8036 -116 8084 -84
rect 8116 -116 8164 -84
rect 8196 -116 8244 -84
rect 8276 -116 8324 -84
rect 8356 -116 8404 -84
rect 8436 -116 8484 -84
rect 8516 -116 8564 -84
rect 8596 -116 8644 -84
rect 8676 -116 8724 -84
rect 8756 -116 8804 -84
rect 8836 -116 8884 -84
rect 8916 -116 8964 -84
rect 8996 -116 9044 -84
rect 9076 -116 9124 -84
rect 9156 -116 9204 -84
rect 9236 -116 9284 -84
rect 9316 -116 9364 -84
rect 9396 -116 9444 -84
rect 9476 -116 9524 -84
rect 9556 -116 9604 -84
rect 9636 -116 9684 -84
rect 9716 -116 9764 -84
rect 9796 -116 9844 -84
rect 9876 -116 9924 -84
rect 9956 -116 10004 -84
rect 10036 -116 10084 -84
rect 10116 -116 10164 -84
rect 10196 -116 10244 -84
rect 10276 -116 10324 -84
rect 10356 -116 10404 -84
rect 10436 -116 10484 -84
rect 10516 -116 10644 -84
rect 10676 -116 10804 -84
rect 10836 -116 10964 -84
rect 10996 -116 11000 -84
rect -720 -120 11000 -116
rect -720 -164 11000 -160
rect -720 -196 -716 -164
rect -684 -196 -556 -164
rect -524 -196 -396 -164
rect -364 -196 -236 -164
rect -204 -196 -156 -164
rect -124 -196 -76 -164
rect -44 -196 4 -164
rect 36 -196 84 -164
rect 116 -196 164 -164
rect 196 -196 244 -164
rect 276 -196 324 -164
rect 356 -196 404 -164
rect 436 -196 484 -164
rect 516 -196 564 -164
rect 596 -196 644 -164
rect 676 -196 724 -164
rect 756 -196 804 -164
rect 836 -196 884 -164
rect 916 -196 964 -164
rect 996 -196 1044 -164
rect 1076 -196 1124 -164
rect 1156 -196 1204 -164
rect 1236 -196 1284 -164
rect 1316 -196 1364 -164
rect 1396 -196 1444 -164
rect 1476 -196 1524 -164
rect 1556 -196 1604 -164
rect 1636 -196 1684 -164
rect 1716 -196 1764 -164
rect 1796 -196 1844 -164
rect 1876 -196 1924 -164
rect 1956 -196 2004 -164
rect 2036 -196 2084 -164
rect 2116 -196 2164 -164
rect 2196 -196 2244 -164
rect 2276 -196 2324 -164
rect 2356 -196 2404 -164
rect 2436 -196 2484 -164
rect 2516 -196 2564 -164
rect 2596 -196 2644 -164
rect 2676 -196 2724 -164
rect 2756 -196 2804 -164
rect 2836 -196 2884 -164
rect 2916 -196 2964 -164
rect 2996 -196 3044 -164
rect 3076 -196 3124 -164
rect 3156 -196 3204 -164
rect 3236 -196 3284 -164
rect 3316 -196 3364 -164
rect 3396 -196 3444 -164
rect 3476 -196 3524 -164
rect 3556 -196 3604 -164
rect 3636 -196 3684 -164
rect 3716 -196 3764 -164
rect 3796 -196 3844 -164
rect 3876 -196 3924 -164
rect 3956 -196 4004 -164
rect 4036 -196 4084 -164
rect 4116 -196 4164 -164
rect 4196 -196 4244 -164
rect 4276 -196 4324 -164
rect 4356 -196 4404 -164
rect 4436 -196 4484 -164
rect 4516 -196 4564 -164
rect 4596 -196 4644 -164
rect 4676 -196 4724 -164
rect 4756 -196 4804 -164
rect 4836 -196 4884 -164
rect 4916 -196 4964 -164
rect 4996 -196 5044 -164
rect 5076 -196 5124 -164
rect 5156 -196 5204 -164
rect 5236 -196 5284 -164
rect 5316 -196 5364 -164
rect 5396 -196 5444 -164
rect 5476 -196 5524 -164
rect 5556 -196 5604 -164
rect 5636 -196 5684 -164
rect 5716 -196 5764 -164
rect 5796 -196 5844 -164
rect 5876 -196 5924 -164
rect 5956 -196 6004 -164
rect 6036 -196 6084 -164
rect 6116 -196 6164 -164
rect 6196 -196 6244 -164
rect 6276 -196 6324 -164
rect 6356 -196 6404 -164
rect 6436 -196 6484 -164
rect 6516 -196 6564 -164
rect 6596 -196 6644 -164
rect 6676 -196 6724 -164
rect 6756 -196 6804 -164
rect 6836 -196 6884 -164
rect 6916 -196 6964 -164
rect 6996 -196 7044 -164
rect 7076 -196 7124 -164
rect 7156 -196 7204 -164
rect 7236 -196 7284 -164
rect 7316 -196 7364 -164
rect 7396 -196 7444 -164
rect 7476 -196 7524 -164
rect 7556 -196 7604 -164
rect 7636 -196 7684 -164
rect 7716 -196 7764 -164
rect 7796 -196 7844 -164
rect 7876 -196 7924 -164
rect 7956 -196 8004 -164
rect 8036 -196 8084 -164
rect 8116 -196 8164 -164
rect 8196 -196 8244 -164
rect 8276 -196 8324 -164
rect 8356 -196 8404 -164
rect 8436 -196 8484 -164
rect 8516 -196 8564 -164
rect 8596 -196 8644 -164
rect 8676 -196 8724 -164
rect 8756 -196 8804 -164
rect 8836 -196 8884 -164
rect 8916 -196 8964 -164
rect 8996 -196 9044 -164
rect 9076 -196 9124 -164
rect 9156 -196 9204 -164
rect 9236 -196 9284 -164
rect 9316 -196 9364 -164
rect 9396 -196 9444 -164
rect 9476 -196 9524 -164
rect 9556 -196 9604 -164
rect 9636 -196 9684 -164
rect 9716 -196 9764 -164
rect 9796 -196 9844 -164
rect 9876 -196 9924 -164
rect 9956 -196 10004 -164
rect 10036 -196 10084 -164
rect 10116 -196 10164 -164
rect 10196 -196 10244 -164
rect 10276 -196 10324 -164
rect 10356 -196 10404 -164
rect 10436 -196 10484 -164
rect 10516 -196 10564 -164
rect 10596 -196 10644 -164
rect 10676 -196 10804 -164
rect 10836 -196 10964 -164
rect 10996 -196 11000 -164
rect -720 -200 11000 -196
rect -720 -244 11000 -240
rect -720 -276 -716 -244
rect -684 -276 -556 -244
rect -524 -276 -396 -244
rect -364 -276 -236 -244
rect -204 -276 -156 -244
rect -124 -276 -76 -244
rect -44 -276 4 -244
rect 36 -276 84 -244
rect 116 -276 164 -244
rect 196 -276 244 -244
rect 276 -276 324 -244
rect 356 -276 404 -244
rect 436 -276 484 -244
rect 516 -276 564 -244
rect 596 -276 644 -244
rect 676 -276 724 -244
rect 756 -276 804 -244
rect 836 -276 884 -244
rect 916 -276 964 -244
rect 996 -276 1044 -244
rect 1076 -276 1124 -244
rect 1156 -276 1204 -244
rect 1236 -276 1284 -244
rect 1316 -276 1364 -244
rect 1396 -276 1444 -244
rect 1476 -276 1524 -244
rect 1556 -276 1604 -244
rect 1636 -276 1684 -244
rect 1716 -276 1764 -244
rect 1796 -276 1844 -244
rect 1876 -276 1924 -244
rect 1956 -276 2004 -244
rect 2036 -276 2084 -244
rect 2116 -276 2164 -244
rect 2196 -276 2244 -244
rect 2276 -276 2324 -244
rect 2356 -276 2404 -244
rect 2436 -276 2484 -244
rect 2516 -276 2564 -244
rect 2596 -276 2644 -244
rect 2676 -276 2724 -244
rect 2756 -276 2804 -244
rect 2836 -276 2884 -244
rect 2916 -276 2964 -244
rect 2996 -276 3044 -244
rect 3076 -276 3124 -244
rect 3156 -276 3204 -244
rect 3236 -276 3284 -244
rect 3316 -276 3364 -244
rect 3396 -276 3444 -244
rect 3476 -276 3524 -244
rect 3556 -276 3604 -244
rect 3636 -276 3684 -244
rect 3716 -276 3764 -244
rect 3796 -276 3844 -244
rect 3876 -276 3924 -244
rect 3956 -276 4004 -244
rect 4036 -276 4084 -244
rect 4116 -276 4164 -244
rect 4196 -276 4244 -244
rect 4276 -276 4324 -244
rect 4356 -276 4404 -244
rect 4436 -276 4484 -244
rect 4516 -276 4564 -244
rect 4596 -276 4644 -244
rect 4676 -276 4724 -244
rect 4756 -276 4804 -244
rect 4836 -276 4884 -244
rect 4916 -276 4964 -244
rect 4996 -276 5044 -244
rect 5076 -276 5124 -244
rect 5156 -276 5204 -244
rect 5236 -276 5284 -244
rect 5316 -276 5364 -244
rect 5396 -276 5444 -244
rect 5476 -276 5524 -244
rect 5556 -276 5604 -244
rect 5636 -276 5684 -244
rect 5716 -276 5764 -244
rect 5796 -276 5844 -244
rect 5876 -276 5924 -244
rect 5956 -276 6004 -244
rect 6036 -276 6084 -244
rect 6116 -276 6164 -244
rect 6196 -276 6244 -244
rect 6276 -276 6324 -244
rect 6356 -276 6404 -244
rect 6436 -276 6484 -244
rect 6516 -276 6564 -244
rect 6596 -276 6644 -244
rect 6676 -276 6724 -244
rect 6756 -276 6804 -244
rect 6836 -276 6884 -244
rect 6916 -276 6964 -244
rect 6996 -276 7044 -244
rect 7076 -276 7124 -244
rect 7156 -276 7204 -244
rect 7236 -276 7284 -244
rect 7316 -276 7364 -244
rect 7396 -276 7444 -244
rect 7476 -276 7524 -244
rect 7556 -276 7604 -244
rect 7636 -276 7684 -244
rect 7716 -276 7764 -244
rect 7796 -276 7844 -244
rect 7876 -276 7924 -244
rect 7956 -276 8004 -244
rect 8036 -276 8084 -244
rect 8116 -276 8164 -244
rect 8196 -276 8244 -244
rect 8276 -276 8324 -244
rect 8356 -276 8404 -244
rect 8436 -276 8484 -244
rect 8516 -276 8564 -244
rect 8596 -276 8644 -244
rect 8676 -276 8724 -244
rect 8756 -276 8804 -244
rect 8836 -276 8884 -244
rect 8916 -276 8964 -244
rect 8996 -276 9044 -244
rect 9076 -276 9124 -244
rect 9156 -276 9204 -244
rect 9236 -276 9284 -244
rect 9316 -276 9364 -244
rect 9396 -276 9444 -244
rect 9476 -276 9524 -244
rect 9556 -276 9604 -244
rect 9636 -276 9684 -244
rect 9716 -276 9764 -244
rect 9796 -276 9844 -244
rect 9876 -276 9924 -244
rect 9956 -276 10004 -244
rect 10036 -276 10084 -244
rect 10116 -276 10164 -244
rect 10196 -276 10244 -244
rect 10276 -276 10324 -244
rect 10356 -276 10404 -244
rect 10436 -276 10484 -244
rect 10516 -276 10564 -244
rect 10596 -276 10644 -244
rect 10676 -276 10804 -244
rect 10836 -276 10964 -244
rect 10996 -276 11000 -244
rect -720 -280 11000 -276
rect -720 -324 11000 -320
rect -720 -356 -716 -324
rect -684 -356 -556 -324
rect -524 -356 -396 -324
rect -364 -356 -236 -324
rect -204 -356 -156 -324
rect -124 -356 -76 -324
rect -44 -356 4 -324
rect 36 -356 84 -324
rect 116 -356 164 -324
rect 196 -356 244 -324
rect 276 -356 324 -324
rect 356 -356 404 -324
rect 436 -356 484 -324
rect 516 -356 564 -324
rect 596 -356 644 -324
rect 676 -356 724 -324
rect 756 -356 804 -324
rect 836 -356 884 -324
rect 916 -356 964 -324
rect 996 -356 1044 -324
rect 1076 -356 1124 -324
rect 1156 -356 1204 -324
rect 1236 -356 1284 -324
rect 1316 -356 1364 -324
rect 1396 -356 1444 -324
rect 1476 -356 1524 -324
rect 1556 -356 1604 -324
rect 1636 -356 1684 -324
rect 1716 -356 1764 -324
rect 1796 -356 1844 -324
rect 1876 -356 1924 -324
rect 1956 -356 2004 -324
rect 2036 -356 2084 -324
rect 2116 -356 2164 -324
rect 2196 -356 2244 -324
rect 2276 -356 2324 -324
rect 2356 -356 2404 -324
rect 2436 -356 2484 -324
rect 2516 -356 2564 -324
rect 2596 -356 2644 -324
rect 2676 -356 2724 -324
rect 2756 -356 2804 -324
rect 2836 -356 2884 -324
rect 2916 -356 2964 -324
rect 2996 -356 3044 -324
rect 3076 -356 3124 -324
rect 3156 -356 3204 -324
rect 3236 -356 3284 -324
rect 3316 -356 3364 -324
rect 3396 -356 3444 -324
rect 3476 -356 3524 -324
rect 3556 -356 3604 -324
rect 3636 -356 3684 -324
rect 3716 -356 3764 -324
rect 3796 -356 3844 -324
rect 3876 -356 3924 -324
rect 3956 -356 4004 -324
rect 4036 -356 4084 -324
rect 4116 -356 4164 -324
rect 4196 -356 4244 -324
rect 4276 -356 4324 -324
rect 4356 -356 4404 -324
rect 4436 -356 4484 -324
rect 4516 -356 4564 -324
rect 4596 -356 4644 -324
rect 4676 -356 4724 -324
rect 4756 -356 4804 -324
rect 4836 -356 4884 -324
rect 4916 -356 4964 -324
rect 4996 -356 5044 -324
rect 5076 -356 5124 -324
rect 5156 -356 5204 -324
rect 5236 -356 5284 -324
rect 5316 -356 5364 -324
rect 5396 -356 5444 -324
rect 5476 -356 5524 -324
rect 5556 -356 5604 -324
rect 5636 -356 5684 -324
rect 5716 -356 5764 -324
rect 5796 -356 5844 -324
rect 5876 -356 5924 -324
rect 5956 -356 6004 -324
rect 6036 -356 6084 -324
rect 6116 -356 6164 -324
rect 6196 -356 6244 -324
rect 6276 -356 6324 -324
rect 6356 -356 6404 -324
rect 6436 -356 6484 -324
rect 6516 -356 6564 -324
rect 6596 -356 6644 -324
rect 6676 -356 6724 -324
rect 6756 -356 6804 -324
rect 6836 -356 6884 -324
rect 6916 -356 6964 -324
rect 6996 -356 7044 -324
rect 7076 -356 7124 -324
rect 7156 -356 7204 -324
rect 7236 -356 7284 -324
rect 7316 -356 7364 -324
rect 7396 -356 7444 -324
rect 7476 -356 7524 -324
rect 7556 -356 7604 -324
rect 7636 -356 7684 -324
rect 7716 -356 7764 -324
rect 7796 -356 7844 -324
rect 7876 -356 7924 -324
rect 7956 -356 8004 -324
rect 8036 -356 8084 -324
rect 8116 -356 8164 -324
rect 8196 -356 8244 -324
rect 8276 -356 8324 -324
rect 8356 -356 8404 -324
rect 8436 -356 8484 -324
rect 8516 -356 8564 -324
rect 8596 -356 8644 -324
rect 8676 -356 8724 -324
rect 8756 -356 8804 -324
rect 8836 -356 8884 -324
rect 8916 -356 8964 -324
rect 8996 -356 9044 -324
rect 9076 -356 9124 -324
rect 9156 -356 9204 -324
rect 9236 -356 9284 -324
rect 9316 -356 9364 -324
rect 9396 -356 9444 -324
rect 9476 -356 9524 -324
rect 9556 -356 9604 -324
rect 9636 -356 9684 -324
rect 9716 -356 9764 -324
rect 9796 -356 9844 -324
rect 9876 -356 9924 -324
rect 9956 -356 10004 -324
rect 10036 -356 10084 -324
rect 10116 -356 10164 -324
rect 10196 -356 10244 -324
rect 10276 -356 10324 -324
rect 10356 -356 10404 -324
rect 10436 -356 10484 -324
rect 10516 -356 10564 -324
rect 10596 -356 10644 -324
rect 10676 -356 10804 -324
rect 10836 -356 10964 -324
rect 10996 -356 11000 -324
rect -720 -360 11000 -356
rect -720 -404 -360 -400
rect -720 -436 -716 -404
rect -684 -436 -556 -404
rect -524 -436 -396 -404
rect -364 -436 -360 -404
rect -720 -440 -360 -436
rect -320 -404 11000 -400
rect -320 -436 -236 -404
rect -204 -436 -156 -404
rect -124 -436 -76 -404
rect -44 -436 4 -404
rect 36 -436 84 -404
rect 116 -436 164 -404
rect 196 -436 244 -404
rect 276 -436 324 -404
rect 356 -436 404 -404
rect 436 -436 484 -404
rect 516 -436 564 -404
rect 596 -436 644 -404
rect 676 -436 724 -404
rect 756 -436 804 -404
rect 836 -436 884 -404
rect 916 -436 964 -404
rect 996 -436 1044 -404
rect 1076 -436 1124 -404
rect 1156 -436 1204 -404
rect 1236 -436 1284 -404
rect 1316 -436 1364 -404
rect 1396 -436 1444 -404
rect 1476 -436 1524 -404
rect 1556 -436 1604 -404
rect 1636 -436 1684 -404
rect 1716 -436 1764 -404
rect 1796 -436 1844 -404
rect 1876 -436 1924 -404
rect 1956 -436 2004 -404
rect 2036 -436 2084 -404
rect 2116 -436 2164 -404
rect 2196 -436 2244 -404
rect 2276 -436 2324 -404
rect 2356 -436 2404 -404
rect 2436 -436 2484 -404
rect 2516 -436 2564 -404
rect 2596 -436 2644 -404
rect 2676 -436 2724 -404
rect 2756 -436 2804 -404
rect 2836 -436 2884 -404
rect 2916 -436 2964 -404
rect 2996 -436 3044 -404
rect 3076 -436 3124 -404
rect 3156 -436 3204 -404
rect 3236 -436 3284 -404
rect 3316 -436 3364 -404
rect 3396 -436 3444 -404
rect 3476 -436 3524 -404
rect 3556 -436 3604 -404
rect 3636 -436 3684 -404
rect 3716 -436 3764 -404
rect 3796 -436 3844 -404
rect 3876 -436 3924 -404
rect 3956 -436 4004 -404
rect 4036 -436 4084 -404
rect 4116 -436 4164 -404
rect 4196 -436 4244 -404
rect 4276 -436 4324 -404
rect 4356 -436 4404 -404
rect 4436 -436 4484 -404
rect 4516 -436 4564 -404
rect 4596 -436 4644 -404
rect 4676 -436 4724 -404
rect 4756 -436 4804 -404
rect 4836 -436 4884 -404
rect 4916 -436 4964 -404
rect 4996 -436 5044 -404
rect 5076 -436 5124 -404
rect 5156 -436 5204 -404
rect 5236 -436 5284 -404
rect 5316 -436 5364 -404
rect 5396 -436 5444 -404
rect 5476 -436 5524 -404
rect 5556 -436 5604 -404
rect 5636 -436 5684 -404
rect 5716 -436 5764 -404
rect 5796 -436 5844 -404
rect 5876 -436 5924 -404
rect 5956 -436 6004 -404
rect 6036 -436 6084 -404
rect 6116 -436 6164 -404
rect 6196 -436 6244 -404
rect 6276 -436 6324 -404
rect 6356 -436 6404 -404
rect 6436 -436 6484 -404
rect 6516 -436 6564 -404
rect 6596 -436 6644 -404
rect 6676 -436 6724 -404
rect 6756 -436 6804 -404
rect 6836 -436 6884 -404
rect 6916 -436 6964 -404
rect 6996 -436 7044 -404
rect 7076 -436 7124 -404
rect 7156 -436 7204 -404
rect 7236 -436 7284 -404
rect 7316 -436 7364 -404
rect 7396 -436 7444 -404
rect 7476 -436 7524 -404
rect 7556 -436 7604 -404
rect 7636 -436 7684 -404
rect 7716 -436 7764 -404
rect 7796 -436 7844 -404
rect 7876 -436 7924 -404
rect 7956 -436 8004 -404
rect 8036 -436 8084 -404
rect 8116 -436 8164 -404
rect 8196 -436 8244 -404
rect 8276 -436 8324 -404
rect 8356 -436 8404 -404
rect 8436 -436 8484 -404
rect 8516 -436 8564 -404
rect 8596 -436 8644 -404
rect 8676 -436 8724 -404
rect 8756 -436 8804 -404
rect 8836 -436 8884 -404
rect 8916 -436 8964 -404
rect 8996 -436 9044 -404
rect 9076 -436 9124 -404
rect 9156 -436 9204 -404
rect 9236 -436 9284 -404
rect 9316 -436 9364 -404
rect 9396 -436 9444 -404
rect 9476 -436 9524 -404
rect 9556 -436 9604 -404
rect 9636 -436 9684 -404
rect 9716 -436 9764 -404
rect 9796 -436 9844 -404
rect 9876 -436 9924 -404
rect 9956 -436 10004 -404
rect 10036 -436 10084 -404
rect 10116 -436 10164 -404
rect 10196 -436 10244 -404
rect 10276 -436 10324 -404
rect 10356 -436 10404 -404
rect 10436 -436 10484 -404
rect 10516 -436 10564 -404
rect 10596 -436 10644 -404
rect 10676 -436 10804 -404
rect 10836 -436 10964 -404
rect 10996 -436 11000 -404
rect -320 -440 11000 -436
rect -720 -484 11000 -480
rect -720 -516 -716 -484
rect -684 -516 -556 -484
rect -524 -516 -396 -484
rect -364 -516 -236 -484
rect -204 -516 -156 -484
rect -124 -516 -76 -484
rect -44 -516 4 -484
rect 36 -516 84 -484
rect 116 -516 164 -484
rect 196 -516 244 -484
rect 276 -516 324 -484
rect 356 -516 404 -484
rect 436 -516 484 -484
rect 516 -516 564 -484
rect 596 -516 644 -484
rect 676 -516 724 -484
rect 756 -516 804 -484
rect 836 -516 884 -484
rect 916 -516 964 -484
rect 996 -516 1044 -484
rect 1076 -516 1124 -484
rect 1156 -516 1204 -484
rect 1236 -516 1284 -484
rect 1316 -516 1364 -484
rect 1396 -516 1444 -484
rect 1476 -516 1524 -484
rect 1556 -516 1604 -484
rect 1636 -516 1684 -484
rect 1716 -516 1764 -484
rect 1796 -516 1844 -484
rect 1876 -516 1924 -484
rect 1956 -516 2004 -484
rect 2036 -516 2084 -484
rect 2116 -516 2164 -484
rect 2196 -516 2244 -484
rect 2276 -516 2324 -484
rect 2356 -516 2404 -484
rect 2436 -516 2484 -484
rect 2516 -516 2564 -484
rect 2596 -516 2644 -484
rect 2676 -516 2724 -484
rect 2756 -516 2804 -484
rect 2836 -516 2884 -484
rect 2916 -516 2964 -484
rect 2996 -516 3044 -484
rect 3076 -516 3124 -484
rect 3156 -516 3204 -484
rect 3236 -516 3284 -484
rect 3316 -516 3364 -484
rect 3396 -516 3444 -484
rect 3476 -516 3524 -484
rect 3556 -516 3604 -484
rect 3636 -516 3684 -484
rect 3716 -516 3764 -484
rect 3796 -516 3844 -484
rect 3876 -516 3924 -484
rect 3956 -516 4004 -484
rect 4036 -516 4084 -484
rect 4116 -516 4164 -484
rect 4196 -516 4244 -484
rect 4276 -516 4324 -484
rect 4356 -516 4404 -484
rect 4436 -516 4484 -484
rect 4516 -516 4564 -484
rect 4596 -516 4644 -484
rect 4676 -516 4724 -484
rect 4756 -516 4804 -484
rect 4836 -516 4884 -484
rect 4916 -516 4964 -484
rect 4996 -516 5044 -484
rect 5076 -516 5124 -484
rect 5156 -516 5204 -484
rect 5236 -516 5284 -484
rect 5316 -516 5364 -484
rect 5396 -516 5444 -484
rect 5476 -516 5524 -484
rect 5556 -516 5604 -484
rect 5636 -516 5684 -484
rect 5716 -516 5764 -484
rect 5796 -516 5844 -484
rect 5876 -516 5924 -484
rect 5956 -516 6004 -484
rect 6036 -516 6084 -484
rect 6116 -516 6164 -484
rect 6196 -516 6244 -484
rect 6276 -516 6324 -484
rect 6356 -516 6404 -484
rect 6436 -516 6484 -484
rect 6516 -516 6564 -484
rect 6596 -516 6644 -484
rect 6676 -516 6724 -484
rect 6756 -516 6804 -484
rect 6836 -516 6884 -484
rect 6916 -516 6964 -484
rect 6996 -516 7044 -484
rect 7076 -516 7124 -484
rect 7156 -516 7204 -484
rect 7236 -516 7284 -484
rect 7316 -516 7364 -484
rect 7396 -516 7444 -484
rect 7476 -516 7524 -484
rect 7556 -516 7604 -484
rect 7636 -516 7684 -484
rect 7716 -516 7764 -484
rect 7796 -516 7844 -484
rect 7876 -516 7924 -484
rect 7956 -516 8004 -484
rect 8036 -516 8084 -484
rect 8116 -516 8164 -484
rect 8196 -516 8244 -484
rect 8276 -516 8324 -484
rect 8356 -516 8404 -484
rect 8436 -516 8484 -484
rect 8516 -516 8564 -484
rect 8596 -516 8644 -484
rect 8676 -516 8724 -484
rect 8756 -516 8804 -484
rect 8836 -516 8884 -484
rect 8916 -516 8964 -484
rect 8996 -516 9044 -484
rect 9076 -516 9124 -484
rect 9156 -516 9204 -484
rect 9236 -516 9284 -484
rect 9316 -516 9364 -484
rect 9396 -516 9444 -484
rect 9476 -516 9524 -484
rect 9556 -516 9604 -484
rect 9636 -516 9684 -484
rect 9716 -516 9764 -484
rect 9796 -516 9844 -484
rect 9876 -516 9924 -484
rect 9956 -516 10004 -484
rect 10036 -516 10084 -484
rect 10116 -516 10164 -484
rect 10196 -516 10244 -484
rect 10276 -516 10324 -484
rect 10356 -516 10404 -484
rect 10436 -516 10484 -484
rect 10516 -516 10564 -484
rect 10596 -516 10644 -484
rect 10676 -516 10804 -484
rect 10836 -516 10964 -484
rect 10996 -516 11000 -484
rect -720 -520 11000 -516
rect -720 -564 -360 -560
rect -720 -596 -716 -564
rect -684 -596 -556 -564
rect -524 -596 -396 -564
rect -364 -596 -360 -564
rect -720 -600 -360 -596
rect -320 -564 11000 -560
rect -320 -596 -236 -564
rect -204 -596 -156 -564
rect -124 -596 -76 -564
rect -44 -596 4 -564
rect 36 -596 84 -564
rect 116 -596 164 -564
rect 196 -596 244 -564
rect 276 -596 324 -564
rect 356 -596 404 -564
rect 436 -596 484 -564
rect 516 -596 564 -564
rect 596 -596 644 -564
rect 676 -596 724 -564
rect 756 -596 804 -564
rect 836 -596 884 -564
rect 916 -596 964 -564
rect 996 -596 1044 -564
rect 1076 -596 1124 -564
rect 1156 -596 1204 -564
rect 1236 -596 1284 -564
rect 1316 -596 1364 -564
rect 1396 -596 1444 -564
rect 1476 -596 1524 -564
rect 1556 -596 1604 -564
rect 1636 -596 1684 -564
rect 1716 -596 1764 -564
rect 1796 -596 1844 -564
rect 1876 -596 1924 -564
rect 1956 -596 2004 -564
rect 2036 -596 2084 -564
rect 2116 -596 2164 -564
rect 2196 -596 2244 -564
rect 2276 -596 2324 -564
rect 2356 -596 2404 -564
rect 2436 -596 2484 -564
rect 2516 -596 2564 -564
rect 2596 -596 2644 -564
rect 2676 -596 2724 -564
rect 2756 -596 2804 -564
rect 2836 -596 2884 -564
rect 2916 -596 2964 -564
rect 2996 -596 3044 -564
rect 3076 -596 3124 -564
rect 3156 -596 3204 -564
rect 3236 -596 3284 -564
rect 3316 -596 3364 -564
rect 3396 -596 3444 -564
rect 3476 -596 3524 -564
rect 3556 -596 3604 -564
rect 3636 -596 3684 -564
rect 3716 -596 3764 -564
rect 3796 -596 3844 -564
rect 3876 -596 3924 -564
rect 3956 -596 4004 -564
rect 4036 -596 4084 -564
rect 4116 -596 4164 -564
rect 4196 -596 4244 -564
rect 4276 -596 4324 -564
rect 4356 -596 4404 -564
rect 4436 -596 4484 -564
rect 4516 -596 4564 -564
rect 4596 -596 4644 -564
rect 4676 -596 4724 -564
rect 4756 -596 4804 -564
rect 4836 -596 4884 -564
rect 4916 -596 4964 -564
rect 4996 -596 5044 -564
rect 5076 -596 5124 -564
rect 5156 -596 5204 -564
rect 5236 -596 5284 -564
rect 5316 -596 5364 -564
rect 5396 -596 5444 -564
rect 5476 -596 5524 -564
rect 5556 -596 5604 -564
rect 5636 -596 5684 -564
rect 5716 -596 5764 -564
rect 5796 -596 5844 -564
rect 5876 -596 5924 -564
rect 5956 -596 6004 -564
rect 6036 -596 6084 -564
rect 6116 -596 6164 -564
rect 6196 -596 6244 -564
rect 6276 -596 6324 -564
rect 6356 -596 6404 -564
rect 6436 -596 6484 -564
rect 6516 -596 6564 -564
rect 6596 -596 6644 -564
rect 6676 -596 6724 -564
rect 6756 -596 6804 -564
rect 6836 -596 6884 -564
rect 6916 -596 6964 -564
rect 6996 -596 7044 -564
rect 7076 -596 7124 -564
rect 7156 -596 7204 -564
rect 7236 -596 7284 -564
rect 7316 -596 7364 -564
rect 7396 -596 7444 -564
rect 7476 -596 7524 -564
rect 7556 -596 7604 -564
rect 7636 -596 7684 -564
rect 7716 -596 7764 -564
rect 7796 -596 7844 -564
rect 7876 -596 7924 -564
rect 7956 -596 8004 -564
rect 8036 -596 8084 -564
rect 8116 -596 8164 -564
rect 8196 -596 8244 -564
rect 8276 -596 8324 -564
rect 8356 -596 8404 -564
rect 8436 -596 8484 -564
rect 8516 -596 8564 -564
rect 8596 -596 8644 -564
rect 8676 -596 8724 -564
rect 8756 -596 8804 -564
rect 8836 -596 8884 -564
rect 8916 -596 8964 -564
rect 8996 -596 9044 -564
rect 9076 -596 9124 -564
rect 9156 -596 9204 -564
rect 9236 -596 9284 -564
rect 9316 -596 9364 -564
rect 9396 -596 9444 -564
rect 9476 -596 9524 -564
rect 9556 -596 9604 -564
rect 9636 -596 9684 -564
rect 9716 -596 9764 -564
rect 9796 -596 9844 -564
rect 9876 -596 9924 -564
rect 9956 -596 10004 -564
rect 10036 -596 10084 -564
rect 10116 -596 10164 -564
rect 10196 -596 10244 -564
rect 10276 -596 10324 -564
rect 10356 -596 10404 -564
rect 10436 -596 10484 -564
rect 10516 -596 10564 -564
rect 10596 -596 10644 -564
rect 10676 -596 10804 -564
rect 10836 -596 10964 -564
rect 10996 -596 11000 -564
rect -320 -600 11000 -596
rect -720 -644 11000 -640
rect -720 -676 -716 -644
rect -684 -676 -556 -644
rect -524 -676 -396 -644
rect -364 -676 -236 -644
rect -204 -676 -156 -644
rect -124 -676 -76 -644
rect -44 -676 4 -644
rect 36 -676 84 -644
rect 116 -676 164 -644
rect 196 -676 244 -644
rect 276 -676 324 -644
rect 356 -676 404 -644
rect 436 -676 484 -644
rect 516 -676 564 -644
rect 596 -676 644 -644
rect 676 -676 724 -644
rect 756 -676 804 -644
rect 836 -676 884 -644
rect 916 -676 964 -644
rect 996 -676 1044 -644
rect 1076 -676 1124 -644
rect 1156 -676 1204 -644
rect 1236 -676 1284 -644
rect 1316 -676 1364 -644
rect 1396 -676 1444 -644
rect 1476 -676 1524 -644
rect 1556 -676 1604 -644
rect 1636 -676 1684 -644
rect 1716 -676 1764 -644
rect 1796 -676 1844 -644
rect 1876 -676 1924 -644
rect 1956 -676 2004 -644
rect 2036 -676 2084 -644
rect 2116 -676 2164 -644
rect 2196 -676 2244 -644
rect 2276 -676 2324 -644
rect 2356 -676 2404 -644
rect 2436 -676 2484 -644
rect 2516 -676 2564 -644
rect 2596 -676 2644 -644
rect 2676 -676 2724 -644
rect 2756 -676 2804 -644
rect 2836 -676 2884 -644
rect 2916 -676 2964 -644
rect 2996 -676 3044 -644
rect 3076 -676 3124 -644
rect 3156 -676 3204 -644
rect 3236 -676 3284 -644
rect 3316 -676 3364 -644
rect 3396 -676 3444 -644
rect 3476 -676 3524 -644
rect 3556 -676 3604 -644
rect 3636 -676 3684 -644
rect 3716 -676 3764 -644
rect 3796 -676 3844 -644
rect 3876 -676 3924 -644
rect 3956 -676 4004 -644
rect 4036 -676 4084 -644
rect 4116 -676 4164 -644
rect 4196 -676 4244 -644
rect 4276 -676 4324 -644
rect 4356 -676 4404 -644
rect 4436 -676 4484 -644
rect 4516 -676 4564 -644
rect 4596 -676 4644 -644
rect 4676 -676 4724 -644
rect 4756 -676 4804 -644
rect 4836 -676 4884 -644
rect 4916 -676 4964 -644
rect 4996 -676 5044 -644
rect 5076 -676 5124 -644
rect 5156 -676 5204 -644
rect 5236 -676 5284 -644
rect 5316 -676 5364 -644
rect 5396 -676 5444 -644
rect 5476 -676 5524 -644
rect 5556 -676 5604 -644
rect 5636 -676 5684 -644
rect 5716 -676 5764 -644
rect 5796 -676 5844 -644
rect 5876 -676 5924 -644
rect 5956 -676 6004 -644
rect 6036 -676 6084 -644
rect 6116 -676 6164 -644
rect 6196 -676 6244 -644
rect 6276 -676 6324 -644
rect 6356 -676 6404 -644
rect 6436 -676 6484 -644
rect 6516 -676 6564 -644
rect 6596 -676 6644 -644
rect 6676 -676 6724 -644
rect 6756 -676 6804 -644
rect 6836 -676 6884 -644
rect 6916 -676 6964 -644
rect 6996 -676 7044 -644
rect 7076 -676 7124 -644
rect 7156 -676 7204 -644
rect 7236 -676 7284 -644
rect 7316 -676 7364 -644
rect 7396 -676 7444 -644
rect 7476 -676 7524 -644
rect 7556 -676 7604 -644
rect 7636 -676 7684 -644
rect 7716 -676 7764 -644
rect 7796 -676 7844 -644
rect 7876 -676 7924 -644
rect 7956 -676 8004 -644
rect 8036 -676 8084 -644
rect 8116 -676 8164 -644
rect 8196 -676 8244 -644
rect 8276 -676 8324 -644
rect 8356 -676 8404 -644
rect 8436 -676 8484 -644
rect 8516 -676 8564 -644
rect 8596 -676 8644 -644
rect 8676 -676 8724 -644
rect 8756 -676 8804 -644
rect 8836 -676 8884 -644
rect 8916 -676 8964 -644
rect 8996 -676 9044 -644
rect 9076 -676 9124 -644
rect 9156 -676 9204 -644
rect 9236 -676 9284 -644
rect 9316 -676 9364 -644
rect 9396 -676 9444 -644
rect 9476 -676 9524 -644
rect 9556 -676 9604 -644
rect 9636 -676 9684 -644
rect 9716 -676 9764 -644
rect 9796 -676 9844 -644
rect 9876 -676 9924 -644
rect 9956 -676 10004 -644
rect 10036 -676 10084 -644
rect 10116 -676 10164 -644
rect 10196 -676 10244 -644
rect 10276 -676 10324 -644
rect 10356 -676 10404 -644
rect 10436 -676 10484 -644
rect 10516 -676 10564 -644
rect 10596 -676 10644 -644
rect 10676 -676 10804 -644
rect 10836 -676 10964 -644
rect 10996 -676 11000 -644
rect -720 -680 11000 -676
rect -720 -724 10600 -720
rect -720 -756 -716 -724
rect -684 -756 -556 -724
rect -524 -756 -396 -724
rect -364 -756 -236 -724
rect -204 -756 -156 -724
rect -124 -756 -76 -724
rect -44 -756 4 -724
rect 36 -756 84 -724
rect 116 -756 164 -724
rect 196 -756 244 -724
rect 276 -756 324 -724
rect 356 -756 404 -724
rect 436 -756 484 -724
rect 516 -756 564 -724
rect 596 -756 644 -724
rect 676 -756 724 -724
rect 756 -756 804 -724
rect 836 -756 884 -724
rect 916 -756 964 -724
rect 996 -756 1044 -724
rect 1076 -756 1124 -724
rect 1156 -756 1204 -724
rect 1236 -756 1284 -724
rect 1316 -756 1364 -724
rect 1396 -756 1444 -724
rect 1476 -756 1524 -724
rect 1556 -756 1604 -724
rect 1636 -756 1684 -724
rect 1716 -756 1764 -724
rect 1796 -756 1844 -724
rect 1876 -756 1924 -724
rect 1956 -756 2004 -724
rect 2036 -756 2084 -724
rect 2116 -756 2164 -724
rect 2196 -756 2244 -724
rect 2276 -756 2324 -724
rect 2356 -756 2404 -724
rect 2436 -756 2484 -724
rect 2516 -756 2564 -724
rect 2596 -756 2644 -724
rect 2676 -756 2724 -724
rect 2756 -756 2804 -724
rect 2836 -756 2884 -724
rect 2916 -756 2964 -724
rect 2996 -756 3044 -724
rect 3076 -756 3124 -724
rect 3156 -756 3204 -724
rect 3236 -756 3284 -724
rect 3316 -756 3364 -724
rect 3396 -756 3444 -724
rect 3476 -756 3524 -724
rect 3556 -756 3604 -724
rect 3636 -756 3684 -724
rect 3716 -756 3764 -724
rect 3796 -756 3844 -724
rect 3876 -756 3924 -724
rect 3956 -756 4004 -724
rect 4036 -756 4084 -724
rect 4116 -756 4164 -724
rect 4196 -756 4244 -724
rect 4276 -756 4324 -724
rect 4356 -756 4404 -724
rect 4436 -756 4484 -724
rect 4516 -756 4564 -724
rect 4596 -756 4644 -724
rect 4676 -756 4724 -724
rect 4756 -756 4804 -724
rect 4836 -756 4884 -724
rect 4916 -756 4964 -724
rect 4996 -756 5044 -724
rect 5076 -756 5124 -724
rect 5156 -756 5204 -724
rect 5236 -756 5284 -724
rect 5316 -756 5364 -724
rect 5396 -756 5444 -724
rect 5476 -756 5524 -724
rect 5556 -756 5604 -724
rect 5636 -756 5684 -724
rect 5716 -756 5764 -724
rect 5796 -756 5844 -724
rect 5876 -756 5924 -724
rect 5956 -756 6004 -724
rect 6036 -756 6084 -724
rect 6116 -756 6164 -724
rect 6196 -756 6244 -724
rect 6276 -756 6324 -724
rect 6356 -756 6404 -724
rect 6436 -756 6484 -724
rect 6516 -756 6564 -724
rect 6596 -756 6644 -724
rect 6676 -756 6724 -724
rect 6756 -756 6804 -724
rect 6836 -756 6884 -724
rect 6916 -756 6964 -724
rect 6996 -756 7044 -724
rect 7076 -756 7124 -724
rect 7156 -756 7204 -724
rect 7236 -756 7284 -724
rect 7316 -756 7364 -724
rect 7396 -756 7444 -724
rect 7476 -756 7524 -724
rect 7556 -756 7604 -724
rect 7636 -756 7684 -724
rect 7716 -756 7764 -724
rect 7796 -756 7844 -724
rect 7876 -756 7924 -724
rect 7956 -756 8004 -724
rect 8036 -756 8084 -724
rect 8116 -756 8164 -724
rect 8196 -756 8244 -724
rect 8276 -756 8324 -724
rect 8356 -756 8404 -724
rect 8436 -756 8484 -724
rect 8516 -756 8564 -724
rect 8596 -756 8644 -724
rect 8676 -756 8724 -724
rect 8756 -756 8804 -724
rect 8836 -756 8884 -724
rect 8916 -756 8964 -724
rect 8996 -756 9044 -724
rect 9076 -756 9124 -724
rect 9156 -756 9204 -724
rect 9236 -756 9284 -724
rect 9316 -756 9364 -724
rect 9396 -756 9444 -724
rect 9476 -756 9524 -724
rect 9556 -756 9604 -724
rect 9636 -756 9684 -724
rect 9716 -756 9764 -724
rect 9796 -756 9844 -724
rect 9876 -756 9924 -724
rect 9956 -756 10004 -724
rect 10036 -756 10084 -724
rect 10116 -756 10164 -724
rect 10196 -756 10244 -724
rect 10276 -756 10324 -724
rect 10356 -756 10404 -724
rect 10436 -756 10484 -724
rect 10516 -756 10564 -724
rect 10596 -756 10600 -724
rect -720 -760 10600 -756
rect 10640 -724 11000 -720
rect 10640 -756 10644 -724
rect 10676 -756 10804 -724
rect 10836 -756 10964 -724
rect 10996 -756 11000 -724
rect 10640 -760 11000 -756
rect -720 -804 11000 -800
rect -720 -836 -716 -804
rect -684 -836 -556 -804
rect -524 -836 -396 -804
rect -364 -836 -236 -804
rect -204 -836 -156 -804
rect -124 -836 -76 -804
rect -44 -836 4 -804
rect 36 -836 84 -804
rect 116 -836 164 -804
rect 196 -836 244 -804
rect 276 -836 324 -804
rect 356 -836 404 -804
rect 436 -836 484 -804
rect 516 -836 564 -804
rect 596 -836 644 -804
rect 676 -836 724 -804
rect 756 -836 804 -804
rect 836 -836 884 -804
rect 916 -836 964 -804
rect 996 -836 1044 -804
rect 1076 -836 1124 -804
rect 1156 -836 1204 -804
rect 1236 -836 1284 -804
rect 1316 -836 1364 -804
rect 1396 -836 1444 -804
rect 1476 -836 1524 -804
rect 1556 -836 1604 -804
rect 1636 -836 1684 -804
rect 1716 -836 1764 -804
rect 1796 -836 1844 -804
rect 1876 -836 1924 -804
rect 1956 -836 2004 -804
rect 2036 -836 2084 -804
rect 2116 -836 2164 -804
rect 2196 -836 2244 -804
rect 2276 -836 2324 -804
rect 2356 -836 2404 -804
rect 2436 -836 2484 -804
rect 2516 -836 2564 -804
rect 2596 -836 2644 -804
rect 2676 -836 2724 -804
rect 2756 -836 2804 -804
rect 2836 -836 2884 -804
rect 2916 -836 2964 -804
rect 2996 -836 3044 -804
rect 3076 -836 3124 -804
rect 3156 -836 3204 -804
rect 3236 -836 3284 -804
rect 3316 -836 3364 -804
rect 3396 -836 3444 -804
rect 3476 -836 3524 -804
rect 3556 -836 3604 -804
rect 3636 -836 3684 -804
rect 3716 -836 3764 -804
rect 3796 -836 3844 -804
rect 3876 -836 3924 -804
rect 3956 -836 4004 -804
rect 4036 -836 4084 -804
rect 4116 -836 4164 -804
rect 4196 -836 4244 -804
rect 4276 -836 4324 -804
rect 4356 -836 4404 -804
rect 4436 -836 4484 -804
rect 4516 -836 4564 -804
rect 4596 -836 4644 -804
rect 4676 -836 4724 -804
rect 4756 -836 4804 -804
rect 4836 -836 4884 -804
rect 4916 -836 4964 -804
rect 4996 -836 5044 -804
rect 5076 -836 5124 -804
rect 5156 -836 5204 -804
rect 5236 -836 5284 -804
rect 5316 -836 5364 -804
rect 5396 -836 5444 -804
rect 5476 -836 5524 -804
rect 5556 -836 5604 -804
rect 5636 -836 5684 -804
rect 5716 -836 5764 -804
rect 5796 -836 5844 -804
rect 5876 -836 5924 -804
rect 5956 -836 6004 -804
rect 6036 -836 6084 -804
rect 6116 -836 6164 -804
rect 6196 -836 6244 -804
rect 6276 -836 6324 -804
rect 6356 -836 6404 -804
rect 6436 -836 6484 -804
rect 6516 -836 6564 -804
rect 6596 -836 6644 -804
rect 6676 -836 6724 -804
rect 6756 -836 6804 -804
rect 6836 -836 6884 -804
rect 6916 -836 6964 -804
rect 6996 -836 7044 -804
rect 7076 -836 7124 -804
rect 7156 -836 7204 -804
rect 7236 -836 7284 -804
rect 7316 -836 7364 -804
rect 7396 -836 7444 -804
rect 7476 -836 7524 -804
rect 7556 -836 7604 -804
rect 7636 -836 7684 -804
rect 7716 -836 7764 -804
rect 7796 -836 7844 -804
rect 7876 -836 7924 -804
rect 7956 -836 8004 -804
rect 8036 -836 8084 -804
rect 8116 -836 8164 -804
rect 8196 -836 8244 -804
rect 8276 -836 8324 -804
rect 8356 -836 8404 -804
rect 8436 -836 8484 -804
rect 8516 -836 8564 -804
rect 8596 -836 8644 -804
rect 8676 -836 8724 -804
rect 8756 -836 8804 -804
rect 8836 -836 8884 -804
rect 8916 -836 8964 -804
rect 8996 -836 9044 -804
rect 9076 -836 9124 -804
rect 9156 -836 9204 -804
rect 9236 -836 9284 -804
rect 9316 -836 9364 -804
rect 9396 -836 9444 -804
rect 9476 -836 9524 -804
rect 9556 -836 9604 -804
rect 9636 -836 9684 -804
rect 9716 -836 9764 -804
rect 9796 -836 9844 -804
rect 9876 -836 9924 -804
rect 9956 -836 10004 -804
rect 10036 -836 10084 -804
rect 10116 -836 10164 -804
rect 10196 -836 10244 -804
rect 10276 -836 10324 -804
rect 10356 -836 10404 -804
rect 10436 -836 10484 -804
rect 10516 -836 10564 -804
rect 10596 -836 10644 -804
rect 10676 -836 10804 -804
rect 10836 -836 10964 -804
rect 10996 -836 11000 -804
rect -720 -840 11000 -836
rect -720 -884 11000 -880
rect -720 -916 -716 -884
rect -684 -916 -556 -884
rect -524 -916 -396 -884
rect -364 -916 -236 -884
rect -204 -916 -156 -884
rect -124 -916 -76 -884
rect -44 -916 4 -884
rect 36 -916 84 -884
rect 116 -916 164 -884
rect 196 -916 244 -884
rect 276 -916 324 -884
rect 356 -916 404 -884
rect 436 -916 484 -884
rect 516 -916 564 -884
rect 596 -916 644 -884
rect 676 -916 724 -884
rect 756 -916 804 -884
rect 836 -916 884 -884
rect 916 -916 964 -884
rect 996 -916 1044 -884
rect 1076 -916 1124 -884
rect 1156 -916 1204 -884
rect 1236 -916 1284 -884
rect 1316 -916 1364 -884
rect 1396 -916 1444 -884
rect 1476 -916 1524 -884
rect 1556 -916 1604 -884
rect 1636 -916 1684 -884
rect 1716 -916 1764 -884
rect 1796 -916 1844 -884
rect 1876 -916 1924 -884
rect 1956 -916 2004 -884
rect 2036 -916 2084 -884
rect 2116 -916 2164 -884
rect 2196 -916 2244 -884
rect 2276 -916 2324 -884
rect 2356 -916 2404 -884
rect 2436 -916 2484 -884
rect 2516 -916 2564 -884
rect 2596 -916 2644 -884
rect 2676 -916 2724 -884
rect 2756 -916 2804 -884
rect 2836 -916 2884 -884
rect 2916 -916 2964 -884
rect 2996 -916 3044 -884
rect 3076 -916 3124 -884
rect 3156 -916 3204 -884
rect 3236 -916 3284 -884
rect 3316 -916 3364 -884
rect 3396 -916 3444 -884
rect 3476 -916 3524 -884
rect 3556 -916 3604 -884
rect 3636 -916 3684 -884
rect 3716 -916 3764 -884
rect 3796 -916 3844 -884
rect 3876 -916 3924 -884
rect 3956 -916 4004 -884
rect 4036 -916 4084 -884
rect 4116 -916 4164 -884
rect 4196 -916 4244 -884
rect 4276 -916 4324 -884
rect 4356 -916 4404 -884
rect 4436 -916 4484 -884
rect 4516 -916 4564 -884
rect 4596 -916 4644 -884
rect 4676 -916 4724 -884
rect 4756 -916 4804 -884
rect 4836 -916 4884 -884
rect 4916 -916 4964 -884
rect 4996 -916 5044 -884
rect 5076 -916 5124 -884
rect 5156 -916 5204 -884
rect 5236 -916 5284 -884
rect 5316 -916 5364 -884
rect 5396 -916 5444 -884
rect 5476 -916 5524 -884
rect 5556 -916 5604 -884
rect 5636 -916 5684 -884
rect 5716 -916 5764 -884
rect 5796 -916 5844 -884
rect 5876 -916 5924 -884
rect 5956 -916 6004 -884
rect 6036 -916 6084 -884
rect 6116 -916 6164 -884
rect 6196 -916 6244 -884
rect 6276 -916 6324 -884
rect 6356 -916 6404 -884
rect 6436 -916 6484 -884
rect 6516 -916 6564 -884
rect 6596 -916 6644 -884
rect 6676 -916 6724 -884
rect 6756 -916 6804 -884
rect 6836 -916 6884 -884
rect 6916 -916 6964 -884
rect 6996 -916 7044 -884
rect 7076 -916 7124 -884
rect 7156 -916 7204 -884
rect 7236 -916 7284 -884
rect 7316 -916 7364 -884
rect 7396 -916 7444 -884
rect 7476 -916 7524 -884
rect 7556 -916 7604 -884
rect 7636 -916 7684 -884
rect 7716 -916 7764 -884
rect 7796 -916 7844 -884
rect 7876 -916 7924 -884
rect 7956 -916 8004 -884
rect 8036 -916 8084 -884
rect 8116 -916 8164 -884
rect 8196 -916 8244 -884
rect 8276 -916 8324 -884
rect 8356 -916 8404 -884
rect 8436 -916 8484 -884
rect 8516 -916 8564 -884
rect 8596 -916 8644 -884
rect 8676 -916 8724 -884
rect 8756 -916 8804 -884
rect 8836 -916 8884 -884
rect 8916 -916 8964 -884
rect 8996 -916 9044 -884
rect 9076 -916 9124 -884
rect 9156 -916 9204 -884
rect 9236 -916 9284 -884
rect 9316 -916 9364 -884
rect 9396 -916 9444 -884
rect 9476 -916 9524 -884
rect 9556 -916 9604 -884
rect 9636 -916 9684 -884
rect 9716 -916 9764 -884
rect 9796 -916 9844 -884
rect 9876 -916 9924 -884
rect 9956 -916 10004 -884
rect 10036 -916 10084 -884
rect 10116 -916 10164 -884
rect 10196 -916 10244 -884
rect 10276 -916 10324 -884
rect 10356 -916 10404 -884
rect 10436 -916 10484 -884
rect 10516 -916 10564 -884
rect 10596 -916 10644 -884
rect 10676 -916 10804 -884
rect 10836 -916 10964 -884
rect 10996 -916 11000 -884
rect -720 -920 11000 -916
rect -720 -964 10600 -960
rect -720 -996 -716 -964
rect -684 -996 -556 -964
rect -524 -996 -396 -964
rect -364 -996 -236 -964
rect -204 -996 -156 -964
rect -124 -996 -76 -964
rect -44 -996 4 -964
rect 36 -996 84 -964
rect 116 -996 164 -964
rect 196 -996 244 -964
rect 276 -996 324 -964
rect 356 -996 404 -964
rect 436 -996 484 -964
rect 516 -996 564 -964
rect 596 -996 644 -964
rect 676 -996 724 -964
rect 756 -996 804 -964
rect 836 -996 884 -964
rect 916 -996 964 -964
rect 996 -996 1044 -964
rect 1076 -996 1124 -964
rect 1156 -996 1204 -964
rect 1236 -996 1284 -964
rect 1316 -996 1364 -964
rect 1396 -996 1444 -964
rect 1476 -996 1524 -964
rect 1556 -996 1604 -964
rect 1636 -996 1684 -964
rect 1716 -996 1764 -964
rect 1796 -996 1844 -964
rect 1876 -996 1924 -964
rect 1956 -996 2004 -964
rect 2036 -996 2084 -964
rect 2116 -996 2164 -964
rect 2196 -996 2244 -964
rect 2276 -996 2324 -964
rect 2356 -996 2404 -964
rect 2436 -996 2484 -964
rect 2516 -996 2564 -964
rect 2596 -996 2644 -964
rect 2676 -996 2724 -964
rect 2756 -996 2804 -964
rect 2836 -996 2884 -964
rect 2916 -996 2964 -964
rect 2996 -996 3044 -964
rect 3076 -996 3124 -964
rect 3156 -996 3204 -964
rect 3236 -996 3284 -964
rect 3316 -996 3364 -964
rect 3396 -996 3444 -964
rect 3476 -996 3524 -964
rect 3556 -996 3604 -964
rect 3636 -996 3684 -964
rect 3716 -996 3764 -964
rect 3796 -996 3844 -964
rect 3876 -996 3924 -964
rect 3956 -996 4004 -964
rect 4036 -996 4084 -964
rect 4116 -996 4164 -964
rect 4196 -996 4244 -964
rect 4276 -996 4324 -964
rect 4356 -996 4404 -964
rect 4436 -996 4484 -964
rect 4516 -996 4564 -964
rect 4596 -996 4644 -964
rect 4676 -996 4724 -964
rect 4756 -996 4804 -964
rect 4836 -996 4884 -964
rect 4916 -996 4964 -964
rect 4996 -996 5044 -964
rect 5076 -996 5124 -964
rect 5156 -996 5204 -964
rect 5236 -996 5284 -964
rect 5316 -996 5364 -964
rect 5396 -996 5444 -964
rect 5476 -996 5524 -964
rect 5556 -996 5604 -964
rect 5636 -996 5684 -964
rect 5716 -996 5764 -964
rect 5796 -996 5844 -964
rect 5876 -996 5924 -964
rect 5956 -996 6004 -964
rect 6036 -996 6084 -964
rect 6116 -996 6164 -964
rect 6196 -996 6244 -964
rect 6276 -996 6324 -964
rect 6356 -996 6404 -964
rect 6436 -996 6484 -964
rect 6516 -996 6564 -964
rect 6596 -996 6644 -964
rect 6676 -996 6724 -964
rect 6756 -996 6804 -964
rect 6836 -996 6884 -964
rect 6916 -996 6964 -964
rect 6996 -996 7044 -964
rect 7076 -996 7124 -964
rect 7156 -996 7204 -964
rect 7236 -996 7284 -964
rect 7316 -996 7364 -964
rect 7396 -996 7444 -964
rect 7476 -996 7524 -964
rect 7556 -996 7604 -964
rect 7636 -996 7684 -964
rect 7716 -996 7764 -964
rect 7796 -996 7844 -964
rect 7876 -996 7924 -964
rect 7956 -996 8004 -964
rect 8036 -996 8084 -964
rect 8116 -996 8164 -964
rect 8196 -996 8244 -964
rect 8276 -996 8324 -964
rect 8356 -996 8404 -964
rect 8436 -996 8484 -964
rect 8516 -996 8564 -964
rect 8596 -996 8644 -964
rect 8676 -996 8724 -964
rect 8756 -996 8804 -964
rect 8836 -996 8884 -964
rect 8916 -996 8964 -964
rect 8996 -996 9044 -964
rect 9076 -996 9124 -964
rect 9156 -996 9204 -964
rect 9236 -996 9284 -964
rect 9316 -996 9364 -964
rect 9396 -996 9444 -964
rect 9476 -996 9524 -964
rect 9556 -996 9604 -964
rect 9636 -996 9684 -964
rect 9716 -996 9764 -964
rect 9796 -996 9844 -964
rect 9876 -996 9924 -964
rect 9956 -996 10004 -964
rect 10036 -996 10084 -964
rect 10116 -996 10164 -964
rect 10196 -996 10244 -964
rect 10276 -996 10324 -964
rect 10356 -996 10404 -964
rect 10436 -996 10484 -964
rect 10516 -996 10564 -964
rect 10596 -996 10600 -964
rect -720 -1000 10600 -996
rect 10640 -964 11000 -960
rect 10640 -996 10644 -964
rect 10676 -996 10804 -964
rect 10836 -996 10964 -964
rect 10996 -996 11000 -964
rect 10640 -1000 11000 -996
rect -720 -1044 10600 -1040
rect -720 -1076 -716 -1044
rect -684 -1076 -556 -1044
rect -524 -1076 -396 -1044
rect -364 -1076 -236 -1044
rect -204 -1076 -156 -1044
rect -124 -1076 -76 -1044
rect -44 -1076 4 -1044
rect 36 -1076 84 -1044
rect 116 -1076 164 -1044
rect 196 -1076 244 -1044
rect 276 -1076 324 -1044
rect 356 -1076 404 -1044
rect 436 -1076 484 -1044
rect 516 -1076 564 -1044
rect 596 -1076 644 -1044
rect 676 -1076 724 -1044
rect 756 -1076 804 -1044
rect 836 -1076 884 -1044
rect 916 -1076 964 -1044
rect 996 -1076 1044 -1044
rect 1076 -1076 1124 -1044
rect 1156 -1076 1204 -1044
rect 1236 -1076 1284 -1044
rect 1316 -1076 1364 -1044
rect 1396 -1076 1444 -1044
rect 1476 -1076 1524 -1044
rect 1556 -1076 1604 -1044
rect 1636 -1076 1684 -1044
rect 1716 -1076 1764 -1044
rect 1796 -1076 1844 -1044
rect 1876 -1076 1924 -1044
rect 1956 -1076 2004 -1044
rect 2036 -1076 2084 -1044
rect 2116 -1076 2164 -1044
rect 2196 -1076 2244 -1044
rect 2276 -1076 2324 -1044
rect 2356 -1076 2404 -1044
rect 2436 -1076 2484 -1044
rect 2516 -1076 2564 -1044
rect 2596 -1076 2644 -1044
rect 2676 -1076 2724 -1044
rect 2756 -1076 2804 -1044
rect 2836 -1076 2884 -1044
rect 2916 -1076 2964 -1044
rect 2996 -1076 3044 -1044
rect 3076 -1076 3124 -1044
rect 3156 -1076 3204 -1044
rect 3236 -1076 3284 -1044
rect 3316 -1076 3364 -1044
rect 3396 -1076 3444 -1044
rect 3476 -1076 3524 -1044
rect 3556 -1076 3604 -1044
rect 3636 -1076 3684 -1044
rect 3716 -1076 3764 -1044
rect 3796 -1076 3844 -1044
rect 3876 -1076 3924 -1044
rect 3956 -1076 4004 -1044
rect 4036 -1076 4084 -1044
rect 4116 -1076 4164 -1044
rect 4196 -1076 4244 -1044
rect 4276 -1076 4324 -1044
rect 4356 -1076 4404 -1044
rect 4436 -1076 4484 -1044
rect 4516 -1076 4564 -1044
rect 4596 -1076 4644 -1044
rect 4676 -1076 4724 -1044
rect 4756 -1076 4804 -1044
rect 4836 -1076 4884 -1044
rect 4916 -1076 4964 -1044
rect 4996 -1076 5044 -1044
rect 5076 -1076 5124 -1044
rect 5156 -1076 5204 -1044
rect 5236 -1076 5284 -1044
rect 5316 -1076 5364 -1044
rect 5396 -1076 5444 -1044
rect 5476 -1076 5524 -1044
rect 5556 -1076 5604 -1044
rect 5636 -1076 5684 -1044
rect 5716 -1076 5764 -1044
rect 5796 -1076 5844 -1044
rect 5876 -1076 5924 -1044
rect 5956 -1076 6004 -1044
rect 6036 -1076 6084 -1044
rect 6116 -1076 6164 -1044
rect 6196 -1076 6244 -1044
rect 6276 -1076 6324 -1044
rect 6356 -1076 6404 -1044
rect 6436 -1076 6484 -1044
rect 6516 -1076 6564 -1044
rect 6596 -1076 6644 -1044
rect 6676 -1076 6724 -1044
rect 6756 -1076 6804 -1044
rect 6836 -1076 6884 -1044
rect 6916 -1076 6964 -1044
rect 6996 -1076 7044 -1044
rect 7076 -1076 7124 -1044
rect 7156 -1076 7204 -1044
rect 7236 -1076 7284 -1044
rect 7316 -1076 7364 -1044
rect 7396 -1076 7444 -1044
rect 7476 -1076 7524 -1044
rect 7556 -1076 7604 -1044
rect 7636 -1076 7684 -1044
rect 7716 -1076 7764 -1044
rect 7796 -1076 7844 -1044
rect 7876 -1076 7924 -1044
rect 7956 -1076 8004 -1044
rect 8036 -1076 8084 -1044
rect 8116 -1076 8164 -1044
rect 8196 -1076 8244 -1044
rect 8276 -1076 8324 -1044
rect 8356 -1076 8404 -1044
rect 8436 -1076 8484 -1044
rect 8516 -1076 8564 -1044
rect 8596 -1076 8644 -1044
rect 8676 -1076 8724 -1044
rect 8756 -1076 8804 -1044
rect 8836 -1076 8884 -1044
rect 8916 -1076 8964 -1044
rect 8996 -1076 9044 -1044
rect 9076 -1076 9124 -1044
rect 9156 -1076 9204 -1044
rect 9236 -1076 9284 -1044
rect 9316 -1076 9364 -1044
rect 9396 -1076 9444 -1044
rect 9476 -1076 9524 -1044
rect 9556 -1076 9604 -1044
rect 9636 -1076 9684 -1044
rect 9716 -1076 9764 -1044
rect 9796 -1076 9844 -1044
rect 9876 -1076 9924 -1044
rect 9956 -1076 10004 -1044
rect 10036 -1076 10084 -1044
rect 10116 -1076 10164 -1044
rect 10196 -1076 10244 -1044
rect 10276 -1076 10324 -1044
rect 10356 -1076 10404 -1044
rect 10436 -1076 10484 -1044
rect 10516 -1076 10564 -1044
rect 10596 -1076 10600 -1044
rect -720 -1080 10600 -1076
rect 10640 -1044 11000 -1040
rect 10640 -1076 10644 -1044
rect 10676 -1076 10804 -1044
rect 10836 -1076 10964 -1044
rect 10996 -1076 11000 -1044
rect 10640 -1080 11000 -1076
rect -720 -1124 11000 -1120
rect -720 -1156 -716 -1124
rect -684 -1156 -556 -1124
rect -524 -1156 -396 -1124
rect -364 -1156 -236 -1124
rect -204 -1156 -156 -1124
rect -124 -1156 -76 -1124
rect -44 -1156 4 -1124
rect 36 -1156 84 -1124
rect 116 -1156 164 -1124
rect 196 -1156 244 -1124
rect 276 -1156 324 -1124
rect 356 -1156 404 -1124
rect 436 -1156 484 -1124
rect 516 -1156 564 -1124
rect 596 -1156 644 -1124
rect 676 -1156 724 -1124
rect 756 -1156 804 -1124
rect 836 -1156 884 -1124
rect 916 -1156 964 -1124
rect 996 -1156 1044 -1124
rect 1076 -1156 1124 -1124
rect 1156 -1156 1204 -1124
rect 1236 -1156 1284 -1124
rect 1316 -1156 1364 -1124
rect 1396 -1156 1444 -1124
rect 1476 -1156 1524 -1124
rect 1556 -1156 1604 -1124
rect 1636 -1156 1684 -1124
rect 1716 -1156 1764 -1124
rect 1796 -1156 1844 -1124
rect 1876 -1156 1924 -1124
rect 1956 -1156 2004 -1124
rect 2036 -1156 2084 -1124
rect 2116 -1156 2164 -1124
rect 2196 -1156 2244 -1124
rect 2276 -1156 2324 -1124
rect 2356 -1156 2404 -1124
rect 2436 -1156 2484 -1124
rect 2516 -1156 2564 -1124
rect 2596 -1156 2644 -1124
rect 2676 -1156 2724 -1124
rect 2756 -1156 2804 -1124
rect 2836 -1156 2884 -1124
rect 2916 -1156 2964 -1124
rect 2996 -1156 3044 -1124
rect 3076 -1156 3124 -1124
rect 3156 -1156 3204 -1124
rect 3236 -1156 3284 -1124
rect 3316 -1156 3364 -1124
rect 3396 -1156 3444 -1124
rect 3476 -1156 3524 -1124
rect 3556 -1156 3604 -1124
rect 3636 -1156 3684 -1124
rect 3716 -1156 3764 -1124
rect 3796 -1156 3844 -1124
rect 3876 -1156 3924 -1124
rect 3956 -1156 4004 -1124
rect 4036 -1156 4084 -1124
rect 4116 -1156 4164 -1124
rect 4196 -1156 4244 -1124
rect 4276 -1156 4324 -1124
rect 4356 -1156 4404 -1124
rect 4436 -1156 4484 -1124
rect 4516 -1156 4564 -1124
rect 4596 -1156 4644 -1124
rect 4676 -1156 4724 -1124
rect 4756 -1156 4804 -1124
rect 4836 -1156 4884 -1124
rect 4916 -1156 4964 -1124
rect 4996 -1156 5044 -1124
rect 5076 -1156 5124 -1124
rect 5156 -1156 5204 -1124
rect 5236 -1156 5284 -1124
rect 5316 -1156 5364 -1124
rect 5396 -1156 5444 -1124
rect 5476 -1156 5524 -1124
rect 5556 -1156 5604 -1124
rect 5636 -1156 5684 -1124
rect 5716 -1156 5764 -1124
rect 5796 -1156 5844 -1124
rect 5876 -1156 5924 -1124
rect 5956 -1156 6004 -1124
rect 6036 -1156 6084 -1124
rect 6116 -1156 6164 -1124
rect 6196 -1156 6244 -1124
rect 6276 -1156 6324 -1124
rect 6356 -1156 6404 -1124
rect 6436 -1156 6484 -1124
rect 6516 -1156 6564 -1124
rect 6596 -1156 6644 -1124
rect 6676 -1156 6724 -1124
rect 6756 -1156 6804 -1124
rect 6836 -1156 6884 -1124
rect 6916 -1156 6964 -1124
rect 6996 -1156 7044 -1124
rect 7076 -1156 7124 -1124
rect 7156 -1156 7204 -1124
rect 7236 -1156 7284 -1124
rect 7316 -1156 7364 -1124
rect 7396 -1156 7444 -1124
rect 7476 -1156 7524 -1124
rect 7556 -1156 7604 -1124
rect 7636 -1156 7684 -1124
rect 7716 -1156 7764 -1124
rect 7796 -1156 7844 -1124
rect 7876 -1156 7924 -1124
rect 7956 -1156 8004 -1124
rect 8036 -1156 8084 -1124
rect 8116 -1156 8164 -1124
rect 8196 -1156 8244 -1124
rect 8276 -1156 8324 -1124
rect 8356 -1156 8404 -1124
rect 8436 -1156 8484 -1124
rect 8516 -1156 8564 -1124
rect 8596 -1156 8644 -1124
rect 8676 -1156 8724 -1124
rect 8756 -1156 8804 -1124
rect 8836 -1156 8884 -1124
rect 8916 -1156 8964 -1124
rect 8996 -1156 9044 -1124
rect 9076 -1156 9124 -1124
rect 9156 -1156 9204 -1124
rect 9236 -1156 9284 -1124
rect 9316 -1156 9364 -1124
rect 9396 -1156 9444 -1124
rect 9476 -1156 9524 -1124
rect 9556 -1156 9604 -1124
rect 9636 -1156 9684 -1124
rect 9716 -1156 9764 -1124
rect 9796 -1156 9844 -1124
rect 9876 -1156 9924 -1124
rect 9956 -1156 10004 -1124
rect 10036 -1156 10084 -1124
rect 10116 -1156 10164 -1124
rect 10196 -1156 10244 -1124
rect 10276 -1156 10324 -1124
rect 10356 -1156 10404 -1124
rect 10436 -1156 10484 -1124
rect 10516 -1156 10564 -1124
rect 10596 -1156 10644 -1124
rect 10676 -1156 10804 -1124
rect 10836 -1156 10964 -1124
rect 10996 -1156 11000 -1124
rect -720 -1160 11000 -1156
rect -720 -1204 11000 -1200
rect -720 -1236 -716 -1204
rect -684 -1236 -556 -1204
rect -524 -1236 -396 -1204
rect -364 -1236 -236 -1204
rect -204 -1236 -156 -1204
rect -124 -1236 -76 -1204
rect -44 -1236 4 -1204
rect 36 -1236 84 -1204
rect 116 -1236 164 -1204
rect 196 -1236 244 -1204
rect 276 -1236 324 -1204
rect 356 -1236 404 -1204
rect 436 -1236 484 -1204
rect 516 -1236 564 -1204
rect 596 -1236 644 -1204
rect 676 -1236 724 -1204
rect 756 -1236 804 -1204
rect 836 -1236 884 -1204
rect 916 -1236 964 -1204
rect 996 -1236 1044 -1204
rect 1076 -1236 1124 -1204
rect 1156 -1236 1204 -1204
rect 1236 -1236 1284 -1204
rect 1316 -1236 1364 -1204
rect 1396 -1236 1444 -1204
rect 1476 -1236 1524 -1204
rect 1556 -1236 1604 -1204
rect 1636 -1236 1684 -1204
rect 1716 -1236 1764 -1204
rect 1796 -1236 1844 -1204
rect 1876 -1236 1924 -1204
rect 1956 -1236 2004 -1204
rect 2036 -1236 2084 -1204
rect 2116 -1236 2164 -1204
rect 2196 -1236 2244 -1204
rect 2276 -1236 2324 -1204
rect 2356 -1236 2404 -1204
rect 2436 -1236 2484 -1204
rect 2516 -1236 2564 -1204
rect 2596 -1236 2644 -1204
rect 2676 -1236 2724 -1204
rect 2756 -1236 2804 -1204
rect 2836 -1236 2884 -1204
rect 2916 -1236 2964 -1204
rect 2996 -1236 3044 -1204
rect 3076 -1236 3124 -1204
rect 3156 -1236 3204 -1204
rect 3236 -1236 3284 -1204
rect 3316 -1236 3364 -1204
rect 3396 -1236 3444 -1204
rect 3476 -1236 3524 -1204
rect 3556 -1236 3604 -1204
rect 3636 -1236 3684 -1204
rect 3716 -1236 3764 -1204
rect 3796 -1236 3844 -1204
rect 3876 -1236 3924 -1204
rect 3956 -1236 4004 -1204
rect 4036 -1236 4084 -1204
rect 4116 -1236 4164 -1204
rect 4196 -1236 4244 -1204
rect 4276 -1236 4324 -1204
rect 4356 -1236 4404 -1204
rect 4436 -1236 4484 -1204
rect 4516 -1236 4564 -1204
rect 4596 -1236 4644 -1204
rect 4676 -1236 4724 -1204
rect 4756 -1236 4804 -1204
rect 4836 -1236 4884 -1204
rect 4916 -1236 4964 -1204
rect 4996 -1236 5044 -1204
rect 5076 -1236 5124 -1204
rect 5156 -1236 5204 -1204
rect 5236 -1236 5284 -1204
rect 5316 -1236 5364 -1204
rect 5396 -1236 5444 -1204
rect 5476 -1236 5524 -1204
rect 5556 -1236 5604 -1204
rect 5636 -1236 5684 -1204
rect 5716 -1236 5764 -1204
rect 5796 -1236 5844 -1204
rect 5876 -1236 5924 -1204
rect 5956 -1236 6004 -1204
rect 6036 -1236 6084 -1204
rect 6116 -1236 6164 -1204
rect 6196 -1236 6244 -1204
rect 6276 -1236 6324 -1204
rect 6356 -1236 6404 -1204
rect 6436 -1236 6484 -1204
rect 6516 -1236 6564 -1204
rect 6596 -1236 6644 -1204
rect 6676 -1236 6724 -1204
rect 6756 -1236 6804 -1204
rect 6836 -1236 6884 -1204
rect 6916 -1236 6964 -1204
rect 6996 -1236 7044 -1204
rect 7076 -1236 7124 -1204
rect 7156 -1236 7204 -1204
rect 7236 -1236 7284 -1204
rect 7316 -1236 7364 -1204
rect 7396 -1236 7444 -1204
rect 7476 -1236 7524 -1204
rect 7556 -1236 7604 -1204
rect 7636 -1236 7684 -1204
rect 7716 -1236 7764 -1204
rect 7796 -1236 7844 -1204
rect 7876 -1236 7924 -1204
rect 7956 -1236 8004 -1204
rect 8036 -1236 8084 -1204
rect 8116 -1236 8164 -1204
rect 8196 -1236 8244 -1204
rect 8276 -1236 8324 -1204
rect 8356 -1236 8404 -1204
rect 8436 -1236 8484 -1204
rect 8516 -1236 8564 -1204
rect 8596 -1236 8644 -1204
rect 8676 -1236 8724 -1204
rect 8756 -1236 8804 -1204
rect 8836 -1236 8884 -1204
rect 8916 -1236 8964 -1204
rect 8996 -1236 9044 -1204
rect 9076 -1236 9124 -1204
rect 9156 -1236 9204 -1204
rect 9236 -1236 9284 -1204
rect 9316 -1236 9364 -1204
rect 9396 -1236 9444 -1204
rect 9476 -1236 9524 -1204
rect 9556 -1236 9604 -1204
rect 9636 -1236 9684 -1204
rect 9716 -1236 9764 -1204
rect 9796 -1236 9844 -1204
rect 9876 -1236 9924 -1204
rect 9956 -1236 10004 -1204
rect 10036 -1236 10084 -1204
rect 10116 -1236 10164 -1204
rect 10196 -1236 10244 -1204
rect 10276 -1236 10324 -1204
rect 10356 -1236 10404 -1204
rect 10436 -1236 10484 -1204
rect 10516 -1236 10564 -1204
rect 10596 -1236 10644 -1204
rect 10676 -1236 10804 -1204
rect 10836 -1236 10964 -1204
rect 10996 -1236 11000 -1204
rect -720 -1240 11000 -1236
rect -720 -1284 11000 -1280
rect -720 -1316 -716 -1284
rect -684 -1316 -556 -1284
rect -524 -1316 -396 -1284
rect -364 -1316 -236 -1284
rect -204 -1316 -156 -1284
rect -124 -1316 -76 -1284
rect -44 -1316 4 -1284
rect 36 -1316 84 -1284
rect 116 -1316 164 -1284
rect 196 -1316 244 -1284
rect 276 -1316 324 -1284
rect 356 -1316 404 -1284
rect 436 -1316 484 -1284
rect 516 -1316 564 -1284
rect 596 -1316 644 -1284
rect 676 -1316 724 -1284
rect 756 -1316 804 -1284
rect 836 -1316 884 -1284
rect 916 -1316 964 -1284
rect 996 -1316 1044 -1284
rect 1076 -1316 1124 -1284
rect 1156 -1316 1204 -1284
rect 1236 -1316 1284 -1284
rect 1316 -1316 1364 -1284
rect 1396 -1316 1444 -1284
rect 1476 -1316 1524 -1284
rect 1556 -1316 1604 -1284
rect 1636 -1316 1684 -1284
rect 1716 -1316 1764 -1284
rect 1796 -1316 1844 -1284
rect 1876 -1316 1924 -1284
rect 1956 -1316 2004 -1284
rect 2036 -1316 2084 -1284
rect 2116 -1316 2164 -1284
rect 2196 -1316 2244 -1284
rect 2276 -1316 2324 -1284
rect 2356 -1316 2404 -1284
rect 2436 -1316 2484 -1284
rect 2516 -1316 2564 -1284
rect 2596 -1316 2644 -1284
rect 2676 -1316 2724 -1284
rect 2756 -1316 2804 -1284
rect 2836 -1316 2884 -1284
rect 2916 -1316 2964 -1284
rect 2996 -1316 3044 -1284
rect 3076 -1316 3124 -1284
rect 3156 -1316 3204 -1284
rect 3236 -1316 3284 -1284
rect 3316 -1316 3364 -1284
rect 3396 -1316 3444 -1284
rect 3476 -1316 3524 -1284
rect 3556 -1316 3604 -1284
rect 3636 -1316 3684 -1284
rect 3716 -1316 3764 -1284
rect 3796 -1316 3844 -1284
rect 3876 -1316 3924 -1284
rect 3956 -1316 4004 -1284
rect 4036 -1316 4084 -1284
rect 4116 -1316 4164 -1284
rect 4196 -1316 4244 -1284
rect 4276 -1316 4324 -1284
rect 4356 -1316 4404 -1284
rect 4436 -1316 4484 -1284
rect 4516 -1316 4564 -1284
rect 4596 -1316 4644 -1284
rect 4676 -1316 4724 -1284
rect 4756 -1316 4804 -1284
rect 4836 -1316 4884 -1284
rect 4916 -1316 4964 -1284
rect 4996 -1316 5044 -1284
rect 5076 -1316 5124 -1284
rect 5156 -1316 5204 -1284
rect 5236 -1316 5284 -1284
rect 5316 -1316 5364 -1284
rect 5396 -1316 5444 -1284
rect 5476 -1316 5524 -1284
rect 5556 -1316 5604 -1284
rect 5636 -1316 5684 -1284
rect 5716 -1316 5764 -1284
rect 5796 -1316 5844 -1284
rect 5876 -1316 5924 -1284
rect 5956 -1316 6004 -1284
rect 6036 -1316 6084 -1284
rect 6116 -1316 6164 -1284
rect 6196 -1316 6244 -1284
rect 6276 -1316 6324 -1284
rect 6356 -1316 6404 -1284
rect 6436 -1316 6484 -1284
rect 6516 -1316 6564 -1284
rect 6596 -1316 6644 -1284
rect 6676 -1316 6724 -1284
rect 6756 -1316 6804 -1284
rect 6836 -1316 6884 -1284
rect 6916 -1316 6964 -1284
rect 6996 -1316 7044 -1284
rect 7076 -1316 7124 -1284
rect 7156 -1316 7204 -1284
rect 7236 -1316 7284 -1284
rect 7316 -1316 7364 -1284
rect 7396 -1316 7444 -1284
rect 7476 -1316 7524 -1284
rect 7556 -1316 7604 -1284
rect 7636 -1316 7684 -1284
rect 7716 -1316 7764 -1284
rect 7796 -1316 7844 -1284
rect 7876 -1316 7924 -1284
rect 7956 -1316 8004 -1284
rect 8036 -1316 8084 -1284
rect 8116 -1316 8164 -1284
rect 8196 -1316 8244 -1284
rect 8276 -1316 8324 -1284
rect 8356 -1316 8404 -1284
rect 8436 -1316 8484 -1284
rect 8516 -1316 8564 -1284
rect 8596 -1316 8644 -1284
rect 8676 -1316 8724 -1284
rect 8756 -1316 8804 -1284
rect 8836 -1316 8884 -1284
rect 8916 -1316 8964 -1284
rect 8996 -1316 9044 -1284
rect 9076 -1316 9124 -1284
rect 9156 -1316 9204 -1284
rect 9236 -1316 9284 -1284
rect 9316 -1316 9364 -1284
rect 9396 -1316 9444 -1284
rect 9476 -1316 9524 -1284
rect 9556 -1316 9604 -1284
rect 9636 -1316 9684 -1284
rect 9716 -1316 9764 -1284
rect 9796 -1316 9844 -1284
rect 9876 -1316 9924 -1284
rect 9956 -1316 10004 -1284
rect 10036 -1316 10084 -1284
rect 10116 -1316 10164 -1284
rect 10196 -1316 10244 -1284
rect 10276 -1316 10324 -1284
rect 10356 -1316 10404 -1284
rect 10436 -1316 10484 -1284
rect 10516 -1316 10564 -1284
rect 10596 -1316 10644 -1284
rect 10676 -1316 10804 -1284
rect 10836 -1316 10964 -1284
rect 10996 -1316 11000 -1284
rect -720 -1320 11000 -1316
rect -720 -1364 11000 -1360
rect -720 -1396 -716 -1364
rect -684 -1396 -556 -1364
rect -524 -1396 -396 -1364
rect -364 -1396 -236 -1364
rect -204 -1396 -156 -1364
rect -124 -1396 -76 -1364
rect -44 -1396 4 -1364
rect 36 -1396 84 -1364
rect 116 -1396 164 -1364
rect 196 -1396 244 -1364
rect 276 -1396 324 -1364
rect 356 -1396 404 -1364
rect 436 -1396 484 -1364
rect 516 -1396 564 -1364
rect 596 -1396 644 -1364
rect 676 -1396 724 -1364
rect 756 -1396 804 -1364
rect 836 -1396 884 -1364
rect 916 -1396 964 -1364
rect 996 -1396 1044 -1364
rect 1076 -1396 1124 -1364
rect 1156 -1396 1204 -1364
rect 1236 -1396 1284 -1364
rect 1316 -1396 1364 -1364
rect 1396 -1396 1444 -1364
rect 1476 -1396 1524 -1364
rect 1556 -1396 1604 -1364
rect 1636 -1396 1684 -1364
rect 1716 -1396 1764 -1364
rect 1796 -1396 1844 -1364
rect 1876 -1396 1924 -1364
rect 1956 -1396 2004 -1364
rect 2036 -1396 2084 -1364
rect 2116 -1396 2164 -1364
rect 2196 -1396 2244 -1364
rect 2276 -1396 2324 -1364
rect 2356 -1396 2404 -1364
rect 2436 -1396 2484 -1364
rect 2516 -1396 2564 -1364
rect 2596 -1396 2644 -1364
rect 2676 -1396 2724 -1364
rect 2756 -1396 2804 -1364
rect 2836 -1396 2884 -1364
rect 2916 -1396 2964 -1364
rect 2996 -1396 3044 -1364
rect 3076 -1396 3124 -1364
rect 3156 -1396 3204 -1364
rect 3236 -1396 3284 -1364
rect 3316 -1396 3364 -1364
rect 3396 -1396 3444 -1364
rect 3476 -1396 3524 -1364
rect 3556 -1396 3604 -1364
rect 3636 -1396 3684 -1364
rect 3716 -1396 3764 -1364
rect 3796 -1396 3844 -1364
rect 3876 -1396 3924 -1364
rect 3956 -1396 4004 -1364
rect 4036 -1396 4084 -1364
rect 4116 -1396 4164 -1364
rect 4196 -1396 4244 -1364
rect 4276 -1396 4324 -1364
rect 4356 -1396 4404 -1364
rect 4436 -1396 4484 -1364
rect 4516 -1396 4564 -1364
rect 4596 -1396 4644 -1364
rect 4676 -1396 4724 -1364
rect 4756 -1396 4804 -1364
rect 4836 -1396 4884 -1364
rect 4916 -1396 4964 -1364
rect 4996 -1396 5044 -1364
rect 5076 -1396 5124 -1364
rect 5156 -1396 5204 -1364
rect 5236 -1396 5284 -1364
rect 5316 -1396 5364 -1364
rect 5396 -1396 5444 -1364
rect 5476 -1396 5524 -1364
rect 5556 -1396 5604 -1364
rect 5636 -1396 5684 -1364
rect 5716 -1396 5764 -1364
rect 5796 -1396 5844 -1364
rect 5876 -1396 5924 -1364
rect 5956 -1396 6004 -1364
rect 6036 -1396 6084 -1364
rect 6116 -1396 6164 -1364
rect 6196 -1396 6244 -1364
rect 6276 -1396 6324 -1364
rect 6356 -1396 6404 -1364
rect 6436 -1396 6484 -1364
rect 6516 -1396 6564 -1364
rect 6596 -1396 6644 -1364
rect 6676 -1396 6724 -1364
rect 6756 -1396 6804 -1364
rect 6836 -1396 6884 -1364
rect 6916 -1396 6964 -1364
rect 6996 -1396 7044 -1364
rect 7076 -1396 7124 -1364
rect 7156 -1396 7204 -1364
rect 7236 -1396 7284 -1364
rect 7316 -1396 7364 -1364
rect 7396 -1396 7444 -1364
rect 7476 -1396 7524 -1364
rect 7556 -1396 7604 -1364
rect 7636 -1396 7684 -1364
rect 7716 -1396 7764 -1364
rect 7796 -1396 7844 -1364
rect 7876 -1396 7924 -1364
rect 7956 -1396 8004 -1364
rect 8036 -1396 8084 -1364
rect 8116 -1396 8164 -1364
rect 8196 -1396 8244 -1364
rect 8276 -1396 8324 -1364
rect 8356 -1396 8404 -1364
rect 8436 -1396 8484 -1364
rect 8516 -1396 8564 -1364
rect 8596 -1396 8644 -1364
rect 8676 -1396 8724 -1364
rect 8756 -1396 8804 -1364
rect 8836 -1396 8884 -1364
rect 8916 -1396 8964 -1364
rect 8996 -1396 9044 -1364
rect 9076 -1396 9124 -1364
rect 9156 -1396 9204 -1364
rect 9236 -1396 9284 -1364
rect 9316 -1396 9364 -1364
rect 9396 -1396 9444 -1364
rect 9476 -1396 9524 -1364
rect 9556 -1396 9604 -1364
rect 9636 -1396 9684 -1364
rect 9716 -1396 9764 -1364
rect 9796 -1396 9844 -1364
rect 9876 -1396 9924 -1364
rect 9956 -1396 10004 -1364
rect 10036 -1396 10084 -1364
rect 10116 -1396 10164 -1364
rect 10196 -1396 10244 -1364
rect 10276 -1396 10324 -1364
rect 10356 -1396 10404 -1364
rect 10436 -1396 10484 -1364
rect 10516 -1396 10564 -1364
rect 10596 -1396 10644 -1364
rect 10676 -1396 10804 -1364
rect 10836 -1396 10964 -1364
rect 10996 -1396 11000 -1364
rect -720 -1400 11000 -1396
rect -720 -1444 11000 -1440
rect -720 -1476 -716 -1444
rect -684 -1476 -556 -1444
rect -524 -1476 -396 -1444
rect -364 -1476 -236 -1444
rect -204 -1476 -156 -1444
rect -124 -1476 -76 -1444
rect -44 -1476 4 -1444
rect 36 -1476 84 -1444
rect 116 -1476 164 -1444
rect 196 -1476 244 -1444
rect 276 -1476 324 -1444
rect 356 -1476 404 -1444
rect 436 -1476 484 -1444
rect 516 -1476 564 -1444
rect 596 -1476 644 -1444
rect 676 -1476 724 -1444
rect 756 -1476 804 -1444
rect 836 -1476 884 -1444
rect 916 -1476 964 -1444
rect 996 -1476 1044 -1444
rect 1076 -1476 1124 -1444
rect 1156 -1476 1204 -1444
rect 1236 -1476 1284 -1444
rect 1316 -1476 1364 -1444
rect 1396 -1476 1444 -1444
rect 1476 -1476 1524 -1444
rect 1556 -1476 1604 -1444
rect 1636 -1476 1684 -1444
rect 1716 -1476 1764 -1444
rect 1796 -1476 1844 -1444
rect 1876 -1476 1924 -1444
rect 1956 -1476 2004 -1444
rect 2036 -1476 2084 -1444
rect 2116 -1476 2164 -1444
rect 2196 -1476 2244 -1444
rect 2276 -1476 2324 -1444
rect 2356 -1476 2404 -1444
rect 2436 -1476 2484 -1444
rect 2516 -1476 2564 -1444
rect 2596 -1476 2644 -1444
rect 2676 -1476 2724 -1444
rect 2756 -1476 2804 -1444
rect 2836 -1476 2884 -1444
rect 2916 -1476 2964 -1444
rect 2996 -1476 3044 -1444
rect 3076 -1476 3124 -1444
rect 3156 -1476 3204 -1444
rect 3236 -1476 3284 -1444
rect 3316 -1476 3364 -1444
rect 3396 -1476 3444 -1444
rect 3476 -1476 3524 -1444
rect 3556 -1476 3604 -1444
rect 3636 -1476 3684 -1444
rect 3716 -1476 3764 -1444
rect 3796 -1476 3844 -1444
rect 3876 -1476 3924 -1444
rect 3956 -1476 4004 -1444
rect 4036 -1476 4084 -1444
rect 4116 -1476 4164 -1444
rect 4196 -1476 4244 -1444
rect 4276 -1476 4324 -1444
rect 4356 -1476 4404 -1444
rect 4436 -1476 4484 -1444
rect 4516 -1476 4564 -1444
rect 4596 -1476 4644 -1444
rect 4676 -1476 4724 -1444
rect 4756 -1476 4804 -1444
rect 4836 -1476 4884 -1444
rect 4916 -1476 4964 -1444
rect 4996 -1476 5044 -1444
rect 5076 -1476 5124 -1444
rect 5156 -1476 5204 -1444
rect 5236 -1476 5284 -1444
rect 5316 -1476 5364 -1444
rect 5396 -1476 5444 -1444
rect 5476 -1476 5524 -1444
rect 5556 -1476 5604 -1444
rect 5636 -1476 5684 -1444
rect 5716 -1476 5764 -1444
rect 5796 -1476 5844 -1444
rect 5876 -1476 5924 -1444
rect 5956 -1476 6004 -1444
rect 6036 -1476 6084 -1444
rect 6116 -1476 6164 -1444
rect 6196 -1476 6244 -1444
rect 6276 -1476 6324 -1444
rect 6356 -1476 6404 -1444
rect 6436 -1476 6484 -1444
rect 6516 -1476 6564 -1444
rect 6596 -1476 6644 -1444
rect 6676 -1476 6724 -1444
rect 6756 -1476 6804 -1444
rect 6836 -1476 6884 -1444
rect 6916 -1476 6964 -1444
rect 6996 -1476 7044 -1444
rect 7076 -1476 7124 -1444
rect 7156 -1476 7204 -1444
rect 7236 -1476 7284 -1444
rect 7316 -1476 7364 -1444
rect 7396 -1476 7444 -1444
rect 7476 -1476 7524 -1444
rect 7556 -1476 7604 -1444
rect 7636 -1476 7684 -1444
rect 7716 -1476 7764 -1444
rect 7796 -1476 7844 -1444
rect 7876 -1476 7924 -1444
rect 7956 -1476 8004 -1444
rect 8036 -1476 8084 -1444
rect 8116 -1476 8164 -1444
rect 8196 -1476 8244 -1444
rect 8276 -1476 8324 -1444
rect 8356 -1476 8404 -1444
rect 8436 -1476 8484 -1444
rect 8516 -1476 8564 -1444
rect 8596 -1476 8644 -1444
rect 8676 -1476 8724 -1444
rect 8756 -1476 8804 -1444
rect 8836 -1476 8884 -1444
rect 8916 -1476 8964 -1444
rect 8996 -1476 9044 -1444
rect 9076 -1476 9124 -1444
rect 9156 -1476 9204 -1444
rect 9236 -1476 9284 -1444
rect 9316 -1476 9364 -1444
rect 9396 -1476 9444 -1444
rect 9476 -1476 9524 -1444
rect 9556 -1476 9604 -1444
rect 9636 -1476 9684 -1444
rect 9716 -1476 9764 -1444
rect 9796 -1476 9844 -1444
rect 9876 -1476 9924 -1444
rect 9956 -1476 10004 -1444
rect 10036 -1476 10084 -1444
rect 10116 -1476 10164 -1444
rect 10196 -1476 10244 -1444
rect 10276 -1476 10324 -1444
rect 10356 -1476 10404 -1444
rect 10436 -1476 10484 -1444
rect 10516 -1476 10564 -1444
rect 10596 -1476 10644 -1444
rect 10676 -1476 10804 -1444
rect 10836 -1476 10964 -1444
rect 10996 -1476 11000 -1444
rect -720 -1480 11000 -1476
rect -720 -1524 11000 -1520
rect -720 -1556 -716 -1524
rect -684 -1556 -556 -1524
rect -524 -1556 -396 -1524
rect -364 -1556 -236 -1524
rect -204 -1556 -156 -1524
rect -124 -1556 -76 -1524
rect -44 -1556 4 -1524
rect 36 -1556 84 -1524
rect 116 -1556 164 -1524
rect 196 -1556 244 -1524
rect 276 -1556 324 -1524
rect 356 -1556 404 -1524
rect 436 -1556 484 -1524
rect 516 -1556 564 -1524
rect 596 -1556 644 -1524
rect 676 -1556 724 -1524
rect 756 -1556 804 -1524
rect 836 -1556 884 -1524
rect 916 -1556 964 -1524
rect 996 -1556 1044 -1524
rect 1076 -1556 1124 -1524
rect 1156 -1556 1204 -1524
rect 1236 -1556 1284 -1524
rect 1316 -1556 1364 -1524
rect 1396 -1556 1444 -1524
rect 1476 -1556 1524 -1524
rect 1556 -1556 1604 -1524
rect 1636 -1556 1684 -1524
rect 1716 -1556 1764 -1524
rect 1796 -1556 1844 -1524
rect 1876 -1556 1924 -1524
rect 1956 -1556 2004 -1524
rect 2036 -1556 2084 -1524
rect 2116 -1556 2164 -1524
rect 2196 -1556 2244 -1524
rect 2276 -1556 2324 -1524
rect 2356 -1556 2404 -1524
rect 2436 -1556 2484 -1524
rect 2516 -1556 2564 -1524
rect 2596 -1556 2644 -1524
rect 2676 -1556 2724 -1524
rect 2756 -1556 2804 -1524
rect 2836 -1556 2884 -1524
rect 2916 -1556 2964 -1524
rect 2996 -1556 3044 -1524
rect 3076 -1556 3124 -1524
rect 3156 -1556 3204 -1524
rect 3236 -1556 3284 -1524
rect 3316 -1556 3364 -1524
rect 3396 -1556 3444 -1524
rect 3476 -1556 3524 -1524
rect 3556 -1556 3604 -1524
rect 3636 -1556 3684 -1524
rect 3716 -1556 3764 -1524
rect 3796 -1556 3844 -1524
rect 3876 -1556 3924 -1524
rect 3956 -1556 4004 -1524
rect 4036 -1556 4084 -1524
rect 4116 -1556 4164 -1524
rect 4196 -1556 4244 -1524
rect 4276 -1556 4324 -1524
rect 4356 -1556 4404 -1524
rect 4436 -1556 4484 -1524
rect 4516 -1556 4564 -1524
rect 4596 -1556 4644 -1524
rect 4676 -1556 4724 -1524
rect 4756 -1556 4804 -1524
rect 4836 -1556 4884 -1524
rect 4916 -1556 4964 -1524
rect 4996 -1556 5044 -1524
rect 5076 -1556 5124 -1524
rect 5156 -1556 5204 -1524
rect 5236 -1556 5284 -1524
rect 5316 -1556 5364 -1524
rect 5396 -1556 5444 -1524
rect 5476 -1556 5524 -1524
rect 5556 -1556 5604 -1524
rect 5636 -1556 5684 -1524
rect 5716 -1556 5764 -1524
rect 5796 -1556 5844 -1524
rect 5876 -1556 5924 -1524
rect 5956 -1556 6004 -1524
rect 6036 -1556 6084 -1524
rect 6116 -1556 6164 -1524
rect 6196 -1556 6244 -1524
rect 6276 -1556 6324 -1524
rect 6356 -1556 6404 -1524
rect 6436 -1556 6484 -1524
rect 6516 -1556 6564 -1524
rect 6596 -1556 6644 -1524
rect 6676 -1556 6724 -1524
rect 6756 -1556 6804 -1524
rect 6836 -1556 6884 -1524
rect 6916 -1556 6964 -1524
rect 6996 -1556 7044 -1524
rect 7076 -1556 7124 -1524
rect 7156 -1556 7204 -1524
rect 7236 -1556 7284 -1524
rect 7316 -1556 7364 -1524
rect 7396 -1556 7444 -1524
rect 7476 -1556 7524 -1524
rect 7556 -1556 7604 -1524
rect 7636 -1556 7684 -1524
rect 7716 -1556 7764 -1524
rect 7796 -1556 7844 -1524
rect 7876 -1556 7924 -1524
rect 7956 -1556 8004 -1524
rect 8036 -1556 8084 -1524
rect 8116 -1556 8164 -1524
rect 8196 -1556 8244 -1524
rect 8276 -1556 8324 -1524
rect 8356 -1556 8404 -1524
rect 8436 -1556 8484 -1524
rect 8516 -1556 8564 -1524
rect 8596 -1556 8644 -1524
rect 8676 -1556 8724 -1524
rect 8756 -1556 8804 -1524
rect 8836 -1556 8884 -1524
rect 8916 -1556 8964 -1524
rect 8996 -1556 9044 -1524
rect 9076 -1556 9124 -1524
rect 9156 -1556 9204 -1524
rect 9236 -1556 9284 -1524
rect 9316 -1556 9364 -1524
rect 9396 -1556 9444 -1524
rect 9476 -1556 9524 -1524
rect 9556 -1556 9604 -1524
rect 9636 -1556 9684 -1524
rect 9716 -1556 9764 -1524
rect 9796 -1556 9844 -1524
rect 9876 -1556 9924 -1524
rect 9956 -1556 10004 -1524
rect 10036 -1556 10084 -1524
rect 10116 -1556 10164 -1524
rect 10196 -1556 10244 -1524
rect 10276 -1556 10324 -1524
rect 10356 -1556 10404 -1524
rect 10436 -1556 10484 -1524
rect 10516 -1556 10564 -1524
rect 10596 -1556 10644 -1524
rect 10676 -1556 10804 -1524
rect 10836 -1556 10964 -1524
rect 10996 -1556 11000 -1524
rect -720 -1560 11000 -1556
rect -720 -1604 10600 -1600
rect -720 -1636 -716 -1604
rect -684 -1636 -556 -1604
rect -524 -1636 -396 -1604
rect -364 -1636 -236 -1604
rect -204 -1636 -156 -1604
rect -124 -1636 -76 -1604
rect -44 -1636 4 -1604
rect 36 -1636 84 -1604
rect 116 -1636 164 -1604
rect 196 -1636 244 -1604
rect 276 -1636 324 -1604
rect 356 -1636 404 -1604
rect 436 -1636 484 -1604
rect 516 -1636 564 -1604
rect 596 -1636 644 -1604
rect 676 -1636 724 -1604
rect 756 -1636 804 -1604
rect 836 -1636 884 -1604
rect 916 -1636 964 -1604
rect 996 -1636 1044 -1604
rect 1076 -1636 1124 -1604
rect 1156 -1636 1204 -1604
rect 1236 -1636 1284 -1604
rect 1316 -1636 1364 -1604
rect 1396 -1636 1444 -1604
rect 1476 -1636 1524 -1604
rect 1556 -1636 1604 -1604
rect 1636 -1636 1684 -1604
rect 1716 -1636 1764 -1604
rect 1796 -1636 1844 -1604
rect 1876 -1636 1924 -1604
rect 1956 -1636 2004 -1604
rect 2036 -1636 2084 -1604
rect 2116 -1636 2164 -1604
rect 2196 -1636 2244 -1604
rect 2276 -1636 2324 -1604
rect 2356 -1636 2404 -1604
rect 2436 -1636 2484 -1604
rect 2516 -1636 2564 -1604
rect 2596 -1636 2644 -1604
rect 2676 -1636 2724 -1604
rect 2756 -1636 2804 -1604
rect 2836 -1636 2884 -1604
rect 2916 -1636 2964 -1604
rect 2996 -1636 3044 -1604
rect 3076 -1636 3124 -1604
rect 3156 -1636 3204 -1604
rect 3236 -1636 3284 -1604
rect 3316 -1636 3364 -1604
rect 3396 -1636 3444 -1604
rect 3476 -1636 3524 -1604
rect 3556 -1636 3604 -1604
rect 3636 -1636 3684 -1604
rect 3716 -1636 3764 -1604
rect 3796 -1636 3844 -1604
rect 3876 -1636 3924 -1604
rect 3956 -1636 4004 -1604
rect 4036 -1636 4084 -1604
rect 4116 -1636 4164 -1604
rect 4196 -1636 4244 -1604
rect 4276 -1636 4324 -1604
rect 4356 -1636 4404 -1604
rect 4436 -1636 4484 -1604
rect 4516 -1636 4564 -1604
rect 4596 -1636 4644 -1604
rect 4676 -1636 4724 -1604
rect 4756 -1636 4804 -1604
rect 4836 -1636 4884 -1604
rect 4916 -1636 4964 -1604
rect 4996 -1636 5044 -1604
rect 5076 -1636 5124 -1604
rect 5156 -1636 5204 -1604
rect 5236 -1636 5284 -1604
rect 5316 -1636 5364 -1604
rect 5396 -1636 5444 -1604
rect 5476 -1636 5524 -1604
rect 5556 -1636 5604 -1604
rect 5636 -1636 5684 -1604
rect 5716 -1636 5764 -1604
rect 5796 -1636 5844 -1604
rect 5876 -1636 5924 -1604
rect 5956 -1636 6004 -1604
rect 6036 -1636 6084 -1604
rect 6116 -1636 6164 -1604
rect 6196 -1636 6244 -1604
rect 6276 -1636 6324 -1604
rect 6356 -1636 6404 -1604
rect 6436 -1636 6484 -1604
rect 6516 -1636 6564 -1604
rect 6596 -1636 6644 -1604
rect 6676 -1636 6724 -1604
rect 6756 -1636 6804 -1604
rect 6836 -1636 6884 -1604
rect 6916 -1636 6964 -1604
rect 6996 -1636 7044 -1604
rect 7076 -1636 7124 -1604
rect 7156 -1636 7204 -1604
rect 7236 -1636 7284 -1604
rect 7316 -1636 7364 -1604
rect 7396 -1636 7444 -1604
rect 7476 -1636 7524 -1604
rect 7556 -1636 7604 -1604
rect 7636 -1636 7684 -1604
rect 7716 -1636 7764 -1604
rect 7796 -1636 7844 -1604
rect 7876 -1636 7924 -1604
rect 7956 -1636 8004 -1604
rect 8036 -1636 8084 -1604
rect 8116 -1636 8164 -1604
rect 8196 -1636 8244 -1604
rect 8276 -1636 8324 -1604
rect 8356 -1636 8404 -1604
rect 8436 -1636 8484 -1604
rect 8516 -1636 8564 -1604
rect 8596 -1636 8644 -1604
rect 8676 -1636 8724 -1604
rect 8756 -1636 8804 -1604
rect 8836 -1636 8884 -1604
rect 8916 -1636 8964 -1604
rect 8996 -1636 9044 -1604
rect 9076 -1636 9124 -1604
rect 9156 -1636 9204 -1604
rect 9236 -1636 9284 -1604
rect 9316 -1636 9364 -1604
rect 9396 -1636 9444 -1604
rect 9476 -1636 9524 -1604
rect 9556 -1636 9604 -1604
rect 9636 -1636 9684 -1604
rect 9716 -1636 9764 -1604
rect 9796 -1636 9844 -1604
rect 9876 -1636 9924 -1604
rect 9956 -1636 10004 -1604
rect 10036 -1636 10084 -1604
rect 10116 -1636 10164 -1604
rect 10196 -1636 10244 -1604
rect 10276 -1636 10324 -1604
rect 10356 -1636 10404 -1604
rect 10436 -1636 10484 -1604
rect 10516 -1636 10564 -1604
rect 10596 -1636 10600 -1604
rect -720 -1640 10600 -1636
rect 10640 -1604 11000 -1600
rect 10640 -1636 10644 -1604
rect 10676 -1636 10804 -1604
rect 10836 -1636 10964 -1604
rect 10996 -1636 11000 -1604
rect 10640 -1640 11000 -1636
rect -720 -1684 10600 -1680
rect -720 -1716 -716 -1684
rect -684 -1716 -556 -1684
rect -524 -1716 -396 -1684
rect -364 -1716 -236 -1684
rect -204 -1716 -156 -1684
rect -124 -1716 -76 -1684
rect -44 -1716 4 -1684
rect 36 -1716 84 -1684
rect 116 -1716 164 -1684
rect 196 -1716 244 -1684
rect 276 -1716 324 -1684
rect 356 -1716 404 -1684
rect 436 -1716 484 -1684
rect 516 -1716 564 -1684
rect 596 -1716 644 -1684
rect 676 -1716 724 -1684
rect 756 -1716 804 -1684
rect 836 -1716 884 -1684
rect 916 -1716 964 -1684
rect 996 -1716 1044 -1684
rect 1076 -1716 1124 -1684
rect 1156 -1716 1204 -1684
rect 1236 -1716 1284 -1684
rect 1316 -1716 1364 -1684
rect 1396 -1716 1444 -1684
rect 1476 -1716 1524 -1684
rect 1556 -1716 1604 -1684
rect 1636 -1716 1684 -1684
rect 1716 -1716 1764 -1684
rect 1796 -1716 1844 -1684
rect 1876 -1716 1924 -1684
rect 1956 -1716 2004 -1684
rect 2036 -1716 2084 -1684
rect 2116 -1716 2164 -1684
rect 2196 -1716 2244 -1684
rect 2276 -1716 2324 -1684
rect 2356 -1716 2404 -1684
rect 2436 -1716 2484 -1684
rect 2516 -1716 2564 -1684
rect 2596 -1716 2644 -1684
rect 2676 -1716 2724 -1684
rect 2756 -1716 2804 -1684
rect 2836 -1716 2884 -1684
rect 2916 -1716 2964 -1684
rect 2996 -1716 3044 -1684
rect 3076 -1716 3124 -1684
rect 3156 -1716 3204 -1684
rect 3236 -1716 3284 -1684
rect 3316 -1716 3364 -1684
rect 3396 -1716 3444 -1684
rect 3476 -1716 3524 -1684
rect 3556 -1716 3604 -1684
rect 3636 -1716 3684 -1684
rect 3716 -1716 3764 -1684
rect 3796 -1716 3844 -1684
rect 3876 -1716 3924 -1684
rect 3956 -1716 4004 -1684
rect 4036 -1716 4084 -1684
rect 4116 -1716 4164 -1684
rect 4196 -1716 4244 -1684
rect 4276 -1716 4324 -1684
rect 4356 -1716 4404 -1684
rect 4436 -1716 4484 -1684
rect 4516 -1716 4564 -1684
rect 4596 -1716 4644 -1684
rect 4676 -1716 4724 -1684
rect 4756 -1716 4804 -1684
rect 4836 -1716 4884 -1684
rect 4916 -1716 4964 -1684
rect 4996 -1716 5044 -1684
rect 5076 -1716 5124 -1684
rect 5156 -1716 5204 -1684
rect 5236 -1716 5284 -1684
rect 5316 -1716 5364 -1684
rect 5396 -1716 5444 -1684
rect 5476 -1716 5524 -1684
rect 5556 -1716 5604 -1684
rect 5636 -1716 5684 -1684
rect 5716 -1716 5764 -1684
rect 5796 -1716 5844 -1684
rect 5876 -1716 5924 -1684
rect 5956 -1716 6004 -1684
rect 6036 -1716 6084 -1684
rect 6116 -1716 6164 -1684
rect 6196 -1716 6244 -1684
rect 6276 -1716 6324 -1684
rect 6356 -1716 6404 -1684
rect 6436 -1716 6484 -1684
rect 6516 -1716 6564 -1684
rect 6596 -1716 6644 -1684
rect 6676 -1716 6724 -1684
rect 6756 -1716 6804 -1684
rect 6836 -1716 6884 -1684
rect 6916 -1716 6964 -1684
rect 6996 -1716 7044 -1684
rect 7076 -1716 7124 -1684
rect 7156 -1716 7204 -1684
rect 7236 -1716 7284 -1684
rect 7316 -1716 7364 -1684
rect 7396 -1716 7444 -1684
rect 7476 -1716 7524 -1684
rect 7556 -1716 7604 -1684
rect 7636 -1716 7684 -1684
rect 7716 -1716 7764 -1684
rect 7796 -1716 7844 -1684
rect 7876 -1716 7924 -1684
rect 7956 -1716 8004 -1684
rect 8036 -1716 8084 -1684
rect 8116 -1716 8164 -1684
rect 8196 -1716 8244 -1684
rect 8276 -1716 8324 -1684
rect 8356 -1716 8404 -1684
rect 8436 -1716 8484 -1684
rect 8516 -1716 8564 -1684
rect 8596 -1716 8644 -1684
rect 8676 -1716 8724 -1684
rect 8756 -1716 8804 -1684
rect 8836 -1716 8884 -1684
rect 8916 -1716 8964 -1684
rect 8996 -1716 9044 -1684
rect 9076 -1716 9124 -1684
rect 9156 -1716 9204 -1684
rect 9236 -1716 9284 -1684
rect 9316 -1716 9364 -1684
rect 9396 -1716 9444 -1684
rect 9476 -1716 9524 -1684
rect 9556 -1716 9604 -1684
rect 9636 -1716 9684 -1684
rect 9716 -1716 9764 -1684
rect 9796 -1716 9844 -1684
rect 9876 -1716 9924 -1684
rect 9956 -1716 10004 -1684
rect 10036 -1716 10084 -1684
rect 10116 -1716 10164 -1684
rect 10196 -1716 10244 -1684
rect 10276 -1716 10324 -1684
rect 10356 -1716 10404 -1684
rect 10436 -1716 10484 -1684
rect 10516 -1716 10564 -1684
rect 10596 -1716 10600 -1684
rect -720 -1720 10600 -1716
rect 10640 -1684 11000 -1680
rect 10640 -1716 10644 -1684
rect 10676 -1716 10804 -1684
rect 10836 -1716 10964 -1684
rect 10996 -1716 11000 -1684
rect 10640 -1720 11000 -1716
rect -720 -1764 11000 -1760
rect -720 -1796 -716 -1764
rect -684 -1796 -556 -1764
rect -524 -1796 -396 -1764
rect -364 -1796 -236 -1764
rect -204 -1796 -156 -1764
rect -124 -1796 -76 -1764
rect -44 -1796 4 -1764
rect 36 -1796 84 -1764
rect 116 -1796 164 -1764
rect 196 -1796 244 -1764
rect 276 -1796 324 -1764
rect 356 -1796 404 -1764
rect 436 -1796 484 -1764
rect 516 -1796 564 -1764
rect 596 -1796 644 -1764
rect 676 -1796 724 -1764
rect 756 -1796 804 -1764
rect 836 -1796 884 -1764
rect 916 -1796 964 -1764
rect 996 -1796 1044 -1764
rect 1076 -1796 1124 -1764
rect 1156 -1796 1204 -1764
rect 1236 -1796 1284 -1764
rect 1316 -1796 1364 -1764
rect 1396 -1796 1444 -1764
rect 1476 -1796 1524 -1764
rect 1556 -1796 1604 -1764
rect 1636 -1796 1684 -1764
rect 1716 -1796 1764 -1764
rect 1796 -1796 1844 -1764
rect 1876 -1796 1924 -1764
rect 1956 -1796 2004 -1764
rect 2036 -1796 2084 -1764
rect 2116 -1796 2164 -1764
rect 2196 -1796 2244 -1764
rect 2276 -1796 2324 -1764
rect 2356 -1796 2404 -1764
rect 2436 -1796 2484 -1764
rect 2516 -1796 2564 -1764
rect 2596 -1796 2644 -1764
rect 2676 -1796 2724 -1764
rect 2756 -1796 2804 -1764
rect 2836 -1796 2884 -1764
rect 2916 -1796 2964 -1764
rect 2996 -1796 3044 -1764
rect 3076 -1796 3124 -1764
rect 3156 -1796 3204 -1764
rect 3236 -1796 3284 -1764
rect 3316 -1796 3364 -1764
rect 3396 -1796 3444 -1764
rect 3476 -1796 3524 -1764
rect 3556 -1796 3604 -1764
rect 3636 -1796 3684 -1764
rect 3716 -1796 3764 -1764
rect 3796 -1796 3844 -1764
rect 3876 -1796 3924 -1764
rect 3956 -1796 4004 -1764
rect 4036 -1796 4084 -1764
rect 4116 -1796 4164 -1764
rect 4196 -1796 4244 -1764
rect 4276 -1796 4324 -1764
rect 4356 -1796 4404 -1764
rect 4436 -1796 4484 -1764
rect 4516 -1796 4564 -1764
rect 4596 -1796 4644 -1764
rect 4676 -1796 4724 -1764
rect 4756 -1796 4804 -1764
rect 4836 -1796 4884 -1764
rect 4916 -1796 4964 -1764
rect 4996 -1796 5044 -1764
rect 5076 -1796 5124 -1764
rect 5156 -1796 5204 -1764
rect 5236 -1796 5284 -1764
rect 5316 -1796 5364 -1764
rect 5396 -1796 5444 -1764
rect 5476 -1796 5524 -1764
rect 5556 -1796 5604 -1764
rect 5636 -1796 5684 -1764
rect 5716 -1796 5764 -1764
rect 5796 -1796 5844 -1764
rect 5876 -1796 5924 -1764
rect 5956 -1796 6004 -1764
rect 6036 -1796 6084 -1764
rect 6116 -1796 6164 -1764
rect 6196 -1796 6244 -1764
rect 6276 -1796 6324 -1764
rect 6356 -1796 6404 -1764
rect 6436 -1796 6484 -1764
rect 6516 -1796 6564 -1764
rect 6596 -1796 6644 -1764
rect 6676 -1796 6724 -1764
rect 6756 -1796 6804 -1764
rect 6836 -1796 6884 -1764
rect 6916 -1796 6964 -1764
rect 6996 -1796 7044 -1764
rect 7076 -1796 7124 -1764
rect 7156 -1796 7204 -1764
rect 7236 -1796 7284 -1764
rect 7316 -1796 7364 -1764
rect 7396 -1796 7444 -1764
rect 7476 -1796 7524 -1764
rect 7556 -1796 7604 -1764
rect 7636 -1796 7684 -1764
rect 7716 -1796 7764 -1764
rect 7796 -1796 7844 -1764
rect 7876 -1796 7924 -1764
rect 7956 -1796 8004 -1764
rect 8036 -1796 8084 -1764
rect 8116 -1796 8164 -1764
rect 8196 -1796 8244 -1764
rect 8276 -1796 8324 -1764
rect 8356 -1796 8404 -1764
rect 8436 -1796 8484 -1764
rect 8516 -1796 8564 -1764
rect 8596 -1796 8644 -1764
rect 8676 -1796 8724 -1764
rect 8756 -1796 8804 -1764
rect 8836 -1796 8884 -1764
rect 8916 -1796 8964 -1764
rect 8996 -1796 9044 -1764
rect 9076 -1796 9124 -1764
rect 9156 -1796 9204 -1764
rect 9236 -1796 9284 -1764
rect 9316 -1796 9364 -1764
rect 9396 -1796 9444 -1764
rect 9476 -1796 9524 -1764
rect 9556 -1796 9604 -1764
rect 9636 -1796 9684 -1764
rect 9716 -1796 9764 -1764
rect 9796 -1796 9844 -1764
rect 9876 -1796 9924 -1764
rect 9956 -1796 10004 -1764
rect 10036 -1796 10084 -1764
rect 10116 -1796 10164 -1764
rect 10196 -1796 10244 -1764
rect 10276 -1796 10324 -1764
rect 10356 -1796 10404 -1764
rect 10436 -1796 10484 -1764
rect 10516 -1796 10564 -1764
rect 10596 -1796 10644 -1764
rect 10676 -1796 10804 -1764
rect 10836 -1796 10964 -1764
rect 10996 -1796 11000 -1764
rect -720 -1800 11000 -1796
rect -720 -1844 11000 -1840
rect -720 -1876 -716 -1844
rect -684 -1876 -556 -1844
rect -524 -1876 -396 -1844
rect -364 -1876 -236 -1844
rect -204 -1876 -156 -1844
rect -124 -1876 -76 -1844
rect -44 -1876 4 -1844
rect 36 -1876 84 -1844
rect 116 -1876 164 -1844
rect 196 -1876 244 -1844
rect 276 -1876 324 -1844
rect 356 -1876 404 -1844
rect 436 -1876 484 -1844
rect 516 -1876 564 -1844
rect 596 -1876 644 -1844
rect 676 -1876 724 -1844
rect 756 -1876 804 -1844
rect 836 -1876 884 -1844
rect 916 -1876 964 -1844
rect 996 -1876 1044 -1844
rect 1076 -1876 1124 -1844
rect 1156 -1876 1204 -1844
rect 1236 -1876 1284 -1844
rect 1316 -1876 1364 -1844
rect 1396 -1876 1444 -1844
rect 1476 -1876 1524 -1844
rect 1556 -1876 1604 -1844
rect 1636 -1876 1684 -1844
rect 1716 -1876 1764 -1844
rect 1796 -1876 1844 -1844
rect 1876 -1876 1924 -1844
rect 1956 -1876 2004 -1844
rect 2036 -1876 2084 -1844
rect 2116 -1876 2164 -1844
rect 2196 -1876 2244 -1844
rect 2276 -1876 2324 -1844
rect 2356 -1876 2404 -1844
rect 2436 -1876 2484 -1844
rect 2516 -1876 2564 -1844
rect 2596 -1876 2644 -1844
rect 2676 -1876 2724 -1844
rect 2756 -1876 2804 -1844
rect 2836 -1876 2884 -1844
rect 2916 -1876 2964 -1844
rect 2996 -1876 3044 -1844
rect 3076 -1876 3124 -1844
rect 3156 -1876 3204 -1844
rect 3236 -1876 3284 -1844
rect 3316 -1876 3364 -1844
rect 3396 -1876 3444 -1844
rect 3476 -1876 3524 -1844
rect 3556 -1876 3604 -1844
rect 3636 -1876 3684 -1844
rect 3716 -1876 3764 -1844
rect 3796 -1876 3844 -1844
rect 3876 -1876 3924 -1844
rect 3956 -1876 4004 -1844
rect 4036 -1876 4084 -1844
rect 4116 -1876 4164 -1844
rect 4196 -1876 4244 -1844
rect 4276 -1876 4324 -1844
rect 4356 -1876 4404 -1844
rect 4436 -1876 4484 -1844
rect 4516 -1876 4564 -1844
rect 4596 -1876 4644 -1844
rect 4676 -1876 4724 -1844
rect 4756 -1876 4804 -1844
rect 4836 -1876 4884 -1844
rect 4916 -1876 4964 -1844
rect 4996 -1876 5044 -1844
rect 5076 -1876 5124 -1844
rect 5156 -1876 5204 -1844
rect 5236 -1876 5284 -1844
rect 5316 -1876 5364 -1844
rect 5396 -1876 5444 -1844
rect 5476 -1876 5524 -1844
rect 5556 -1876 5604 -1844
rect 5636 -1876 5684 -1844
rect 5716 -1876 5764 -1844
rect 5796 -1876 5844 -1844
rect 5876 -1876 5924 -1844
rect 5956 -1876 6004 -1844
rect 6036 -1876 6084 -1844
rect 6116 -1876 6164 -1844
rect 6196 -1876 6244 -1844
rect 6276 -1876 6324 -1844
rect 6356 -1876 6404 -1844
rect 6436 -1876 6484 -1844
rect 6516 -1876 6564 -1844
rect 6596 -1876 6644 -1844
rect 6676 -1876 6724 -1844
rect 6756 -1876 6804 -1844
rect 6836 -1876 6884 -1844
rect 6916 -1876 6964 -1844
rect 6996 -1876 7044 -1844
rect 7076 -1876 7124 -1844
rect 7156 -1876 7204 -1844
rect 7236 -1876 7284 -1844
rect 7316 -1876 7364 -1844
rect 7396 -1876 7444 -1844
rect 7476 -1876 7524 -1844
rect 7556 -1876 7604 -1844
rect 7636 -1876 7684 -1844
rect 7716 -1876 7764 -1844
rect 7796 -1876 7844 -1844
rect 7876 -1876 7924 -1844
rect 7956 -1876 8004 -1844
rect 8036 -1876 8084 -1844
rect 8116 -1876 8164 -1844
rect 8196 -1876 8244 -1844
rect 8276 -1876 8324 -1844
rect 8356 -1876 8404 -1844
rect 8436 -1876 8484 -1844
rect 8516 -1876 8564 -1844
rect 8596 -1876 8644 -1844
rect 8676 -1876 8724 -1844
rect 8756 -1876 8804 -1844
rect 8836 -1876 8884 -1844
rect 8916 -1876 8964 -1844
rect 8996 -1876 9044 -1844
rect 9076 -1876 9124 -1844
rect 9156 -1876 9204 -1844
rect 9236 -1876 9284 -1844
rect 9316 -1876 9364 -1844
rect 9396 -1876 9444 -1844
rect 9476 -1876 9524 -1844
rect 9556 -1876 9604 -1844
rect 9636 -1876 9684 -1844
rect 9716 -1876 9764 -1844
rect 9796 -1876 9844 -1844
rect 9876 -1876 9924 -1844
rect 9956 -1876 10004 -1844
rect 10036 -1876 10084 -1844
rect 10116 -1876 10164 -1844
rect 10196 -1876 10244 -1844
rect 10276 -1876 10324 -1844
rect 10356 -1876 10404 -1844
rect 10436 -1876 10484 -1844
rect 10516 -1876 10564 -1844
rect 10596 -1876 10644 -1844
rect 10676 -1876 10804 -1844
rect 10836 -1876 10964 -1844
rect 10996 -1876 11000 -1844
rect -720 -1880 11000 -1876
rect -720 -1924 10600 -1920
rect -720 -1956 -716 -1924
rect -684 -1956 -556 -1924
rect -524 -1956 -396 -1924
rect -364 -1956 -236 -1924
rect -204 -1956 -156 -1924
rect -124 -1956 -76 -1924
rect -44 -1956 4 -1924
rect 36 -1956 84 -1924
rect 116 -1956 164 -1924
rect 196 -1956 244 -1924
rect 276 -1956 324 -1924
rect 356 -1956 404 -1924
rect 436 -1956 484 -1924
rect 516 -1956 564 -1924
rect 596 -1956 644 -1924
rect 676 -1956 724 -1924
rect 756 -1956 804 -1924
rect 836 -1956 884 -1924
rect 916 -1956 964 -1924
rect 996 -1956 1044 -1924
rect 1076 -1956 1124 -1924
rect 1156 -1956 1204 -1924
rect 1236 -1956 1284 -1924
rect 1316 -1956 1364 -1924
rect 1396 -1956 1444 -1924
rect 1476 -1956 1524 -1924
rect 1556 -1956 1604 -1924
rect 1636 -1956 1684 -1924
rect 1716 -1956 1764 -1924
rect 1796 -1956 1844 -1924
rect 1876 -1956 1924 -1924
rect 1956 -1956 2004 -1924
rect 2036 -1956 2084 -1924
rect 2116 -1956 2164 -1924
rect 2196 -1956 2244 -1924
rect 2276 -1956 2324 -1924
rect 2356 -1956 2404 -1924
rect 2436 -1956 2484 -1924
rect 2516 -1956 2564 -1924
rect 2596 -1956 2644 -1924
rect 2676 -1956 2724 -1924
rect 2756 -1956 2804 -1924
rect 2836 -1956 2884 -1924
rect 2916 -1956 2964 -1924
rect 2996 -1956 3044 -1924
rect 3076 -1956 3124 -1924
rect 3156 -1956 3204 -1924
rect 3236 -1956 3284 -1924
rect 3316 -1956 3364 -1924
rect 3396 -1956 3444 -1924
rect 3476 -1956 3524 -1924
rect 3556 -1956 3604 -1924
rect 3636 -1956 3684 -1924
rect 3716 -1956 3764 -1924
rect 3796 -1956 3844 -1924
rect 3876 -1956 3924 -1924
rect 3956 -1956 4004 -1924
rect 4036 -1956 4084 -1924
rect 4116 -1956 4164 -1924
rect 4196 -1956 4244 -1924
rect 4276 -1956 4324 -1924
rect 4356 -1956 4404 -1924
rect 4436 -1956 4484 -1924
rect 4516 -1956 4564 -1924
rect 4596 -1956 4644 -1924
rect 4676 -1956 4724 -1924
rect 4756 -1956 4804 -1924
rect 4836 -1956 4884 -1924
rect 4916 -1956 4964 -1924
rect 4996 -1956 5044 -1924
rect 5076 -1956 5124 -1924
rect 5156 -1956 5204 -1924
rect 5236 -1956 5284 -1924
rect 5316 -1956 5364 -1924
rect 5396 -1956 5444 -1924
rect 5476 -1956 5524 -1924
rect 5556 -1956 5604 -1924
rect 5636 -1956 5684 -1924
rect 5716 -1956 5764 -1924
rect 5796 -1956 5844 -1924
rect 5876 -1956 5924 -1924
rect 5956 -1956 6004 -1924
rect 6036 -1956 6084 -1924
rect 6116 -1956 6164 -1924
rect 6196 -1956 6244 -1924
rect 6276 -1956 6324 -1924
rect 6356 -1956 6404 -1924
rect 6436 -1956 6484 -1924
rect 6516 -1956 6564 -1924
rect 6596 -1956 6644 -1924
rect 6676 -1956 6724 -1924
rect 6756 -1956 6804 -1924
rect 6836 -1956 6884 -1924
rect 6916 -1956 6964 -1924
rect 6996 -1956 7044 -1924
rect 7076 -1956 7124 -1924
rect 7156 -1956 7204 -1924
rect 7236 -1956 7284 -1924
rect 7316 -1956 7364 -1924
rect 7396 -1956 7444 -1924
rect 7476 -1956 7524 -1924
rect 7556 -1956 7604 -1924
rect 7636 -1956 7684 -1924
rect 7716 -1956 7764 -1924
rect 7796 -1956 7844 -1924
rect 7876 -1956 7924 -1924
rect 7956 -1956 8004 -1924
rect 8036 -1956 8084 -1924
rect 8116 -1956 8164 -1924
rect 8196 -1956 8244 -1924
rect 8276 -1956 8324 -1924
rect 8356 -1956 8404 -1924
rect 8436 -1956 8484 -1924
rect 8516 -1956 8564 -1924
rect 8596 -1956 8644 -1924
rect 8676 -1956 8724 -1924
rect 8756 -1956 8804 -1924
rect 8836 -1956 8884 -1924
rect 8916 -1956 8964 -1924
rect 8996 -1956 9044 -1924
rect 9076 -1956 9124 -1924
rect 9156 -1956 9204 -1924
rect 9236 -1956 9284 -1924
rect 9316 -1956 9364 -1924
rect 9396 -1956 9444 -1924
rect 9476 -1956 9524 -1924
rect 9556 -1956 9604 -1924
rect 9636 -1956 9684 -1924
rect 9716 -1956 9764 -1924
rect 9796 -1956 9844 -1924
rect 9876 -1956 9924 -1924
rect 9956 -1956 10004 -1924
rect 10036 -1956 10084 -1924
rect 10116 -1956 10164 -1924
rect 10196 -1956 10244 -1924
rect 10276 -1956 10324 -1924
rect 10356 -1956 10404 -1924
rect 10436 -1956 10484 -1924
rect 10516 -1956 10564 -1924
rect 10596 -1956 10600 -1924
rect -720 -1960 10600 -1956
rect 10640 -1924 11000 -1920
rect 10640 -1956 10644 -1924
rect 10676 -1956 10804 -1924
rect 10836 -1956 10964 -1924
rect 10996 -1956 11000 -1924
rect 10640 -1960 11000 -1956
rect -720 -2004 11000 -2000
rect -720 -2036 -716 -2004
rect -684 -2036 -556 -2004
rect -524 -2036 -396 -2004
rect -364 -2036 -236 -2004
rect -204 -2036 -156 -2004
rect -124 -2036 -76 -2004
rect -44 -2036 4 -2004
rect 36 -2036 84 -2004
rect 116 -2036 164 -2004
rect 196 -2036 244 -2004
rect 276 -2036 324 -2004
rect 356 -2036 404 -2004
rect 436 -2036 484 -2004
rect 516 -2036 564 -2004
rect 596 -2036 644 -2004
rect 676 -2036 724 -2004
rect 756 -2036 804 -2004
rect 836 -2036 884 -2004
rect 916 -2036 964 -2004
rect 996 -2036 1044 -2004
rect 1076 -2036 1124 -2004
rect 1156 -2036 1204 -2004
rect 1236 -2036 1284 -2004
rect 1316 -2036 1364 -2004
rect 1396 -2036 1444 -2004
rect 1476 -2036 1524 -2004
rect 1556 -2036 1604 -2004
rect 1636 -2036 1684 -2004
rect 1716 -2036 1764 -2004
rect 1796 -2036 1844 -2004
rect 1876 -2036 1924 -2004
rect 1956 -2036 2004 -2004
rect 2036 -2036 2084 -2004
rect 2116 -2036 2164 -2004
rect 2196 -2036 2244 -2004
rect 2276 -2036 2324 -2004
rect 2356 -2036 2404 -2004
rect 2436 -2036 2484 -2004
rect 2516 -2036 2564 -2004
rect 2596 -2036 2644 -2004
rect 2676 -2036 2724 -2004
rect 2756 -2036 2804 -2004
rect 2836 -2036 2884 -2004
rect 2916 -2036 2964 -2004
rect 2996 -2036 3044 -2004
rect 3076 -2036 3124 -2004
rect 3156 -2036 3204 -2004
rect 3236 -2036 3284 -2004
rect 3316 -2036 3364 -2004
rect 3396 -2036 3444 -2004
rect 3476 -2036 3524 -2004
rect 3556 -2036 3604 -2004
rect 3636 -2036 3684 -2004
rect 3716 -2036 3764 -2004
rect 3796 -2036 3844 -2004
rect 3876 -2036 3924 -2004
rect 3956 -2036 4004 -2004
rect 4036 -2036 4084 -2004
rect 4116 -2036 4164 -2004
rect 4196 -2036 4244 -2004
rect 4276 -2036 4324 -2004
rect 4356 -2036 4404 -2004
rect 4436 -2036 4484 -2004
rect 4516 -2036 4564 -2004
rect 4596 -2036 4644 -2004
rect 4676 -2036 4724 -2004
rect 4756 -2036 4804 -2004
rect 4836 -2036 4884 -2004
rect 4916 -2036 4964 -2004
rect 4996 -2036 5044 -2004
rect 5076 -2036 5124 -2004
rect 5156 -2036 5204 -2004
rect 5236 -2036 5284 -2004
rect 5316 -2036 5364 -2004
rect 5396 -2036 5444 -2004
rect 5476 -2036 5524 -2004
rect 5556 -2036 5604 -2004
rect 5636 -2036 5684 -2004
rect 5716 -2036 5764 -2004
rect 5796 -2036 5844 -2004
rect 5876 -2036 5924 -2004
rect 5956 -2036 6004 -2004
rect 6036 -2036 6084 -2004
rect 6116 -2036 6164 -2004
rect 6196 -2036 6244 -2004
rect 6276 -2036 6324 -2004
rect 6356 -2036 6404 -2004
rect 6436 -2036 6484 -2004
rect 6516 -2036 6564 -2004
rect 6596 -2036 6644 -2004
rect 6676 -2036 6724 -2004
rect 6756 -2036 6804 -2004
rect 6836 -2036 6884 -2004
rect 6916 -2036 6964 -2004
rect 6996 -2036 7044 -2004
rect 7076 -2036 7124 -2004
rect 7156 -2036 7204 -2004
rect 7236 -2036 7284 -2004
rect 7316 -2036 7364 -2004
rect 7396 -2036 7444 -2004
rect 7476 -2036 7524 -2004
rect 7556 -2036 7604 -2004
rect 7636 -2036 7684 -2004
rect 7716 -2036 7764 -2004
rect 7796 -2036 7844 -2004
rect 7876 -2036 7924 -2004
rect 7956 -2036 8004 -2004
rect 8036 -2036 8084 -2004
rect 8116 -2036 8164 -2004
rect 8196 -2036 8244 -2004
rect 8276 -2036 8324 -2004
rect 8356 -2036 8404 -2004
rect 8436 -2036 8484 -2004
rect 8516 -2036 8564 -2004
rect 8596 -2036 8644 -2004
rect 8676 -2036 8724 -2004
rect 8756 -2036 8804 -2004
rect 8836 -2036 8884 -2004
rect 8916 -2036 8964 -2004
rect 8996 -2036 9044 -2004
rect 9076 -2036 9124 -2004
rect 9156 -2036 9204 -2004
rect 9236 -2036 9284 -2004
rect 9316 -2036 9364 -2004
rect 9396 -2036 9444 -2004
rect 9476 -2036 9524 -2004
rect 9556 -2036 9604 -2004
rect 9636 -2036 9684 -2004
rect 9716 -2036 9764 -2004
rect 9796 -2036 9844 -2004
rect 9876 -2036 9924 -2004
rect 9956 -2036 10004 -2004
rect 10036 -2036 10084 -2004
rect 10116 -2036 10164 -2004
rect 10196 -2036 10244 -2004
rect 10276 -2036 10324 -2004
rect 10356 -2036 10404 -2004
rect 10436 -2036 10484 -2004
rect 10516 -2036 10564 -2004
rect 10596 -2036 10644 -2004
rect 10676 -2036 10804 -2004
rect 10836 -2036 10964 -2004
rect 10996 -2036 11000 -2004
rect -720 -2040 11000 -2036
rect -720 -2084 -360 -2080
rect -720 -2116 -716 -2084
rect -684 -2116 -556 -2084
rect -524 -2116 -396 -2084
rect -364 -2116 -360 -2084
rect -720 -2120 -360 -2116
rect -320 -2084 11000 -2080
rect -320 -2116 -236 -2084
rect -204 -2116 -156 -2084
rect -124 -2116 -76 -2084
rect -44 -2116 4 -2084
rect 36 -2116 84 -2084
rect 116 -2116 164 -2084
rect 196 -2116 244 -2084
rect 276 -2116 324 -2084
rect 356 -2116 404 -2084
rect 436 -2116 484 -2084
rect 516 -2116 564 -2084
rect 596 -2116 644 -2084
rect 676 -2116 724 -2084
rect 756 -2116 804 -2084
rect 836 -2116 884 -2084
rect 916 -2116 964 -2084
rect 996 -2116 1044 -2084
rect 1076 -2116 1124 -2084
rect 1156 -2116 1204 -2084
rect 1236 -2116 1284 -2084
rect 1316 -2116 1364 -2084
rect 1396 -2116 1444 -2084
rect 1476 -2116 1524 -2084
rect 1556 -2116 1604 -2084
rect 1636 -2116 1684 -2084
rect 1716 -2116 1764 -2084
rect 1796 -2116 1844 -2084
rect 1876 -2116 1924 -2084
rect 1956 -2116 2004 -2084
rect 2036 -2116 2084 -2084
rect 2116 -2116 2164 -2084
rect 2196 -2116 2244 -2084
rect 2276 -2116 2324 -2084
rect 2356 -2116 2404 -2084
rect 2436 -2116 2484 -2084
rect 2516 -2116 2564 -2084
rect 2596 -2116 2644 -2084
rect 2676 -2116 2724 -2084
rect 2756 -2116 2804 -2084
rect 2836 -2116 2884 -2084
rect 2916 -2116 2964 -2084
rect 2996 -2116 3044 -2084
rect 3076 -2116 3124 -2084
rect 3156 -2116 3204 -2084
rect 3236 -2116 3284 -2084
rect 3316 -2116 3364 -2084
rect 3396 -2116 3444 -2084
rect 3476 -2116 3524 -2084
rect 3556 -2116 3604 -2084
rect 3636 -2116 3684 -2084
rect 3716 -2116 3764 -2084
rect 3796 -2116 3844 -2084
rect 3876 -2116 3924 -2084
rect 3956 -2116 4004 -2084
rect 4036 -2116 4084 -2084
rect 4116 -2116 4164 -2084
rect 4196 -2116 4244 -2084
rect 4276 -2116 4324 -2084
rect 4356 -2116 4404 -2084
rect 4436 -2116 4484 -2084
rect 4516 -2116 4564 -2084
rect 4596 -2116 4644 -2084
rect 4676 -2116 4724 -2084
rect 4756 -2116 4804 -2084
rect 4836 -2116 4884 -2084
rect 4916 -2116 4964 -2084
rect 4996 -2116 5044 -2084
rect 5076 -2116 5124 -2084
rect 5156 -2116 5204 -2084
rect 5236 -2116 5284 -2084
rect 5316 -2116 5364 -2084
rect 5396 -2116 5444 -2084
rect 5476 -2116 5524 -2084
rect 5556 -2116 5604 -2084
rect 5636 -2116 5684 -2084
rect 5716 -2116 5764 -2084
rect 5796 -2116 5844 -2084
rect 5876 -2116 5924 -2084
rect 5956 -2116 6004 -2084
rect 6036 -2116 6084 -2084
rect 6116 -2116 6164 -2084
rect 6196 -2116 6244 -2084
rect 6276 -2116 6324 -2084
rect 6356 -2116 6404 -2084
rect 6436 -2116 6484 -2084
rect 6516 -2116 6564 -2084
rect 6596 -2116 6644 -2084
rect 6676 -2116 6724 -2084
rect 6756 -2116 6804 -2084
rect 6836 -2116 6884 -2084
rect 6916 -2116 6964 -2084
rect 6996 -2116 7044 -2084
rect 7076 -2116 7124 -2084
rect 7156 -2116 7204 -2084
rect 7236 -2116 7284 -2084
rect 7316 -2116 7364 -2084
rect 7396 -2116 7444 -2084
rect 7476 -2116 7524 -2084
rect 7556 -2116 7604 -2084
rect 7636 -2116 7684 -2084
rect 7716 -2116 7764 -2084
rect 7796 -2116 7844 -2084
rect 7876 -2116 7924 -2084
rect 7956 -2116 8004 -2084
rect 8036 -2116 8084 -2084
rect 8116 -2116 8164 -2084
rect 8196 -2116 8244 -2084
rect 8276 -2116 8324 -2084
rect 8356 -2116 8404 -2084
rect 8436 -2116 8484 -2084
rect 8516 -2116 8564 -2084
rect 8596 -2116 8644 -2084
rect 8676 -2116 8724 -2084
rect 8756 -2116 8804 -2084
rect 8836 -2116 8884 -2084
rect 8916 -2116 8964 -2084
rect 8996 -2116 9044 -2084
rect 9076 -2116 9124 -2084
rect 9156 -2116 9204 -2084
rect 9236 -2116 9284 -2084
rect 9316 -2116 9364 -2084
rect 9396 -2116 9444 -2084
rect 9476 -2116 9524 -2084
rect 9556 -2116 9604 -2084
rect 9636 -2116 9684 -2084
rect 9716 -2116 9764 -2084
rect 9796 -2116 9844 -2084
rect 9876 -2116 9924 -2084
rect 9956 -2116 10004 -2084
rect 10036 -2116 10084 -2084
rect 10116 -2116 10164 -2084
rect 10196 -2116 10244 -2084
rect 10276 -2116 10324 -2084
rect 10356 -2116 10404 -2084
rect 10436 -2116 10484 -2084
rect 10516 -2116 10564 -2084
rect 10596 -2116 10644 -2084
rect 10676 -2116 10804 -2084
rect 10836 -2116 10964 -2084
rect 10996 -2116 11000 -2084
rect -320 -2120 11000 -2116
rect -720 -2164 11000 -2160
rect -720 -2196 -716 -2164
rect -684 -2196 -556 -2164
rect -524 -2196 -396 -2164
rect -364 -2196 -236 -2164
rect -204 -2196 -156 -2164
rect -124 -2196 -76 -2164
rect -44 -2196 4 -2164
rect 36 -2196 84 -2164
rect 116 -2196 164 -2164
rect 196 -2196 244 -2164
rect 276 -2196 324 -2164
rect 356 -2196 404 -2164
rect 436 -2196 484 -2164
rect 516 -2196 564 -2164
rect 596 -2196 644 -2164
rect 676 -2196 724 -2164
rect 756 -2196 804 -2164
rect 836 -2196 884 -2164
rect 916 -2196 964 -2164
rect 996 -2196 1044 -2164
rect 1076 -2196 1124 -2164
rect 1156 -2196 1204 -2164
rect 1236 -2196 1284 -2164
rect 1316 -2196 1364 -2164
rect 1396 -2196 1444 -2164
rect 1476 -2196 1524 -2164
rect 1556 -2196 1604 -2164
rect 1636 -2196 1684 -2164
rect 1716 -2196 1764 -2164
rect 1796 -2196 1844 -2164
rect 1876 -2196 1924 -2164
rect 1956 -2196 2004 -2164
rect 2036 -2196 2084 -2164
rect 2116 -2196 2164 -2164
rect 2196 -2196 2244 -2164
rect 2276 -2196 2324 -2164
rect 2356 -2196 2404 -2164
rect 2436 -2196 2484 -2164
rect 2516 -2196 2564 -2164
rect 2596 -2196 2644 -2164
rect 2676 -2196 2724 -2164
rect 2756 -2196 2804 -2164
rect 2836 -2196 2884 -2164
rect 2916 -2196 2964 -2164
rect 2996 -2196 3044 -2164
rect 3076 -2196 3124 -2164
rect 3156 -2196 3204 -2164
rect 3236 -2196 3284 -2164
rect 3316 -2196 3364 -2164
rect 3396 -2196 3444 -2164
rect 3476 -2196 3524 -2164
rect 3556 -2196 3604 -2164
rect 3636 -2196 3684 -2164
rect 3716 -2196 3764 -2164
rect 3796 -2196 3844 -2164
rect 3876 -2196 3924 -2164
rect 3956 -2196 4004 -2164
rect 4036 -2196 4084 -2164
rect 4116 -2196 4164 -2164
rect 4196 -2196 4244 -2164
rect 4276 -2196 4324 -2164
rect 4356 -2196 4404 -2164
rect 4436 -2196 4484 -2164
rect 4516 -2196 4564 -2164
rect 4596 -2196 4644 -2164
rect 4676 -2196 4724 -2164
rect 4756 -2196 4804 -2164
rect 4836 -2196 4884 -2164
rect 4916 -2196 4964 -2164
rect 4996 -2196 5044 -2164
rect 5076 -2196 5124 -2164
rect 5156 -2196 5204 -2164
rect 5236 -2196 5284 -2164
rect 5316 -2196 5364 -2164
rect 5396 -2196 5444 -2164
rect 5476 -2196 5524 -2164
rect 5556 -2196 5604 -2164
rect 5636 -2196 5684 -2164
rect 5716 -2196 5764 -2164
rect 5796 -2196 5844 -2164
rect 5876 -2196 5924 -2164
rect 5956 -2196 6004 -2164
rect 6036 -2196 6084 -2164
rect 6116 -2196 6164 -2164
rect 6196 -2196 6244 -2164
rect 6276 -2196 6324 -2164
rect 6356 -2196 6404 -2164
rect 6436 -2196 6484 -2164
rect 6516 -2196 6564 -2164
rect 6596 -2196 6644 -2164
rect 6676 -2196 6724 -2164
rect 6756 -2196 6804 -2164
rect 6836 -2196 6884 -2164
rect 6916 -2196 6964 -2164
rect 6996 -2196 7044 -2164
rect 7076 -2196 7124 -2164
rect 7156 -2196 7204 -2164
rect 7236 -2196 7284 -2164
rect 7316 -2196 7364 -2164
rect 7396 -2196 7444 -2164
rect 7476 -2196 7524 -2164
rect 7556 -2196 7604 -2164
rect 7636 -2196 7684 -2164
rect 7716 -2196 7764 -2164
rect 7796 -2196 7844 -2164
rect 7876 -2196 7924 -2164
rect 7956 -2196 8004 -2164
rect 8036 -2196 8084 -2164
rect 8116 -2196 8164 -2164
rect 8196 -2196 8244 -2164
rect 8276 -2196 8324 -2164
rect 8356 -2196 8404 -2164
rect 8436 -2196 8484 -2164
rect 8516 -2196 8564 -2164
rect 8596 -2196 8644 -2164
rect 8676 -2196 8724 -2164
rect 8756 -2196 8804 -2164
rect 8836 -2196 8884 -2164
rect 8916 -2196 8964 -2164
rect 8996 -2196 9044 -2164
rect 9076 -2196 9124 -2164
rect 9156 -2196 9204 -2164
rect 9236 -2196 9284 -2164
rect 9316 -2196 9364 -2164
rect 9396 -2196 9444 -2164
rect 9476 -2196 9524 -2164
rect 9556 -2196 9604 -2164
rect 9636 -2196 9684 -2164
rect 9716 -2196 9764 -2164
rect 9796 -2196 9844 -2164
rect 9876 -2196 9924 -2164
rect 9956 -2196 10004 -2164
rect 10036 -2196 10084 -2164
rect 10116 -2196 10164 -2164
rect 10196 -2196 10244 -2164
rect 10276 -2196 10324 -2164
rect 10356 -2196 10404 -2164
rect 10436 -2196 10484 -2164
rect 10516 -2196 10564 -2164
rect 10596 -2196 10644 -2164
rect 10676 -2196 10804 -2164
rect 10836 -2196 10964 -2164
rect 10996 -2196 11000 -2164
rect -720 -2200 11000 -2196
rect -720 -2244 -360 -2240
rect -720 -2276 -716 -2244
rect -684 -2276 -556 -2244
rect -524 -2276 -396 -2244
rect -364 -2276 -360 -2244
rect -720 -2280 -360 -2276
rect -320 -2244 11000 -2240
rect -320 -2276 -236 -2244
rect -204 -2276 -156 -2244
rect -124 -2276 -76 -2244
rect -44 -2276 4 -2244
rect 36 -2276 84 -2244
rect 116 -2276 164 -2244
rect 196 -2276 244 -2244
rect 276 -2276 324 -2244
rect 356 -2276 404 -2244
rect 436 -2276 484 -2244
rect 516 -2276 564 -2244
rect 596 -2276 644 -2244
rect 676 -2276 724 -2244
rect 756 -2276 804 -2244
rect 836 -2276 884 -2244
rect 916 -2276 964 -2244
rect 996 -2276 1044 -2244
rect 1076 -2276 1124 -2244
rect 1156 -2276 1204 -2244
rect 1236 -2276 1284 -2244
rect 1316 -2276 1364 -2244
rect 1396 -2276 1444 -2244
rect 1476 -2276 1524 -2244
rect 1556 -2276 1604 -2244
rect 1636 -2276 1684 -2244
rect 1716 -2276 1764 -2244
rect 1796 -2276 1844 -2244
rect 1876 -2276 1924 -2244
rect 1956 -2276 2004 -2244
rect 2036 -2276 2084 -2244
rect 2116 -2276 2164 -2244
rect 2196 -2276 2244 -2244
rect 2276 -2276 2324 -2244
rect 2356 -2276 2404 -2244
rect 2436 -2276 2484 -2244
rect 2516 -2276 2564 -2244
rect 2596 -2276 2644 -2244
rect 2676 -2276 2724 -2244
rect 2756 -2276 2804 -2244
rect 2836 -2276 2884 -2244
rect 2916 -2276 2964 -2244
rect 2996 -2276 3044 -2244
rect 3076 -2276 3124 -2244
rect 3156 -2276 3204 -2244
rect 3236 -2276 3284 -2244
rect 3316 -2276 3364 -2244
rect 3396 -2276 3444 -2244
rect 3476 -2276 3524 -2244
rect 3556 -2276 3604 -2244
rect 3636 -2276 3684 -2244
rect 3716 -2276 3764 -2244
rect 3796 -2276 3844 -2244
rect 3876 -2276 3924 -2244
rect 3956 -2276 4004 -2244
rect 4036 -2276 4084 -2244
rect 4116 -2276 4164 -2244
rect 4196 -2276 4244 -2244
rect 4276 -2276 4324 -2244
rect 4356 -2276 4404 -2244
rect 4436 -2276 4484 -2244
rect 4516 -2276 4564 -2244
rect 4596 -2276 4644 -2244
rect 4676 -2276 4724 -2244
rect 4756 -2276 4804 -2244
rect 4836 -2276 4884 -2244
rect 4916 -2276 4964 -2244
rect 4996 -2276 5044 -2244
rect 5076 -2276 5124 -2244
rect 5156 -2276 5204 -2244
rect 5236 -2276 5284 -2244
rect 5316 -2276 5364 -2244
rect 5396 -2276 5444 -2244
rect 5476 -2276 5524 -2244
rect 5556 -2276 5604 -2244
rect 5636 -2276 5684 -2244
rect 5716 -2276 5764 -2244
rect 5796 -2276 5844 -2244
rect 5876 -2276 5924 -2244
rect 5956 -2276 6004 -2244
rect 6036 -2276 6084 -2244
rect 6116 -2276 6164 -2244
rect 6196 -2276 6244 -2244
rect 6276 -2276 6324 -2244
rect 6356 -2276 6404 -2244
rect 6436 -2276 6484 -2244
rect 6516 -2276 6564 -2244
rect 6596 -2276 6644 -2244
rect 6676 -2276 6724 -2244
rect 6756 -2276 6804 -2244
rect 6836 -2276 6884 -2244
rect 6916 -2276 6964 -2244
rect 6996 -2276 7044 -2244
rect 7076 -2276 7124 -2244
rect 7156 -2276 7204 -2244
rect 7236 -2276 7284 -2244
rect 7316 -2276 7364 -2244
rect 7396 -2276 7444 -2244
rect 7476 -2276 7524 -2244
rect 7556 -2276 7604 -2244
rect 7636 -2276 7684 -2244
rect 7716 -2276 7764 -2244
rect 7796 -2276 7844 -2244
rect 7876 -2276 7924 -2244
rect 7956 -2276 8004 -2244
rect 8036 -2276 8084 -2244
rect 8116 -2276 8164 -2244
rect 8196 -2276 8244 -2244
rect 8276 -2276 8324 -2244
rect 8356 -2276 8404 -2244
rect 8436 -2276 8484 -2244
rect 8516 -2276 8564 -2244
rect 8596 -2276 8644 -2244
rect 8676 -2276 8724 -2244
rect 8756 -2276 8804 -2244
rect 8836 -2276 8884 -2244
rect 8916 -2276 8964 -2244
rect 8996 -2276 9044 -2244
rect 9076 -2276 9124 -2244
rect 9156 -2276 9204 -2244
rect 9236 -2276 9284 -2244
rect 9316 -2276 9364 -2244
rect 9396 -2276 9444 -2244
rect 9476 -2276 9524 -2244
rect 9556 -2276 9604 -2244
rect 9636 -2276 9684 -2244
rect 9716 -2276 9764 -2244
rect 9796 -2276 9844 -2244
rect 9876 -2276 9924 -2244
rect 9956 -2276 10004 -2244
rect 10036 -2276 10084 -2244
rect 10116 -2276 10164 -2244
rect 10196 -2276 10244 -2244
rect 10276 -2276 10324 -2244
rect 10356 -2276 10404 -2244
rect 10436 -2276 10484 -2244
rect 10516 -2276 10564 -2244
rect 10596 -2276 10644 -2244
rect 10676 -2276 10804 -2244
rect 10836 -2276 10964 -2244
rect 10996 -2276 11000 -2244
rect -320 -2280 11000 -2276
rect -720 -2324 11000 -2320
rect -720 -2356 -716 -2324
rect -684 -2356 -556 -2324
rect -524 -2356 -396 -2324
rect -364 -2356 -236 -2324
rect -204 -2356 -156 -2324
rect -124 -2356 -76 -2324
rect -44 -2356 4 -2324
rect 36 -2356 84 -2324
rect 116 -2356 164 -2324
rect 196 -2356 244 -2324
rect 276 -2356 324 -2324
rect 356 -2356 404 -2324
rect 436 -2356 484 -2324
rect 516 -2356 564 -2324
rect 596 -2356 644 -2324
rect 676 -2356 724 -2324
rect 756 -2356 804 -2324
rect 836 -2356 884 -2324
rect 916 -2356 964 -2324
rect 996 -2356 1044 -2324
rect 1076 -2356 1124 -2324
rect 1156 -2356 1204 -2324
rect 1236 -2356 1284 -2324
rect 1316 -2356 1364 -2324
rect 1396 -2356 1444 -2324
rect 1476 -2356 1524 -2324
rect 1556 -2356 1604 -2324
rect 1636 -2356 1684 -2324
rect 1716 -2356 1764 -2324
rect 1796 -2356 1844 -2324
rect 1876 -2356 1924 -2324
rect 1956 -2356 2004 -2324
rect 2036 -2356 2084 -2324
rect 2116 -2356 2164 -2324
rect 2196 -2356 2244 -2324
rect 2276 -2356 2324 -2324
rect 2356 -2356 2404 -2324
rect 2436 -2356 2484 -2324
rect 2516 -2356 2564 -2324
rect 2596 -2356 2644 -2324
rect 2676 -2356 2724 -2324
rect 2756 -2356 2804 -2324
rect 2836 -2356 2884 -2324
rect 2916 -2356 2964 -2324
rect 2996 -2356 3044 -2324
rect 3076 -2356 3124 -2324
rect 3156 -2356 3204 -2324
rect 3236 -2356 3284 -2324
rect 3316 -2356 3364 -2324
rect 3396 -2356 3444 -2324
rect 3476 -2356 3524 -2324
rect 3556 -2356 3604 -2324
rect 3636 -2356 3684 -2324
rect 3716 -2356 3764 -2324
rect 3796 -2356 3844 -2324
rect 3876 -2356 3924 -2324
rect 3956 -2356 4004 -2324
rect 4036 -2356 4084 -2324
rect 4116 -2356 4164 -2324
rect 4196 -2356 4244 -2324
rect 4276 -2356 4324 -2324
rect 4356 -2356 4404 -2324
rect 4436 -2356 4484 -2324
rect 4516 -2356 4564 -2324
rect 4596 -2356 4644 -2324
rect 4676 -2356 4724 -2324
rect 4756 -2356 4804 -2324
rect 4836 -2356 4884 -2324
rect 4916 -2356 4964 -2324
rect 4996 -2356 5044 -2324
rect 5076 -2356 5124 -2324
rect 5156 -2356 5204 -2324
rect 5236 -2356 5284 -2324
rect 5316 -2356 5364 -2324
rect 5396 -2356 5444 -2324
rect 5476 -2356 5524 -2324
rect 5556 -2356 5604 -2324
rect 5636 -2356 5684 -2324
rect 5716 -2356 5764 -2324
rect 5796 -2356 5844 -2324
rect 5876 -2356 5924 -2324
rect 5956 -2356 6004 -2324
rect 6036 -2356 6084 -2324
rect 6116 -2356 6164 -2324
rect 6196 -2356 6244 -2324
rect 6276 -2356 6324 -2324
rect 6356 -2356 6404 -2324
rect 6436 -2356 6484 -2324
rect 6516 -2356 6564 -2324
rect 6596 -2356 6644 -2324
rect 6676 -2356 6724 -2324
rect 6756 -2356 6804 -2324
rect 6836 -2356 6884 -2324
rect 6916 -2356 6964 -2324
rect 6996 -2356 7044 -2324
rect 7076 -2356 7124 -2324
rect 7156 -2356 7204 -2324
rect 7236 -2356 7284 -2324
rect 7316 -2356 7364 -2324
rect 7396 -2356 7444 -2324
rect 7476 -2356 7524 -2324
rect 7556 -2356 7604 -2324
rect 7636 -2356 7684 -2324
rect 7716 -2356 7764 -2324
rect 7796 -2356 7844 -2324
rect 7876 -2356 7924 -2324
rect 7956 -2356 8004 -2324
rect 8036 -2356 8084 -2324
rect 8116 -2356 8164 -2324
rect 8196 -2356 8244 -2324
rect 8276 -2356 8324 -2324
rect 8356 -2356 8404 -2324
rect 8436 -2356 8484 -2324
rect 8516 -2356 8564 -2324
rect 8596 -2356 8644 -2324
rect 8676 -2356 8724 -2324
rect 8756 -2356 8804 -2324
rect 8836 -2356 8884 -2324
rect 8916 -2356 8964 -2324
rect 8996 -2356 9044 -2324
rect 9076 -2356 9124 -2324
rect 9156 -2356 9204 -2324
rect 9236 -2356 9284 -2324
rect 9316 -2356 9364 -2324
rect 9396 -2356 9444 -2324
rect 9476 -2356 9524 -2324
rect 9556 -2356 9604 -2324
rect 9636 -2356 9684 -2324
rect 9716 -2356 9764 -2324
rect 9796 -2356 9844 -2324
rect 9876 -2356 9924 -2324
rect 9956 -2356 10004 -2324
rect 10036 -2356 10084 -2324
rect 10116 -2356 10164 -2324
rect 10196 -2356 10244 -2324
rect 10276 -2356 10324 -2324
rect 10356 -2356 10404 -2324
rect 10436 -2356 10484 -2324
rect 10516 -2356 10564 -2324
rect 10596 -2356 10644 -2324
rect 10676 -2356 10804 -2324
rect 10836 -2356 10964 -2324
rect 10996 -2356 11000 -2324
rect -720 -2360 11000 -2356
rect -720 -2404 11000 -2400
rect -720 -2436 -716 -2404
rect -684 -2436 -556 -2404
rect -524 -2436 -396 -2404
rect -364 -2436 -236 -2404
rect -204 -2436 -156 -2404
rect -124 -2436 -76 -2404
rect -44 -2436 4 -2404
rect 36 -2436 84 -2404
rect 116 -2436 164 -2404
rect 196 -2436 244 -2404
rect 276 -2436 324 -2404
rect 356 -2436 404 -2404
rect 436 -2436 484 -2404
rect 516 -2436 564 -2404
rect 596 -2436 644 -2404
rect 676 -2436 724 -2404
rect 756 -2436 804 -2404
rect 836 -2436 884 -2404
rect 916 -2436 964 -2404
rect 996 -2436 1044 -2404
rect 1076 -2436 1124 -2404
rect 1156 -2436 1204 -2404
rect 1236 -2436 1284 -2404
rect 1316 -2436 1364 -2404
rect 1396 -2436 1444 -2404
rect 1476 -2436 1524 -2404
rect 1556 -2436 1604 -2404
rect 1636 -2436 1684 -2404
rect 1716 -2436 1764 -2404
rect 1796 -2436 1844 -2404
rect 1876 -2436 1924 -2404
rect 1956 -2436 2004 -2404
rect 2036 -2436 2084 -2404
rect 2116 -2436 2164 -2404
rect 2196 -2436 2244 -2404
rect 2276 -2436 2324 -2404
rect 2356 -2436 2404 -2404
rect 2436 -2436 2484 -2404
rect 2516 -2436 2564 -2404
rect 2596 -2436 2644 -2404
rect 2676 -2436 2724 -2404
rect 2756 -2436 2804 -2404
rect 2836 -2436 2884 -2404
rect 2916 -2436 2964 -2404
rect 2996 -2436 3044 -2404
rect 3076 -2436 3124 -2404
rect 3156 -2436 3204 -2404
rect 3236 -2436 3284 -2404
rect 3316 -2436 3364 -2404
rect 3396 -2436 3444 -2404
rect 3476 -2436 3524 -2404
rect 3556 -2436 3604 -2404
rect 3636 -2436 3684 -2404
rect 3716 -2436 3764 -2404
rect 3796 -2436 3844 -2404
rect 3876 -2436 3924 -2404
rect 3956 -2436 4004 -2404
rect 4036 -2436 4084 -2404
rect 4116 -2436 4164 -2404
rect 4196 -2436 4244 -2404
rect 4276 -2436 4324 -2404
rect 4356 -2436 4404 -2404
rect 4436 -2436 4484 -2404
rect 4516 -2436 4564 -2404
rect 4596 -2436 4644 -2404
rect 4676 -2436 4724 -2404
rect 4756 -2436 4804 -2404
rect 4836 -2436 4884 -2404
rect 4916 -2436 4964 -2404
rect 4996 -2436 5044 -2404
rect 5076 -2436 5124 -2404
rect 5156 -2436 5204 -2404
rect 5236 -2436 5284 -2404
rect 5316 -2436 5364 -2404
rect 5396 -2436 5444 -2404
rect 5476 -2436 5524 -2404
rect 5556 -2436 5604 -2404
rect 5636 -2436 5684 -2404
rect 5716 -2436 5764 -2404
rect 5796 -2436 5844 -2404
rect 5876 -2436 5924 -2404
rect 5956 -2436 6004 -2404
rect 6036 -2436 6084 -2404
rect 6116 -2436 6164 -2404
rect 6196 -2436 6244 -2404
rect 6276 -2436 6324 -2404
rect 6356 -2436 6404 -2404
rect 6436 -2436 6484 -2404
rect 6516 -2436 6564 -2404
rect 6596 -2436 6644 -2404
rect 6676 -2436 6724 -2404
rect 6756 -2436 6804 -2404
rect 6836 -2436 6884 -2404
rect 6916 -2436 6964 -2404
rect 6996 -2436 7044 -2404
rect 7076 -2436 7124 -2404
rect 7156 -2436 7204 -2404
rect 7236 -2436 7284 -2404
rect 7316 -2436 7364 -2404
rect 7396 -2436 7444 -2404
rect 7476 -2436 7524 -2404
rect 7556 -2436 7604 -2404
rect 7636 -2436 7684 -2404
rect 7716 -2436 7764 -2404
rect 7796 -2436 7844 -2404
rect 7876 -2436 7924 -2404
rect 7956 -2436 8004 -2404
rect 8036 -2436 8084 -2404
rect 8116 -2436 8164 -2404
rect 8196 -2436 8244 -2404
rect 8276 -2436 8324 -2404
rect 8356 -2436 8404 -2404
rect 8436 -2436 8484 -2404
rect 8516 -2436 8564 -2404
rect 8596 -2436 8644 -2404
rect 8676 -2436 8724 -2404
rect 8756 -2436 8804 -2404
rect 8836 -2436 8884 -2404
rect 8916 -2436 8964 -2404
rect 8996 -2436 9044 -2404
rect 9076 -2436 9124 -2404
rect 9156 -2436 9204 -2404
rect 9236 -2436 9284 -2404
rect 9316 -2436 9364 -2404
rect 9396 -2436 9444 -2404
rect 9476 -2436 9524 -2404
rect 9556 -2436 9604 -2404
rect 9636 -2436 9684 -2404
rect 9716 -2436 9764 -2404
rect 9796 -2436 9844 -2404
rect 9876 -2436 9924 -2404
rect 9956 -2436 10004 -2404
rect 10036 -2436 10084 -2404
rect 10116 -2436 10164 -2404
rect 10196 -2436 10244 -2404
rect 10276 -2436 10324 -2404
rect 10356 -2436 10404 -2404
rect 10436 -2436 10484 -2404
rect 10516 -2436 10564 -2404
rect 10596 -2436 10644 -2404
rect 10676 -2436 10804 -2404
rect 10836 -2436 10964 -2404
rect 10996 -2436 11000 -2404
rect -720 -2440 11000 -2436
rect -720 -2484 11000 -2480
rect -720 -2516 -716 -2484
rect -684 -2516 -556 -2484
rect -524 -2516 -396 -2484
rect -364 -2516 -236 -2484
rect -204 -2516 -156 -2484
rect -124 -2516 -76 -2484
rect -44 -2516 4 -2484
rect 36 -2516 84 -2484
rect 116 -2516 164 -2484
rect 196 -2516 244 -2484
rect 276 -2516 324 -2484
rect 356 -2516 404 -2484
rect 436 -2516 484 -2484
rect 516 -2516 564 -2484
rect 596 -2516 644 -2484
rect 676 -2516 724 -2484
rect 756 -2516 804 -2484
rect 836 -2516 884 -2484
rect 916 -2516 964 -2484
rect 996 -2516 1044 -2484
rect 1076 -2516 1124 -2484
rect 1156 -2516 1204 -2484
rect 1236 -2516 1284 -2484
rect 1316 -2516 1364 -2484
rect 1396 -2516 1444 -2484
rect 1476 -2516 1524 -2484
rect 1556 -2516 1604 -2484
rect 1636 -2516 1684 -2484
rect 1716 -2516 1764 -2484
rect 1796 -2516 1844 -2484
rect 1876 -2516 1924 -2484
rect 1956 -2516 2004 -2484
rect 2036 -2516 2084 -2484
rect 2116 -2516 2164 -2484
rect 2196 -2516 2244 -2484
rect 2276 -2516 2324 -2484
rect 2356 -2516 2404 -2484
rect 2436 -2516 2484 -2484
rect 2516 -2516 2564 -2484
rect 2596 -2516 2644 -2484
rect 2676 -2516 2724 -2484
rect 2756 -2516 2804 -2484
rect 2836 -2516 2884 -2484
rect 2916 -2516 2964 -2484
rect 2996 -2516 3044 -2484
rect 3076 -2516 3124 -2484
rect 3156 -2516 3204 -2484
rect 3236 -2516 3284 -2484
rect 3316 -2516 3364 -2484
rect 3396 -2516 3444 -2484
rect 3476 -2516 3524 -2484
rect 3556 -2516 3604 -2484
rect 3636 -2516 3684 -2484
rect 3716 -2516 3764 -2484
rect 3796 -2516 3844 -2484
rect 3876 -2516 3924 -2484
rect 3956 -2516 4004 -2484
rect 4036 -2516 4084 -2484
rect 4116 -2516 4164 -2484
rect 4196 -2516 4244 -2484
rect 4276 -2516 4324 -2484
rect 4356 -2516 4404 -2484
rect 4436 -2516 4484 -2484
rect 4516 -2516 4564 -2484
rect 4596 -2516 4644 -2484
rect 4676 -2516 4724 -2484
rect 4756 -2516 4804 -2484
rect 4836 -2516 4884 -2484
rect 4916 -2516 4964 -2484
rect 4996 -2516 5044 -2484
rect 5076 -2516 5124 -2484
rect 5156 -2516 5204 -2484
rect 5236 -2516 5284 -2484
rect 5316 -2516 5364 -2484
rect 5396 -2516 5444 -2484
rect 5476 -2516 5524 -2484
rect 5556 -2516 5604 -2484
rect 5636 -2516 5684 -2484
rect 5716 -2516 5764 -2484
rect 5796 -2516 5844 -2484
rect 5876 -2516 5924 -2484
rect 5956 -2516 6004 -2484
rect 6036 -2516 6084 -2484
rect 6116 -2516 6164 -2484
rect 6196 -2516 6244 -2484
rect 6276 -2516 6324 -2484
rect 6356 -2516 6404 -2484
rect 6436 -2516 6484 -2484
rect 6516 -2516 6564 -2484
rect 6596 -2516 6644 -2484
rect 6676 -2516 6724 -2484
rect 6756 -2516 6804 -2484
rect 6836 -2516 6884 -2484
rect 6916 -2516 6964 -2484
rect 6996 -2516 7044 -2484
rect 7076 -2516 7124 -2484
rect 7156 -2516 7204 -2484
rect 7236 -2516 7284 -2484
rect 7316 -2516 7364 -2484
rect 7396 -2516 7444 -2484
rect 7476 -2516 7524 -2484
rect 7556 -2516 7604 -2484
rect 7636 -2516 7684 -2484
rect 7716 -2516 7764 -2484
rect 7796 -2516 7844 -2484
rect 7876 -2516 7924 -2484
rect 7956 -2516 8004 -2484
rect 8036 -2516 8084 -2484
rect 8116 -2516 8164 -2484
rect 8196 -2516 8244 -2484
rect 8276 -2516 8324 -2484
rect 8356 -2516 8404 -2484
rect 8436 -2516 8484 -2484
rect 8516 -2516 8564 -2484
rect 8596 -2516 8644 -2484
rect 8676 -2516 8724 -2484
rect 8756 -2516 8804 -2484
rect 8836 -2516 8884 -2484
rect 8916 -2516 8964 -2484
rect 8996 -2516 9044 -2484
rect 9076 -2516 9124 -2484
rect 9156 -2516 9204 -2484
rect 9236 -2516 9284 -2484
rect 9316 -2516 9364 -2484
rect 9396 -2516 9444 -2484
rect 9476 -2516 9524 -2484
rect 9556 -2516 9604 -2484
rect 9636 -2516 9684 -2484
rect 9716 -2516 9764 -2484
rect 9796 -2516 9844 -2484
rect 9876 -2516 9924 -2484
rect 9956 -2516 10004 -2484
rect 10036 -2516 10084 -2484
rect 10116 -2516 10164 -2484
rect 10196 -2516 10244 -2484
rect 10276 -2516 10324 -2484
rect 10356 -2516 10404 -2484
rect 10436 -2516 10484 -2484
rect 10516 -2516 10564 -2484
rect 10596 -2516 10644 -2484
rect 10676 -2516 10804 -2484
rect 10836 -2516 10964 -2484
rect 10996 -2516 11000 -2484
rect -720 -2520 11000 -2516
rect -720 -2564 11000 -2560
rect -720 -2596 -716 -2564
rect -684 -2596 -556 -2564
rect -524 -2596 -396 -2564
rect -364 -2596 -316 -2564
rect -284 -2596 -236 -2564
rect -204 -2596 -156 -2564
rect -124 -2596 -76 -2564
rect -44 -2596 4 -2564
rect 36 -2596 84 -2564
rect 116 -2596 164 -2564
rect 196 -2596 244 -2564
rect 276 -2596 324 -2564
rect 356 -2596 404 -2564
rect 436 -2596 484 -2564
rect 516 -2596 564 -2564
rect 596 -2596 644 -2564
rect 676 -2596 724 -2564
rect 756 -2596 804 -2564
rect 836 -2596 884 -2564
rect 916 -2596 964 -2564
rect 996 -2596 1044 -2564
rect 1076 -2596 1124 -2564
rect 1156 -2596 1204 -2564
rect 1236 -2596 1284 -2564
rect 1316 -2596 1364 -2564
rect 1396 -2596 1444 -2564
rect 1476 -2596 1524 -2564
rect 1556 -2596 1604 -2564
rect 1636 -2596 1684 -2564
rect 1716 -2596 1764 -2564
rect 1796 -2596 1844 -2564
rect 1876 -2596 1924 -2564
rect 1956 -2596 2004 -2564
rect 2036 -2596 2084 -2564
rect 2116 -2596 2164 -2564
rect 2196 -2596 2244 -2564
rect 2276 -2596 2324 -2564
rect 2356 -2596 2404 -2564
rect 2436 -2596 2484 -2564
rect 2516 -2596 2564 -2564
rect 2596 -2596 2644 -2564
rect 2676 -2596 2724 -2564
rect 2756 -2596 2804 -2564
rect 2836 -2596 2884 -2564
rect 2916 -2596 2964 -2564
rect 2996 -2596 3044 -2564
rect 3076 -2596 3124 -2564
rect 3156 -2596 3204 -2564
rect 3236 -2596 3284 -2564
rect 3316 -2596 3364 -2564
rect 3396 -2596 3444 -2564
rect 3476 -2596 3524 -2564
rect 3556 -2596 3604 -2564
rect 3636 -2596 3684 -2564
rect 3716 -2596 3764 -2564
rect 3796 -2596 3844 -2564
rect 3876 -2596 3924 -2564
rect 3956 -2596 4004 -2564
rect 4036 -2596 4084 -2564
rect 4116 -2596 4164 -2564
rect 4196 -2596 4244 -2564
rect 4276 -2596 4324 -2564
rect 4356 -2596 4404 -2564
rect 4436 -2596 4484 -2564
rect 4516 -2596 4564 -2564
rect 4596 -2596 4644 -2564
rect 4676 -2596 4724 -2564
rect 4756 -2596 4804 -2564
rect 4836 -2596 4884 -2564
rect 4916 -2596 4964 -2564
rect 4996 -2596 5044 -2564
rect 5076 -2596 5124 -2564
rect 5156 -2596 5204 -2564
rect 5236 -2596 5284 -2564
rect 5316 -2596 5364 -2564
rect 5396 -2596 5444 -2564
rect 5476 -2596 5524 -2564
rect 5556 -2596 5604 -2564
rect 5636 -2596 5684 -2564
rect 5716 -2596 5764 -2564
rect 5796 -2596 5844 -2564
rect 5876 -2596 5924 -2564
rect 5956 -2596 6004 -2564
rect 6036 -2596 6084 -2564
rect 6116 -2596 6164 -2564
rect 6196 -2596 6244 -2564
rect 6276 -2596 6324 -2564
rect 6356 -2596 6404 -2564
rect 6436 -2596 6484 -2564
rect 6516 -2596 6564 -2564
rect 6596 -2596 6644 -2564
rect 6676 -2596 6724 -2564
rect 6756 -2596 6804 -2564
rect 6836 -2596 6884 -2564
rect 6916 -2596 6964 -2564
rect 6996 -2596 7044 -2564
rect 7076 -2596 7124 -2564
rect 7156 -2596 7204 -2564
rect 7236 -2596 7284 -2564
rect 7316 -2596 7364 -2564
rect 7396 -2596 7444 -2564
rect 7476 -2596 7524 -2564
rect 7556 -2596 7604 -2564
rect 7636 -2596 7684 -2564
rect 7716 -2596 7764 -2564
rect 7796 -2596 7844 -2564
rect 7876 -2596 7924 -2564
rect 7956 -2596 8004 -2564
rect 8036 -2596 8084 -2564
rect 8116 -2596 8164 -2564
rect 8196 -2596 8244 -2564
rect 8276 -2596 8324 -2564
rect 8356 -2596 8404 -2564
rect 8436 -2596 8484 -2564
rect 8516 -2596 8564 -2564
rect 8596 -2596 8644 -2564
rect 8676 -2596 8724 -2564
rect 8756 -2596 8804 -2564
rect 8836 -2596 8884 -2564
rect 8916 -2596 8964 -2564
rect 8996 -2596 9044 -2564
rect 9076 -2596 9124 -2564
rect 9156 -2596 9204 -2564
rect 9236 -2596 9284 -2564
rect 9316 -2596 9364 -2564
rect 9396 -2596 9444 -2564
rect 9476 -2596 9524 -2564
rect 9556 -2596 9604 -2564
rect 9636 -2596 9684 -2564
rect 9716 -2596 9764 -2564
rect 9796 -2596 9844 -2564
rect 9876 -2596 9924 -2564
rect 9956 -2596 10004 -2564
rect 10036 -2596 10084 -2564
rect 10116 -2596 10164 -2564
rect 10196 -2596 10244 -2564
rect 10276 -2596 10324 -2564
rect 10356 -2596 10404 -2564
rect 10436 -2596 10484 -2564
rect 10516 -2596 10644 -2564
rect 10676 -2596 10804 -2564
rect 10836 -2596 10964 -2564
rect 10996 -2596 11000 -2564
rect -720 -2600 11000 -2596
rect -720 -2644 11000 -2640
rect -720 -2676 -716 -2644
rect -684 -2676 -556 -2644
rect -524 -2676 -396 -2644
rect -364 -2676 -316 -2644
rect -284 -2676 -236 -2644
rect -204 -2676 -156 -2644
rect -124 -2676 -76 -2644
rect -44 -2676 4 -2644
rect 36 -2676 84 -2644
rect 116 -2676 164 -2644
rect 196 -2676 244 -2644
rect 276 -2676 324 -2644
rect 356 -2676 404 -2644
rect 436 -2676 484 -2644
rect 516 -2676 564 -2644
rect 596 -2676 644 -2644
rect 676 -2676 724 -2644
rect 756 -2676 804 -2644
rect 836 -2676 884 -2644
rect 916 -2676 964 -2644
rect 996 -2676 1044 -2644
rect 1076 -2676 1124 -2644
rect 1156 -2676 1204 -2644
rect 1236 -2676 1284 -2644
rect 1316 -2676 1364 -2644
rect 1396 -2676 1444 -2644
rect 1476 -2676 1524 -2644
rect 1556 -2676 1604 -2644
rect 1636 -2676 1684 -2644
rect 1716 -2676 1764 -2644
rect 1796 -2676 1844 -2644
rect 1876 -2676 1924 -2644
rect 1956 -2676 2004 -2644
rect 2036 -2676 2084 -2644
rect 2116 -2676 2164 -2644
rect 2196 -2676 2244 -2644
rect 2276 -2676 2324 -2644
rect 2356 -2676 2404 -2644
rect 2436 -2676 2484 -2644
rect 2516 -2676 2564 -2644
rect 2596 -2676 2644 -2644
rect 2676 -2676 2724 -2644
rect 2756 -2676 2804 -2644
rect 2836 -2676 2884 -2644
rect 2916 -2676 2964 -2644
rect 2996 -2676 3044 -2644
rect 3076 -2676 3124 -2644
rect 3156 -2676 3204 -2644
rect 3236 -2676 3284 -2644
rect 3316 -2676 3364 -2644
rect 3396 -2676 3444 -2644
rect 3476 -2676 3524 -2644
rect 3556 -2676 3604 -2644
rect 3636 -2676 3684 -2644
rect 3716 -2676 3764 -2644
rect 3796 -2676 3844 -2644
rect 3876 -2676 3924 -2644
rect 3956 -2676 4004 -2644
rect 4036 -2676 4084 -2644
rect 4116 -2676 4164 -2644
rect 4196 -2676 4244 -2644
rect 4276 -2676 4324 -2644
rect 4356 -2676 4404 -2644
rect 4436 -2676 4484 -2644
rect 4516 -2676 4564 -2644
rect 4596 -2676 4644 -2644
rect 4676 -2676 4724 -2644
rect 4756 -2676 4804 -2644
rect 4836 -2676 4884 -2644
rect 4916 -2676 4964 -2644
rect 4996 -2676 5044 -2644
rect 5076 -2676 5124 -2644
rect 5156 -2676 5204 -2644
rect 5236 -2676 5284 -2644
rect 5316 -2676 5364 -2644
rect 5396 -2676 5444 -2644
rect 5476 -2676 5524 -2644
rect 5556 -2676 5604 -2644
rect 5636 -2676 5684 -2644
rect 5716 -2676 5764 -2644
rect 5796 -2676 5844 -2644
rect 5876 -2676 5924 -2644
rect 5956 -2676 6004 -2644
rect 6036 -2676 6084 -2644
rect 6116 -2676 6164 -2644
rect 6196 -2676 6244 -2644
rect 6276 -2676 6324 -2644
rect 6356 -2676 6404 -2644
rect 6436 -2676 6484 -2644
rect 6516 -2676 6564 -2644
rect 6596 -2676 6644 -2644
rect 6676 -2676 6724 -2644
rect 6756 -2676 6804 -2644
rect 6836 -2676 6884 -2644
rect 6916 -2676 6964 -2644
rect 6996 -2676 7044 -2644
rect 7076 -2676 7124 -2644
rect 7156 -2676 7204 -2644
rect 7236 -2676 7284 -2644
rect 7316 -2676 7364 -2644
rect 7396 -2676 7444 -2644
rect 7476 -2676 7524 -2644
rect 7556 -2676 7604 -2644
rect 7636 -2676 7684 -2644
rect 7716 -2676 7764 -2644
rect 7796 -2676 7844 -2644
rect 7876 -2676 7924 -2644
rect 7956 -2676 8004 -2644
rect 8036 -2676 8084 -2644
rect 8116 -2676 8164 -2644
rect 8196 -2676 8244 -2644
rect 8276 -2676 8324 -2644
rect 8356 -2676 8404 -2644
rect 8436 -2676 8484 -2644
rect 8516 -2676 8564 -2644
rect 8596 -2676 8644 -2644
rect 8676 -2676 8724 -2644
rect 8756 -2676 8804 -2644
rect 8836 -2676 8884 -2644
rect 8916 -2676 8964 -2644
rect 8996 -2676 9044 -2644
rect 9076 -2676 9124 -2644
rect 9156 -2676 9204 -2644
rect 9236 -2676 9284 -2644
rect 9316 -2676 9364 -2644
rect 9396 -2676 9444 -2644
rect 9476 -2676 9524 -2644
rect 9556 -2676 9604 -2644
rect 9636 -2676 9684 -2644
rect 9716 -2676 9764 -2644
rect 9796 -2676 9844 -2644
rect 9876 -2676 9924 -2644
rect 9956 -2676 10004 -2644
rect 10036 -2676 10084 -2644
rect 10116 -2676 10164 -2644
rect 10196 -2676 10244 -2644
rect 10276 -2676 10324 -2644
rect 10356 -2676 10404 -2644
rect 10436 -2676 10484 -2644
rect 10516 -2676 10644 -2644
rect 10676 -2676 10804 -2644
rect 10836 -2676 10964 -2644
rect 10996 -2676 11000 -2644
rect -720 -2680 11000 -2676
rect -720 -2724 11000 -2720
rect -720 -2756 -716 -2724
rect -684 -2756 -556 -2724
rect -524 -2756 -396 -2724
rect -364 -2756 -316 -2724
rect -284 -2756 -236 -2724
rect -204 -2756 -156 -2724
rect -124 -2756 -76 -2724
rect -44 -2756 4 -2724
rect 36 -2756 84 -2724
rect 116 -2756 164 -2724
rect 196 -2756 244 -2724
rect 276 -2756 324 -2724
rect 356 -2756 404 -2724
rect 436 -2756 484 -2724
rect 516 -2756 564 -2724
rect 596 -2756 644 -2724
rect 676 -2756 724 -2724
rect 756 -2756 804 -2724
rect 836 -2756 884 -2724
rect 916 -2756 964 -2724
rect 996 -2756 1044 -2724
rect 1076 -2756 1124 -2724
rect 1156 -2756 1204 -2724
rect 1236 -2756 1284 -2724
rect 1316 -2756 1364 -2724
rect 1396 -2756 1444 -2724
rect 1476 -2756 1524 -2724
rect 1556 -2756 1604 -2724
rect 1636 -2756 1684 -2724
rect 1716 -2756 1764 -2724
rect 1796 -2756 1844 -2724
rect 1876 -2756 1924 -2724
rect 1956 -2756 2004 -2724
rect 2036 -2756 2084 -2724
rect 2116 -2756 2164 -2724
rect 2196 -2756 2244 -2724
rect 2276 -2756 2324 -2724
rect 2356 -2756 2404 -2724
rect 2436 -2756 2484 -2724
rect 2516 -2756 2564 -2724
rect 2596 -2756 2644 -2724
rect 2676 -2756 2724 -2724
rect 2756 -2756 2804 -2724
rect 2836 -2756 2884 -2724
rect 2916 -2756 2964 -2724
rect 2996 -2756 3044 -2724
rect 3076 -2756 3124 -2724
rect 3156 -2756 3204 -2724
rect 3236 -2756 3284 -2724
rect 3316 -2756 3364 -2724
rect 3396 -2756 3444 -2724
rect 3476 -2756 3524 -2724
rect 3556 -2756 3604 -2724
rect 3636 -2756 3684 -2724
rect 3716 -2756 3764 -2724
rect 3796 -2756 3844 -2724
rect 3876 -2756 3924 -2724
rect 3956 -2756 4004 -2724
rect 4036 -2756 4084 -2724
rect 4116 -2756 4164 -2724
rect 4196 -2756 4244 -2724
rect 4276 -2756 4324 -2724
rect 4356 -2756 4404 -2724
rect 4436 -2756 4484 -2724
rect 4516 -2756 4564 -2724
rect 4596 -2756 4644 -2724
rect 4676 -2756 4724 -2724
rect 4756 -2756 4804 -2724
rect 4836 -2756 4884 -2724
rect 4916 -2756 4964 -2724
rect 4996 -2756 5044 -2724
rect 5076 -2756 5124 -2724
rect 5156 -2756 5204 -2724
rect 5236 -2756 5284 -2724
rect 5316 -2756 5364 -2724
rect 5396 -2756 5444 -2724
rect 5476 -2756 5524 -2724
rect 5556 -2756 5604 -2724
rect 5636 -2756 5684 -2724
rect 5716 -2756 5764 -2724
rect 5796 -2756 5844 -2724
rect 5876 -2756 5924 -2724
rect 5956 -2756 6004 -2724
rect 6036 -2756 6084 -2724
rect 6116 -2756 6164 -2724
rect 6196 -2756 6244 -2724
rect 6276 -2756 6324 -2724
rect 6356 -2756 6404 -2724
rect 6436 -2756 6484 -2724
rect 6516 -2756 6564 -2724
rect 6596 -2756 6644 -2724
rect 6676 -2756 6724 -2724
rect 6756 -2756 6804 -2724
rect 6836 -2756 6884 -2724
rect 6916 -2756 6964 -2724
rect 6996 -2756 7044 -2724
rect 7076 -2756 7124 -2724
rect 7156 -2756 7204 -2724
rect 7236 -2756 7284 -2724
rect 7316 -2756 7364 -2724
rect 7396 -2756 7444 -2724
rect 7476 -2756 7524 -2724
rect 7556 -2756 7604 -2724
rect 7636 -2756 7684 -2724
rect 7716 -2756 7764 -2724
rect 7796 -2756 7844 -2724
rect 7876 -2756 7924 -2724
rect 7956 -2756 8004 -2724
rect 8036 -2756 8084 -2724
rect 8116 -2756 8164 -2724
rect 8196 -2756 8244 -2724
rect 8276 -2756 8324 -2724
rect 8356 -2756 8404 -2724
rect 8436 -2756 8484 -2724
rect 8516 -2756 8564 -2724
rect 8596 -2756 8644 -2724
rect 8676 -2756 8724 -2724
rect 8756 -2756 8804 -2724
rect 8836 -2756 8884 -2724
rect 8916 -2756 8964 -2724
rect 8996 -2756 9044 -2724
rect 9076 -2756 9124 -2724
rect 9156 -2756 9204 -2724
rect 9236 -2756 9284 -2724
rect 9316 -2756 9364 -2724
rect 9396 -2756 9444 -2724
rect 9476 -2756 9524 -2724
rect 9556 -2756 9604 -2724
rect 9636 -2756 9684 -2724
rect 9716 -2756 9764 -2724
rect 9796 -2756 9844 -2724
rect 9876 -2756 9924 -2724
rect 9956 -2756 10004 -2724
rect 10036 -2756 10084 -2724
rect 10116 -2756 10164 -2724
rect 10196 -2756 10244 -2724
rect 10276 -2756 10324 -2724
rect 10356 -2756 10404 -2724
rect 10436 -2756 10484 -2724
rect 10516 -2756 10644 -2724
rect 10676 -2756 10804 -2724
rect 10836 -2756 10964 -2724
rect 10996 -2756 11000 -2724
rect -720 -2760 11000 -2756
rect -720 -2804 -360 -2800
rect -720 -2836 -716 -2804
rect -684 -2836 -556 -2804
rect -524 -2836 -396 -2804
rect -364 -2836 -360 -2804
rect -720 -2840 -360 -2836
rect -320 -2804 11000 -2800
rect -320 -2836 -316 -2804
rect -284 -2836 -236 -2804
rect -204 -2836 -156 -2804
rect -124 -2836 -76 -2804
rect -44 -2836 4 -2804
rect 36 -2836 84 -2804
rect 116 -2836 164 -2804
rect 196 -2836 244 -2804
rect 276 -2836 324 -2804
rect 356 -2836 404 -2804
rect 436 -2836 484 -2804
rect 516 -2836 564 -2804
rect 596 -2836 644 -2804
rect 676 -2836 724 -2804
rect 756 -2836 804 -2804
rect 836 -2836 884 -2804
rect 916 -2836 964 -2804
rect 996 -2836 1044 -2804
rect 1076 -2836 1124 -2804
rect 1156 -2836 1204 -2804
rect 1236 -2836 1284 -2804
rect 1316 -2836 1364 -2804
rect 1396 -2836 1444 -2804
rect 1476 -2836 1524 -2804
rect 1556 -2836 1604 -2804
rect 1636 -2836 1684 -2804
rect 1716 -2836 1764 -2804
rect 1796 -2836 1844 -2804
rect 1876 -2836 1924 -2804
rect 1956 -2836 2004 -2804
rect 2036 -2836 2084 -2804
rect 2116 -2836 2164 -2804
rect 2196 -2836 2244 -2804
rect 2276 -2836 2324 -2804
rect 2356 -2836 2404 -2804
rect 2436 -2836 2484 -2804
rect 2516 -2836 2564 -2804
rect 2596 -2836 2644 -2804
rect 2676 -2836 2724 -2804
rect 2756 -2836 2804 -2804
rect 2836 -2836 2884 -2804
rect 2916 -2836 2964 -2804
rect 2996 -2836 3044 -2804
rect 3076 -2836 3124 -2804
rect 3156 -2836 3204 -2804
rect 3236 -2836 3284 -2804
rect 3316 -2836 3364 -2804
rect 3396 -2836 3444 -2804
rect 3476 -2836 3524 -2804
rect 3556 -2836 3604 -2804
rect 3636 -2836 3684 -2804
rect 3716 -2836 3764 -2804
rect 3796 -2836 3844 -2804
rect 3876 -2836 3924 -2804
rect 3956 -2836 4004 -2804
rect 4036 -2836 4084 -2804
rect 4116 -2836 4164 -2804
rect 4196 -2836 4244 -2804
rect 4276 -2836 4324 -2804
rect 4356 -2836 4404 -2804
rect 4436 -2836 4484 -2804
rect 4516 -2836 4564 -2804
rect 4596 -2836 4644 -2804
rect 4676 -2836 4724 -2804
rect 4756 -2836 4804 -2804
rect 4836 -2836 4884 -2804
rect 4916 -2836 4964 -2804
rect 4996 -2836 5044 -2804
rect 5076 -2836 5124 -2804
rect 5156 -2836 5204 -2804
rect 5236 -2836 5284 -2804
rect 5316 -2836 5364 -2804
rect 5396 -2836 5444 -2804
rect 5476 -2836 5524 -2804
rect 5556 -2836 5604 -2804
rect 5636 -2836 5684 -2804
rect 5716 -2836 5764 -2804
rect 5796 -2836 5844 -2804
rect 5876 -2836 5924 -2804
rect 5956 -2836 6004 -2804
rect 6036 -2836 6084 -2804
rect 6116 -2836 6164 -2804
rect 6196 -2836 6244 -2804
rect 6276 -2836 6324 -2804
rect 6356 -2836 6404 -2804
rect 6436 -2836 6484 -2804
rect 6516 -2836 6564 -2804
rect 6596 -2836 6644 -2804
rect 6676 -2836 6724 -2804
rect 6756 -2836 6804 -2804
rect 6836 -2836 6884 -2804
rect 6916 -2836 6964 -2804
rect 6996 -2836 7044 -2804
rect 7076 -2836 7124 -2804
rect 7156 -2836 7204 -2804
rect 7236 -2836 7284 -2804
rect 7316 -2836 7364 -2804
rect 7396 -2836 7444 -2804
rect 7476 -2836 7524 -2804
rect 7556 -2836 7604 -2804
rect 7636 -2836 7684 -2804
rect 7716 -2836 7764 -2804
rect 7796 -2836 7844 -2804
rect 7876 -2836 7924 -2804
rect 7956 -2836 8004 -2804
rect 8036 -2836 8084 -2804
rect 8116 -2836 8164 -2804
rect 8196 -2836 8244 -2804
rect 8276 -2836 8324 -2804
rect 8356 -2836 8404 -2804
rect 8436 -2836 8484 -2804
rect 8516 -2836 8564 -2804
rect 8596 -2836 8644 -2804
rect 8676 -2836 8724 -2804
rect 8756 -2836 8804 -2804
rect 8836 -2836 8884 -2804
rect 8916 -2836 8964 -2804
rect 8996 -2836 9044 -2804
rect 9076 -2836 9124 -2804
rect 9156 -2836 9204 -2804
rect 9236 -2836 9284 -2804
rect 9316 -2836 9364 -2804
rect 9396 -2836 9444 -2804
rect 9476 -2836 9524 -2804
rect 9556 -2836 9604 -2804
rect 9636 -2836 9684 -2804
rect 9716 -2836 9764 -2804
rect 9796 -2836 9844 -2804
rect 9876 -2836 9924 -2804
rect 9956 -2836 10004 -2804
rect 10036 -2836 10084 -2804
rect 10116 -2836 10164 -2804
rect 10196 -2836 10244 -2804
rect 10276 -2836 10324 -2804
rect 10356 -2836 10404 -2804
rect 10436 -2836 10484 -2804
rect 10516 -2836 10644 -2804
rect 10676 -2836 10804 -2804
rect 10836 -2836 10964 -2804
rect 10996 -2836 11000 -2804
rect -320 -2840 11000 -2836
rect -720 -2884 11000 -2880
rect -720 -2916 -716 -2884
rect -684 -2916 -556 -2884
rect -524 -2916 -396 -2884
rect -364 -2916 -316 -2884
rect -284 -2916 -236 -2884
rect -204 -2916 -156 -2884
rect -124 -2916 -76 -2884
rect -44 -2916 4 -2884
rect 36 -2916 84 -2884
rect 116 -2916 164 -2884
rect 196 -2916 244 -2884
rect 276 -2916 324 -2884
rect 356 -2916 404 -2884
rect 436 -2916 484 -2884
rect 516 -2916 564 -2884
rect 596 -2916 644 -2884
rect 676 -2916 724 -2884
rect 756 -2916 804 -2884
rect 836 -2916 884 -2884
rect 916 -2916 964 -2884
rect 996 -2916 1044 -2884
rect 1076 -2916 1124 -2884
rect 1156 -2916 1204 -2884
rect 1236 -2916 1284 -2884
rect 1316 -2916 1364 -2884
rect 1396 -2916 1444 -2884
rect 1476 -2916 1524 -2884
rect 1556 -2916 1604 -2884
rect 1636 -2916 1684 -2884
rect 1716 -2916 1764 -2884
rect 1796 -2916 1844 -2884
rect 1876 -2916 1924 -2884
rect 1956 -2916 2004 -2884
rect 2036 -2916 2084 -2884
rect 2116 -2916 2164 -2884
rect 2196 -2916 2244 -2884
rect 2276 -2916 2324 -2884
rect 2356 -2916 2404 -2884
rect 2436 -2916 2484 -2884
rect 2516 -2916 2564 -2884
rect 2596 -2916 2644 -2884
rect 2676 -2916 2724 -2884
rect 2756 -2916 2804 -2884
rect 2836 -2916 2884 -2884
rect 2916 -2916 2964 -2884
rect 2996 -2916 3044 -2884
rect 3076 -2916 3124 -2884
rect 3156 -2916 3204 -2884
rect 3236 -2916 3284 -2884
rect 3316 -2916 3364 -2884
rect 3396 -2916 3444 -2884
rect 3476 -2916 3524 -2884
rect 3556 -2916 3604 -2884
rect 3636 -2916 3684 -2884
rect 3716 -2916 3764 -2884
rect 3796 -2916 3844 -2884
rect 3876 -2916 3924 -2884
rect 3956 -2916 4004 -2884
rect 4036 -2916 4084 -2884
rect 4116 -2916 4164 -2884
rect 4196 -2916 4244 -2884
rect 4276 -2916 4324 -2884
rect 4356 -2916 4404 -2884
rect 4436 -2916 4484 -2884
rect 4516 -2916 4564 -2884
rect 4596 -2916 4644 -2884
rect 4676 -2916 4724 -2884
rect 4756 -2916 4804 -2884
rect 4836 -2916 4884 -2884
rect 4916 -2916 4964 -2884
rect 4996 -2916 5044 -2884
rect 5076 -2916 5124 -2884
rect 5156 -2916 5204 -2884
rect 5236 -2916 5284 -2884
rect 5316 -2916 5364 -2884
rect 5396 -2916 5444 -2884
rect 5476 -2916 5524 -2884
rect 5556 -2916 5604 -2884
rect 5636 -2916 5684 -2884
rect 5716 -2916 5764 -2884
rect 5796 -2916 5844 -2884
rect 5876 -2916 5924 -2884
rect 5956 -2916 6004 -2884
rect 6036 -2916 6084 -2884
rect 6116 -2916 6164 -2884
rect 6196 -2916 6244 -2884
rect 6276 -2916 6324 -2884
rect 6356 -2916 6404 -2884
rect 6436 -2916 6484 -2884
rect 6516 -2916 6564 -2884
rect 6596 -2916 6644 -2884
rect 6676 -2916 6724 -2884
rect 6756 -2916 6804 -2884
rect 6836 -2916 6884 -2884
rect 6916 -2916 6964 -2884
rect 6996 -2916 7044 -2884
rect 7076 -2916 7124 -2884
rect 7156 -2916 7204 -2884
rect 7236 -2916 7284 -2884
rect 7316 -2916 7364 -2884
rect 7396 -2916 7444 -2884
rect 7476 -2916 7524 -2884
rect 7556 -2916 7604 -2884
rect 7636 -2916 7684 -2884
rect 7716 -2916 7764 -2884
rect 7796 -2916 7844 -2884
rect 7876 -2916 7924 -2884
rect 7956 -2916 8004 -2884
rect 8036 -2916 8084 -2884
rect 8116 -2916 8164 -2884
rect 8196 -2916 8244 -2884
rect 8276 -2916 8324 -2884
rect 8356 -2916 8404 -2884
rect 8436 -2916 8484 -2884
rect 8516 -2916 8564 -2884
rect 8596 -2916 8644 -2884
rect 8676 -2916 8724 -2884
rect 8756 -2916 8804 -2884
rect 8836 -2916 8884 -2884
rect 8916 -2916 8964 -2884
rect 8996 -2916 9044 -2884
rect 9076 -2916 9124 -2884
rect 9156 -2916 9204 -2884
rect 9236 -2916 9284 -2884
rect 9316 -2916 9364 -2884
rect 9396 -2916 9444 -2884
rect 9476 -2916 9524 -2884
rect 9556 -2916 9604 -2884
rect 9636 -2916 9684 -2884
rect 9716 -2916 9764 -2884
rect 9796 -2916 9844 -2884
rect 9876 -2916 9924 -2884
rect 9956 -2916 10004 -2884
rect 10036 -2916 10084 -2884
rect 10116 -2916 10164 -2884
rect 10196 -2916 10244 -2884
rect 10276 -2916 10324 -2884
rect 10356 -2916 10404 -2884
rect 10436 -2916 10484 -2884
rect 10516 -2916 10644 -2884
rect 10676 -2916 10804 -2884
rect 10836 -2916 10964 -2884
rect 10996 -2916 11000 -2884
rect -720 -2920 11000 -2916
rect -720 -2964 -360 -2960
rect -720 -2996 -716 -2964
rect -684 -2996 -556 -2964
rect -524 -2996 -396 -2964
rect -364 -2996 -360 -2964
rect -720 -3000 -360 -2996
rect -320 -2964 11000 -2960
rect -320 -2996 -316 -2964
rect -284 -2996 -236 -2964
rect -204 -2996 -156 -2964
rect -124 -2996 -76 -2964
rect -44 -2996 4 -2964
rect 36 -2996 84 -2964
rect 116 -2996 164 -2964
rect 196 -2996 244 -2964
rect 276 -2996 324 -2964
rect 356 -2996 404 -2964
rect 436 -2996 484 -2964
rect 516 -2996 564 -2964
rect 596 -2996 644 -2964
rect 676 -2996 724 -2964
rect 756 -2996 804 -2964
rect 836 -2996 884 -2964
rect 916 -2996 964 -2964
rect 996 -2996 1044 -2964
rect 1076 -2996 1124 -2964
rect 1156 -2996 1204 -2964
rect 1236 -2996 1284 -2964
rect 1316 -2996 1364 -2964
rect 1396 -2996 1444 -2964
rect 1476 -2996 1524 -2964
rect 1556 -2996 1604 -2964
rect 1636 -2996 1684 -2964
rect 1716 -2996 1764 -2964
rect 1796 -2996 1844 -2964
rect 1876 -2996 1924 -2964
rect 1956 -2996 2004 -2964
rect 2036 -2996 2084 -2964
rect 2116 -2996 2164 -2964
rect 2196 -2996 2244 -2964
rect 2276 -2996 2324 -2964
rect 2356 -2996 2404 -2964
rect 2436 -2996 2484 -2964
rect 2516 -2996 2564 -2964
rect 2596 -2996 2644 -2964
rect 2676 -2996 2724 -2964
rect 2756 -2996 2804 -2964
rect 2836 -2996 2884 -2964
rect 2916 -2996 2964 -2964
rect 2996 -2996 3044 -2964
rect 3076 -2996 3124 -2964
rect 3156 -2996 3204 -2964
rect 3236 -2996 3284 -2964
rect 3316 -2996 3364 -2964
rect 3396 -2996 3444 -2964
rect 3476 -2996 3524 -2964
rect 3556 -2996 3604 -2964
rect 3636 -2996 3684 -2964
rect 3716 -2996 3764 -2964
rect 3796 -2996 3844 -2964
rect 3876 -2996 3924 -2964
rect 3956 -2996 4004 -2964
rect 4036 -2996 4084 -2964
rect 4116 -2996 4164 -2964
rect 4196 -2996 4244 -2964
rect 4276 -2996 4324 -2964
rect 4356 -2996 4404 -2964
rect 4436 -2996 4484 -2964
rect 4516 -2996 4564 -2964
rect 4596 -2996 4644 -2964
rect 4676 -2996 4724 -2964
rect 4756 -2996 4804 -2964
rect 4836 -2996 4884 -2964
rect 4916 -2996 4964 -2964
rect 4996 -2996 5044 -2964
rect 5076 -2996 5124 -2964
rect 5156 -2996 5204 -2964
rect 5236 -2996 5284 -2964
rect 5316 -2996 5364 -2964
rect 5396 -2996 5444 -2964
rect 5476 -2996 5524 -2964
rect 5556 -2996 5604 -2964
rect 5636 -2996 5684 -2964
rect 5716 -2996 5764 -2964
rect 5796 -2996 5844 -2964
rect 5876 -2996 5924 -2964
rect 5956 -2996 6004 -2964
rect 6036 -2996 6084 -2964
rect 6116 -2996 6164 -2964
rect 6196 -2996 6244 -2964
rect 6276 -2996 6324 -2964
rect 6356 -2996 6404 -2964
rect 6436 -2996 6484 -2964
rect 6516 -2996 6564 -2964
rect 6596 -2996 6644 -2964
rect 6676 -2996 6724 -2964
rect 6756 -2996 6804 -2964
rect 6836 -2996 6884 -2964
rect 6916 -2996 6964 -2964
rect 6996 -2996 7044 -2964
rect 7076 -2996 7124 -2964
rect 7156 -2996 7204 -2964
rect 7236 -2996 7284 -2964
rect 7316 -2996 7364 -2964
rect 7396 -2996 7444 -2964
rect 7476 -2996 7524 -2964
rect 7556 -2996 7604 -2964
rect 7636 -2996 7684 -2964
rect 7716 -2996 7764 -2964
rect 7796 -2996 7844 -2964
rect 7876 -2996 7924 -2964
rect 7956 -2996 8004 -2964
rect 8036 -2996 8084 -2964
rect 8116 -2996 8164 -2964
rect 8196 -2996 8244 -2964
rect 8276 -2996 8324 -2964
rect 8356 -2996 8404 -2964
rect 8436 -2996 8484 -2964
rect 8516 -2996 8564 -2964
rect 8596 -2996 8644 -2964
rect 8676 -2996 8724 -2964
rect 8756 -2996 8804 -2964
rect 8836 -2996 8884 -2964
rect 8916 -2996 8964 -2964
rect 8996 -2996 9044 -2964
rect 9076 -2996 9124 -2964
rect 9156 -2996 9204 -2964
rect 9236 -2996 9284 -2964
rect 9316 -2996 9364 -2964
rect 9396 -2996 9444 -2964
rect 9476 -2996 9524 -2964
rect 9556 -2996 9604 -2964
rect 9636 -2996 9684 -2964
rect 9716 -2996 9764 -2964
rect 9796 -2996 9844 -2964
rect 9876 -2996 9924 -2964
rect 9956 -2996 10004 -2964
rect 10036 -2996 10084 -2964
rect 10116 -2996 10164 -2964
rect 10196 -2996 10244 -2964
rect 10276 -2996 10324 -2964
rect 10356 -2996 10404 -2964
rect 10436 -2996 10484 -2964
rect 10516 -2996 10644 -2964
rect 10676 -2996 10804 -2964
rect 10836 -2996 10964 -2964
rect 10996 -2996 11000 -2964
rect -320 -3000 11000 -2996
rect -720 -3044 11000 -3040
rect -720 -3076 -716 -3044
rect -684 -3076 -556 -3044
rect -524 -3076 -396 -3044
rect -364 -3076 -316 -3044
rect -284 -3076 -236 -3044
rect -204 -3076 -156 -3044
rect -124 -3076 -76 -3044
rect -44 -3076 4 -3044
rect 36 -3076 84 -3044
rect 116 -3076 164 -3044
rect 196 -3076 244 -3044
rect 276 -3076 324 -3044
rect 356 -3076 404 -3044
rect 436 -3076 484 -3044
rect 516 -3076 564 -3044
rect 596 -3076 644 -3044
rect 676 -3076 724 -3044
rect 756 -3076 804 -3044
rect 836 -3076 884 -3044
rect 916 -3076 964 -3044
rect 996 -3076 1044 -3044
rect 1076 -3076 1124 -3044
rect 1156 -3076 1204 -3044
rect 1236 -3076 1284 -3044
rect 1316 -3076 1364 -3044
rect 1396 -3076 1444 -3044
rect 1476 -3076 1524 -3044
rect 1556 -3076 1604 -3044
rect 1636 -3076 1684 -3044
rect 1716 -3076 1764 -3044
rect 1796 -3076 1844 -3044
rect 1876 -3076 1924 -3044
rect 1956 -3076 2004 -3044
rect 2036 -3076 2084 -3044
rect 2116 -3076 2164 -3044
rect 2196 -3076 2244 -3044
rect 2276 -3076 2324 -3044
rect 2356 -3076 2404 -3044
rect 2436 -3076 2484 -3044
rect 2516 -3076 2564 -3044
rect 2596 -3076 2644 -3044
rect 2676 -3076 2724 -3044
rect 2756 -3076 2804 -3044
rect 2836 -3076 2884 -3044
rect 2916 -3076 2964 -3044
rect 2996 -3076 3044 -3044
rect 3076 -3076 3124 -3044
rect 3156 -3076 3204 -3044
rect 3236 -3076 3284 -3044
rect 3316 -3076 3364 -3044
rect 3396 -3076 3444 -3044
rect 3476 -3076 3524 -3044
rect 3556 -3076 3604 -3044
rect 3636 -3076 3684 -3044
rect 3716 -3076 3764 -3044
rect 3796 -3076 3844 -3044
rect 3876 -3076 3924 -3044
rect 3956 -3076 4004 -3044
rect 4036 -3076 4084 -3044
rect 4116 -3076 4164 -3044
rect 4196 -3076 4244 -3044
rect 4276 -3076 4324 -3044
rect 4356 -3076 4404 -3044
rect 4436 -3076 4484 -3044
rect 4516 -3076 4564 -3044
rect 4596 -3076 4644 -3044
rect 4676 -3076 4724 -3044
rect 4756 -3076 4804 -3044
rect 4836 -3076 4884 -3044
rect 4916 -3076 4964 -3044
rect 4996 -3076 5044 -3044
rect 5076 -3076 5124 -3044
rect 5156 -3076 5204 -3044
rect 5236 -3076 5284 -3044
rect 5316 -3076 5364 -3044
rect 5396 -3076 5444 -3044
rect 5476 -3076 5524 -3044
rect 5556 -3076 5604 -3044
rect 5636 -3076 5684 -3044
rect 5716 -3076 5764 -3044
rect 5796 -3076 5844 -3044
rect 5876 -3076 5924 -3044
rect 5956 -3076 6004 -3044
rect 6036 -3076 6084 -3044
rect 6116 -3076 6164 -3044
rect 6196 -3076 6244 -3044
rect 6276 -3076 6324 -3044
rect 6356 -3076 6404 -3044
rect 6436 -3076 6484 -3044
rect 6516 -3076 6564 -3044
rect 6596 -3076 6644 -3044
rect 6676 -3076 6724 -3044
rect 6756 -3076 6804 -3044
rect 6836 -3076 6884 -3044
rect 6916 -3076 6964 -3044
rect 6996 -3076 7044 -3044
rect 7076 -3076 7124 -3044
rect 7156 -3076 7204 -3044
rect 7236 -3076 7284 -3044
rect 7316 -3076 7364 -3044
rect 7396 -3076 7444 -3044
rect 7476 -3076 7524 -3044
rect 7556 -3076 7604 -3044
rect 7636 -3076 7684 -3044
rect 7716 -3076 7764 -3044
rect 7796 -3076 7844 -3044
rect 7876 -3076 7924 -3044
rect 7956 -3076 8004 -3044
rect 8036 -3076 8084 -3044
rect 8116 -3076 8164 -3044
rect 8196 -3076 8244 -3044
rect 8276 -3076 8324 -3044
rect 8356 -3076 8404 -3044
rect 8436 -3076 8484 -3044
rect 8516 -3076 8564 -3044
rect 8596 -3076 8644 -3044
rect 8676 -3076 8724 -3044
rect 8756 -3076 8804 -3044
rect 8836 -3076 8884 -3044
rect 8916 -3076 8964 -3044
rect 8996 -3076 9044 -3044
rect 9076 -3076 9124 -3044
rect 9156 -3076 9204 -3044
rect 9236 -3076 9284 -3044
rect 9316 -3076 9364 -3044
rect 9396 -3076 9444 -3044
rect 9476 -3076 9524 -3044
rect 9556 -3076 9604 -3044
rect 9636 -3076 9684 -3044
rect 9716 -3076 9764 -3044
rect 9796 -3076 9844 -3044
rect 9876 -3076 9924 -3044
rect 9956 -3076 10004 -3044
rect 10036 -3076 10084 -3044
rect 10116 -3076 10164 -3044
rect 10196 -3076 10244 -3044
rect 10276 -3076 10324 -3044
rect 10356 -3076 10404 -3044
rect 10436 -3076 10484 -3044
rect 10516 -3076 10644 -3044
rect 10676 -3076 10804 -3044
rect 10836 -3076 10964 -3044
rect 10996 -3076 11000 -3044
rect -720 -3080 11000 -3076
rect -720 -3124 10600 -3120
rect -720 -3156 -716 -3124
rect -684 -3156 -556 -3124
rect -524 -3156 -396 -3124
rect -364 -3156 -316 -3124
rect -284 -3156 -236 -3124
rect -204 -3156 -156 -3124
rect -124 -3156 -76 -3124
rect -44 -3156 4 -3124
rect 36 -3156 84 -3124
rect 116 -3156 164 -3124
rect 196 -3156 244 -3124
rect 276 -3156 324 -3124
rect 356 -3156 404 -3124
rect 436 -3156 484 -3124
rect 516 -3156 564 -3124
rect 596 -3156 644 -3124
rect 676 -3156 724 -3124
rect 756 -3156 804 -3124
rect 836 -3156 884 -3124
rect 916 -3156 964 -3124
rect 996 -3156 1044 -3124
rect 1076 -3156 1124 -3124
rect 1156 -3156 1204 -3124
rect 1236 -3156 1284 -3124
rect 1316 -3156 1364 -3124
rect 1396 -3156 1444 -3124
rect 1476 -3156 1524 -3124
rect 1556 -3156 1604 -3124
rect 1636 -3156 1684 -3124
rect 1716 -3156 1764 -3124
rect 1796 -3156 1844 -3124
rect 1876 -3156 1924 -3124
rect 1956 -3156 2004 -3124
rect 2036 -3156 2084 -3124
rect 2116 -3156 2164 -3124
rect 2196 -3156 2244 -3124
rect 2276 -3156 2324 -3124
rect 2356 -3156 2404 -3124
rect 2436 -3156 2484 -3124
rect 2516 -3156 2564 -3124
rect 2596 -3156 2644 -3124
rect 2676 -3156 2724 -3124
rect 2756 -3156 2804 -3124
rect 2836 -3156 2884 -3124
rect 2916 -3156 2964 -3124
rect 2996 -3156 3044 -3124
rect 3076 -3156 3124 -3124
rect 3156 -3156 3204 -3124
rect 3236 -3156 3284 -3124
rect 3316 -3156 3364 -3124
rect 3396 -3156 3444 -3124
rect 3476 -3156 3524 -3124
rect 3556 -3156 3604 -3124
rect 3636 -3156 3684 -3124
rect 3716 -3156 3764 -3124
rect 3796 -3156 3844 -3124
rect 3876 -3156 3924 -3124
rect 3956 -3156 4004 -3124
rect 4036 -3156 4084 -3124
rect 4116 -3156 4164 -3124
rect 4196 -3156 4244 -3124
rect 4276 -3156 4324 -3124
rect 4356 -3156 4404 -3124
rect 4436 -3156 4484 -3124
rect 4516 -3156 4564 -3124
rect 4596 -3156 4644 -3124
rect 4676 -3156 4724 -3124
rect 4756 -3156 4804 -3124
rect 4836 -3156 4884 -3124
rect 4916 -3156 4964 -3124
rect 4996 -3156 5044 -3124
rect 5076 -3156 5124 -3124
rect 5156 -3156 5204 -3124
rect 5236 -3156 5284 -3124
rect 5316 -3156 5364 -3124
rect 5396 -3156 5444 -3124
rect 5476 -3156 5524 -3124
rect 5556 -3156 5604 -3124
rect 5636 -3156 5684 -3124
rect 5716 -3156 5764 -3124
rect 5796 -3156 5844 -3124
rect 5876 -3156 5924 -3124
rect 5956 -3156 6004 -3124
rect 6036 -3156 6084 -3124
rect 6116 -3156 6164 -3124
rect 6196 -3156 6244 -3124
rect 6276 -3156 6324 -3124
rect 6356 -3156 6404 -3124
rect 6436 -3156 6484 -3124
rect 6516 -3156 6564 -3124
rect 6596 -3156 6644 -3124
rect 6676 -3156 6724 -3124
rect 6756 -3156 6804 -3124
rect 6836 -3156 6884 -3124
rect 6916 -3156 6964 -3124
rect 6996 -3156 7044 -3124
rect 7076 -3156 7124 -3124
rect 7156 -3156 7204 -3124
rect 7236 -3156 7284 -3124
rect 7316 -3156 7364 -3124
rect 7396 -3156 7444 -3124
rect 7476 -3156 7524 -3124
rect 7556 -3156 7604 -3124
rect 7636 -3156 7684 -3124
rect 7716 -3156 7764 -3124
rect 7796 -3156 7844 -3124
rect 7876 -3156 7924 -3124
rect 7956 -3156 8004 -3124
rect 8036 -3156 8084 -3124
rect 8116 -3156 8164 -3124
rect 8196 -3156 8244 -3124
rect 8276 -3156 8324 -3124
rect 8356 -3156 8404 -3124
rect 8436 -3156 8484 -3124
rect 8516 -3156 8564 -3124
rect 8596 -3156 8644 -3124
rect 8676 -3156 8724 -3124
rect 8756 -3156 8804 -3124
rect 8836 -3156 8884 -3124
rect 8916 -3156 8964 -3124
rect 8996 -3156 9044 -3124
rect 9076 -3156 9124 -3124
rect 9156 -3156 9204 -3124
rect 9236 -3156 9284 -3124
rect 9316 -3156 9364 -3124
rect 9396 -3156 9444 -3124
rect 9476 -3156 9524 -3124
rect 9556 -3156 9604 -3124
rect 9636 -3156 9684 -3124
rect 9716 -3156 9764 -3124
rect 9796 -3156 9844 -3124
rect 9876 -3156 9924 -3124
rect 9956 -3156 10004 -3124
rect 10036 -3156 10084 -3124
rect 10116 -3156 10164 -3124
rect 10196 -3156 10244 -3124
rect 10276 -3156 10324 -3124
rect 10356 -3156 10404 -3124
rect 10436 -3156 10484 -3124
rect 10516 -3156 10600 -3124
rect -720 -3160 10600 -3156
rect 10640 -3124 11000 -3120
rect 10640 -3156 10644 -3124
rect 10676 -3156 10804 -3124
rect 10836 -3156 10964 -3124
rect 10996 -3156 11000 -3124
rect 10640 -3160 11000 -3156
rect -720 -3204 11000 -3200
rect -720 -3236 -716 -3204
rect -684 -3236 -556 -3204
rect -524 -3236 -396 -3204
rect -364 -3236 -316 -3204
rect -284 -3236 -236 -3204
rect -204 -3236 -156 -3204
rect -124 -3236 -76 -3204
rect -44 -3236 4 -3204
rect 36 -3236 84 -3204
rect 116 -3236 164 -3204
rect 196 -3236 244 -3204
rect 276 -3236 324 -3204
rect 356 -3236 404 -3204
rect 436 -3236 484 -3204
rect 516 -3236 564 -3204
rect 596 -3236 644 -3204
rect 676 -3236 724 -3204
rect 756 -3236 804 -3204
rect 836 -3236 884 -3204
rect 916 -3236 964 -3204
rect 996 -3236 1044 -3204
rect 1076 -3236 1124 -3204
rect 1156 -3236 1204 -3204
rect 1236 -3236 1284 -3204
rect 1316 -3236 1364 -3204
rect 1396 -3236 1444 -3204
rect 1476 -3236 1524 -3204
rect 1556 -3236 1604 -3204
rect 1636 -3236 1684 -3204
rect 1716 -3236 1764 -3204
rect 1796 -3236 1844 -3204
rect 1876 -3236 1924 -3204
rect 1956 -3236 2004 -3204
rect 2036 -3236 2084 -3204
rect 2116 -3236 2164 -3204
rect 2196 -3236 2244 -3204
rect 2276 -3236 2324 -3204
rect 2356 -3236 2404 -3204
rect 2436 -3236 2484 -3204
rect 2516 -3236 2564 -3204
rect 2596 -3236 2644 -3204
rect 2676 -3236 2724 -3204
rect 2756 -3236 2804 -3204
rect 2836 -3236 2884 -3204
rect 2916 -3236 2964 -3204
rect 2996 -3236 3044 -3204
rect 3076 -3236 3124 -3204
rect 3156 -3236 3204 -3204
rect 3236 -3236 3284 -3204
rect 3316 -3236 3364 -3204
rect 3396 -3236 3444 -3204
rect 3476 -3236 3524 -3204
rect 3556 -3236 3604 -3204
rect 3636 -3236 3684 -3204
rect 3716 -3236 3764 -3204
rect 3796 -3236 3844 -3204
rect 3876 -3236 3924 -3204
rect 3956 -3236 4004 -3204
rect 4036 -3236 4084 -3204
rect 4116 -3236 4164 -3204
rect 4196 -3236 4244 -3204
rect 4276 -3236 4324 -3204
rect 4356 -3236 4404 -3204
rect 4436 -3236 4484 -3204
rect 4516 -3236 4564 -3204
rect 4596 -3236 4644 -3204
rect 4676 -3236 4724 -3204
rect 4756 -3236 4804 -3204
rect 4836 -3236 4884 -3204
rect 4916 -3236 4964 -3204
rect 4996 -3236 5044 -3204
rect 5076 -3236 5124 -3204
rect 5156 -3236 5204 -3204
rect 5236 -3236 5284 -3204
rect 5316 -3236 5364 -3204
rect 5396 -3236 5444 -3204
rect 5476 -3236 5524 -3204
rect 5556 -3236 5604 -3204
rect 5636 -3236 5684 -3204
rect 5716 -3236 5764 -3204
rect 5796 -3236 5844 -3204
rect 5876 -3236 5924 -3204
rect 5956 -3236 6004 -3204
rect 6036 -3236 6084 -3204
rect 6116 -3236 6164 -3204
rect 6196 -3236 6244 -3204
rect 6276 -3236 6324 -3204
rect 6356 -3236 6404 -3204
rect 6436 -3236 6484 -3204
rect 6516 -3236 6564 -3204
rect 6596 -3236 6644 -3204
rect 6676 -3236 6724 -3204
rect 6756 -3236 6804 -3204
rect 6836 -3236 6884 -3204
rect 6916 -3236 6964 -3204
rect 6996 -3236 7044 -3204
rect 7076 -3236 7124 -3204
rect 7156 -3236 7204 -3204
rect 7236 -3236 7284 -3204
rect 7316 -3236 7364 -3204
rect 7396 -3236 7444 -3204
rect 7476 -3236 7524 -3204
rect 7556 -3236 7604 -3204
rect 7636 -3236 7684 -3204
rect 7716 -3236 7764 -3204
rect 7796 -3236 7844 -3204
rect 7876 -3236 7924 -3204
rect 7956 -3236 8004 -3204
rect 8036 -3236 8084 -3204
rect 8116 -3236 8164 -3204
rect 8196 -3236 8244 -3204
rect 8276 -3236 8324 -3204
rect 8356 -3236 8404 -3204
rect 8436 -3236 8484 -3204
rect 8516 -3236 8564 -3204
rect 8596 -3236 8644 -3204
rect 8676 -3236 8724 -3204
rect 8756 -3236 8804 -3204
rect 8836 -3236 8884 -3204
rect 8916 -3236 8964 -3204
rect 8996 -3236 9044 -3204
rect 9076 -3236 9124 -3204
rect 9156 -3236 9204 -3204
rect 9236 -3236 9284 -3204
rect 9316 -3236 9364 -3204
rect 9396 -3236 9444 -3204
rect 9476 -3236 9524 -3204
rect 9556 -3236 9604 -3204
rect 9636 -3236 9684 -3204
rect 9716 -3236 9764 -3204
rect 9796 -3236 9844 -3204
rect 9876 -3236 9924 -3204
rect 9956 -3236 10004 -3204
rect 10036 -3236 10084 -3204
rect 10116 -3236 10164 -3204
rect 10196 -3236 10244 -3204
rect 10276 -3236 10324 -3204
rect 10356 -3236 10404 -3204
rect 10436 -3236 10484 -3204
rect 10516 -3236 10644 -3204
rect 10676 -3236 10804 -3204
rect 10836 -3236 10964 -3204
rect 10996 -3236 11000 -3204
rect -720 -3240 11000 -3236
rect -720 -3284 11000 -3280
rect -720 -3316 -716 -3284
rect -684 -3316 -556 -3284
rect -524 -3316 -396 -3284
rect -364 -3316 -316 -3284
rect -284 -3316 -236 -3284
rect -204 -3316 -156 -3284
rect -124 -3316 -76 -3284
rect -44 -3316 4 -3284
rect 36 -3316 84 -3284
rect 116 -3316 164 -3284
rect 196 -3316 244 -3284
rect 276 -3316 324 -3284
rect 356 -3316 404 -3284
rect 436 -3316 484 -3284
rect 516 -3316 564 -3284
rect 596 -3316 644 -3284
rect 676 -3316 724 -3284
rect 756 -3316 804 -3284
rect 836 -3316 884 -3284
rect 916 -3316 964 -3284
rect 996 -3316 1044 -3284
rect 1076 -3316 1124 -3284
rect 1156 -3316 1204 -3284
rect 1236 -3316 1284 -3284
rect 1316 -3316 1364 -3284
rect 1396 -3316 1444 -3284
rect 1476 -3316 1524 -3284
rect 1556 -3316 1604 -3284
rect 1636 -3316 1684 -3284
rect 1716 -3316 1764 -3284
rect 1796 -3316 1844 -3284
rect 1876 -3316 1924 -3284
rect 1956 -3316 2004 -3284
rect 2036 -3316 2084 -3284
rect 2116 -3316 2164 -3284
rect 2196 -3316 2244 -3284
rect 2276 -3316 2324 -3284
rect 2356 -3316 2404 -3284
rect 2436 -3316 2484 -3284
rect 2516 -3316 2564 -3284
rect 2596 -3316 2644 -3284
rect 2676 -3316 2724 -3284
rect 2756 -3316 2804 -3284
rect 2836 -3316 2884 -3284
rect 2916 -3316 2964 -3284
rect 2996 -3316 3044 -3284
rect 3076 -3316 3124 -3284
rect 3156 -3316 3204 -3284
rect 3236 -3316 3284 -3284
rect 3316 -3316 3364 -3284
rect 3396 -3316 3444 -3284
rect 3476 -3316 3524 -3284
rect 3556 -3316 3604 -3284
rect 3636 -3316 3684 -3284
rect 3716 -3316 3764 -3284
rect 3796 -3316 3844 -3284
rect 3876 -3316 3924 -3284
rect 3956 -3316 4004 -3284
rect 4036 -3316 4084 -3284
rect 4116 -3316 4164 -3284
rect 4196 -3316 4244 -3284
rect 4276 -3316 4324 -3284
rect 4356 -3316 4404 -3284
rect 4436 -3316 4484 -3284
rect 4516 -3316 4564 -3284
rect 4596 -3316 4644 -3284
rect 4676 -3316 4724 -3284
rect 4756 -3316 4804 -3284
rect 4836 -3316 4884 -3284
rect 4916 -3316 4964 -3284
rect 4996 -3316 5044 -3284
rect 5076 -3316 5124 -3284
rect 5156 -3316 5204 -3284
rect 5236 -3316 5284 -3284
rect 5316 -3316 5364 -3284
rect 5396 -3316 5444 -3284
rect 5476 -3316 5524 -3284
rect 5556 -3316 5604 -3284
rect 5636 -3316 5684 -3284
rect 5716 -3316 5764 -3284
rect 5796 -3316 5844 -3284
rect 5876 -3316 5924 -3284
rect 5956 -3316 6004 -3284
rect 6036 -3316 6084 -3284
rect 6116 -3316 6164 -3284
rect 6196 -3316 6244 -3284
rect 6276 -3316 6324 -3284
rect 6356 -3316 6404 -3284
rect 6436 -3316 6484 -3284
rect 6516 -3316 6564 -3284
rect 6596 -3316 6644 -3284
rect 6676 -3316 6724 -3284
rect 6756 -3316 6804 -3284
rect 6836 -3316 6884 -3284
rect 6916 -3316 6964 -3284
rect 6996 -3316 7044 -3284
rect 7076 -3316 7124 -3284
rect 7156 -3316 7204 -3284
rect 7236 -3316 7284 -3284
rect 7316 -3316 7364 -3284
rect 7396 -3316 7444 -3284
rect 7476 -3316 7524 -3284
rect 7556 -3316 7604 -3284
rect 7636 -3316 7684 -3284
rect 7716 -3316 7764 -3284
rect 7796 -3316 7844 -3284
rect 7876 -3316 7924 -3284
rect 7956 -3316 8004 -3284
rect 8036 -3316 8084 -3284
rect 8116 -3316 8164 -3284
rect 8196 -3316 8244 -3284
rect 8276 -3316 8324 -3284
rect 8356 -3316 8404 -3284
rect 8436 -3316 8484 -3284
rect 8516 -3316 8564 -3284
rect 8596 -3316 8644 -3284
rect 8676 -3316 8724 -3284
rect 8756 -3316 8804 -3284
rect 8836 -3316 8884 -3284
rect 8916 -3316 8964 -3284
rect 8996 -3316 9044 -3284
rect 9076 -3316 9124 -3284
rect 9156 -3316 9204 -3284
rect 9236 -3316 9284 -3284
rect 9316 -3316 9364 -3284
rect 9396 -3316 9444 -3284
rect 9476 -3316 9524 -3284
rect 9556 -3316 9604 -3284
rect 9636 -3316 9684 -3284
rect 9716 -3316 9764 -3284
rect 9796 -3316 9844 -3284
rect 9876 -3316 9924 -3284
rect 9956 -3316 10004 -3284
rect 10036 -3316 10084 -3284
rect 10116 -3316 10164 -3284
rect 10196 -3316 10244 -3284
rect 10276 -3316 10324 -3284
rect 10356 -3316 10404 -3284
rect 10436 -3316 10484 -3284
rect 10516 -3316 10644 -3284
rect 10676 -3316 10804 -3284
rect 10836 -3316 10964 -3284
rect 10996 -3316 11000 -3284
rect -720 -3320 11000 -3316
rect -720 -3364 10600 -3360
rect -720 -3396 -716 -3364
rect -684 -3396 -556 -3364
rect -524 -3396 -396 -3364
rect -364 -3396 -316 -3364
rect -284 -3396 -236 -3364
rect -204 -3396 -156 -3364
rect -124 -3396 -76 -3364
rect -44 -3396 4 -3364
rect 36 -3396 84 -3364
rect 116 -3396 164 -3364
rect 196 -3396 244 -3364
rect 276 -3396 324 -3364
rect 356 -3396 404 -3364
rect 436 -3396 484 -3364
rect 516 -3396 564 -3364
rect 596 -3396 644 -3364
rect 676 -3396 724 -3364
rect 756 -3396 804 -3364
rect 836 -3396 884 -3364
rect 916 -3396 964 -3364
rect 996 -3396 1044 -3364
rect 1076 -3396 1124 -3364
rect 1156 -3396 1204 -3364
rect 1236 -3396 1284 -3364
rect 1316 -3396 1364 -3364
rect 1396 -3396 1444 -3364
rect 1476 -3396 1524 -3364
rect 1556 -3396 1604 -3364
rect 1636 -3396 1684 -3364
rect 1716 -3396 1764 -3364
rect 1796 -3396 1844 -3364
rect 1876 -3396 1924 -3364
rect 1956 -3396 2004 -3364
rect 2036 -3396 2084 -3364
rect 2116 -3396 2164 -3364
rect 2196 -3396 2244 -3364
rect 2276 -3396 2324 -3364
rect 2356 -3396 2404 -3364
rect 2436 -3396 2484 -3364
rect 2516 -3396 2564 -3364
rect 2596 -3396 2644 -3364
rect 2676 -3396 2724 -3364
rect 2756 -3396 2804 -3364
rect 2836 -3396 2884 -3364
rect 2916 -3396 2964 -3364
rect 2996 -3396 3044 -3364
rect 3076 -3396 3124 -3364
rect 3156 -3396 3204 -3364
rect 3236 -3396 3284 -3364
rect 3316 -3396 3364 -3364
rect 3396 -3396 3444 -3364
rect 3476 -3396 3524 -3364
rect 3556 -3396 3604 -3364
rect 3636 -3396 3684 -3364
rect 3716 -3396 3764 -3364
rect 3796 -3396 3844 -3364
rect 3876 -3396 3924 -3364
rect 3956 -3396 4004 -3364
rect 4036 -3396 4084 -3364
rect 4116 -3396 4164 -3364
rect 4196 -3396 4244 -3364
rect 4276 -3396 4324 -3364
rect 4356 -3396 4404 -3364
rect 4436 -3396 4484 -3364
rect 4516 -3396 4564 -3364
rect 4596 -3396 4644 -3364
rect 4676 -3396 4724 -3364
rect 4756 -3396 4804 -3364
rect 4836 -3396 4884 -3364
rect 4916 -3396 4964 -3364
rect 4996 -3396 5044 -3364
rect 5076 -3396 5124 -3364
rect 5156 -3396 5204 -3364
rect 5236 -3396 5284 -3364
rect 5316 -3396 5364 -3364
rect 5396 -3396 5444 -3364
rect 5476 -3396 5524 -3364
rect 5556 -3396 5604 -3364
rect 5636 -3396 5684 -3364
rect 5716 -3396 5764 -3364
rect 5796 -3396 5844 -3364
rect 5876 -3396 5924 -3364
rect 5956 -3396 6004 -3364
rect 6036 -3396 6084 -3364
rect 6116 -3396 6164 -3364
rect 6196 -3396 6244 -3364
rect 6276 -3396 6324 -3364
rect 6356 -3396 6404 -3364
rect 6436 -3396 6484 -3364
rect 6516 -3396 6564 -3364
rect 6596 -3396 6644 -3364
rect 6676 -3396 6724 -3364
rect 6756 -3396 6804 -3364
rect 6836 -3396 6884 -3364
rect 6916 -3396 6964 -3364
rect 6996 -3396 7044 -3364
rect 7076 -3396 7124 -3364
rect 7156 -3396 7204 -3364
rect 7236 -3396 7284 -3364
rect 7316 -3396 7364 -3364
rect 7396 -3396 7444 -3364
rect 7476 -3396 7524 -3364
rect 7556 -3396 7604 -3364
rect 7636 -3396 7684 -3364
rect 7716 -3396 7764 -3364
rect 7796 -3396 7844 -3364
rect 7876 -3396 7924 -3364
rect 7956 -3396 8004 -3364
rect 8036 -3396 8084 -3364
rect 8116 -3396 8164 -3364
rect 8196 -3396 8244 -3364
rect 8276 -3396 8324 -3364
rect 8356 -3396 8404 -3364
rect 8436 -3396 8484 -3364
rect 8516 -3396 8564 -3364
rect 8596 -3396 8644 -3364
rect 8676 -3396 8724 -3364
rect 8756 -3396 8804 -3364
rect 8836 -3396 8884 -3364
rect 8916 -3396 8964 -3364
rect 8996 -3396 9044 -3364
rect 9076 -3396 9124 -3364
rect 9156 -3396 9204 -3364
rect 9236 -3396 9284 -3364
rect 9316 -3396 9364 -3364
rect 9396 -3396 9444 -3364
rect 9476 -3396 9524 -3364
rect 9556 -3396 9604 -3364
rect 9636 -3396 9684 -3364
rect 9716 -3396 9764 -3364
rect 9796 -3396 9844 -3364
rect 9876 -3396 9924 -3364
rect 9956 -3396 10004 -3364
rect 10036 -3396 10084 -3364
rect 10116 -3396 10164 -3364
rect 10196 -3396 10244 -3364
rect 10276 -3396 10324 -3364
rect 10356 -3396 10404 -3364
rect 10436 -3396 10484 -3364
rect 10516 -3396 10600 -3364
rect -720 -3400 10600 -3396
rect 10640 -3364 11000 -3360
rect 10640 -3396 10644 -3364
rect 10676 -3396 10804 -3364
rect 10836 -3396 10964 -3364
rect 10996 -3396 11000 -3364
rect 10640 -3400 11000 -3396
rect -720 -3444 10600 -3440
rect -720 -3476 -716 -3444
rect -684 -3476 -556 -3444
rect -524 -3476 -396 -3444
rect -364 -3476 -316 -3444
rect -284 -3476 -236 -3444
rect -204 -3476 -156 -3444
rect -124 -3476 -76 -3444
rect -44 -3476 4 -3444
rect 36 -3476 84 -3444
rect 116 -3476 164 -3444
rect 196 -3476 244 -3444
rect 276 -3476 324 -3444
rect 356 -3476 404 -3444
rect 436 -3476 484 -3444
rect 516 -3476 564 -3444
rect 596 -3476 644 -3444
rect 676 -3476 724 -3444
rect 756 -3476 804 -3444
rect 836 -3476 884 -3444
rect 916 -3476 964 -3444
rect 996 -3476 1044 -3444
rect 1076 -3476 1124 -3444
rect 1156 -3476 1204 -3444
rect 1236 -3476 1284 -3444
rect 1316 -3476 1364 -3444
rect 1396 -3476 1444 -3444
rect 1476 -3476 1524 -3444
rect 1556 -3476 1604 -3444
rect 1636 -3476 1684 -3444
rect 1716 -3476 1764 -3444
rect 1796 -3476 1844 -3444
rect 1876 -3476 1924 -3444
rect 1956 -3476 2004 -3444
rect 2036 -3476 2084 -3444
rect 2116 -3476 2164 -3444
rect 2196 -3476 2244 -3444
rect 2276 -3476 2324 -3444
rect 2356 -3476 2404 -3444
rect 2436 -3476 2484 -3444
rect 2516 -3476 2564 -3444
rect 2596 -3476 2644 -3444
rect 2676 -3476 2724 -3444
rect 2756 -3476 2804 -3444
rect 2836 -3476 2884 -3444
rect 2916 -3476 2964 -3444
rect 2996 -3476 3044 -3444
rect 3076 -3476 3124 -3444
rect 3156 -3476 3204 -3444
rect 3236 -3476 3284 -3444
rect 3316 -3476 3364 -3444
rect 3396 -3476 3444 -3444
rect 3476 -3476 3524 -3444
rect 3556 -3476 3604 -3444
rect 3636 -3476 3684 -3444
rect 3716 -3476 3764 -3444
rect 3796 -3476 3844 -3444
rect 3876 -3476 3924 -3444
rect 3956 -3476 4004 -3444
rect 4036 -3476 4084 -3444
rect 4116 -3476 4164 -3444
rect 4196 -3476 4244 -3444
rect 4276 -3476 4324 -3444
rect 4356 -3476 4404 -3444
rect 4436 -3476 4484 -3444
rect 4516 -3476 4564 -3444
rect 4596 -3476 4644 -3444
rect 4676 -3476 4724 -3444
rect 4756 -3476 4804 -3444
rect 4836 -3476 4884 -3444
rect 4916 -3476 4964 -3444
rect 4996 -3476 5044 -3444
rect 5076 -3476 5124 -3444
rect 5156 -3476 5204 -3444
rect 5236 -3476 5284 -3444
rect 5316 -3476 5364 -3444
rect 5396 -3476 5444 -3444
rect 5476 -3476 5524 -3444
rect 5556 -3476 5604 -3444
rect 5636 -3476 5684 -3444
rect 5716 -3476 5764 -3444
rect 5796 -3476 5844 -3444
rect 5876 -3476 5924 -3444
rect 5956 -3476 6004 -3444
rect 6036 -3476 6084 -3444
rect 6116 -3476 6164 -3444
rect 6196 -3476 6244 -3444
rect 6276 -3476 6324 -3444
rect 6356 -3476 6404 -3444
rect 6436 -3476 6484 -3444
rect 6516 -3476 6564 -3444
rect 6596 -3476 6644 -3444
rect 6676 -3476 6724 -3444
rect 6756 -3476 6804 -3444
rect 6836 -3476 6884 -3444
rect 6916 -3476 6964 -3444
rect 6996 -3476 7044 -3444
rect 7076 -3476 7124 -3444
rect 7156 -3476 7204 -3444
rect 7236 -3476 7284 -3444
rect 7316 -3476 7364 -3444
rect 7396 -3476 7444 -3444
rect 7476 -3476 7524 -3444
rect 7556 -3476 7604 -3444
rect 7636 -3476 7684 -3444
rect 7716 -3476 7764 -3444
rect 7796 -3476 7844 -3444
rect 7876 -3476 7924 -3444
rect 7956 -3476 8004 -3444
rect 8036 -3476 8084 -3444
rect 8116 -3476 8164 -3444
rect 8196 -3476 8244 -3444
rect 8276 -3476 8324 -3444
rect 8356 -3476 8404 -3444
rect 8436 -3476 8484 -3444
rect 8516 -3476 8564 -3444
rect 8596 -3476 8644 -3444
rect 8676 -3476 8724 -3444
rect 8756 -3476 8804 -3444
rect 8836 -3476 8884 -3444
rect 8916 -3476 8964 -3444
rect 8996 -3476 9044 -3444
rect 9076 -3476 9124 -3444
rect 9156 -3476 9204 -3444
rect 9236 -3476 9284 -3444
rect 9316 -3476 9364 -3444
rect 9396 -3476 9444 -3444
rect 9476 -3476 9524 -3444
rect 9556 -3476 9604 -3444
rect 9636 -3476 9684 -3444
rect 9716 -3476 9764 -3444
rect 9796 -3476 9844 -3444
rect 9876 -3476 9924 -3444
rect 9956 -3476 10004 -3444
rect 10036 -3476 10084 -3444
rect 10116 -3476 10164 -3444
rect 10196 -3476 10244 -3444
rect 10276 -3476 10324 -3444
rect 10356 -3476 10404 -3444
rect 10436 -3476 10484 -3444
rect 10516 -3476 10600 -3444
rect -720 -3480 10600 -3476
rect 10640 -3444 11000 -3440
rect 10640 -3476 10644 -3444
rect 10676 -3476 10804 -3444
rect 10836 -3476 10964 -3444
rect 10996 -3476 11000 -3444
rect 10640 -3480 11000 -3476
rect -720 -3524 11000 -3520
rect -720 -3556 -716 -3524
rect -684 -3556 -556 -3524
rect -524 -3556 -396 -3524
rect -364 -3556 -316 -3524
rect -284 -3556 -236 -3524
rect -204 -3556 -156 -3524
rect -124 -3556 -76 -3524
rect -44 -3556 4 -3524
rect 36 -3556 84 -3524
rect 116 -3556 164 -3524
rect 196 -3556 244 -3524
rect 276 -3556 324 -3524
rect 356 -3556 404 -3524
rect 436 -3556 484 -3524
rect 516 -3556 564 -3524
rect 596 -3556 644 -3524
rect 676 -3556 724 -3524
rect 756 -3556 804 -3524
rect 836 -3556 884 -3524
rect 916 -3556 964 -3524
rect 996 -3556 1044 -3524
rect 1076 -3556 1124 -3524
rect 1156 -3556 1204 -3524
rect 1236 -3556 1284 -3524
rect 1316 -3556 1364 -3524
rect 1396 -3556 1444 -3524
rect 1476 -3556 1524 -3524
rect 1556 -3556 1604 -3524
rect 1636 -3556 1684 -3524
rect 1716 -3556 1764 -3524
rect 1796 -3556 1844 -3524
rect 1876 -3556 1924 -3524
rect 1956 -3556 2004 -3524
rect 2036 -3556 2084 -3524
rect 2116 -3556 2164 -3524
rect 2196 -3556 2244 -3524
rect 2276 -3556 2324 -3524
rect 2356 -3556 2404 -3524
rect 2436 -3556 2484 -3524
rect 2516 -3556 2564 -3524
rect 2596 -3556 2644 -3524
rect 2676 -3556 2724 -3524
rect 2756 -3556 2804 -3524
rect 2836 -3556 2884 -3524
rect 2916 -3556 2964 -3524
rect 2996 -3556 3044 -3524
rect 3076 -3556 3124 -3524
rect 3156 -3556 3204 -3524
rect 3236 -3556 3284 -3524
rect 3316 -3556 3364 -3524
rect 3396 -3556 3444 -3524
rect 3476 -3556 3524 -3524
rect 3556 -3556 3604 -3524
rect 3636 -3556 3684 -3524
rect 3716 -3556 3764 -3524
rect 3796 -3556 3844 -3524
rect 3876 -3556 3924 -3524
rect 3956 -3556 4004 -3524
rect 4036 -3556 4084 -3524
rect 4116 -3556 4164 -3524
rect 4196 -3556 4244 -3524
rect 4276 -3556 4324 -3524
rect 4356 -3556 4404 -3524
rect 4436 -3556 4484 -3524
rect 4516 -3556 4564 -3524
rect 4596 -3556 4644 -3524
rect 4676 -3556 4724 -3524
rect 4756 -3556 4804 -3524
rect 4836 -3556 4884 -3524
rect 4916 -3556 4964 -3524
rect 4996 -3556 5044 -3524
rect 5076 -3556 5124 -3524
rect 5156 -3556 5204 -3524
rect 5236 -3556 5284 -3524
rect 5316 -3556 5364 -3524
rect 5396 -3556 5444 -3524
rect 5476 -3556 5524 -3524
rect 5556 -3556 5604 -3524
rect 5636 -3556 5684 -3524
rect 5716 -3556 5764 -3524
rect 5796 -3556 5844 -3524
rect 5876 -3556 5924 -3524
rect 5956 -3556 6004 -3524
rect 6036 -3556 6084 -3524
rect 6116 -3556 6164 -3524
rect 6196 -3556 6244 -3524
rect 6276 -3556 6324 -3524
rect 6356 -3556 6404 -3524
rect 6436 -3556 6484 -3524
rect 6516 -3556 6564 -3524
rect 6596 -3556 6644 -3524
rect 6676 -3556 6724 -3524
rect 6756 -3556 6804 -3524
rect 6836 -3556 6884 -3524
rect 6916 -3556 6964 -3524
rect 6996 -3556 7044 -3524
rect 7076 -3556 7124 -3524
rect 7156 -3556 7204 -3524
rect 7236 -3556 7284 -3524
rect 7316 -3556 7364 -3524
rect 7396 -3556 7444 -3524
rect 7476 -3556 7524 -3524
rect 7556 -3556 7604 -3524
rect 7636 -3556 7684 -3524
rect 7716 -3556 7764 -3524
rect 7796 -3556 7844 -3524
rect 7876 -3556 7924 -3524
rect 7956 -3556 8004 -3524
rect 8036 -3556 8084 -3524
rect 8116 -3556 8164 -3524
rect 8196 -3556 8244 -3524
rect 8276 -3556 8324 -3524
rect 8356 -3556 8404 -3524
rect 8436 -3556 8484 -3524
rect 8516 -3556 8564 -3524
rect 8596 -3556 8644 -3524
rect 8676 -3556 8724 -3524
rect 8756 -3556 8804 -3524
rect 8836 -3556 8884 -3524
rect 8916 -3556 8964 -3524
rect 8996 -3556 9044 -3524
rect 9076 -3556 9124 -3524
rect 9156 -3556 9204 -3524
rect 9236 -3556 9284 -3524
rect 9316 -3556 9364 -3524
rect 9396 -3556 9444 -3524
rect 9476 -3556 9524 -3524
rect 9556 -3556 9604 -3524
rect 9636 -3556 9684 -3524
rect 9716 -3556 9764 -3524
rect 9796 -3556 9844 -3524
rect 9876 -3556 9924 -3524
rect 9956 -3556 10004 -3524
rect 10036 -3556 10084 -3524
rect 10116 -3556 10164 -3524
rect 10196 -3556 10244 -3524
rect 10276 -3556 10324 -3524
rect 10356 -3556 10404 -3524
rect 10436 -3556 10484 -3524
rect 10516 -3556 10644 -3524
rect 10676 -3556 10804 -3524
rect 10836 -3556 10964 -3524
rect 10996 -3556 11000 -3524
rect -720 -3560 11000 -3556
rect -720 -3604 11000 -3600
rect -720 -3636 -716 -3604
rect -684 -3636 -556 -3604
rect -524 -3636 -396 -3604
rect -364 -3636 -316 -3604
rect -284 -3636 -236 -3604
rect -204 -3636 -156 -3604
rect -124 -3636 -76 -3604
rect -44 -3636 4 -3604
rect 36 -3636 84 -3604
rect 116 -3636 164 -3604
rect 196 -3636 244 -3604
rect 276 -3636 324 -3604
rect 356 -3636 404 -3604
rect 436 -3636 484 -3604
rect 516 -3636 564 -3604
rect 596 -3636 644 -3604
rect 676 -3636 724 -3604
rect 756 -3636 804 -3604
rect 836 -3636 884 -3604
rect 916 -3636 964 -3604
rect 996 -3636 1044 -3604
rect 1076 -3636 1124 -3604
rect 1156 -3636 1204 -3604
rect 1236 -3636 1284 -3604
rect 1316 -3636 1364 -3604
rect 1396 -3636 1444 -3604
rect 1476 -3636 1524 -3604
rect 1556 -3636 1604 -3604
rect 1636 -3636 1684 -3604
rect 1716 -3636 1764 -3604
rect 1796 -3636 1844 -3604
rect 1876 -3636 1924 -3604
rect 1956 -3636 2004 -3604
rect 2036 -3636 2084 -3604
rect 2116 -3636 2164 -3604
rect 2196 -3636 2244 -3604
rect 2276 -3636 2324 -3604
rect 2356 -3636 2404 -3604
rect 2436 -3636 2484 -3604
rect 2516 -3636 2564 -3604
rect 2596 -3636 2644 -3604
rect 2676 -3636 2724 -3604
rect 2756 -3636 2804 -3604
rect 2836 -3636 2884 -3604
rect 2916 -3636 2964 -3604
rect 2996 -3636 3044 -3604
rect 3076 -3636 3124 -3604
rect 3156 -3636 3204 -3604
rect 3236 -3636 3284 -3604
rect 3316 -3636 3364 -3604
rect 3396 -3636 3444 -3604
rect 3476 -3636 3524 -3604
rect 3556 -3636 3604 -3604
rect 3636 -3636 3684 -3604
rect 3716 -3636 3764 -3604
rect 3796 -3636 3844 -3604
rect 3876 -3636 3924 -3604
rect 3956 -3636 4004 -3604
rect 4036 -3636 4084 -3604
rect 4116 -3636 4164 -3604
rect 4196 -3636 4244 -3604
rect 4276 -3636 4324 -3604
rect 4356 -3636 4404 -3604
rect 4436 -3636 4484 -3604
rect 4516 -3636 4564 -3604
rect 4596 -3636 4644 -3604
rect 4676 -3636 4724 -3604
rect 4756 -3636 4804 -3604
rect 4836 -3636 4884 -3604
rect 4916 -3636 4964 -3604
rect 4996 -3636 5044 -3604
rect 5076 -3636 5124 -3604
rect 5156 -3636 5204 -3604
rect 5236 -3636 5284 -3604
rect 5316 -3636 5364 -3604
rect 5396 -3636 5444 -3604
rect 5476 -3636 5524 -3604
rect 5556 -3636 5604 -3604
rect 5636 -3636 5684 -3604
rect 5716 -3636 5764 -3604
rect 5796 -3636 5844 -3604
rect 5876 -3636 5924 -3604
rect 5956 -3636 6004 -3604
rect 6036 -3636 6084 -3604
rect 6116 -3636 6164 -3604
rect 6196 -3636 6244 -3604
rect 6276 -3636 6324 -3604
rect 6356 -3636 6404 -3604
rect 6436 -3636 6484 -3604
rect 6516 -3636 6564 -3604
rect 6596 -3636 6644 -3604
rect 6676 -3636 6724 -3604
rect 6756 -3636 6804 -3604
rect 6836 -3636 6884 -3604
rect 6916 -3636 6964 -3604
rect 6996 -3636 7044 -3604
rect 7076 -3636 7124 -3604
rect 7156 -3636 7204 -3604
rect 7236 -3636 7284 -3604
rect 7316 -3636 7364 -3604
rect 7396 -3636 7444 -3604
rect 7476 -3636 7524 -3604
rect 7556 -3636 7604 -3604
rect 7636 -3636 7684 -3604
rect 7716 -3636 7764 -3604
rect 7796 -3636 7844 -3604
rect 7876 -3636 7924 -3604
rect 7956 -3636 8004 -3604
rect 8036 -3636 8084 -3604
rect 8116 -3636 8164 -3604
rect 8196 -3636 8244 -3604
rect 8276 -3636 8324 -3604
rect 8356 -3636 8404 -3604
rect 8436 -3636 8484 -3604
rect 8516 -3636 8564 -3604
rect 8596 -3636 8644 -3604
rect 8676 -3636 8724 -3604
rect 8756 -3636 8804 -3604
rect 8836 -3636 8884 -3604
rect 8916 -3636 8964 -3604
rect 8996 -3636 9044 -3604
rect 9076 -3636 9124 -3604
rect 9156 -3636 9204 -3604
rect 9236 -3636 9284 -3604
rect 9316 -3636 9364 -3604
rect 9396 -3636 9444 -3604
rect 9476 -3636 9524 -3604
rect 9556 -3636 9604 -3604
rect 9636 -3636 9684 -3604
rect 9716 -3636 9764 -3604
rect 9796 -3636 9844 -3604
rect 9876 -3636 9924 -3604
rect 9956 -3636 10004 -3604
rect 10036 -3636 10084 -3604
rect 10116 -3636 10164 -3604
rect 10196 -3636 10244 -3604
rect 10276 -3636 10324 -3604
rect 10356 -3636 10404 -3604
rect 10436 -3636 10484 -3604
rect 10516 -3636 10644 -3604
rect 10676 -3636 10804 -3604
rect 10836 -3636 10964 -3604
rect 10996 -3636 11000 -3604
rect -720 -3640 11000 -3636
rect -720 -3684 11000 -3680
rect -720 -3716 -716 -3684
rect -684 -3716 -556 -3684
rect -524 -3716 -396 -3684
rect -364 -3716 -316 -3684
rect -284 -3716 -236 -3684
rect -204 -3716 -156 -3684
rect -124 -3716 -76 -3684
rect -44 -3716 4 -3684
rect 36 -3716 84 -3684
rect 116 -3716 164 -3684
rect 196 -3716 244 -3684
rect 276 -3716 324 -3684
rect 356 -3716 404 -3684
rect 436 -3716 484 -3684
rect 516 -3716 564 -3684
rect 596 -3716 644 -3684
rect 676 -3716 724 -3684
rect 756 -3716 804 -3684
rect 836 -3716 884 -3684
rect 916 -3716 964 -3684
rect 996 -3716 1044 -3684
rect 1076 -3716 1124 -3684
rect 1156 -3716 1204 -3684
rect 1236 -3716 1284 -3684
rect 1316 -3716 1364 -3684
rect 1396 -3716 1444 -3684
rect 1476 -3716 1524 -3684
rect 1556 -3716 1604 -3684
rect 1636 -3716 1684 -3684
rect 1716 -3716 1764 -3684
rect 1796 -3716 1844 -3684
rect 1876 -3716 1924 -3684
rect 1956 -3716 2004 -3684
rect 2036 -3716 2084 -3684
rect 2116 -3716 2164 -3684
rect 2196 -3716 2244 -3684
rect 2276 -3716 2324 -3684
rect 2356 -3716 2404 -3684
rect 2436 -3716 2484 -3684
rect 2516 -3716 2564 -3684
rect 2596 -3716 2644 -3684
rect 2676 -3716 2724 -3684
rect 2756 -3716 2804 -3684
rect 2836 -3716 2884 -3684
rect 2916 -3716 2964 -3684
rect 2996 -3716 3044 -3684
rect 3076 -3716 3124 -3684
rect 3156 -3716 3204 -3684
rect 3236 -3716 3284 -3684
rect 3316 -3716 3364 -3684
rect 3396 -3716 3444 -3684
rect 3476 -3716 3524 -3684
rect 3556 -3716 3604 -3684
rect 3636 -3716 3684 -3684
rect 3716 -3716 3764 -3684
rect 3796 -3716 3844 -3684
rect 3876 -3716 3924 -3684
rect 3956 -3716 4004 -3684
rect 4036 -3716 4084 -3684
rect 4116 -3716 4164 -3684
rect 4196 -3716 4244 -3684
rect 4276 -3716 4324 -3684
rect 4356 -3716 4404 -3684
rect 4436 -3716 4484 -3684
rect 4516 -3716 4564 -3684
rect 4596 -3716 4644 -3684
rect 4676 -3716 4724 -3684
rect 4756 -3716 4804 -3684
rect 4836 -3716 4884 -3684
rect 4916 -3716 4964 -3684
rect 4996 -3716 5044 -3684
rect 5076 -3716 5124 -3684
rect 5156 -3716 5204 -3684
rect 5236 -3716 5284 -3684
rect 5316 -3716 5364 -3684
rect 5396 -3716 5444 -3684
rect 5476 -3716 5524 -3684
rect 5556 -3716 5604 -3684
rect 5636 -3716 5684 -3684
rect 5716 -3716 5764 -3684
rect 5796 -3716 5844 -3684
rect 5876 -3716 5924 -3684
rect 5956 -3716 6004 -3684
rect 6036 -3716 6084 -3684
rect 6116 -3716 6164 -3684
rect 6196 -3716 6244 -3684
rect 6276 -3716 6324 -3684
rect 6356 -3716 6404 -3684
rect 6436 -3716 6484 -3684
rect 6516 -3716 6564 -3684
rect 6596 -3716 6644 -3684
rect 6676 -3716 6724 -3684
rect 6756 -3716 6804 -3684
rect 6836 -3716 6884 -3684
rect 6916 -3716 6964 -3684
rect 6996 -3716 7044 -3684
rect 7076 -3716 7124 -3684
rect 7156 -3716 7204 -3684
rect 7236 -3716 7284 -3684
rect 7316 -3716 7364 -3684
rect 7396 -3716 7444 -3684
rect 7476 -3716 7524 -3684
rect 7556 -3716 7604 -3684
rect 7636 -3716 7684 -3684
rect 7716 -3716 7764 -3684
rect 7796 -3716 7844 -3684
rect 7876 -3716 7924 -3684
rect 7956 -3716 8004 -3684
rect 8036 -3716 8084 -3684
rect 8116 -3716 8164 -3684
rect 8196 -3716 8244 -3684
rect 8276 -3716 8324 -3684
rect 8356 -3716 8404 -3684
rect 8436 -3716 8484 -3684
rect 8516 -3716 8564 -3684
rect 8596 -3716 8644 -3684
rect 8676 -3716 8724 -3684
rect 8756 -3716 8804 -3684
rect 8836 -3716 8884 -3684
rect 8916 -3716 8964 -3684
rect 8996 -3716 9044 -3684
rect 9076 -3716 9124 -3684
rect 9156 -3716 9204 -3684
rect 9236 -3716 9284 -3684
rect 9316 -3716 9364 -3684
rect 9396 -3716 9444 -3684
rect 9476 -3716 9524 -3684
rect 9556 -3716 9604 -3684
rect 9636 -3716 9684 -3684
rect 9716 -3716 9764 -3684
rect 9796 -3716 9844 -3684
rect 9876 -3716 9924 -3684
rect 9956 -3716 10004 -3684
rect 10036 -3716 10084 -3684
rect 10116 -3716 10164 -3684
rect 10196 -3716 10244 -3684
rect 10276 -3716 10324 -3684
rect 10356 -3716 10404 -3684
rect 10436 -3716 10484 -3684
rect 10516 -3716 10644 -3684
rect 10676 -3716 10804 -3684
rect 10836 -3716 10964 -3684
rect 10996 -3716 11000 -3684
rect -720 -3720 11000 -3716
<< labels >>
rlabel metal3 -640 1040 -600 1080 0 ii
port 1 nsew
rlabel metal3 -480 1040 -440 1080 0 vi
port 2 nsew
rlabel metal3 10720 1040 10760 1080 0 n
rlabel metal3 10880 1040 10920 1080 0 vo
port 3 nsew
rlabel metal3 10960 1040 11000 1080 0 vssa
port 4 nsew
<< end >>
