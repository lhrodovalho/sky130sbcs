* Self-biased current source testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0

.include "../mag/sbcs1v8.spice"

* supply voltages
vdda	vdda 0 1.8
vssa	vssa 0 0.0

.subckt p1_2 d g s b
xd d g x b sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=4
xs x g s b sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=4
.ends

.subckt p1_4 d g s b
xd d g x b p1_2
xs x g s b p1_2
.ends

.subckt p1_8 d g s b
xd d g x b p1_4
xs x g s b p1_4
.ends

.subckt p1_16 d g s b
xd d g x b p1_8
xs x g s b p1_8
.ends

.subckt p1_32 d g s b
xd d g x b p1_16
xs x g s b p1_16
.ends

.subckt p1_64 d g s b
xd d g x b p1_32
xs x g s b p1_32
.ends

.subckt p2_2 d g s b
xl d g s b p1_2
xr d g s b p1_2
.ends

.subckt p4_2 d g s b
xl d g s b p2_2
xr d g s b p2_2
.ends

.subckt p8_2 d g s b
xl d g s b p4_2
xr d g s b p4_2
.ends

.subckt p2_4 d g s b
xl d g s b p1_4
xr d g s b p1_4
.ends

.subckt p4_4 d g s b
xl d g s b p2_4
xr d g s b p2_4
.ends

.subckt p2_8 d g s b
xl d g s b p1_8
xr d g s b p1_8
.ends

.subckt buffer in out vdda vssa
xpa  n   p   out  in    p1_16
xpb  p   p   out  out   p1_16
xna  n   n   vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=8
xnb  p   n   vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=8
is vdda out 100n
.ends

* DUT
x0 io vdda vssa x sbcs1v8
vo io y 0.0

xpa  n   x   y    y    p1_16
xpb1 ref ref y    y    sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=64
xna  n   n   vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=8
xnb  ref n   vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u m=8

x1 ref ref0 vdda vssa buffer

.option gmin=1e-13
.control
  dc vdda 10m 1.95 10m
  plot x ref
  plot i(vo)
  plot abs(deriv(ref)/ref) ylog
  
  dc temp -40 125 1
  meas dc r27 find ref at=27
  let refN = ref/r27
  plot refN
  
.endc

.end
