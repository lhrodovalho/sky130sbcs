* NGSPICE file created from sbcs1v8.ext - technology: sky130A

.subckt sbcs1v8 io vdda vssa x
X0 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X1 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X2 a_11920_2720# p1 a_11360_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X3 a_15440_3840# y a_14800_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X4 p0 y a_1680_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X5 io p2 a_14800_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X6 a_13200_6560# p0 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X7 a_10320_n10720# s a_9680_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X8 a_400_n7320# p0 a_n160_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X9 a_4560_n3480# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X10 a_9680_n7320# p2 a_9040_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X11 a_4560_9960# s a_3920_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X12 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X13 p2 n a_6160_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X14 a_6160_9960# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X15 a_11920_n760# y y vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X16 x p2 a_n160_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X17 a_4560_6120# p2 p1 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X18 x p2 a_15440_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X19 a_6160_6120# p2 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X20 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X21 a_11920_10400# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X22 a_6160_7680# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X23 vdda p1 a_n160_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X24 a_15440_n3480# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X25 vdda p1 a_15440_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X26 a_n960_3800# a_n960_3800# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X27 a_10960_n3480# p1 a_10320_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X28 a_16080_n7320# p0 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X29 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X30 a_400_n760# x vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X31 vdda p0 a_400_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X32 vdda s a_11920_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X33 a_16080_n760# x z vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X34 vssa a_17120_0# a_17120_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X35 vssa n a_10320_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X36 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X37 a_16720_n7320# p0 a_16080_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X38 a_9680_6560# p2 a_9040_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X39 a_6160_n10720# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X40 a_12560_9960# s a_11920_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X41 a_14800_n11160# p1 a_14240_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X42 vdda p1 a_1040_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X43 a_14800_3840# y p0 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X44 a_1040_n8440# s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X45 p1 p2 a_11920_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X46 a_3920_9960# s a_3280_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X47 a_9040_n3480# p1 a_8480_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X48 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X49 vssa x a_16080_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X50 a_13840_2280# p2 a_13200_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X51 p1 p2 a_3280_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X52 a_4560_n10720# s a_3920_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X53 vdda p1 a_11920_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X54 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X55 vdda a_17120_n7320# a_17120_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X56 a_13840_2280# p1 a_13200_2720# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X57 p2 p2 a_7440_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X58 a_7440_n7320# p2 a_6800_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X59 a_5200_2280# p2 a_4560_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X60 vdda p1 a_400_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X61 a_3280_n11160# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X62 a_8080_n3480# p2 a_7440_n3040# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X63 a_5200_2280# p1 a_4560_2720# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X64 vdda s a_7440_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X65 vdda a_17120_n11160# a_17120_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X66 vssa x a_13200_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X67 n n a_7440_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X68 vssa n a_7440_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X69 x p2 a_1040_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X70 a_10320_3840# n p2 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X71 a_5200_n3480# p1 a_4560_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X72 a_10320_n7320# p2 a_9680_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X73 a_3280_2280# p2 a_2720_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X74 a_6800_n10720# s a_6160_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X75 p2 p2 a_7440_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X76 y y a_4560_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X77 vdda p1 a_1040_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X78 s n a_7440_7680# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X79 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X80 a_3280_2720# p1 a_2720_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X81 vdda a_17120_6120# a_17120_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X82 a_13840_n7320# p0 a_13200_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X83 vdda s a_10320_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X84 a_7440_6560# p2 a_6800_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X85 a_1680_n760# x z vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X86 a_1680_n11160# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X87 a_9040_6560# p2 p2 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X88 a_3280_n760# x vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X89 a_11920_9960# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X90 a_6160_n3480# p1 a_5600_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X91 a_11920_6120# p2 a_11360_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X92 a_400_n6880# p2 a_n160_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X93 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X94 a_13200_n10720# s a_12560_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X95 z x a_400_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X96 a_9680_n6880# p2 a_9040_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X97 a_13200_2280# p2 y vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X98 vdda s a_3280_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X99 x p2 a_n160_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X100 a_4560_n7320# p0 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X101 a_400_n4600# y vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X102 n p2 a_9040_n3040# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X103 a_400_9960# p2 a_n160_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X104 vssa y a_16080_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X105 a_400_n10720# p2 a_n160_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X106 a_13200_2720# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X107 a_16080_9960# p2 io vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X108 p2 n a_9040_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X109 vdda s a_7440_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X110 vdda p1 a_6160_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X111 a_400_6120# p2 a_n160_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X112 a_2320_n3480# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X113 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X114 vdda s a_7440_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X115 a_16080_6120# p2 p0 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X116 a_13200_n760# x z vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X117 vdda p2 a_10320_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X118 p1 s a_15440_7680# vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X119 a_n960_n3600# a_n960_n3600# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X120 a_16080_n6880# p2 p0 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X121 vdda p0 a_14800_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X122 vdda p2 a_10320_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X123 a_4560_3840# n a_3920_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X124 vdda p0 a_14800_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X125 a_2320_6120# p0 a_1680_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X126 x p2 a_15440_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X127 a_6160_3840# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X128 a_16080_n4600# y a_15440_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X129 a_1040_2280# p2 x vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X130 a_13200_n3480# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X131 a_6800_6560# p2 a_6160_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X132 vdda p1 a_14800_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X133 a_10320_n11160# s a_9680_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X134 a_1040_2280# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X135 a_16720_n7320# p2 a_16080_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X136 a_3280_n3480# p1 a_2720_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X137 a_16720_n3480# p2 x vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X138 z x a_400_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X139 a_n960_6000# a_n960_6000# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X140 n p2 a_9040_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X141 vssa y a_16080_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X142 a_6800_0# n a_6160_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X143 a_400_10400# p1 a_n160_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X144 a_9040_n10720# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X145 a_1680_n7320# p0 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X146 a_1680_0# x z vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X147 a_9680_10400# s a_9040_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X148 vdda p1 a_9040_2720# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X149 a_400_0# x vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X150 vdda s a_13200_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X151 vdda p1 a_3280_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X152 a_9040_n7320# p2 p2 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X153 vdda a_17120_n7320# a_17120_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X154 a_9680_n760# n a_9040_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X155 a_2320_n11160# p2 a_1680_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X156 a_11920_0# y y vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X157 a_13840_6120# p2 a_13200_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X158 a_7440_n6880# p2 a_6800_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X159 vdda s a_4560_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X160 a_12560_3840# n a_11920_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X161 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X162 vdda p0 a_11920_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X163 vdda a_17120_n3480# a_17120_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X164 a_7440_n10720# s a_6800_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X165 vssa a_17120_n4600# a_17120_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X166 a_7440_n3040# p2 n vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X167 a_16080_10400# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X168 vdda p1 a_14240_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X169 a_5200_6120# p2 a_4560_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X170 a_1680_9960# p2 io vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X171 a_7440_n4600# n p2 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X172 a_3920_3840# n a_3280_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X173 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X174 a_14800_6560# p0 a_14240_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X175 a_3280_9960# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X176 a_10320_n6880# p2 a_9680_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X177 a_7440_0# n a_6800_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X178 s n a_7440_n8440# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X179 a_6160_n11160# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X180 a_1680_6120# p2 p0 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X181 a_5200_n7320# p0 a_4560_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X182 a_1040_n3480# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X183 a_3280_0# x vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X184 a_10320_n3040# p2 n vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X185 a_3280_6120# p2 a_2720_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X186 p1 s a_1040_7680# vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X187 a_13840_n7320# p2 a_13200_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X188 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X189 a_10320_n4600# n p2 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X190 vdda a_17120_2280# a_17120_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X191 a_16720_9960# p1 a_16080_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X192 a_13840_n3480# p2 a_13200_n3040# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X193 z y a_11920_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X194 vssa n a_13200_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X195 vdda s a_13200_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X196 vdda a_17120_2280# a_17120_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X197 a_7440_2280# p2 n vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X198 vssa n a_7440_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X199 a_9040_2280# p2 a_8480_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X200 a_4560_n11160# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X201 a_7440_2720# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X202 a_9040_2720# p1 a_8480_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X203 a_10320_6560# p2 a_9680_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X204 a_6160_n7320# p2 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X205 vssa a_17120_n760# a_17120_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X206 a_9040_0# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X207 x x a_1680_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X208 a_13200_9960# s a_12560_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X209 a_7440_n760# n a_6800_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X210 a_4560_n6880# p2 p1 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X211 vdda a_17120_n11160# a_17120_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X212 a_9040_n760# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X213 vdda a_17120_9960# a_17120_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X214 a_13200_6120# p2 p1 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X215 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X216 a_11920_3840# n p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X217 a_7440_10400# s a_6800_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X218 a_4560_n3040# p2 y vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X219 a_6800_n11160# s a_6160_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X220 a_11920_n3480# p1 a_11360_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X221 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X222 a_4560_n4600# n a_3920_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X223 a_9680_n8440# n a_9040_n8440# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X224 a_6800_n7320# p2 a_6160_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X225 vdda s a_10320_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X226 p0 p2 a_14800_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X227 a_2320_n7320# p0 a_1680_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X228 a_10320_10400# s a_9680_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X229 a_10960_2280# p2 a_10320_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X230 vdda p2 a_10320_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X231 a_n960_n7440# a_n960_n7440# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X232 a_15440_n3480# p2 x vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X233 a_400_3840# y vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X234 io p2 a_400_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X235 a_15440_n4600# y a_14800_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X236 a_10960_2280# p1 a_10320_2720# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X237 a_9680_0# n a_9040_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X238 vdda s a_13200_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X239 a_10960_n3480# p2 a_10320_n3040# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X240 a_15440_2280# p2 x vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X241 a_2320_2280# p2 x vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X242 a_16080_3840# y a_15440_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X243 vssa n a_10320_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X244 p1 s a_15440_n8440# vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X245 p0 p2 a_400_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X246 a_13200_n7320# p0 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X247 a_15440_2280# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X248 a_13200_n11160# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X249 a_2320_2280# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X250 a_16720_6120# p0 a_16080_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X251 a_1040_7680# s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X252 vssa n a_10320_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X253 n p2 a_6160_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X254 a_9680_n10720# s a_9040_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X255 a_13200_0# x z vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X256 a_3280_n7320# p0 a_2720_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X257 vdda p1 a_6160_2720# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X258 a_9680_9960# s a_9040_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X259 z x a_14800_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X260 x x a_1680_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X261 a_400_n11160# p1 a_n160_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X262 a_1680_n6880# p2 p0 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X263 a_n960_2160# a_n960_2160# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X264 a_9680_6120# p2 a_9040_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X265 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X266 a_11920_n10720# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X267 a_6800_n760# n a_6160_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X268 a_4560_6560# p0 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X269 a_9680_7680# n a_9040_7680# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X270 a_6160_6560# p2 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X271 a_4560_10400# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X272 x p2 a_1040_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X273 a_9040_n6880# p2 p2 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X274 a_n960_2160# a_n960_2160# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X275 a_1680_n4600# y a_1040_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X276 vdda p0 a_3280_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X277 a_9040_n3040# p2 a_8480_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X278 p1 p2 a_11920_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X279 a_16080_n10720# p2 io vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X280 a_9040_n4600# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X281 a_n960_n880# a_n960_n880# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X282 vssa x a_13200_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X283 y p2 a_11920_n3040# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X284 vdda p1 a_14800_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X285 vdda s a_4560_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X286 a_12560_n4600# n a_11920_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X287 vdda s a_10320_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X288 vssa a_17120_n8440# a_17120_n8440# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X289 a_14800_n7320# p0 a_14240_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X290 vssa n a_13200_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X291 a_7440_n8440# n a_6800_n8440# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X292 a_5200_n7320# p2 a_4560_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X293 x p2 a_14240_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X294 a_10320_0# n a_9680_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X295 vdda p1 a_14240_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X296 p1 n a_4560_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X297 a_5200_n3480# p2 a_4560_n3040# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X298 vdda a_17120_9960# a_17120_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X299 vdda p0 a_400_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X300 a_9040_n11160# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X301 p1 n a_4560_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X302 a_10320_n8440# n a_9680_n8440# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X303 a_n960_n11280# a_n960_n11280# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X304 a_7440_9960# s a_6800_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X305 a_1680_3840# y a_1040_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X306 vdda a_17120_6120# a_17120_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X307 a_14800_n760# x x vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X308 vdda p0 a_11920_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X309 a_9040_9960# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X310 vssa a_17120_7680# a_17120_7680# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X311 a_3280_3840# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X312 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X313 a_7440_6120# p2 a_6800_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X314 a_2320_n11160# p1 a_1680_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X315 a_1680_10400# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X316 a_7440_7680# n a_6800_7680# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X317 a_9040_6120# p2 p2 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X318 a_16720_n11160# p2 a_16080_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X319 a_6160_n6880# p2 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X320 vdda p0 a_3280_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X321 a_9040_7680# n s vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X322 a_7440_n11160# s a_6800_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X323 a_10320_2280# p2 n vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X324 a_9040_10400# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X325 a_6160_n3040# p2 a_5600_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X326 a_6160_n4600# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X327 a_8080_n3480# p1 a_7440_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X328 a_10320_2720# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X329 vdda s a_11920_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X330 a_6800_n6880# p2 a_6160_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X331 p2 p2 a_7440_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X332 a_11920_n7320# p0 a_11360_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X333 a_10320_n760# n a_9680_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X334 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X335 a_2320_n7320# p2 a_1680_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X336 vdda s a_10320_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X337 a_13200_3840# n a_12560_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X338 n p2 a_6160_n3040# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X339 a_n960_n7440# a_n960_n7440# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X340 a_16080_0# x z vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X341 p2 n a_6160_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X342 vdda s a_4560_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X343 a_2320_n3480# p2 x vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X344 vdda s a_13200_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X345 vdda p2 a_10320_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X346 io p2 a_14800_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X347 p0 y a_1680_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X348 a_2320_9960# p2 a_1680_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X349 a_n960_n3600# a_n960_n3600# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X350 vssa n a_10320_7680# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X351 a_n960_n4720# a_n960_n4720# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X352 a_15440_n8440# s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X353 a_13200_n6880# p2 p1 vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X354 p0 p2 a_14800_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X355 a_2320_6120# p2 a_1680_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X356 a_6800_9960# s a_6160_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X357 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X358 a_15440_7680# s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X359 vssa n a_10320_n8440# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X360 a_11920_6560# p0 a_11360_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X361 a_13200_n3040# p2 y vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X362 a_12560_n10720# s a_11920_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X363 a_16720_2280# p2 x vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X364 a_3280_n6880# p2 a_2720_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X365 a_13200_n4600# n a_12560_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X366 a_6800_6120# p2 a_6160_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X367 a_6800_7680# n a_6160_7680# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X368 vdda p1 a_n160_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X369 a_16720_2280# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X370 a_6160_10400# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X371 vdda p1 a_9040_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X372 a_3280_n3040# p2 a_2720_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X373 a_1040_3840# y a_400_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X374 a_n960_9840# a_n960_9840# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X375 a_3280_n4600# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X376 a_400_6560# p0 a_n160_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X377 vssa x a_16080_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X378 a_n960_6000# a_n960_6000# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X379 a_4560_2280# p2 y vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X380 a_16080_6560# p0 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X381 a_n960_7640# a_n960_7640# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X382 a_6160_2280# p2 a_5600_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X383 a_14800_n10720# p2 a_14240_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X384 p1 p2 a_3280_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X385 z x a_3280_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X386 p1 s a_1040_n8440# vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X387 a_4560_2720# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X388 a_6160_2720# p1 a_5600_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X389 p2 n a_9040_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X390 a_6800_10400# s a_6160_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X391 y p2 a_3280_n3040# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X392 vdda p1 a_15440_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X393 a_3920_n4600# n a_3280_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X394 a_2320_9960# p1 a_1680_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X395 a_9040_n8440# n s vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X396 a_4560_n760# y z vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X397 a_n960_9840# a_n960_9840# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X398 a_6160_n760# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X399 a_14800_n6880# p2 a_14240_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X400 a_9680_n11160# s a_9040_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X401 a_14800_9960# p2 a_14240_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X402 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X403 x p2 a_14240_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X404 a_14800_6120# p2 a_14240_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X405 p0 p2 a_400_n6880# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X406 a_14800_n4600# y p0 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X407 io p2 a_400_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X408 a_3280_n10720# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X409 a_13200_10400# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X410 p1 s n vssa sky130_fd_pr__nfet_01v8_lvt ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X411 a_16720_n3480# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X412 a_11920_n11160# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X413 a_4560_0# y z vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X414 a_1040_n3480# p2 x vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X415 a_n960_n40# a_n960_n40# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X416 a_3280_10400# s vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X417 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X418 a_1040_n4600# y a_400_n4600# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X419 y p2 a_11920_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X420 a_16080_n11160# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X421 a_14800_0# x x vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X422 a_1680_n10720# p2 io vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X423 vdda p1 a_11920_2720# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X424 a_13840_6120# p0 a_13200_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X425 a_10320_9960# s a_9680_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X426 y p2 a_3280_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X427 vssa a_17120_3840# a_17120_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X428 vdda s a_4560_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X429 vdda a_17120_n3480# a_17120_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X430 vdda s a_3280_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X431 a_7440_n3480# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X432 vdda p1 a_3280_2720# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X433 a_7440_3840# n p2 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X434 a_10320_6120# p2 a_9680_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X435 z y a_11920_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X436 a_5200_6120# p0 a_4560_6560# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X437 a_9040_3840# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X438 a_10320_7680# n a_9680_7680# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X439 a_6160_n8440# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X440 p2 p2 a_7440_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X441 a_6160_0# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X442 a_11920_n6880# p2 a_11360_n7320# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X443 a_1680_6560# p0 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X444 z x a_3280_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X445 a_3920_n10720# s a_3280_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X446 a_3280_6560# p0 a_2720_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X447 a_10320_n3480# p1 vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X448 a_14800_10400# p1 a_14240_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X449 a_n960_n11280# a_n960_n11280# vdda vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X450 a_11920_n3040# p2 a_11360_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X451 a_8080_2280# p2 a_7440_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X452 a_11920_n4600# n p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X453 z x a_14800_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X454 a_13840_n3480# p1 a_13200_n3480# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X455 a_8080_2280# p1 a_7440_2720# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X456 a_6800_n8440# n a_6160_n8440# vssa sky130_fd_pr__nfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X457 vdda p1 a_400_10400# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X458 vdda s a_7440_n10720# vdda sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X459 n s p1 vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X460 a_16720_n11160# p1 a_16080_n11160# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X461 a_n960_n8560# a_n960_n8560# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X462 n n a_7440_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=7.42857e+11p pd=3.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X463 a_16720_9960# p2 a_16080_9960# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X464 y y a_4560_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X465 vssa n a_10320_3840# vssa sky130_fd_pr__nfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X466 a_11920_2280# p2 a_11360_2280# vdda sky130_fd_pr__pfet_01v8_lvt ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X467 a_16720_6120# p2 a_16080_6120# vdda sky130_fd_pr__pfet_01v8_lvt ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
.ends

