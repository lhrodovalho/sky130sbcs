* NGSPICE file created from vref1v8.ext - technology: sky130A

.subckt vref1v8 ii vi vo vssa
X0 n vi a_9360_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=3.2e+12p pd=1.44e+07u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X1 a_1680_n4800# n a_1040_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X2 a_19280_n4800# n a_18640_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X3 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=4.32e+13p pd=1.664e+08u as=3.12e+13p ps=1.144e+08u w=1e+06u l=2e+06u
X4 a_13520_n6880# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X5 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6 a_14800_n5560# n a_14160_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X7 n n a_17360_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=9.6e+12p pd=3.52e+07u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X8 a_15440_n3480# vi a_14800_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X9 a_12240_1320# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X10 a_10960_n3480# vi n ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X11 vssa n a_4240_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=2.24e+13p pd=9.28e+07u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X12 a_19920_n4800# n a_19280_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X13 a_400_n760# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X14 a_1040_n5560# n a_400_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X15 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X16 a_16080_n760# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X17 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X18 vssa n a_19920_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X19 a_10960_0# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X20 a_11600_n3480# vi a_10960_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X21 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X22 a_5520_n5560# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X23 a_6160_1320# vi a_5520_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X24 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X25 vssa n a_19920_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X26 a_16080_n2080# vi a_15440_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X27 a_19280_n3480# vi a_18640_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X28 a_6160_n4800# n a_5520_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X29 a_16720_0# n a_16080_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X30 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X31 a_19280_0# n a_18640_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X32 a_16720_n2080# vi a_16080_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X33 a_19920_n3480# vi a_19280_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X34 a_8080_n6880# vi a_7440_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X35 a_6800_n4800# n a_6160_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X36 a_5520_0# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X37 a_12240_n2080# vi a_11600_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X38 a_9360_n5560# n a_8720_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X39 vo n a_1680_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=9.6e+12p pd=3.52e+07u as=0p ps=0u w=1e+06u l=2e+06u
X40 a_8080_0# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X41 a_3600_n760# n a_2960_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X42 a_19920_n760# n a_19280_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X43 vo n a_12240_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X44 ii vo a_13520_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X45 a_8720_n6880# vi a_8080_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X46 a_1680_n760# n a_1040_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X47 a_4240_n6880# vi a_3600_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X48 vssa n a_9360_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X49 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X50 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X51 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X52 n vi a_9360_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X53 a_9360_n760# n a_8720_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X54 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X55 a_13520_n5560# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X56 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X57 a_1040_0# n a_400_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X58 a_400_n6880# vi ii ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X59 a_18640_n4800# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X60 a_14160_n4800# n a_13520_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X61 a_8080_1320# vi a_7440_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X62 a_12240_0# n a_11600_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X63 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X64 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X65 a_11600_n760# n a_10960_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X66 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X67 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X68 a_14800_n4800# n a_14160_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X69 a_17360_n5560# n a_16720_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X70 vssa n a_4240_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X71 a_1040_n4800# n a_400_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X72 vo n a_17360_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X73 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X74 vo n a_12240_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X75 a_17360_n760# n a_16720_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X76 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X77 vssa n a_19920_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X78 a_5520_n760# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X79 a_12240_n6880# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X80 a_400_1320# vi ii ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X81 a_6800_0# n a_6160_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X82 a_1040_n760# n a_400_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X83 a_15440_n2080# vi a_14800_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X84 vo n a_17360_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X85 a_5520_n4800# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X86 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X87 a_1680_0# n a_1040_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X88 a_10960_n2080# vi n ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X89 a_18640_n3480# vi a_18000_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X90 a_400_0# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X91 a_9360_0# n a_8720_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X92 a_14160_n3480# vi a_13520_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X93 a_8080_n5560# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X94 a_18640_0# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X95 a_7440_n6880# vi a_6800_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X96 a_11600_n2080# vi a_10960_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X97 a_2960_n6880# vi a_2320_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X98 a_14800_n3480# vi a_14160_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X99 a_8720_n5560# n a_8080_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X100 n n a_6800_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X101 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X102 a_4240_n5560# n a_3600_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X103 a_19280_n2080# vi a_18640_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X104 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X105 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X106 a_9360_n4800# n a_8720_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X107 a_13520_n760# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X108 a_3600_n6880# vi a_2960_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X109 ii vi a_19920_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X110 a_400_n5560# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X111 n n a_12240_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X112 a_19920_n2080# vi a_19280_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X113 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X114 vssa n a_9360_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X115 a_3600_1320# vi a_2960_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X116 a_2960_n760# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X117 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X118 n n a_1680_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X119 a_19280_n760# n a_18640_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X120 vo n a_6800_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X121 a_13520_n4800# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X122 a_1680_1320# vi a_1040_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X123 a_16080_n5560# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X124 a_11600_0# n a_10960_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X125 a_14160_0# n a_13520_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X126 a_9360_1320# vi a_8720_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X127 ii vo a_14800_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X128 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X129 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X130 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X131 a_16720_n5560# n a_16080_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X132 a_2960_0# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X133 a_12240_n5560# n a_11600_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X134 a_12880_n3480# vi a_12240_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X135 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X136 a_10960_n760# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X137 a_17360_n4800# n a_16720_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X138 a_19920_0# n a_19280_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X139 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X140 vo n a_1680_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X141 vssa n a_14800_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X142 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X143 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X144 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X145 a_1680_n6880# vi a_1040_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X146 a_6800_n760# n a_6160_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X147 a_13520_n3480# vi a_12880_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X148 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X149 n n a_6800_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X150 a_8720_0# n a_8080_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X151 a_2960_n5560# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X152 n n a_17360_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X153 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X154 a_5520_1320# vi a_4880_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X155 vssa n a_4240_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X156 a_8080_n4800# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X157 a_1040_1320# vi a_400_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X158 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X159 a_3600_n5560# n a_2960_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X160 a_18640_n2080# vi a_18000_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X161 a_8720_n4800# n a_8080_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X162 a_14160_n2080# vi a_13520_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X163 a_4240_n4800# n a_3600_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X164 a_17360_n3480# vi a_16720_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X165 a_14800_n760# n a_14160_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X166 a_400_n4800# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X167 a_13520_1320# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X168 n n a_12240_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X169 a_14800_n2080# vi a_14160_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X170 a_18000_n3480# vi a_17360_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X171 a_6160_n6880# vi a_5520_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X172 a_4240_0# n a_3600_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X173 a_4240_n760# n a_3600_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X174 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X175 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X176 vssa n a_14800_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X177 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X178 a_8720_n760# n a_8080_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X179 a_10960_n5560# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X180 a_2960_1320# vi a_2320_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X181 ii vi a_19920_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X182 a_6800_n6880# vi a_6160_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X183 a_16080_n4800# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X184 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X185 a_13520_0# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X186 a_2320_n6880# vi a_1680_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X187 a_7440_1320# vi a_6800_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X188 a_16080_0# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X189 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X190 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X191 vssa n a_9360_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X192 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X193 a_11600_n5560# n a_10960_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X194 vssa n a_4240_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X195 a_16720_n4800# n a_16080_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X196 a_1680_n5560# n a_1040_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X197 a_12240_n4800# n a_11600_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X198 a_19280_n5560# n a_18640_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X199 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X200 a_12240_n760# n a_11600_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X201 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X202 a_16720_n760# n a_16080_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X203 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X204 ii vo a_13520_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X205 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X206 a_19920_n5560# n a_19280_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X207 vo n a_6800_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X208 a_12880_n2080# vi a_12240_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X209 a_2960_n4800# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X210 a_2320_1320# vi a_1680_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X211 ii vo a_14800_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X212 a_16080_n3480# vi a_15440_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X213 a_6800_1320# vi a_6160_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X214 a_6160_n760# n a_5520_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X215 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X216 a_14800_n6880# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X217 a_13520_n2080# vi a_12880_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X218 a_4880_n6880# vi a_4240_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X219 a_1040_n6880# vi a_400_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X220 a_3600_n4800# n a_2960_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X221 a_4880_1320# vi a_4240_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.2e+12p ps=4.4e+06u w=1e+06u l=2e+06u
X222 a_16720_n3480# vi a_16080_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X223 a_12240_n3480# vi a_11600_n3480# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X224 a_6160_n5560# n a_5520_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X225 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X226 a_14800_0# n a_14160_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X227 a_5520_n6880# vi a_4880_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X228 a_17360_0# n a_16720_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X229 a_6800_n5560# n a_6160_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X230 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X231 n n a_1680_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X232 a_14800_1320# vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X233 a_3600_0# n a_2960_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X234 a_14160_n760# n a_13520_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X235 a_17360_n2080# vi a_16720_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X236 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X237 a_6160_0# n a_5520_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X238 a_18640_n760# n n vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X239 vssa n a_14800_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X240 ii vo a_12240_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X241 a_10960_n4800# n vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=4.4e+06u as=0p ps=0u w=1e+06u l=2e+06u
X242 vssa n a_14800_0# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X243 vssa n a_9360_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X244 a_4240_1320# vi a_3600_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X245 vssa n a_19920_n760# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X246 a_18000_n2080# vi a_17360_n2080# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X247 ii vo vo ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X248 a_9360_n6880# vi a_8720_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X249 a_8720_1320# vi a_8080_1320# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X250 a_8080_n760# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X251 vo vo ii ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X252 ii vo a_12240_n6880# ii sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X253 a_18640_n5560# n vo vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X254 a_11600_n4800# n a_10960_n4800# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X255 a_14160_n5560# n a_13520_n5560# vssa sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
.ends

