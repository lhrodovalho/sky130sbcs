magic
tech sky130A
timestamp 1640909703
<< nwell >>
rect -200 920 320 1440
rect 520 920 1040 1440
<< mvpsubdiff >>
rect -320 1520 -240 1560
rect 1080 1520 1160 1560
rect -320 1480 -280 1520
rect 400 1480 440 1520
rect 1120 1480 1160 1520
rect 400 840 440 880
rect -280 800 -240 840
rect -160 800 280 840
rect 560 800 1000 840
rect 1080 800 1120 840
rect -160 480 280 520
rect -160 440 -120 480
rect 240 440 280 480
rect -160 120 -120 160
rect 240 120 280 160
rect 560 480 1000 520
rect 560 440 600 480
rect 960 440 1000 480
rect 560 120 600 160
rect 960 120 1000 160
rect -320 80 -240 120
rect 1080 80 1160 120
<< mvnsubdiff >>
rect -160 1360 -80 1400
rect 200 1360 280 1400
rect -160 1320 -120 1360
rect 240 1320 280 1360
rect -160 1000 -120 1040
rect 240 1000 280 1040
rect -160 960 280 1000
rect 560 1360 640 1400
rect 920 1360 1000 1400
rect 560 1320 600 1360
rect 960 1320 1000 1360
rect 560 1000 600 1040
rect 960 1000 1000 1040
rect 560 960 1000 1000
<< mvpsubdiffcont >>
rect -240 1520 1080 1560
rect -320 120 -280 1480
rect 400 880 440 1480
rect -240 800 -160 840
rect 280 800 560 840
rect 1000 800 1080 840
rect -160 160 -120 440
rect 240 160 280 440
rect 560 160 600 440
rect 960 160 1000 440
rect 1120 120 1160 1480
rect -240 80 1080 120
<< mvnsubdiffcont >>
rect -80 1360 200 1400
rect -160 1040 -120 1320
rect 240 1040 280 1320
rect 640 1360 920 1400
rect 560 1040 600 1320
rect 960 1040 1000 1320
<< xpolycontact >>
rect -80 600 200 720
rect 640 600 920 720
<< ppolyres >>
rect 200 600 640 720
<< pdiode >>
rect -80 1280 200 1320
rect -80 1080 -40 1280
rect 160 1080 200 1280
rect -80 1040 200 1080
rect 640 1280 920 1320
rect 640 1080 680 1280
rect 880 1080 920 1280
rect 640 1040 920 1080
<< ndiode >>
rect -80 400 200 440
rect -80 200 -40 400
rect 160 200 200 400
rect -80 160 200 200
rect 640 400 920 440
rect 640 200 680 400
rect 880 200 920 400
rect 640 160 920 200
<< pdiodec >>
rect -40 1080 160 1280
rect 680 1080 880 1280
<< ndiodec >>
rect -40 200 160 400
rect 680 200 880 400
<< locali >>
rect -320 1520 -240 1560
rect 1080 1520 1160 1560
rect -320 1480 -280 1520
rect -400 750 -360 760
rect -400 730 -390 750
rect -370 730 -360 750
rect -400 590 -360 730
rect -400 570 -390 590
rect -370 570 -360 590
rect -400 560 -360 570
rect 400 1480 440 1520
rect -160 1360 -80 1400
rect 200 1360 280 1400
rect -160 1320 -120 1360
rect 240 1320 280 1360
rect -160 960 -120 1040
rect -80 1280 200 1320
rect -80 1080 -40 1280
rect 160 1080 200 1280
rect -280 800 -240 840
rect -160 800 -120 840
rect -240 750 -200 760
rect -240 730 -230 750
rect -210 730 -200 750
rect -240 590 -200 730
rect -240 570 -230 590
rect -210 570 -200 590
rect -240 560 -200 570
rect -160 750 -120 760
rect -160 730 -150 750
rect -130 730 -120 750
rect -160 590 -120 730
rect -160 570 -150 590
rect -130 570 -120 590
rect -160 560 -120 570
rect -80 720 200 1080
rect 240 960 280 1040
rect 1120 1480 1160 1520
rect 560 1360 640 1400
rect 920 1360 1000 1400
rect 560 1320 600 1360
rect 960 1320 1000 1360
rect 560 960 600 1040
rect 640 1280 920 1320
rect 640 1080 680 1280
rect 880 1080 920 1280
rect 400 840 440 880
rect 240 800 280 840
rect 560 800 600 840
rect -160 440 -120 520
rect -80 400 200 600
rect 640 720 920 1080
rect 960 960 1000 1040
rect 960 800 1000 840
rect 1080 800 1120 840
rect -80 200 -40 400
rect 160 200 200 400
rect -80 160 200 200
rect 240 440 280 520
rect -160 120 -120 160
rect 240 120 280 160
rect 560 440 600 520
rect 640 400 920 600
rect 960 750 1000 760
rect 960 730 970 750
rect 990 730 1000 750
rect 960 590 1000 730
rect 960 570 970 590
rect 990 570 1000 590
rect 960 560 1000 570
rect 1040 750 1080 760
rect 1040 730 1050 750
rect 1070 730 1080 750
rect 1040 590 1080 730
rect 1040 570 1050 590
rect 1070 570 1080 590
rect 1040 560 1080 570
rect 640 200 680 400
rect 880 200 920 400
rect 640 160 920 200
rect 960 440 1000 520
rect 560 120 600 160
rect 960 120 1000 160
rect 1200 750 1240 760
rect 1200 730 1210 750
rect 1230 730 1240 750
rect 1200 590 1240 730
rect 1200 570 1210 590
rect 1230 570 1240 590
rect 1200 560 1240 570
rect -320 80 -240 120
rect 1080 80 1160 120
<< viali >>
rect -390 730 -370 750
rect -390 570 -370 590
rect -70 1365 190 1395
rect -310 730 -290 750
rect -310 570 -290 590
rect -230 730 -210 750
rect -230 570 -210 590
rect -150 730 -130 750
rect -150 570 -130 590
rect 650 1365 910 1395
rect -70 645 190 675
rect 650 645 910 675
rect 970 730 990 750
rect 970 570 990 590
rect 1050 730 1070 750
rect 1050 570 1070 590
rect 1130 730 1150 750
rect 1130 570 1150 590
rect 1210 730 1230 750
rect 1210 570 1230 590
rect -70 85 190 115
rect 650 85 910 115
<< metal1 >>
rect -80 1395 200 1400
rect -80 1365 -70 1395
rect 190 1365 200 1395
rect -80 1360 200 1365
rect 640 1395 920 1400
rect 640 1365 650 1395
rect 910 1365 920 1395
rect 640 1360 920 1365
rect -400 755 -360 760
rect -400 725 -395 755
rect -365 725 -360 755
rect -400 720 -360 725
rect -320 755 -280 760
rect -320 725 -315 755
rect -285 725 -280 755
rect -320 720 -280 725
rect -240 755 -200 760
rect -240 725 -235 755
rect -205 725 -200 755
rect -240 720 -200 725
rect -160 755 -120 760
rect -160 725 -155 755
rect -125 725 -120 755
rect -160 720 -120 725
rect 960 755 1000 760
rect 960 725 965 755
rect 995 725 1000 755
rect 960 720 1000 725
rect 1040 755 1080 760
rect 1040 725 1045 755
rect 1075 725 1080 755
rect 1040 720 1080 725
rect 1120 755 1160 760
rect 1120 725 1125 755
rect 1155 725 1160 755
rect 1120 720 1160 725
rect 1200 755 1240 760
rect 1200 725 1205 755
rect 1235 725 1240 755
rect 1200 720 1240 725
rect -80 675 200 680
rect -80 645 -70 675
rect 190 645 200 675
rect -80 640 200 645
rect 640 675 920 680
rect 640 645 650 675
rect 910 645 920 675
rect 640 640 920 645
rect -400 595 -360 600
rect -400 565 -395 595
rect -365 565 -360 595
rect -400 560 -360 565
rect -320 595 -280 600
rect -320 565 -315 595
rect -285 565 -280 595
rect -320 560 -280 565
rect -240 595 -200 600
rect -240 565 -235 595
rect -205 565 -200 595
rect -240 560 -200 565
rect -160 595 -120 600
rect -160 565 -155 595
rect -125 565 -120 595
rect -160 560 -120 565
rect 960 595 1000 600
rect 960 565 965 595
rect 995 565 1000 595
rect 960 560 1000 565
rect 1040 595 1080 600
rect 1040 565 1045 595
rect 1075 565 1080 595
rect 1040 560 1080 565
rect 1120 595 1160 600
rect 1120 565 1125 595
rect 1155 565 1160 595
rect 1120 560 1160 565
rect 1200 595 1240 600
rect 1200 565 1205 595
rect 1235 565 1240 595
rect 1200 560 1240 565
rect -80 115 200 120
rect -80 85 -70 115
rect 190 85 200 115
rect -80 80 200 85
rect 640 115 920 120
rect 640 85 650 115
rect 910 85 920 115
rect 640 80 920 85
<< via1 >>
rect -70 1365 190 1395
rect 650 1365 910 1395
rect -395 750 -365 755
rect -395 730 -390 750
rect -390 730 -370 750
rect -370 730 -365 750
rect -395 725 -365 730
rect -315 750 -285 755
rect -315 730 -310 750
rect -310 730 -290 750
rect -290 730 -285 750
rect -315 725 -285 730
rect -235 750 -205 755
rect -235 730 -230 750
rect -230 730 -210 750
rect -210 730 -205 750
rect -235 725 -205 730
rect -155 750 -125 755
rect -155 730 -150 750
rect -150 730 -130 750
rect -130 730 -125 750
rect -155 725 -125 730
rect 965 750 995 755
rect 965 730 970 750
rect 970 730 990 750
rect 990 730 995 750
rect 965 725 995 730
rect 1045 750 1075 755
rect 1045 730 1050 750
rect 1050 730 1070 750
rect 1070 730 1075 750
rect 1045 725 1075 730
rect 1125 750 1155 755
rect 1125 730 1130 750
rect 1130 730 1150 750
rect 1150 730 1155 750
rect 1125 725 1155 730
rect 1205 750 1235 755
rect 1205 730 1210 750
rect 1210 730 1230 750
rect 1230 730 1235 750
rect 1205 725 1235 730
rect -70 645 190 675
rect 650 645 910 675
rect -395 590 -365 595
rect -395 570 -390 590
rect -390 570 -370 590
rect -370 570 -365 590
rect -395 565 -365 570
rect -315 590 -285 595
rect -315 570 -310 590
rect -310 570 -290 590
rect -290 570 -285 590
rect -315 565 -285 570
rect -235 590 -205 595
rect -235 570 -230 590
rect -230 570 -210 590
rect -210 570 -205 590
rect -235 565 -205 570
rect -155 590 -125 595
rect -155 570 -150 590
rect -150 570 -130 590
rect -130 570 -125 590
rect -155 565 -125 570
rect 965 590 995 595
rect 965 570 970 590
rect 970 570 990 590
rect 990 570 995 590
rect 965 565 995 570
rect 1045 590 1075 595
rect 1045 570 1050 590
rect 1050 570 1070 590
rect 1070 570 1075 590
rect 1045 565 1075 570
rect 1125 590 1155 595
rect 1125 570 1130 590
rect 1130 570 1150 590
rect 1150 570 1155 590
rect 1125 565 1155 570
rect 1205 590 1235 595
rect 1205 570 1210 590
rect 1210 570 1230 590
rect 1230 570 1235 590
rect 1205 565 1235 570
rect -70 85 190 115
rect 650 85 910 115
<< metal2 >>
rect -80 1395 200 1400
rect -80 1365 -70 1395
rect 190 1365 200 1395
rect -80 1360 200 1365
rect 640 1395 920 1400
rect 640 1365 650 1395
rect 910 1365 920 1395
rect 640 1360 920 1365
rect -440 755 1280 760
rect -440 725 -395 755
rect -365 725 -315 755
rect -285 725 -235 755
rect -205 725 -155 755
rect -125 725 965 755
rect 995 725 1045 755
rect 1075 725 1125 755
rect 1155 725 1205 755
rect 1235 725 1280 755
rect -440 720 1280 725
rect -440 675 200 680
rect -440 645 -70 675
rect 190 645 200 675
rect -440 640 200 645
rect 640 675 1280 680
rect 640 645 650 675
rect 910 645 1280 675
rect 640 640 1280 645
rect -440 595 1280 600
rect -440 565 -395 595
rect -365 565 -315 595
rect -285 565 -235 595
rect -205 565 -155 595
rect -125 565 965 595
rect 995 565 1045 595
rect 1075 565 1125 595
rect 1155 565 1205 595
rect 1235 565 1280 595
rect -440 560 1280 565
rect -80 115 200 120
rect -80 85 -70 115
rect 190 85 200 115
rect -80 80 200 85
rect 640 115 920 120
rect 640 85 650 115
rect 910 85 920 115
rect 640 80 920 85
<< via2 >>
rect -70 1365 190 1395
rect 650 1365 910 1395
rect -395 725 -365 755
rect -315 725 -285 755
rect -235 725 -205 755
rect -155 725 -125 755
rect 965 725 995 755
rect 1045 725 1075 755
rect 1125 725 1155 755
rect 1205 725 1235 755
rect -395 565 -365 595
rect -315 565 -285 595
rect -235 565 -205 595
rect -155 565 -125 595
rect 965 565 995 595
rect 1045 565 1075 595
rect 1125 565 1155 595
rect 1205 565 1235 595
rect -70 85 190 115
rect 650 85 910 115
<< metal3 >>
rect -80 1396 200 1400
rect -80 1364 -71 1396
rect 191 1364 200 1396
rect -80 1360 200 1364
rect 640 1396 920 1400
rect 640 1364 649 1396
rect 911 1364 920 1396
rect 640 1360 920 1364
rect -400 755 -360 760
rect -400 725 -395 755
rect -365 725 -360 755
rect -400 595 -360 725
rect -400 565 -395 595
rect -365 565 -360 595
rect -400 560 -360 565
rect -320 755 -280 760
rect -320 725 -315 755
rect -285 725 -280 755
rect -320 595 -280 725
rect -320 565 -315 595
rect -285 565 -280 595
rect -320 560 -280 565
rect -240 755 -200 760
rect -240 725 -235 755
rect -205 725 -200 755
rect -240 595 -200 725
rect -240 565 -235 595
rect -205 565 -200 595
rect -240 560 -200 565
rect -160 755 -120 760
rect -160 725 -155 755
rect -125 725 -120 755
rect -160 595 -120 725
rect -160 565 -155 595
rect -125 565 -120 595
rect -160 560 -120 565
rect 960 755 1000 760
rect 960 725 965 755
rect 995 725 1000 755
rect 960 595 1000 725
rect 960 565 965 595
rect 995 565 1000 595
rect 960 560 1000 565
rect 1040 755 1080 760
rect 1040 725 1045 755
rect 1075 725 1080 755
rect 1040 595 1080 725
rect 1040 565 1045 595
rect 1075 565 1080 595
rect 1040 560 1080 565
rect 1120 755 1160 760
rect 1120 725 1125 755
rect 1155 725 1160 755
rect 1120 595 1160 725
rect 1120 565 1125 595
rect 1155 565 1160 595
rect 1120 560 1160 565
rect 1200 755 1240 760
rect 1200 725 1205 755
rect 1235 725 1240 755
rect 1200 595 1240 725
rect 1200 565 1205 595
rect 1235 565 1240 595
rect 1200 560 1240 565
rect -80 116 200 120
rect -80 84 -71 116
rect 191 84 200 116
rect -80 80 200 84
rect 640 116 920 120
rect 640 84 649 116
rect 911 84 920 116
rect 640 80 920 84
<< via3 >>
rect -71 1395 191 1396
rect -71 1365 -70 1395
rect -70 1365 190 1395
rect 190 1365 191 1395
rect -71 1364 191 1365
rect 649 1395 911 1396
rect 649 1365 650 1395
rect 650 1365 910 1395
rect 910 1365 911 1395
rect 649 1364 911 1365
rect -71 115 191 116
rect -71 85 -70 115
rect -70 85 190 115
rect 190 85 191 115
rect -71 84 191 85
rect 649 115 911 116
rect 649 85 650 115
rect 650 85 910 115
rect 910 85 911 115
rect 649 84 911 85
<< metal4 >>
rect -400 1396 1280 1560
rect -400 1364 -71 1396
rect 191 1364 649 1396
rect 911 1364 1280 1396
rect -400 1360 1280 1364
rect -440 116 1240 280
rect -440 84 -71 116
rect 191 84 649 116
rect 911 84 1240 116
rect -440 80 1240 84
<< labels >>
rlabel metal2 -440 640 -400 680 0 a
port 1 nsew
rlabel metal2 1240 640 1280 680 0 b
port 2 nsew
rlabel metal4 -400 1360 1280 1560 0 vdda
port 3 nsew
rlabel metal4 -440 80 1240 280 0 vssa
port 4 nsew
<< end >>
