magic
tech sky130A
timestamp 1640954171
<< nwell >>
rect -200 480 10520 920
<< pmoslvt >>
rect 0 660 200 760
rect 320 660 520 760
rect 640 660 840 760
rect 960 660 1160 760
rect 1280 660 1480 760
rect 1600 660 1800 760
rect 1920 660 2120 760
rect 2240 660 2440 760
rect 2560 660 2760 760
rect 2880 660 3080 760
rect 3200 660 3400 760
rect 3520 660 3720 760
rect 3840 660 4040 760
rect 4160 660 4360 760
rect 4480 660 4680 760
rect 4800 660 5000 760
rect 5280 660 5480 760
rect 5600 660 5800 760
rect 5920 660 6120 760
rect 6240 660 6440 760
rect 6560 660 6760 760
rect 6880 660 7080 760
rect 7200 660 7400 760
rect 7520 660 7720 760
rect 7840 660 8040 760
rect 8160 660 8360 760
rect 8480 660 8680 760
rect 8800 660 9000 760
rect 9120 660 9320 760
rect 9440 660 9640 760
rect 9760 660 9960 760
rect 10080 660 10280 760
<< nmoslvt >>
rect 0 0 200 100
rect 320 0 520 100
rect 640 0 840 100
rect 960 0 1160 100
rect 1280 0 1480 100
rect 1600 0 1800 100
rect 1920 0 2120 100
rect 2240 0 2440 100
rect 2560 0 2760 100
rect 2880 0 3080 100
rect 3200 0 3400 100
rect 3520 0 3720 100
rect 3840 0 4040 100
rect 4160 0 4360 100
rect 4480 0 4680 100
rect 4800 0 5000 100
rect 5280 0 5480 100
rect 5600 0 5800 100
rect 5920 0 6120 100
rect 6240 0 6440 100
rect 6560 0 6760 100
rect 6880 0 7080 100
rect 7200 0 7400 100
rect 7520 0 7720 100
rect 7840 0 8040 100
rect 8160 0 8360 100
rect 8480 0 8680 100
rect 8800 0 9000 100
rect 9120 0 9320 100
rect 9440 0 9640 100
rect 9760 0 9960 100
rect 10080 0 10280 100
<< ndiff >>
rect -80 90 0 100
rect -80 10 -75 90
rect -45 10 0 90
rect -80 0 0 10
rect 200 90 320 100
rect 200 10 245 90
rect 275 10 320 90
rect 200 0 320 10
rect 520 90 640 100
rect 520 10 565 90
rect 595 10 640 90
rect 520 0 640 10
rect 840 90 960 100
rect 840 10 885 90
rect 915 10 960 90
rect 840 0 960 10
rect 1160 90 1280 100
rect 1160 10 1205 90
rect 1235 10 1280 90
rect 1160 0 1280 10
rect 1480 90 1600 100
rect 1480 10 1525 90
rect 1555 10 1600 90
rect 1480 0 1600 10
rect 1800 90 1920 100
rect 1800 10 1845 90
rect 1875 10 1920 90
rect 1800 0 1920 10
rect 2120 90 2240 100
rect 2120 10 2165 90
rect 2195 10 2240 90
rect 2120 0 2240 10
rect 2440 90 2560 100
rect 2440 10 2485 90
rect 2515 10 2560 90
rect 2440 0 2560 10
rect 2760 90 2880 100
rect 2760 10 2805 90
rect 2835 10 2880 90
rect 2760 0 2880 10
rect 3080 90 3200 100
rect 3080 10 3125 90
rect 3155 10 3200 90
rect 3080 0 3200 10
rect 3400 90 3520 100
rect 3400 10 3445 90
rect 3475 10 3520 90
rect 3400 0 3520 10
rect 3720 90 3840 100
rect 3720 10 3765 90
rect 3795 10 3840 90
rect 3720 0 3840 10
rect 4040 90 4160 100
rect 4040 10 4085 90
rect 4115 10 4160 90
rect 4040 0 4160 10
rect 4360 90 4480 100
rect 4360 10 4405 90
rect 4435 10 4480 90
rect 4360 0 4480 10
rect 4680 90 4800 100
rect 4680 10 4725 90
rect 4755 10 4800 90
rect 4680 0 4800 10
rect 5000 90 5080 100
rect 5000 10 5045 90
rect 5075 10 5080 90
rect 5000 0 5080 10
rect 5200 90 5280 100
rect 5200 10 5205 90
rect 5235 10 5280 90
rect 5200 0 5280 10
rect 5480 90 5600 100
rect 5480 10 5525 90
rect 5555 10 5600 90
rect 5480 0 5600 10
rect 5800 90 5920 100
rect 5800 10 5845 90
rect 5875 10 5920 90
rect 5800 0 5920 10
rect 6120 90 6240 100
rect 6120 10 6165 90
rect 6195 10 6240 90
rect 6120 0 6240 10
rect 6440 90 6560 100
rect 6440 10 6485 90
rect 6515 10 6560 90
rect 6440 0 6560 10
rect 6760 90 6880 100
rect 6760 10 6805 90
rect 6835 10 6880 90
rect 6760 0 6880 10
rect 7080 90 7200 100
rect 7080 10 7125 90
rect 7155 10 7200 90
rect 7080 0 7200 10
rect 7400 90 7520 100
rect 7400 10 7445 90
rect 7475 10 7520 90
rect 7400 0 7520 10
rect 7720 90 7840 100
rect 7720 10 7765 90
rect 7795 10 7840 90
rect 7720 0 7840 10
rect 8040 90 8160 100
rect 8040 10 8085 90
rect 8115 10 8160 90
rect 8040 0 8160 10
rect 8360 90 8480 100
rect 8360 10 8405 90
rect 8435 10 8480 90
rect 8360 0 8480 10
rect 8680 90 8800 100
rect 8680 10 8725 90
rect 8755 10 8800 90
rect 8680 0 8800 10
rect 9000 90 9120 100
rect 9000 10 9045 90
rect 9075 10 9120 90
rect 9000 0 9120 10
rect 9320 90 9440 100
rect 9320 10 9365 90
rect 9395 10 9440 90
rect 9320 0 9440 10
rect 9640 90 9760 100
rect 9640 10 9685 90
rect 9715 10 9760 90
rect 9640 0 9760 10
rect 9960 90 10080 100
rect 9960 10 10005 90
rect 10035 10 10080 90
rect 9960 0 10080 10
rect 10280 90 10360 100
rect 10280 10 10325 90
rect 10355 10 10360 90
rect 10280 0 10360 10
<< pdiff >>
rect -80 750 0 760
rect -80 670 -75 750
rect -45 670 0 750
rect -80 660 0 670
rect 200 750 320 760
rect 200 670 245 750
rect 275 670 320 750
rect 200 660 320 670
rect 520 750 640 760
rect 520 670 565 750
rect 595 670 640 750
rect 520 660 640 670
rect 840 750 960 760
rect 840 670 885 750
rect 915 670 960 750
rect 840 660 960 670
rect 1160 750 1280 760
rect 1160 670 1205 750
rect 1235 670 1280 750
rect 1160 660 1280 670
rect 1480 750 1600 760
rect 1480 670 1525 750
rect 1555 670 1600 750
rect 1480 660 1600 670
rect 1800 750 1920 760
rect 1800 670 1845 750
rect 1875 670 1920 750
rect 1800 660 1920 670
rect 2120 750 2240 760
rect 2120 670 2165 750
rect 2195 670 2240 750
rect 2120 660 2240 670
rect 2440 750 2560 760
rect 2440 670 2485 750
rect 2515 670 2560 750
rect 2440 660 2560 670
rect 2760 750 2880 760
rect 2760 670 2805 750
rect 2835 670 2880 750
rect 2760 660 2880 670
rect 3080 750 3200 760
rect 3080 670 3125 750
rect 3155 670 3200 750
rect 3080 660 3200 670
rect 3400 750 3520 760
rect 3400 670 3445 750
rect 3475 670 3520 750
rect 3400 660 3520 670
rect 3720 750 3840 760
rect 3720 670 3765 750
rect 3795 670 3840 750
rect 3720 660 3840 670
rect 4040 750 4160 760
rect 4040 670 4085 750
rect 4115 670 4160 750
rect 4040 660 4160 670
rect 4360 750 4480 760
rect 4360 670 4405 750
rect 4435 670 4480 750
rect 4360 660 4480 670
rect 4680 750 4800 760
rect 4680 670 4725 750
rect 4755 670 4800 750
rect 4680 660 4800 670
rect 5000 750 5080 760
rect 5000 670 5045 750
rect 5075 670 5080 750
rect 5000 660 5080 670
rect 5200 750 5280 760
rect 5200 670 5205 750
rect 5235 670 5280 750
rect 5200 660 5280 670
rect 5480 750 5600 760
rect 5480 670 5525 750
rect 5555 670 5600 750
rect 5480 660 5600 670
rect 5800 750 5920 760
rect 5800 670 5845 750
rect 5875 670 5920 750
rect 5800 660 5920 670
rect 6120 750 6240 760
rect 6120 670 6165 750
rect 6195 670 6240 750
rect 6120 660 6240 670
rect 6440 750 6560 760
rect 6440 670 6485 750
rect 6515 670 6560 750
rect 6440 660 6560 670
rect 6760 750 6880 760
rect 6760 670 6805 750
rect 6835 670 6880 750
rect 6760 660 6880 670
rect 7080 750 7200 760
rect 7080 670 7125 750
rect 7155 670 7200 750
rect 7080 660 7200 670
rect 7400 750 7520 760
rect 7400 670 7445 750
rect 7475 670 7520 750
rect 7400 660 7520 670
rect 7720 750 7840 760
rect 7720 670 7765 750
rect 7795 670 7840 750
rect 7720 660 7840 670
rect 8040 750 8160 760
rect 8040 670 8085 750
rect 8115 670 8160 750
rect 8040 660 8160 670
rect 8360 750 8480 760
rect 8360 670 8405 750
rect 8435 670 8480 750
rect 8360 660 8480 670
rect 8680 750 8800 760
rect 8680 670 8725 750
rect 8755 670 8800 750
rect 8680 660 8800 670
rect 9000 750 9120 760
rect 9000 670 9045 750
rect 9075 670 9120 750
rect 9000 660 9120 670
rect 9320 750 9440 760
rect 9320 670 9365 750
rect 9395 670 9440 750
rect 9320 660 9440 670
rect 9640 750 9760 760
rect 9640 670 9685 750
rect 9715 670 9760 750
rect 9640 660 9760 670
rect 9960 750 10080 760
rect 9960 670 10005 750
rect 10035 670 10080 750
rect 9960 660 10080 670
rect 10280 750 10360 760
rect 10280 670 10325 750
rect 10355 670 10360 750
rect 10280 660 10360 670
<< ndiffc >>
rect -75 10 -45 90
rect 245 10 275 90
rect 565 10 595 90
rect 885 10 915 90
rect 1205 10 1235 90
rect 1525 10 1555 90
rect 1845 10 1875 90
rect 2165 10 2195 90
rect 2485 10 2515 90
rect 2805 10 2835 90
rect 3125 10 3155 90
rect 3445 10 3475 90
rect 3765 10 3795 90
rect 4085 10 4115 90
rect 4405 10 4435 90
rect 4725 10 4755 90
rect 5045 10 5075 90
rect 5205 10 5235 90
rect 5525 10 5555 90
rect 5845 10 5875 90
rect 6165 10 6195 90
rect 6485 10 6515 90
rect 6805 10 6835 90
rect 7125 10 7155 90
rect 7445 10 7475 90
rect 7765 10 7795 90
rect 8085 10 8115 90
rect 8405 10 8435 90
rect 8725 10 8755 90
rect 9045 10 9075 90
rect 9365 10 9395 90
rect 9685 10 9715 90
rect 10005 10 10035 90
rect 10325 10 10355 90
<< pdiffc >>
rect -75 670 -45 750
rect 245 670 275 750
rect 565 670 595 750
rect 885 670 915 750
rect 1205 670 1235 750
rect 1525 670 1555 750
rect 1845 670 1875 750
rect 2165 670 2195 750
rect 2485 670 2515 750
rect 2805 670 2835 750
rect 3125 670 3155 750
rect 3445 670 3475 750
rect 3765 670 3795 750
rect 4085 670 4115 750
rect 4405 670 4435 750
rect 4725 670 4755 750
rect 5045 670 5075 750
rect 5205 670 5235 750
rect 5525 670 5555 750
rect 5845 670 5875 750
rect 6165 670 6195 750
rect 6485 670 6515 750
rect 6805 670 6835 750
rect 7125 670 7155 750
rect 7445 670 7475 750
rect 7765 670 7795 750
rect 8085 670 8115 750
rect 8405 670 8435 750
rect 8725 670 8755 750
rect 9045 670 9075 750
rect 9365 670 9395 750
rect 9685 670 9715 750
rect 10005 670 10035 750
rect 10325 670 10355 750
<< psubdiff >>
rect -320 1000 -40 1040
rect 240 1000 280 1040
rect 560 1000 600 1040
rect 880 1000 920 1040
rect 1200 1000 1240 1040
rect 1520 1000 1560 1040
rect 1840 1000 1880 1040
rect 2160 1000 2200 1040
rect 2480 1000 2520 1040
rect 2800 1000 2840 1040
rect 3120 1000 3160 1040
rect 3440 1000 3480 1040
rect 3760 1000 3800 1040
rect 4080 1000 4120 1040
rect 4400 1000 4440 1040
rect 4720 1000 4760 1040
rect 5040 1000 5240 1040
rect 5520 1000 5560 1040
rect 5840 1000 5880 1040
rect 6160 1000 6200 1040
rect 6480 1000 6520 1040
rect 6800 1000 6840 1040
rect 7120 1000 7160 1040
rect 7440 1000 7480 1040
rect 7760 1000 7800 1040
rect 8080 1000 8120 1040
rect 8400 1000 8440 1040
rect 8720 1000 8760 1040
rect 9040 1000 9080 1040
rect 9360 1000 9400 1040
rect 9680 1000 9720 1040
rect 10000 1000 10040 1040
rect 10320 1000 10640 1040
rect -320 960 -280 1000
rect 10600 960 10640 1000
rect -280 360 -40 400
rect 240 360 280 400
rect 560 360 600 400
rect 880 360 920 400
rect 1200 360 1240 400
rect 1520 360 1560 400
rect 1840 360 1880 400
rect 2160 360 2200 400
rect 2480 360 2520 400
rect 2800 360 2840 400
rect 3120 360 3160 400
rect 3440 360 3480 400
rect 3760 360 3800 400
rect 4080 360 4120 400
rect 4400 360 4440 400
rect 4720 360 4760 400
rect 5040 360 5240 400
rect 5520 360 5560 400
rect 5840 360 5880 400
rect 6160 360 6200 400
rect 6480 360 6520 400
rect 6800 360 6840 400
rect 7120 360 7160 400
rect 7440 360 7480 400
rect 7760 360 7800 400
rect 8080 360 8120 400
rect 8400 360 8440 400
rect 8720 360 8760 400
rect 9040 360 9080 400
rect 9360 360 9400 400
rect 9680 360 9720 400
rect 10000 360 10040 400
rect 10320 360 10600 400
rect -320 -80 -280 -40
rect -160 200 -40 240
rect 240 200 280 240
rect 560 200 600 240
rect 880 200 920 240
rect 1200 200 1240 240
rect 1520 200 1560 240
rect 1840 200 1880 240
rect 2160 200 2200 240
rect 2480 200 2520 240
rect 2800 200 2840 240
rect 3120 200 3160 240
rect 3440 200 3480 240
rect 3760 200 3800 240
rect 4080 200 4120 240
rect 4400 200 4440 240
rect 4720 200 4760 240
rect 5040 200 5240 240
rect 5520 200 5560 240
rect 5840 200 5880 240
rect 6160 200 6200 240
rect 6480 200 6520 240
rect 6800 200 6840 240
rect 7120 200 7160 240
rect 7440 200 7480 240
rect 7760 200 7800 240
rect 8080 200 8120 240
rect 8400 200 8440 240
rect 8720 200 8760 240
rect 9040 200 9080 240
rect 9360 200 9400 240
rect 9680 200 9720 240
rect 10000 200 10040 240
rect 10320 200 10480 240
rect -160 160 -120 200
rect 5120 160 5160 200
rect 10400 160 10440 200
rect -160 -80 -120 -40
rect 5120 -80 5160 -40
rect 10400 -80 10440 -40
rect 10600 -80 10640 -40
rect -320 -120 -40 -80
rect 240 -120 280 -80
rect 560 -120 600 -80
rect 880 -120 920 -80
rect 1200 -120 1240 -80
rect 1520 -120 1560 -80
rect 1840 -120 1880 -80
rect 2160 -120 2200 -80
rect 2480 -120 2520 -80
rect 2800 -120 2840 -80
rect 3120 -120 3160 -80
rect 3440 -120 3480 -80
rect 3760 -120 3800 -80
rect 4080 -120 4120 -80
rect 4400 -120 4440 -80
rect 4720 -120 4760 -80
rect 5040 -120 5240 -80
rect 5520 -120 5560 -80
rect 5840 -120 5880 -80
rect 6160 -120 6200 -80
rect 6480 -120 6520 -80
rect 6800 -120 6840 -80
rect 7120 -120 7160 -80
rect 7440 -120 7480 -80
rect 7760 -120 7800 -80
rect 8080 -120 8120 -80
rect 8400 -120 8440 -80
rect 8720 -120 8760 -80
rect 9040 -120 9080 -80
rect 9360 -120 9400 -80
rect 9680 -120 9720 -80
rect 10000 -120 10040 -80
rect 10320 -120 10640 -80
<< nsubdiff >>
rect -160 840 -40 880
rect 240 840 280 880
rect 560 840 600 880
rect 880 840 920 880
rect 1200 840 1240 880
rect 1520 840 1560 880
rect 1840 840 1880 880
rect 2160 840 2200 880
rect 2480 840 2520 880
rect 2800 840 2840 880
rect 3120 840 3160 880
rect 3440 840 3480 880
rect 3760 840 3800 880
rect 4080 840 4120 880
rect 4400 840 4440 880
rect 4720 840 4760 880
rect 5040 840 5240 880
rect 5520 840 5560 880
rect 5840 840 5880 880
rect 6160 840 6200 880
rect 6480 840 6520 880
rect 6800 840 6840 880
rect 7120 840 7160 880
rect 7440 840 7480 880
rect 7760 840 7800 880
rect 8080 840 8120 880
rect 8400 840 8440 880
rect 8720 840 8760 880
rect 9040 840 9080 880
rect 9360 840 9400 880
rect 9680 840 9720 880
rect 10000 840 10040 880
rect 10320 840 10480 880
rect -160 800 -120 840
rect 5120 800 5160 840
rect 10400 800 10440 840
rect -160 560 -120 600
rect 5120 560 5160 600
rect 10400 560 10440 600
rect -160 520 -40 560
rect 240 520 280 560
rect 560 520 600 560
rect 880 520 920 560
rect 1200 520 1240 560
rect 1520 520 1560 560
rect 1840 520 1880 560
rect 2160 520 2200 560
rect 2480 520 2520 560
rect 2800 520 2840 560
rect 3120 520 3160 560
rect 3440 520 3480 560
rect 3760 520 3800 560
rect 4080 520 4120 560
rect 4400 520 4440 560
rect 4720 520 4760 560
rect 5040 520 5240 560
rect 5520 520 5560 560
rect 5840 520 5880 560
rect 6160 520 6200 560
rect 6480 520 6520 560
rect 6800 520 6840 560
rect 7120 520 7160 560
rect 7440 520 7480 560
rect 7760 520 7800 560
rect 8080 520 8120 560
rect 8400 520 8440 560
rect 8720 520 8760 560
rect 9040 520 9080 560
rect 9360 520 9400 560
rect 9680 520 9720 560
rect 10000 520 10040 560
rect 10320 520 10480 560
<< psubdiffcont >>
rect -40 1000 240 1040
rect 280 1000 560 1040
rect 600 1000 880 1040
rect 920 1000 1200 1040
rect 1240 1000 1520 1040
rect 1560 1000 1840 1040
rect 1880 1000 2160 1040
rect 2200 1000 2480 1040
rect 2520 1000 2800 1040
rect 2840 1000 3120 1040
rect 3160 1000 3440 1040
rect 3480 1000 3760 1040
rect 3800 1000 4080 1040
rect 4120 1000 4400 1040
rect 4440 1000 4720 1040
rect 4760 1000 5040 1040
rect 5240 1000 5520 1040
rect 5560 1000 5840 1040
rect 5880 1000 6160 1040
rect 6200 1000 6480 1040
rect 6520 1000 6800 1040
rect 6840 1000 7120 1040
rect 7160 1000 7440 1040
rect 7480 1000 7760 1040
rect 7800 1000 8080 1040
rect 8120 1000 8400 1040
rect 8440 1000 8720 1040
rect 8760 1000 9040 1040
rect 9080 1000 9360 1040
rect 9400 1000 9680 1040
rect 9720 1000 10000 1040
rect 10040 1000 10320 1040
rect -320 -40 -280 960
rect -40 360 240 400
rect 280 360 560 400
rect 600 360 880 400
rect 920 360 1200 400
rect 1240 360 1520 400
rect 1560 360 1840 400
rect 1880 360 2160 400
rect 2200 360 2480 400
rect 2520 360 2800 400
rect 2840 360 3120 400
rect 3160 360 3440 400
rect 3480 360 3760 400
rect 3800 360 4080 400
rect 4120 360 4400 400
rect 4440 360 4720 400
rect 4760 360 5040 400
rect 5240 360 5520 400
rect 5560 360 5840 400
rect 5880 360 6160 400
rect 6200 360 6480 400
rect 6520 360 6800 400
rect 6840 360 7120 400
rect 7160 360 7440 400
rect 7480 360 7760 400
rect 7800 360 8080 400
rect 8120 360 8400 400
rect 8440 360 8720 400
rect 8760 360 9040 400
rect 9080 360 9360 400
rect 9400 360 9680 400
rect 9720 360 10000 400
rect 10040 360 10320 400
rect -40 200 240 240
rect 280 200 560 240
rect 600 200 880 240
rect 920 200 1200 240
rect 1240 200 1520 240
rect 1560 200 1840 240
rect 1880 200 2160 240
rect 2200 200 2480 240
rect 2520 200 2800 240
rect 2840 200 3120 240
rect 3160 200 3440 240
rect 3480 200 3760 240
rect 3800 200 4080 240
rect 4120 200 4400 240
rect 4440 200 4720 240
rect 4760 200 5040 240
rect 5240 200 5520 240
rect 5560 200 5840 240
rect 5880 200 6160 240
rect 6200 200 6480 240
rect 6520 200 6800 240
rect 6840 200 7120 240
rect 7160 200 7440 240
rect 7480 200 7760 240
rect 7800 200 8080 240
rect 8120 200 8400 240
rect 8440 200 8720 240
rect 8760 200 9040 240
rect 9080 200 9360 240
rect 9400 200 9680 240
rect 9720 200 10000 240
rect 10040 200 10320 240
rect -160 -40 -120 160
rect 5120 -40 5160 160
rect 10400 -40 10440 160
rect 10600 -40 10640 960
rect -40 -120 240 -80
rect 280 -120 560 -80
rect 600 -120 880 -80
rect 920 -120 1200 -80
rect 1240 -120 1520 -80
rect 1560 -120 1840 -80
rect 1880 -120 2160 -80
rect 2200 -120 2480 -80
rect 2520 -120 2800 -80
rect 2840 -120 3120 -80
rect 3160 -120 3440 -80
rect 3480 -120 3760 -80
rect 3800 -120 4080 -80
rect 4120 -120 4400 -80
rect 4440 -120 4720 -80
rect 4760 -120 5040 -80
rect 5240 -120 5520 -80
rect 5560 -120 5840 -80
rect 5880 -120 6160 -80
rect 6200 -120 6480 -80
rect 6520 -120 6800 -80
rect 6840 -120 7120 -80
rect 7160 -120 7440 -80
rect 7480 -120 7760 -80
rect 7800 -120 8080 -80
rect 8120 -120 8400 -80
rect 8440 -120 8720 -80
rect 8760 -120 9040 -80
rect 9080 -120 9360 -80
rect 9400 -120 9680 -80
rect 9720 -120 10000 -80
rect 10040 -120 10320 -80
<< nsubdiffcont >>
rect -40 840 240 880
rect 280 840 560 880
rect 600 840 880 880
rect 920 840 1200 880
rect 1240 840 1520 880
rect 1560 840 1840 880
rect 1880 840 2160 880
rect 2200 840 2480 880
rect 2520 840 2800 880
rect 2840 840 3120 880
rect 3160 840 3440 880
rect 3480 840 3760 880
rect 3800 840 4080 880
rect 4120 840 4400 880
rect 4440 840 4720 880
rect 4760 840 5040 880
rect 5240 840 5520 880
rect 5560 840 5840 880
rect 5880 840 6160 880
rect 6200 840 6480 880
rect 6520 840 6800 880
rect 6840 840 7120 880
rect 7160 840 7440 880
rect 7480 840 7760 880
rect 7800 840 8080 880
rect 8120 840 8400 880
rect 8440 840 8720 880
rect 8760 840 9040 880
rect 9080 840 9360 880
rect 9400 840 9680 880
rect 9720 840 10000 880
rect 10040 840 10320 880
rect -160 600 -120 800
rect 5120 600 5160 800
rect 10400 600 10440 800
rect -40 520 240 560
rect 280 520 560 560
rect 600 520 880 560
rect 920 520 1200 560
rect 1240 520 1520 560
rect 1560 520 1840 560
rect 1880 520 2160 560
rect 2200 520 2480 560
rect 2520 520 2800 560
rect 2840 520 3120 560
rect 3160 520 3440 560
rect 3480 520 3760 560
rect 3800 520 4080 560
rect 4120 520 4400 560
rect 4440 520 4720 560
rect 4760 520 5040 560
rect 5240 520 5520 560
rect 5560 520 5840 560
rect 5880 520 6160 560
rect 6200 520 6480 560
rect 6520 520 6800 560
rect 6840 520 7120 560
rect 7160 520 7440 560
rect 7480 520 7760 560
rect 7800 520 8080 560
rect 8120 520 8400 560
rect 8440 520 8720 560
rect 8760 520 9040 560
rect 9080 520 9360 560
rect 9400 520 9680 560
rect 9720 520 10000 560
rect 10040 520 10320 560
<< poly >>
rect 0 760 200 780
rect 320 760 520 780
rect 640 760 840 780
rect 960 760 1160 780
rect 1280 760 1480 780
rect 1600 760 1800 780
rect 1920 760 2120 780
rect 2240 760 2440 780
rect 2560 760 2760 780
rect 2880 760 3080 780
rect 3200 760 3400 780
rect 3520 760 3720 780
rect 3840 760 4040 780
rect 4160 760 4360 780
rect 4480 760 4680 780
rect 4800 760 5000 780
rect 0 635 200 660
rect 0 605 10 635
rect 190 605 200 635
rect 0 600 200 605
rect 320 635 520 660
rect 320 605 330 635
rect 510 605 520 635
rect 320 600 520 605
rect 640 635 840 660
rect 640 605 650 635
rect 830 605 840 635
rect 640 600 840 605
rect 960 635 1160 660
rect 960 605 970 635
rect 1150 605 1160 635
rect 960 600 1160 605
rect 1280 635 1480 660
rect 1280 605 1290 635
rect 1470 605 1480 635
rect 1280 600 1480 605
rect 1600 635 1800 660
rect 1600 605 1610 635
rect 1790 605 1800 635
rect 1600 600 1800 605
rect 1920 635 2120 660
rect 1920 605 1930 635
rect 2110 605 2120 635
rect 1920 600 2120 605
rect 2240 635 2440 660
rect 2240 605 2250 635
rect 2430 605 2440 635
rect 2240 600 2440 605
rect 2560 635 2760 660
rect 2560 605 2570 635
rect 2750 605 2760 635
rect 2560 600 2760 605
rect 2880 635 3080 660
rect 2880 605 2890 635
rect 3070 605 3080 635
rect 2880 600 3080 605
rect 3200 635 3400 660
rect 3200 605 3210 635
rect 3390 605 3400 635
rect 3200 600 3400 605
rect 3520 635 3720 660
rect 3520 605 3530 635
rect 3710 605 3720 635
rect 3520 600 3720 605
rect 3840 635 4040 660
rect 3840 605 3850 635
rect 4030 605 4040 635
rect 3840 600 4040 605
rect 4160 635 4360 660
rect 4160 605 4170 635
rect 4350 605 4360 635
rect 4160 600 4360 605
rect 4480 635 4680 660
rect 4480 605 4490 635
rect 4670 605 4680 635
rect 4480 600 4680 605
rect 4800 635 5000 660
rect 4800 605 4810 635
rect 4990 605 5000 635
rect 4800 600 5000 605
rect 5280 760 5480 780
rect 5600 760 5800 780
rect 5920 760 6120 780
rect 6240 760 6440 780
rect 6560 760 6760 780
rect 6880 760 7080 780
rect 7200 760 7400 780
rect 7520 760 7720 780
rect 7840 760 8040 780
rect 8160 760 8360 780
rect 8480 760 8680 780
rect 8800 760 9000 780
rect 9120 760 9320 780
rect 9440 760 9640 780
rect 9760 760 9960 780
rect 10080 760 10280 780
rect 5280 635 5480 660
rect 5280 605 5290 635
rect 5470 605 5480 635
rect 5280 600 5480 605
rect 5600 635 5800 660
rect 5600 605 5610 635
rect 5790 605 5800 635
rect 5600 600 5800 605
rect 5920 635 6120 660
rect 5920 605 5930 635
rect 6110 605 6120 635
rect 5920 600 6120 605
rect 6240 635 6440 660
rect 6240 605 6250 635
rect 6430 605 6440 635
rect 6240 600 6440 605
rect 6560 635 6760 660
rect 6560 605 6570 635
rect 6750 605 6760 635
rect 6560 600 6760 605
rect 6880 635 7080 660
rect 6880 605 6890 635
rect 7070 605 7080 635
rect 6880 600 7080 605
rect 7200 635 7400 660
rect 7200 605 7210 635
rect 7390 605 7400 635
rect 7200 600 7400 605
rect 7520 635 7720 660
rect 7520 605 7530 635
rect 7710 605 7720 635
rect 7520 600 7720 605
rect 7840 635 8040 660
rect 7840 605 7850 635
rect 8030 605 8040 635
rect 7840 600 8040 605
rect 8160 635 8360 660
rect 8160 605 8170 635
rect 8350 605 8360 635
rect 8160 600 8360 605
rect 8480 635 8680 660
rect 8480 605 8490 635
rect 8670 605 8680 635
rect 8480 600 8680 605
rect 8800 635 9000 660
rect 8800 605 8810 635
rect 8990 605 9000 635
rect 8800 600 9000 605
rect 9120 635 9320 660
rect 9120 605 9130 635
rect 9310 605 9320 635
rect 9120 600 9320 605
rect 9440 635 9640 660
rect 9440 605 9450 635
rect 9630 605 9640 635
rect 9440 600 9640 605
rect 9760 635 9960 660
rect 9760 605 9770 635
rect 9950 605 9960 635
rect 9760 600 9960 605
rect 10080 635 10280 660
rect 10080 605 10090 635
rect 10270 605 10280 635
rect 10080 600 10280 605
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 100 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 100 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 100 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 100 1160 125
rect 1280 155 1480 160
rect 1280 125 1290 155
rect 1470 125 1480 155
rect 1280 100 1480 125
rect 1600 155 1800 160
rect 1600 125 1610 155
rect 1790 125 1800 155
rect 1600 100 1800 125
rect 1920 155 2120 160
rect 1920 125 1930 155
rect 2110 125 2120 155
rect 1920 100 2120 125
rect 2240 155 2440 160
rect 2240 125 2250 155
rect 2430 125 2440 155
rect 2240 100 2440 125
rect 2560 155 2760 160
rect 2560 125 2570 155
rect 2750 125 2760 155
rect 2560 100 2760 125
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 100 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 100 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 100 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 100 4040 125
rect 4160 155 4360 160
rect 4160 125 4170 155
rect 4350 125 4360 155
rect 4160 100 4360 125
rect 4480 155 4680 160
rect 4480 125 4490 155
rect 4670 125 4680 155
rect 4480 100 4680 125
rect 4800 155 5000 160
rect 4800 125 4810 155
rect 4990 125 5000 155
rect 4800 100 5000 125
rect 0 -20 200 0
rect 320 -20 520 0
rect 640 -20 840 0
rect 960 -20 1160 0
rect 1280 -20 1480 0
rect 1600 -20 1800 0
rect 1920 -20 2120 0
rect 2240 -20 2440 0
rect 2560 -20 2760 0
rect 2880 -20 3080 0
rect 3200 -20 3400 0
rect 3520 -20 3720 0
rect 3840 -20 4040 0
rect 4160 -20 4360 0
rect 4480 -20 4680 0
rect 4800 -20 5000 0
rect 5280 155 5480 160
rect 5280 125 5290 155
rect 5470 125 5480 155
rect 5280 100 5480 125
rect 5600 155 5800 160
rect 5600 125 5610 155
rect 5790 125 5800 155
rect 5600 100 5800 125
rect 5920 155 6120 160
rect 5920 125 5930 155
rect 6110 125 6120 155
rect 5920 100 6120 125
rect 6240 155 6440 160
rect 6240 125 6250 155
rect 6430 125 6440 155
rect 6240 100 6440 125
rect 6560 155 6760 160
rect 6560 125 6570 155
rect 6750 125 6760 155
rect 6560 100 6760 125
rect 6880 155 7080 160
rect 6880 125 6890 155
rect 7070 125 7080 155
rect 6880 100 7080 125
rect 7200 155 7400 160
rect 7200 125 7210 155
rect 7390 125 7400 155
rect 7200 100 7400 125
rect 7520 155 7720 160
rect 7520 125 7530 155
rect 7710 125 7720 155
rect 7520 100 7720 125
rect 7840 155 8040 160
rect 7840 125 7850 155
rect 8030 125 8040 155
rect 7840 100 8040 125
rect 8160 155 8360 160
rect 8160 125 8170 155
rect 8350 125 8360 155
rect 8160 100 8360 125
rect 8480 155 8680 160
rect 8480 125 8490 155
rect 8670 125 8680 155
rect 8480 100 8680 125
rect 8800 155 9000 160
rect 8800 125 8810 155
rect 8990 125 9000 155
rect 8800 100 9000 125
rect 9120 155 9320 160
rect 9120 125 9130 155
rect 9310 125 9320 155
rect 9120 100 9320 125
rect 9440 155 9640 160
rect 9440 125 9450 155
rect 9630 125 9640 155
rect 9440 100 9640 125
rect 9760 155 9960 160
rect 9760 125 9770 155
rect 9950 125 9960 155
rect 9760 100 9960 125
rect 10080 155 10280 160
rect 10080 125 10090 155
rect 10270 125 10280 155
rect 10080 100 10280 125
rect 5280 -20 5480 0
rect 5600 -20 5800 0
rect 5920 -20 6120 0
rect 6240 -20 6440 0
rect 6560 -20 6760 0
rect 6880 -20 7080 0
rect 7200 -20 7400 0
rect 7520 -20 7720 0
rect 7840 -20 8040 0
rect 8160 -20 8360 0
rect 8480 -20 8680 0
rect 8800 -20 9000 0
rect 9120 -20 9320 0
rect 9440 -20 9640 0
rect 9760 -20 9960 0
rect 10080 -20 10280 0
<< polycont >>
rect 10 605 190 635
rect 330 605 510 635
rect 650 605 830 635
rect 970 605 1150 635
rect 1290 605 1470 635
rect 1610 605 1790 635
rect 1930 605 2110 635
rect 2250 605 2430 635
rect 2570 605 2750 635
rect 2890 605 3070 635
rect 3210 605 3390 635
rect 3530 605 3710 635
rect 3850 605 4030 635
rect 4170 605 4350 635
rect 4490 605 4670 635
rect 4810 605 4990 635
rect 5290 605 5470 635
rect 5610 605 5790 635
rect 5930 605 6110 635
rect 6250 605 6430 635
rect 6570 605 6750 635
rect 6890 605 7070 635
rect 7210 605 7390 635
rect 7530 605 7710 635
rect 7850 605 8030 635
rect 8170 605 8350 635
rect 8490 605 8670 635
rect 8810 605 8990 635
rect 9130 605 9310 635
rect 9450 605 9630 635
rect 9770 605 9950 635
rect 10090 605 10270 635
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect 1290 125 1470 155
rect 1610 125 1790 155
rect 1930 125 2110 155
rect 2250 125 2430 155
rect 2570 125 2750 155
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3850 125 4030 155
rect 4170 125 4350 155
rect 4490 125 4670 155
rect 4810 125 4990 155
rect 5290 125 5470 155
rect 5610 125 5790 155
rect 5930 125 6110 155
rect 6250 125 6430 155
rect 6570 125 6750 155
rect 6890 125 7070 155
rect 7210 125 7390 155
rect 7530 125 7710 155
rect 7850 125 8030 155
rect 8170 125 8350 155
rect 8490 125 8670 155
rect 8810 125 8990 155
rect 9130 125 9310 155
rect 9450 125 9630 155
rect 9770 125 9950 155
rect 10090 125 10270 155
<< locali >>
rect -320 1000 -40 1040
rect 240 1000 280 1040
rect 560 1000 600 1040
rect 880 1000 920 1040
rect 1200 1000 1240 1040
rect 1520 1000 1560 1040
rect 1840 1000 1880 1040
rect 2160 1000 2200 1040
rect 2480 1000 2520 1040
rect 2800 1000 2840 1040
rect 3120 1000 3160 1040
rect 3440 1000 3480 1040
rect 3760 1000 3800 1040
rect 4080 1000 4120 1040
rect 4400 1000 4440 1040
rect 4720 1000 4760 1040
rect 5040 1000 5240 1040
rect 5520 1000 5560 1040
rect 5840 1000 5880 1040
rect 6160 1000 6200 1040
rect 6480 1000 6520 1040
rect 6800 1000 6840 1040
rect 7120 1000 7160 1040
rect 7440 1000 7480 1040
rect 7760 1000 7800 1040
rect 8080 1000 8120 1040
rect 8400 1000 8440 1040
rect 8720 1000 8760 1040
rect 9040 1000 9080 1040
rect 9360 1000 9400 1040
rect 9680 1000 9720 1040
rect 10000 1000 10040 1040
rect 10320 1000 10640 1040
rect -320 960 -280 1000
rect 10600 960 10640 1000
rect -160 840 -40 880
rect 240 840 280 880
rect 560 840 600 880
rect 880 840 920 880
rect 1200 840 1240 880
rect 1520 840 1560 880
rect 1840 840 1880 880
rect 2160 840 2200 880
rect 2480 840 2520 880
rect 2800 840 2840 880
rect 3120 840 3160 880
rect 3440 840 3480 880
rect 3760 840 3800 880
rect 4080 840 4120 880
rect 4400 840 4440 880
rect 4720 840 4760 880
rect 5040 840 5240 880
rect 5520 840 5560 880
rect -160 800 -120 840
rect -160 560 -120 600
rect -80 750 -40 840
rect 5120 800 5160 840
rect -80 670 -75 750
rect -45 670 -40 750
rect -80 560 -40 670
rect 240 750 280 760
rect 240 670 245 750
rect 275 670 280 750
rect 240 660 280 670
rect 560 750 600 760
rect 560 670 565 750
rect 595 670 600 750
rect 560 660 600 670
rect 880 750 920 760
rect 880 670 885 750
rect 915 670 920 750
rect 880 660 920 670
rect 1200 750 1240 760
rect 1200 670 1205 750
rect 1235 670 1240 750
rect 1200 660 1240 670
rect 1520 750 1560 760
rect 1520 670 1525 750
rect 1555 670 1560 750
rect 1520 660 1560 670
rect 1840 750 1880 760
rect 1840 670 1845 750
rect 1875 670 1880 750
rect 1840 660 1880 670
rect 2160 750 2200 760
rect 2160 670 2165 750
rect 2195 670 2200 750
rect 2160 660 2200 670
rect 2480 750 2520 760
rect 2480 670 2485 750
rect 2515 670 2520 750
rect 2480 660 2520 670
rect 2800 750 2840 760
rect 2800 670 2805 750
rect 2835 670 2840 750
rect 2800 660 2840 670
rect 3120 750 3160 760
rect 3120 670 3125 750
rect 3155 670 3160 750
rect 3120 660 3160 670
rect 3440 750 3480 760
rect 3440 670 3445 750
rect 3475 670 3480 750
rect 3440 660 3480 670
rect 3760 750 3800 760
rect 3760 670 3765 750
rect 3795 670 3800 750
rect 3760 660 3800 670
rect 4080 750 4120 760
rect 4080 670 4085 750
rect 4115 670 4120 750
rect 4080 660 4120 670
rect 4400 750 4440 760
rect 4400 670 4405 750
rect 4435 670 4440 750
rect 4400 660 4440 670
rect 4720 750 4760 760
rect 4720 670 4725 750
rect 4755 670 4760 750
rect 4720 660 4760 670
rect 5040 750 5080 760
rect 5040 670 5045 750
rect 5075 670 5080 750
rect 5040 660 5080 670
rect 0 635 200 640
rect 0 605 10 635
rect 190 605 200 635
rect 0 600 200 605
rect 320 635 520 640
rect 320 605 330 635
rect 510 605 520 635
rect 320 600 520 605
rect 640 635 840 640
rect 640 605 650 635
rect 830 605 840 635
rect 640 600 840 605
rect 960 635 1160 640
rect 960 605 970 635
rect 1150 605 1160 635
rect 960 600 1160 605
rect 1280 635 1480 640
rect 1280 605 1290 635
rect 1470 605 1480 635
rect 1280 600 1480 605
rect 1600 635 1800 640
rect 1600 605 1610 635
rect 1790 605 1800 635
rect 1600 600 1800 605
rect 1920 635 2120 640
rect 1920 605 1930 635
rect 2110 605 2120 635
rect 1920 600 2120 605
rect 2240 635 2440 640
rect 2240 605 2250 635
rect 2430 605 2440 635
rect 2240 600 2440 605
rect 2560 635 2760 640
rect 2560 605 2570 635
rect 2750 605 2760 635
rect 2560 600 2760 605
rect 2880 635 3080 640
rect 2880 605 2890 635
rect 3070 605 3080 635
rect 2880 600 3080 605
rect 3200 635 3400 640
rect 3200 605 3210 635
rect 3390 605 3400 635
rect 3200 600 3400 605
rect 3520 635 3720 640
rect 3520 605 3530 635
rect 3710 605 3720 635
rect 3520 600 3720 605
rect 3840 635 4040 640
rect 3840 605 3850 635
rect 4030 605 4040 635
rect 3840 600 4040 605
rect 4160 635 4360 640
rect 4160 605 4170 635
rect 4350 605 4360 635
rect 4160 600 4360 605
rect 4480 635 4680 640
rect 4480 605 4490 635
rect 4670 605 4680 635
rect 4480 600 4680 605
rect 4800 635 5000 640
rect 4800 605 4810 635
rect 4990 605 5000 635
rect 4800 600 5000 605
rect 5120 560 5160 600
rect 5200 750 5240 840
rect 5200 670 5205 750
rect 5235 670 5240 750
rect 5200 560 5240 670
rect 5520 750 5560 760
rect 5520 670 5525 750
rect 5555 670 5560 750
rect 5520 660 5560 670
rect 5840 750 5880 880
rect 6160 840 6200 880
rect 5840 670 5845 750
rect 5875 670 5880 750
rect 5280 635 5480 640
rect 5280 605 5290 635
rect 5470 605 5480 635
rect 5280 600 5480 605
rect 5600 635 5800 640
rect 5600 605 5610 635
rect 5790 605 5800 635
rect 5600 600 5800 605
rect -160 520 -40 560
rect 240 520 280 560
rect 560 520 600 560
rect 880 520 920 560
rect 1200 520 1240 560
rect 1520 520 1560 560
rect 1840 520 1880 560
rect 2160 520 2200 560
rect 2480 520 2520 560
rect 2800 520 2840 560
rect 3120 520 3160 560
rect 3440 520 3480 560
rect 3760 520 3800 560
rect 4080 520 4120 560
rect 4400 520 4440 560
rect 4720 520 4760 560
rect 5040 520 5240 560
rect 5520 520 5560 560
rect 5840 520 5880 670
rect 6160 750 6200 760
rect 6160 670 6165 750
rect 6195 670 6200 750
rect 6160 660 6200 670
rect 6480 750 6520 880
rect 6800 840 6840 880
rect 6480 670 6485 750
rect 6515 670 6520 750
rect 5920 635 6120 640
rect 5920 605 5930 635
rect 6110 605 6120 635
rect 5920 600 6120 605
rect 6240 635 6440 640
rect 6240 605 6250 635
rect 6430 605 6440 635
rect 6240 600 6440 605
rect 6160 520 6200 560
rect 6480 520 6520 670
rect 6800 750 6840 760
rect 6800 670 6805 750
rect 6835 670 6840 750
rect 6800 660 6840 670
rect 7120 750 7160 880
rect 7440 840 7480 880
rect 7120 670 7125 750
rect 7155 670 7160 750
rect 6560 635 6760 640
rect 6560 605 6570 635
rect 6750 605 6760 635
rect 6560 600 6760 605
rect 6880 635 7080 640
rect 6880 605 6890 635
rect 7070 605 7080 635
rect 6880 600 7080 605
rect 6800 520 6840 560
rect 7120 520 7160 670
rect 7440 750 7480 760
rect 7440 670 7445 750
rect 7475 670 7480 750
rect 7440 660 7480 670
rect 7760 750 7800 880
rect 8080 840 8120 880
rect 7760 670 7765 750
rect 7795 670 7800 750
rect 7200 635 7400 640
rect 7200 605 7210 635
rect 7390 605 7400 635
rect 7200 600 7400 605
rect 7520 635 7720 640
rect 7520 605 7530 635
rect 7710 605 7720 635
rect 7520 600 7720 605
rect 7440 520 7480 560
rect 7760 520 7800 670
rect 8080 750 8120 760
rect 8080 670 8085 750
rect 8115 670 8120 750
rect 8080 660 8120 670
rect 8400 750 8440 880
rect 8720 840 8760 880
rect 8400 670 8405 750
rect 8435 670 8440 750
rect 7840 635 8040 640
rect 7840 605 7850 635
rect 8030 605 8040 635
rect 7840 600 8040 605
rect 8160 635 8360 640
rect 8160 605 8170 635
rect 8350 605 8360 635
rect 8160 600 8360 605
rect 8080 520 8120 560
rect 8400 520 8440 670
rect 8720 750 8760 760
rect 8720 670 8725 750
rect 8755 670 8760 750
rect 8720 660 8760 670
rect 9040 750 9080 880
rect 9360 840 9400 880
rect 9040 670 9045 750
rect 9075 670 9080 750
rect 8480 635 8680 640
rect 8480 605 8490 635
rect 8670 605 8680 635
rect 8480 600 8680 605
rect 8800 635 9000 640
rect 8800 605 8810 635
rect 8990 605 9000 635
rect 8800 600 9000 605
rect 8720 520 8760 560
rect 9040 520 9080 670
rect 9360 750 9400 760
rect 9360 670 9365 750
rect 9395 670 9400 750
rect 9360 660 9400 670
rect 9680 750 9720 880
rect 10000 840 10040 880
rect 10320 840 10480 880
rect 9680 670 9685 750
rect 9715 670 9720 750
rect 9120 635 9320 640
rect 9120 605 9130 635
rect 9310 605 9320 635
rect 9120 600 9320 605
rect 9440 635 9640 640
rect 9440 605 9450 635
rect 9630 605 9640 635
rect 9440 600 9640 605
rect 9360 520 9400 560
rect 9680 520 9720 670
rect 10000 750 10040 760
rect 10000 670 10005 750
rect 10035 670 10040 750
rect 10000 660 10040 670
rect 10320 750 10360 840
rect 10320 670 10325 750
rect 10355 670 10360 750
rect 9760 635 9960 640
rect 9760 605 9770 635
rect 9950 605 9960 635
rect 9760 600 9960 605
rect 10080 635 10280 640
rect 10080 605 10090 635
rect 10270 605 10280 635
rect 10080 600 10280 605
rect 10320 560 10360 670
rect 10400 800 10440 840
rect 10400 560 10440 600
rect 10000 520 10040 560
rect 10320 520 10480 560
rect -280 360 -40 400
rect 240 360 280 400
rect 560 360 600 400
rect 880 360 920 400
rect 1200 360 1240 400
rect 1520 360 1560 400
rect 1840 360 1880 400
rect 2160 360 2200 400
rect 2480 360 2520 400
rect 2800 360 2840 400
rect 3120 360 3160 400
rect 3440 360 3480 400
rect 3760 360 3800 400
rect 4080 360 4120 400
rect 4400 360 4440 400
rect 4720 360 4760 400
rect 5040 360 5240 400
rect 5520 360 5560 400
rect 5840 360 5880 400
rect 6160 360 6200 400
rect 6480 360 6520 400
rect 6800 360 6840 400
rect 7120 360 7160 400
rect 7440 360 7480 400
rect 7760 360 7800 400
rect 8080 360 8120 400
rect 8400 360 8440 400
rect 8720 360 8760 400
rect 9040 360 9080 400
rect 9360 360 9400 400
rect 9680 360 9720 400
rect 10000 360 10040 400
rect 10320 360 10600 400
rect -320 -80 -280 -40
rect -160 200 -40 240
rect 240 200 280 240
rect 560 200 600 240
rect 880 200 920 240
rect 1200 200 1240 240
rect 1520 200 1560 240
rect 1840 200 1880 240
rect 2160 200 2200 240
rect -160 160 -120 200
rect -160 -80 -120 -40
rect -80 90 -40 200
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 120 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 120 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 120 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 120 1160 125
rect 1280 155 1480 160
rect 1280 125 1290 155
rect 1470 125 1480 155
rect 1280 120 1480 125
rect 1600 155 1800 160
rect 1600 125 1610 155
rect 1790 125 1800 155
rect 1600 120 1800 125
rect 1920 155 2120 160
rect 1920 125 1930 155
rect 2110 125 2120 155
rect 1920 120 2120 125
rect 2240 155 2440 160
rect 2240 125 2250 155
rect 2430 125 2440 155
rect 2240 120 2440 125
rect -80 10 -75 90
rect -45 10 -40 90
rect -80 -80 -40 10
rect 240 90 280 100
rect 240 10 245 90
rect 275 10 280 90
rect 240 0 280 10
rect 560 90 600 100
rect 560 10 565 90
rect 595 10 600 90
rect 560 0 600 10
rect 880 90 920 100
rect 880 10 885 90
rect 915 10 920 90
rect 880 0 920 10
rect 1200 90 1240 100
rect 1200 10 1205 90
rect 1235 10 1240 90
rect 1200 0 1240 10
rect 1520 90 1560 100
rect 1520 10 1525 90
rect 1555 10 1560 90
rect 1520 0 1560 10
rect 1840 90 1880 100
rect 1840 10 1845 90
rect 1875 10 1880 90
rect 1840 0 1880 10
rect 2160 90 2200 100
rect 2160 10 2165 90
rect 2195 10 2200 90
rect 2160 0 2200 10
rect 2480 90 2520 240
rect 2800 200 2840 240
rect 3120 200 3160 240
rect 3440 200 3480 240
rect 3760 200 3800 240
rect 4080 200 4120 240
rect 4400 200 4440 240
rect 4720 200 4760 240
rect 5040 200 5240 240
rect 5520 200 5560 240
rect 5840 200 5880 240
rect 6160 200 6200 240
rect 6480 200 6520 240
rect 6800 200 6840 240
rect 7120 200 7160 240
rect 7440 200 7480 240
rect 2560 155 2760 160
rect 2560 125 2570 155
rect 2750 125 2760 155
rect 2560 120 2760 125
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 120 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 120 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 120 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 120 4040 125
rect 4160 155 4360 160
rect 4160 125 4170 155
rect 4350 125 4360 155
rect 4160 120 4360 125
rect 4480 155 4680 160
rect 4480 125 4490 155
rect 4670 125 4680 155
rect 4480 120 4680 125
rect 4800 155 5000 160
rect 4800 125 4810 155
rect 4990 125 5000 155
rect 4800 120 5000 125
rect 2480 10 2485 90
rect 2515 10 2520 90
rect -320 -120 -40 -80
rect 240 -120 280 -80
rect 560 -120 600 -80
rect 880 -120 920 -80
rect 1200 -120 1240 -80
rect 1520 -120 1560 -80
rect 1840 -120 1880 -80
rect 2160 -120 2200 -80
rect 2480 -120 2520 10
rect 2800 90 2840 100
rect 2800 10 2805 90
rect 2835 10 2840 90
rect 2800 0 2840 10
rect 3120 90 3160 100
rect 3120 10 3125 90
rect 3155 10 3160 90
rect 3120 0 3160 10
rect 3440 90 3480 100
rect 3440 10 3445 90
rect 3475 10 3480 90
rect 3440 0 3480 10
rect 3760 90 3800 100
rect 3760 10 3765 90
rect 3795 10 3800 90
rect 3760 0 3800 10
rect 4080 90 4120 100
rect 4080 10 4085 90
rect 4115 10 4120 90
rect 4080 0 4120 10
rect 4400 90 4440 100
rect 4400 10 4405 90
rect 4435 10 4440 90
rect 4400 0 4440 10
rect 4720 90 4760 100
rect 4720 10 4725 90
rect 4755 10 4760 90
rect 4720 0 4760 10
rect 5040 90 5080 200
rect 5040 10 5045 90
rect 5075 10 5080 90
rect 5040 -80 5080 10
rect 5120 160 5160 200
rect 5120 -80 5160 -40
rect 5200 90 5240 200
rect 5280 155 5480 160
rect 5280 125 5290 155
rect 5470 125 5480 155
rect 5280 120 5480 125
rect 5600 155 5800 160
rect 5600 125 5610 155
rect 5790 125 5800 155
rect 5600 120 5800 125
rect 5920 155 6120 160
rect 5920 125 5930 155
rect 6110 125 6120 155
rect 5920 120 6120 125
rect 6240 155 6440 160
rect 6240 125 6250 155
rect 6430 125 6440 155
rect 6240 120 6440 125
rect 6560 155 6760 160
rect 6560 125 6570 155
rect 6750 125 6760 155
rect 6560 120 6760 125
rect 6880 155 7080 160
rect 6880 125 6890 155
rect 7070 125 7080 155
rect 6880 120 7080 125
rect 7200 155 7400 160
rect 7200 125 7210 155
rect 7390 125 7400 155
rect 7200 120 7400 125
rect 7520 155 7720 160
rect 7520 125 7530 155
rect 7710 125 7720 155
rect 7520 120 7720 125
rect 5200 10 5205 90
rect 5235 10 5240 90
rect 5200 -80 5240 10
rect 5520 90 5560 100
rect 5520 10 5525 90
rect 5555 10 5560 90
rect 5520 0 5560 10
rect 5840 90 5880 100
rect 5840 10 5845 90
rect 5875 10 5880 90
rect 5840 0 5880 10
rect 6160 90 6200 100
rect 6160 10 6165 90
rect 6195 10 6200 90
rect 6160 0 6200 10
rect 6480 90 6520 100
rect 6480 10 6485 90
rect 6515 10 6520 90
rect 6480 0 6520 10
rect 6800 90 6840 100
rect 6800 10 6805 90
rect 6835 10 6840 90
rect 6800 0 6840 10
rect 7120 90 7160 100
rect 7120 10 7125 90
rect 7155 10 7160 90
rect 7120 0 7160 10
rect 7440 90 7480 100
rect 7440 10 7445 90
rect 7475 10 7480 90
rect 7440 0 7480 10
rect 7760 90 7800 240
rect 8080 200 8120 240
rect 8400 200 8440 240
rect 8720 200 8760 240
rect 9040 200 9080 240
rect 9360 200 9400 240
rect 9680 200 9720 240
rect 10000 200 10040 240
rect 10320 200 10480 240
rect 7840 155 8040 160
rect 7840 125 7850 155
rect 8030 125 8040 155
rect 7840 120 8040 125
rect 8160 155 8360 160
rect 8160 125 8170 155
rect 8350 125 8360 155
rect 8160 120 8360 125
rect 8480 155 8680 160
rect 8480 125 8490 155
rect 8670 125 8680 155
rect 8480 120 8680 125
rect 8800 155 9000 160
rect 8800 125 8810 155
rect 8990 125 9000 155
rect 8800 120 9000 125
rect 9120 155 9320 160
rect 9120 125 9130 155
rect 9310 125 9320 155
rect 9120 120 9320 125
rect 9440 155 9640 160
rect 9440 125 9450 155
rect 9630 125 9640 155
rect 9440 120 9640 125
rect 9760 155 9960 160
rect 9760 125 9770 155
rect 9950 125 9960 155
rect 9760 120 9960 125
rect 10080 155 10280 160
rect 10080 125 10090 155
rect 10270 125 10280 155
rect 10080 120 10280 125
rect 7760 10 7765 90
rect 7795 10 7800 90
rect 2800 -120 2840 -80
rect 3120 -120 3160 -80
rect 3440 -120 3480 -80
rect 3760 -120 3800 -80
rect 4080 -120 4120 -80
rect 4400 -120 4440 -80
rect 4720 -120 4760 -80
rect 5040 -120 5240 -80
rect 5520 -120 5560 -80
rect 5840 -120 5880 -80
rect 6160 -120 6200 -80
rect 6480 -120 6520 -80
rect 6800 -120 6840 -80
rect 7120 -120 7160 -80
rect 7440 -120 7480 -80
rect 7760 -120 7800 10
rect 8080 90 8120 100
rect 8080 10 8085 90
rect 8115 10 8120 90
rect 8080 0 8120 10
rect 8400 90 8440 100
rect 8400 10 8405 90
rect 8435 10 8440 90
rect 8400 0 8440 10
rect 8720 90 8760 100
rect 8720 10 8725 90
rect 8755 10 8760 90
rect 8720 0 8760 10
rect 9040 90 9080 100
rect 9040 10 9045 90
rect 9075 10 9080 90
rect 9040 0 9080 10
rect 9360 90 9400 100
rect 9360 10 9365 90
rect 9395 10 9400 90
rect 9360 0 9400 10
rect 9680 90 9720 100
rect 9680 10 9685 90
rect 9715 10 9720 90
rect 9680 0 9720 10
rect 10000 90 10040 100
rect 10000 10 10005 90
rect 10035 10 10040 90
rect 10000 0 10040 10
rect 10320 90 10360 200
rect 10320 10 10325 90
rect 10355 10 10360 90
rect 10320 -80 10360 10
rect 10400 160 10440 200
rect 10400 -80 10440 -40
rect 10600 -80 10640 -40
rect 8080 -120 8120 -80
rect 8400 -120 8440 -80
rect 8720 -120 8760 -80
rect 9040 -120 9080 -80
rect 9360 -120 9400 -80
rect 9680 -120 9720 -80
rect 10000 -120 10040 -80
rect 10320 -120 10640 -80
<< viali >>
rect -75 670 -45 750
rect 245 670 275 750
rect 565 670 595 750
rect 885 670 915 750
rect 1205 670 1235 750
rect 1525 670 1555 750
rect 1845 670 1875 750
rect 2165 670 2195 750
rect 2485 670 2515 750
rect 2805 670 2835 750
rect 3125 670 3155 750
rect 3445 670 3475 750
rect 3765 670 3795 750
rect 4085 670 4115 750
rect 4405 670 4435 750
rect 4725 670 4755 750
rect 5045 670 5075 750
rect 10 605 190 635
rect 330 605 510 635
rect 650 605 830 635
rect 970 605 1150 635
rect 1290 605 1470 635
rect 1610 605 1790 635
rect 1930 605 2110 635
rect 2250 605 2430 635
rect 2570 605 2750 635
rect 2890 605 3070 635
rect 3210 605 3390 635
rect 3530 605 3710 635
rect 3850 605 4030 635
rect 4170 605 4350 635
rect 4490 605 4670 635
rect 4810 605 4990 635
rect 5205 670 5235 750
rect 5525 670 5555 750
rect 5845 670 5875 750
rect 5290 605 5470 635
rect 5610 605 5790 635
rect 6165 670 6195 750
rect 6485 670 6515 750
rect 5930 605 6110 635
rect 6250 605 6430 635
rect 6805 670 6835 750
rect 7125 670 7155 750
rect 6570 605 6750 635
rect 6890 605 7070 635
rect 7445 670 7475 750
rect 7765 670 7795 750
rect 7210 605 7390 635
rect 7530 605 7710 635
rect 8085 670 8115 750
rect 8405 670 8435 750
rect 7850 605 8030 635
rect 8170 605 8350 635
rect 8725 670 8755 750
rect 9045 670 9075 750
rect 8490 605 8670 635
rect 8810 605 8990 635
rect 9365 670 9395 750
rect 9685 670 9715 750
rect 9130 605 9310 635
rect 9450 605 9630 635
rect 10005 670 10035 750
rect 10325 670 10355 750
rect 9770 605 9950 635
rect 10090 605 10270 635
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect 1290 125 1470 155
rect 1610 125 1790 155
rect 1930 125 2110 155
rect 2250 125 2430 155
rect -75 10 -45 90
rect 245 10 275 90
rect 565 10 595 90
rect 885 10 915 90
rect 1205 10 1235 90
rect 1525 10 1555 90
rect 1845 10 1875 90
rect 2165 10 2195 90
rect 2570 125 2750 155
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3850 125 4030 155
rect 4170 125 4350 155
rect 4490 125 4670 155
rect 4810 125 4990 155
rect 2485 10 2515 90
rect 2805 10 2835 90
rect 3125 10 3155 90
rect 3445 10 3475 90
rect 3765 10 3795 90
rect 4085 10 4115 90
rect 4405 10 4435 90
rect 4725 10 4755 90
rect 5045 10 5075 90
rect 5290 125 5470 155
rect 5610 125 5790 155
rect 5930 125 6110 155
rect 6250 125 6430 155
rect 6570 125 6750 155
rect 6890 125 7070 155
rect 7210 125 7390 155
rect 7530 125 7710 155
rect 5205 10 5235 90
rect 5525 10 5555 90
rect 5845 10 5875 90
rect 6165 10 6195 90
rect 6485 10 6515 90
rect 6805 10 6835 90
rect 7125 10 7155 90
rect 7445 10 7475 90
rect 7850 125 8030 155
rect 8170 125 8350 155
rect 8490 125 8670 155
rect 8810 125 8990 155
rect 9130 125 9310 155
rect 9450 125 9630 155
rect 9770 125 9950 155
rect 10090 125 10270 155
rect 7765 10 7795 90
rect 8085 10 8115 90
rect 8405 10 8435 90
rect 8725 10 8755 90
rect 9045 10 9075 90
rect 9365 10 9395 90
rect 9685 10 9715 90
rect 10005 10 10035 90
rect 10325 10 10355 90
<< metal1 >>
rect -80 795 -40 800
rect -80 765 -75 795
rect -45 765 -40 795
rect -80 750 -40 765
rect 5200 795 5240 800
rect 5200 765 5205 795
rect 5235 765 5240 795
rect -80 670 -75 750
rect -45 670 -40 750
rect -80 660 -40 670
rect 240 750 280 760
rect 240 670 245 750
rect 275 670 280 750
rect 240 660 280 670
rect 560 750 600 760
rect 560 670 565 750
rect 595 670 600 750
rect 560 660 600 670
rect 880 750 920 760
rect 880 670 885 750
rect 915 670 920 750
rect 880 660 920 670
rect 1200 750 1240 760
rect 1200 670 1205 750
rect 1235 670 1240 750
rect 1200 660 1240 670
rect 1520 750 1560 760
rect 1520 670 1525 750
rect 1555 670 1560 750
rect 1520 660 1560 670
rect 1840 750 1880 760
rect 1840 670 1845 750
rect 1875 670 1880 750
rect 1840 660 1880 670
rect 2160 750 2200 760
rect 2160 670 2165 750
rect 2195 670 2200 750
rect 2160 660 2200 670
rect 2480 750 2520 760
rect 2480 670 2485 750
rect 2515 670 2520 750
rect 2480 660 2520 670
rect 2800 750 2840 760
rect 2800 670 2805 750
rect 2835 670 2840 750
rect 2800 660 2840 670
rect 3120 750 3160 760
rect 3120 670 3125 750
rect 3155 670 3160 750
rect 3120 660 3160 670
rect 3440 750 3480 760
rect 3440 670 3445 750
rect 3475 670 3480 750
rect 3440 660 3480 670
rect 3760 750 3800 760
rect 3760 670 3765 750
rect 3795 670 3800 750
rect 3760 660 3800 670
rect 4080 750 4120 760
rect 4080 670 4085 750
rect 4115 670 4120 750
rect 4080 660 4120 670
rect 4400 750 4440 760
rect 4400 670 4405 750
rect 4435 670 4440 750
rect 4400 660 4440 670
rect 4720 750 4760 760
rect 4720 670 4725 750
rect 4755 670 4760 750
rect 4720 660 4760 670
rect 5040 750 5080 760
rect 5040 670 5045 750
rect 5075 670 5080 750
rect 0 635 200 640
rect 0 605 10 635
rect 190 605 200 635
rect 0 600 200 605
rect 320 635 520 640
rect 320 605 330 635
rect 510 605 520 635
rect 320 600 520 605
rect 640 635 840 640
rect 640 605 650 635
rect 830 605 840 635
rect 640 600 840 605
rect 960 635 1160 640
rect 960 605 970 635
rect 1150 605 1160 635
rect 960 600 1160 605
rect 1280 635 1480 640
rect 1280 605 1290 635
rect 1470 605 1480 635
rect 1280 600 1480 605
rect 1600 635 1800 640
rect 1600 605 1610 635
rect 1790 605 1800 635
rect 1600 600 1800 605
rect 1920 635 2120 640
rect 1920 605 1930 635
rect 2110 605 2120 635
rect 1920 600 2120 605
rect 2240 635 2440 640
rect 2240 605 2250 635
rect 2430 605 2440 635
rect 2240 600 2440 605
rect 2560 635 2760 640
rect 2560 605 2570 635
rect 2750 605 2760 635
rect 2560 600 2760 605
rect 2880 635 3080 640
rect 2880 605 2890 635
rect 3070 605 3080 635
rect 2880 600 3080 605
rect 3200 635 3400 640
rect 3200 605 3210 635
rect 3390 605 3400 635
rect 3200 600 3400 605
rect 3520 635 3720 640
rect 3520 605 3530 635
rect 3710 605 3720 635
rect 3520 600 3720 605
rect 3840 635 4040 640
rect 3840 605 3850 635
rect 4030 605 4040 635
rect 3840 600 4040 605
rect 4160 635 4360 640
rect 4160 605 4170 635
rect 4350 605 4360 635
rect 4160 600 4360 605
rect 4480 635 4680 640
rect 4480 605 4490 635
rect 4670 605 4680 635
rect 4480 600 4680 605
rect 4800 635 5000 640
rect 4800 605 4810 635
rect 4990 605 5000 635
rect 4800 600 5000 605
rect 80 475 120 600
rect 80 445 85 475
rect 115 445 120 475
rect 80 440 120 445
rect 400 475 440 600
rect 400 445 405 475
rect 435 445 440 475
rect 400 440 440 445
rect 720 475 760 600
rect 720 445 725 475
rect 755 445 760 475
rect 720 440 760 445
rect 1040 475 1080 600
rect 1040 445 1045 475
rect 1075 445 1080 475
rect 1040 440 1080 445
rect 1360 475 1400 600
rect 1360 445 1365 475
rect 1395 445 1400 475
rect 1360 440 1400 445
rect 1680 475 1720 600
rect 1680 445 1685 475
rect 1715 445 1720 475
rect 1680 440 1720 445
rect 2000 475 2040 600
rect 2000 445 2005 475
rect 2035 445 2040 475
rect 2000 440 2040 445
rect 2320 475 2360 600
rect 2320 445 2325 475
rect 2355 445 2360 475
rect 2320 440 2360 445
rect 2640 475 2680 600
rect 2640 445 2645 475
rect 2675 445 2680 475
rect 2640 440 2680 445
rect 2960 475 3000 600
rect 2960 445 2965 475
rect 2995 445 3000 475
rect 2960 440 3000 445
rect 3280 475 3320 600
rect 3280 445 3285 475
rect 3315 445 3320 475
rect 3280 440 3320 445
rect 3600 475 3640 600
rect 3600 445 3605 475
rect 3635 445 3640 475
rect 3600 440 3640 445
rect 3920 475 3960 600
rect 3920 445 3925 475
rect 3955 445 3960 475
rect 3920 440 3960 445
rect 4240 475 4280 600
rect 4240 445 4245 475
rect 4275 445 4280 475
rect 4240 440 4280 445
rect 4560 475 4600 600
rect 4560 445 4565 475
rect 4595 445 4600 475
rect 4560 440 4600 445
rect 4880 475 4920 600
rect 4880 445 4885 475
rect 4915 445 4920 475
rect 4880 440 4920 445
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 120 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 120 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 120 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 120 1160 125
rect 1200 155 1240 160
rect 1200 125 1205 155
rect 1235 125 1240 155
rect -80 90 -40 100
rect -80 10 -75 90
rect -45 10 -40 90
rect -80 -5 -40 10
rect 240 90 280 100
rect 240 10 245 90
rect 275 10 280 90
rect 240 0 280 10
rect 560 90 600 100
rect 560 10 565 90
rect 595 10 600 90
rect 560 0 600 10
rect 880 90 920 100
rect 880 10 885 90
rect 915 10 920 90
rect 880 0 920 10
rect 1200 90 1240 125
rect 1280 155 1480 160
rect 1280 125 1290 155
rect 1470 125 1480 155
rect 1280 120 1480 125
rect 1600 155 1800 160
rect 1600 125 1610 155
rect 1790 125 1800 155
rect 1600 120 1800 125
rect 1920 155 2120 160
rect 1920 125 1930 155
rect 2110 125 2120 155
rect 1920 120 2120 125
rect 2240 155 2440 160
rect 2240 125 2250 155
rect 2430 125 2440 155
rect 2240 120 2440 125
rect 2560 155 2760 160
rect 2560 125 2570 155
rect 2750 125 2760 155
rect 2560 120 2760 125
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 120 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 120 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 120 3720 125
rect 3760 155 3800 160
rect 3760 125 3765 155
rect 3795 125 3800 155
rect 1200 10 1205 90
rect 1235 10 1240 90
rect 1200 0 1240 10
rect 1520 90 1560 100
rect 1520 10 1525 90
rect 1555 10 1560 90
rect 1520 0 1560 10
rect 1840 90 1880 100
rect 1840 10 1845 90
rect 1875 10 1880 90
rect 1840 0 1880 10
rect 2160 90 2200 100
rect 2160 10 2165 90
rect 2195 10 2200 90
rect 2160 0 2200 10
rect 2480 90 2520 100
rect 2480 10 2485 90
rect 2515 10 2520 90
rect -80 -35 -75 -5
rect -45 -35 -40 -5
rect -80 -40 -40 -35
rect 2480 -5 2520 10
rect 2800 90 2840 100
rect 2800 10 2805 90
rect 2835 10 2840 90
rect 2800 0 2840 10
rect 3120 90 3160 100
rect 3120 10 3125 90
rect 3155 10 3160 90
rect 3120 0 3160 10
rect 3440 90 3480 100
rect 3440 10 3445 90
rect 3475 10 3480 90
rect 3440 0 3480 10
rect 3760 90 3800 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 120 4040 125
rect 4160 155 4360 160
rect 4160 125 4170 155
rect 4350 125 4360 155
rect 4160 120 4360 125
rect 4480 155 4680 160
rect 4480 125 4490 155
rect 4670 125 4680 155
rect 4480 120 4680 125
rect 4800 155 5000 160
rect 4800 125 4810 155
rect 4990 125 5000 155
rect 4800 120 5000 125
rect 5040 155 5080 670
rect 5200 750 5240 765
rect 5840 795 5880 800
rect 5840 765 5845 795
rect 5875 765 5880 795
rect 5200 670 5205 750
rect 5235 670 5240 750
rect 5200 660 5240 670
rect 5520 750 5560 760
rect 5520 670 5525 750
rect 5555 670 5560 750
rect 5280 635 5480 640
rect 5280 605 5290 635
rect 5470 605 5480 635
rect 5280 600 5480 605
rect 5360 315 5400 600
rect 5360 285 5365 315
rect 5395 285 5400 315
rect 5360 280 5400 285
rect 5520 315 5560 670
rect 5840 750 5880 765
rect 6480 795 6520 800
rect 6480 765 6485 795
rect 6515 765 6520 795
rect 5840 670 5845 750
rect 5875 670 5880 750
rect 5840 660 5880 670
rect 6160 750 6200 760
rect 6160 670 6165 750
rect 6195 670 6200 750
rect 6160 660 6200 670
rect 6480 750 6520 765
rect 7120 795 7160 800
rect 7120 765 7125 795
rect 7155 765 7160 795
rect 6480 670 6485 750
rect 6515 670 6520 750
rect 6480 660 6520 670
rect 6800 750 6840 760
rect 6800 670 6805 750
rect 6835 670 6840 750
rect 6800 660 6840 670
rect 7120 750 7160 765
rect 7760 795 7800 800
rect 7760 765 7765 795
rect 7795 765 7800 795
rect 7120 670 7125 750
rect 7155 670 7160 750
rect 7120 660 7160 670
rect 7440 750 7480 760
rect 7440 670 7445 750
rect 7475 670 7480 750
rect 7440 660 7480 670
rect 7760 750 7800 765
rect 8400 795 8440 800
rect 8400 765 8405 795
rect 8435 765 8440 795
rect 7760 670 7765 750
rect 7795 670 7800 750
rect 7760 660 7800 670
rect 8080 750 8120 760
rect 8080 670 8085 750
rect 8115 670 8120 750
rect 8080 660 8120 670
rect 8400 750 8440 765
rect 9040 795 9080 800
rect 9040 765 9045 795
rect 9075 765 9080 795
rect 8400 670 8405 750
rect 8435 670 8440 750
rect 8400 660 8440 670
rect 8720 750 8760 760
rect 8720 670 8725 750
rect 8755 670 8760 750
rect 8720 660 8760 670
rect 9040 750 9080 765
rect 9680 795 9720 800
rect 9680 765 9685 795
rect 9715 765 9720 795
rect 9040 670 9045 750
rect 9075 670 9080 750
rect 9040 660 9080 670
rect 9360 750 9400 760
rect 9360 670 9365 750
rect 9395 670 9400 750
rect 9360 660 9400 670
rect 9680 750 9720 765
rect 10320 795 10360 800
rect 10320 765 10325 795
rect 10355 765 10360 795
rect 9680 670 9685 750
rect 9715 670 9720 750
rect 9680 660 9720 670
rect 10000 750 10040 760
rect 10000 670 10005 750
rect 10035 670 10040 750
rect 10000 660 10040 670
rect 10320 750 10360 765
rect 10320 670 10325 750
rect 10355 670 10360 750
rect 10320 660 10360 670
rect 5600 635 5800 640
rect 5600 605 5610 635
rect 5790 605 5800 635
rect 5600 600 5800 605
rect 5920 635 6120 640
rect 5920 605 5930 635
rect 6110 605 6120 635
rect 5920 600 6120 605
rect 6240 635 6440 640
rect 6240 605 6250 635
rect 6430 605 6440 635
rect 6240 600 6440 605
rect 6560 635 6760 640
rect 6560 605 6570 635
rect 6750 605 6760 635
rect 6560 600 6760 605
rect 6880 635 7080 640
rect 6880 605 6890 635
rect 7070 605 7080 635
rect 6880 600 7080 605
rect 7200 635 7400 640
rect 7200 605 7210 635
rect 7390 605 7400 635
rect 7200 600 7400 605
rect 7520 635 7720 640
rect 7520 605 7530 635
rect 7710 605 7720 635
rect 7520 600 7720 605
rect 7840 635 8040 640
rect 7840 605 7850 635
rect 8030 605 8040 635
rect 7840 600 8040 605
rect 8160 635 8360 640
rect 8160 605 8170 635
rect 8350 605 8360 635
rect 8160 600 8360 605
rect 8480 635 8680 640
rect 8480 605 8490 635
rect 8670 605 8680 635
rect 8480 600 8680 605
rect 8800 635 9000 640
rect 8800 605 8810 635
rect 8990 605 9000 635
rect 8800 600 9000 605
rect 9120 635 9320 640
rect 9120 605 9130 635
rect 9310 605 9320 635
rect 9120 600 9320 605
rect 9440 635 9640 640
rect 9440 605 9450 635
rect 9630 605 9640 635
rect 9440 600 9640 605
rect 9760 635 9960 640
rect 9760 605 9770 635
rect 9950 605 9960 635
rect 9760 600 9960 605
rect 10080 635 10280 640
rect 10080 605 10090 635
rect 10270 605 10280 635
rect 10080 600 10280 605
rect 5520 285 5525 315
rect 5555 285 5560 315
rect 5520 280 5560 285
rect 5680 315 5720 600
rect 5680 285 5685 315
rect 5715 285 5720 315
rect 5680 280 5720 285
rect 6000 315 6040 600
rect 6000 285 6005 315
rect 6035 285 6040 315
rect 6000 280 6040 285
rect 6160 315 6200 600
rect 6160 285 6165 315
rect 6195 285 6200 315
rect 6160 280 6200 285
rect 6320 315 6360 600
rect 6320 285 6325 315
rect 6355 285 6360 315
rect 6320 280 6360 285
rect 6480 315 6520 320
rect 6480 285 6485 315
rect 6515 285 6520 315
rect 5040 125 5045 155
rect 5075 125 5080 155
rect 5040 120 5080 125
rect 5280 155 5480 160
rect 5280 125 5290 155
rect 5470 125 5480 155
rect 5280 120 5480 125
rect 5600 155 5800 160
rect 5600 125 5610 155
rect 5790 125 5800 155
rect 5600 120 5800 125
rect 5920 155 6120 160
rect 5920 125 5930 155
rect 6110 125 6120 155
rect 5920 120 6120 125
rect 6240 155 6440 160
rect 6240 125 6250 155
rect 6430 125 6440 155
rect 6240 120 6440 125
rect 3760 10 3765 90
rect 3795 10 3800 90
rect 3760 0 3800 10
rect 4080 90 4120 100
rect 4080 10 4085 90
rect 4115 10 4120 90
rect 4080 0 4120 10
rect 4400 90 4440 100
rect 4400 10 4405 90
rect 4435 10 4440 90
rect 4400 0 4440 10
rect 4720 90 4760 100
rect 4720 10 4725 90
rect 4755 10 4760 90
rect 4720 0 4760 10
rect 5040 90 5080 100
rect 5040 10 5045 90
rect 5075 10 5080 90
rect 2480 -35 2485 -5
rect 2515 -35 2520 -5
rect 2480 -40 2520 -35
rect 5040 -5 5080 10
rect 5040 -35 5045 -5
rect 5075 -35 5080 -5
rect 5040 -40 5080 -35
rect 5200 90 5240 100
rect 5200 10 5205 90
rect 5235 10 5240 90
rect 5200 -5 5240 10
rect 5520 90 5560 100
rect 5520 10 5525 90
rect 5555 10 5560 90
rect 5520 0 5560 10
rect 5840 90 5880 100
rect 5840 10 5845 90
rect 5875 10 5880 90
rect 5840 0 5880 10
rect 6160 90 6200 100
rect 6160 10 6165 90
rect 6195 10 6200 90
rect 6160 0 6200 10
rect 6480 90 6520 285
rect 6640 315 6680 600
rect 6640 285 6645 315
rect 6675 285 6680 315
rect 6640 280 6680 285
rect 6800 315 6840 600
rect 6800 285 6805 315
rect 6835 285 6840 315
rect 6800 280 6840 285
rect 6960 315 7000 600
rect 6960 285 6965 315
rect 6995 285 7000 315
rect 6960 280 7000 285
rect 7280 315 7320 600
rect 7280 285 7285 315
rect 7315 285 7320 315
rect 7280 280 7320 285
rect 7440 315 7480 600
rect 7440 285 7445 315
rect 7475 285 7480 315
rect 7440 280 7480 285
rect 7600 315 7640 600
rect 7600 285 7605 315
rect 7635 285 7640 315
rect 7600 280 7640 285
rect 7920 315 7960 600
rect 7920 285 7925 315
rect 7955 285 7960 315
rect 7920 280 7960 285
rect 8080 315 8120 600
rect 8080 285 8085 315
rect 8115 285 8120 315
rect 8080 280 8120 285
rect 8240 315 8280 600
rect 8240 285 8245 315
rect 8275 285 8280 315
rect 8240 280 8280 285
rect 8560 315 8600 600
rect 8560 285 8565 315
rect 8595 285 8600 315
rect 8560 280 8600 285
rect 8720 315 8760 600
rect 8720 285 8725 315
rect 8755 285 8760 315
rect 8720 280 8760 285
rect 8880 315 8920 600
rect 8880 285 8885 315
rect 8915 285 8920 315
rect 8880 280 8920 285
rect 9040 315 9080 320
rect 9040 285 9045 315
rect 9075 285 9080 315
rect 6560 155 6760 160
rect 6560 125 6570 155
rect 6750 125 6760 155
rect 6560 120 6760 125
rect 6880 155 7080 160
rect 6880 125 6890 155
rect 7070 125 7080 155
rect 6880 120 7080 125
rect 7200 155 7400 160
rect 7200 125 7210 155
rect 7390 125 7400 155
rect 7200 120 7400 125
rect 7520 155 7720 160
rect 7520 125 7530 155
rect 7710 125 7720 155
rect 7520 120 7720 125
rect 7840 155 8040 160
rect 7840 125 7850 155
rect 8030 125 8040 155
rect 7840 120 8040 125
rect 8160 155 8360 160
rect 8160 125 8170 155
rect 8350 125 8360 155
rect 8160 120 8360 125
rect 8480 155 8680 160
rect 8480 125 8490 155
rect 8670 125 8680 155
rect 8480 120 8680 125
rect 8800 155 9000 160
rect 8800 125 8810 155
rect 8990 125 9000 155
rect 8800 120 9000 125
rect 6480 10 6485 90
rect 6515 10 6520 90
rect 6480 0 6520 10
rect 6800 90 6840 100
rect 6800 10 6805 90
rect 6835 10 6840 90
rect 6800 0 6840 10
rect 7120 90 7160 100
rect 7120 10 7125 90
rect 7155 10 7160 90
rect 7120 0 7160 10
rect 7440 90 7480 100
rect 7440 10 7445 90
rect 7475 10 7480 90
rect 7440 0 7480 10
rect 7760 90 7800 100
rect 7760 10 7765 90
rect 7795 10 7800 90
rect 5200 -35 5205 -5
rect 5235 -35 5240 -5
rect 5200 -40 5240 -35
rect 7760 -5 7800 10
rect 8080 90 8120 100
rect 8080 10 8085 90
rect 8115 10 8120 90
rect 8080 0 8120 10
rect 8400 90 8440 100
rect 8400 10 8405 90
rect 8435 10 8440 90
rect 8400 0 8440 10
rect 8720 90 8760 100
rect 8720 10 8725 90
rect 8755 10 8760 90
rect 8720 0 8760 10
rect 9040 90 9080 285
rect 9200 315 9240 600
rect 9200 285 9205 315
rect 9235 285 9240 315
rect 9200 280 9240 285
rect 9360 315 9400 600
rect 9360 285 9365 315
rect 9395 285 9400 315
rect 9360 280 9400 285
rect 9520 315 9560 600
rect 9520 285 9525 315
rect 9555 285 9560 315
rect 9520 280 9560 285
rect 9840 315 9880 600
rect 9840 285 9845 315
rect 9875 285 9880 315
rect 9840 280 9880 285
rect 10000 315 10040 600
rect 10000 285 10005 315
rect 10035 285 10040 315
rect 10000 280 10040 285
rect 10160 315 10200 600
rect 10160 285 10165 315
rect 10195 285 10200 315
rect 10160 280 10200 285
rect 9120 155 9320 160
rect 9120 125 9130 155
rect 9310 125 9320 155
rect 9120 120 9320 125
rect 9440 155 9640 160
rect 9440 125 9450 155
rect 9630 125 9640 155
rect 9440 120 9640 125
rect 9760 155 9960 160
rect 9760 125 9770 155
rect 9950 125 9960 155
rect 9760 120 9960 125
rect 10080 155 10280 160
rect 10080 125 10090 155
rect 10270 125 10280 155
rect 10080 120 10280 125
rect 9040 10 9045 90
rect 9075 10 9080 90
rect 9040 0 9080 10
rect 9360 90 9400 100
rect 9360 10 9365 90
rect 9395 10 9400 90
rect 9360 0 9400 10
rect 9680 90 9720 100
rect 9680 10 9685 90
rect 9715 10 9720 90
rect 9680 0 9720 10
rect 10000 90 10040 100
rect 10000 10 10005 90
rect 10035 10 10040 90
rect 10000 0 10040 10
rect 10320 90 10360 100
rect 10320 10 10325 90
rect 10355 10 10360 90
rect 7760 -35 7765 -5
rect 7795 -35 7800 -5
rect 7760 -40 7800 -35
rect 10320 -5 10360 10
rect 10320 -35 10325 -5
rect 10355 -35 10360 -5
rect 10320 -40 10360 -35
<< via1 >>
rect -75 765 -45 795
rect 5205 765 5235 795
rect -75 685 -45 715
rect 85 445 115 475
rect 405 445 435 475
rect 725 445 755 475
rect 1045 445 1075 475
rect 1365 445 1395 475
rect 1685 445 1715 475
rect 2005 445 2035 475
rect 2325 445 2355 475
rect 2645 445 2675 475
rect 2965 445 2995 475
rect 3285 445 3315 475
rect 3605 445 3635 475
rect 3925 445 3955 475
rect 4245 445 4275 475
rect 4565 445 4595 475
rect 4885 445 4915 475
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect 1205 125 1235 155
rect -75 45 -45 75
rect 1290 125 1470 155
rect 1610 125 1790 155
rect 1930 125 2110 155
rect 2250 125 2430 155
rect 2570 125 2750 155
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3765 125 3795 155
rect 2485 45 2515 75
rect -75 -35 -45 -5
rect 3850 125 4030 155
rect 4170 125 4350 155
rect 4490 125 4670 155
rect 4810 125 4990 155
rect 5845 765 5875 795
rect 5205 685 5235 715
rect 5365 285 5395 315
rect 6485 765 6515 795
rect 5845 685 5875 715
rect 7125 765 7155 795
rect 6485 685 6515 715
rect 7765 765 7795 795
rect 7125 685 7155 715
rect 8405 765 8435 795
rect 7765 685 7795 715
rect 9045 765 9075 795
rect 8405 685 8435 715
rect 9685 765 9715 795
rect 9045 685 9075 715
rect 10325 765 10355 795
rect 9685 685 9715 715
rect 10325 685 10355 715
rect 5525 285 5555 315
rect 5685 285 5715 315
rect 6005 285 6035 315
rect 6165 285 6195 315
rect 6325 285 6355 315
rect 6485 285 6515 315
rect 5045 125 5075 155
rect 5290 125 5470 155
rect 5610 125 5790 155
rect 5930 125 6110 155
rect 6250 125 6430 155
rect 5045 45 5075 75
rect 2485 -35 2515 -5
rect 5045 -35 5075 -5
rect 5205 45 5235 75
rect 6645 285 6675 315
rect 6805 285 6835 315
rect 6965 285 6995 315
rect 7285 285 7315 315
rect 7445 285 7475 315
rect 7605 285 7635 315
rect 7925 285 7955 315
rect 8085 285 8115 315
rect 8245 285 8275 315
rect 8565 285 8595 315
rect 8725 285 8755 315
rect 8885 285 8915 315
rect 9045 285 9075 315
rect 6570 125 6750 155
rect 6890 125 7070 155
rect 7210 125 7390 155
rect 7530 125 7710 155
rect 7850 125 8030 155
rect 8170 125 8350 155
rect 8490 125 8670 155
rect 8810 125 8990 155
rect 7765 45 7795 75
rect 5205 -35 5235 -5
rect 9205 285 9235 315
rect 9365 285 9395 315
rect 9525 285 9555 315
rect 9845 285 9875 315
rect 10005 285 10035 315
rect 10165 285 10195 315
rect 9130 125 9310 155
rect 9450 125 9630 155
rect 9770 125 9950 155
rect 10090 125 10270 155
rect 10325 45 10355 75
rect 7765 -35 7795 -5
rect 10325 -35 10355 -5
<< metal2 >>
rect -720 1035 10640 1040
rect -720 1005 -715 1035
rect -685 1005 10640 1035
rect -720 1000 10640 1005
rect -320 920 10640 960
rect -320 840 10640 880
rect -640 795 10640 800
rect -640 765 -635 795
rect -605 765 -75 795
rect -45 765 5205 795
rect 5235 765 5845 795
rect 5875 765 6485 795
rect 6515 765 7125 795
rect 7155 765 7765 795
rect 7795 765 8405 795
rect 8435 765 9045 795
rect 9075 765 9685 795
rect 9715 765 10325 795
rect 10355 765 10640 795
rect -640 760 10640 765
rect -640 715 10640 720
rect -640 685 -635 715
rect -605 685 -75 715
rect -45 685 5205 715
rect 5235 685 5845 715
rect 5875 685 6485 715
rect 6515 685 7125 715
rect 7155 685 7765 715
rect 7795 685 8405 715
rect 8435 685 9045 715
rect 9075 685 9685 715
rect 9715 685 10325 715
rect 10355 685 10640 715
rect -640 680 10640 685
rect -320 600 10640 640
rect -320 520 10640 560
rect -480 475 10640 480
rect -480 445 -475 475
rect -445 445 85 475
rect 115 445 405 475
rect 435 445 725 475
rect 755 445 1045 475
rect 1075 445 1365 475
rect 1395 445 1685 475
rect 1715 445 2005 475
rect 2035 445 2325 475
rect 2355 445 2645 475
rect 2675 445 2965 475
rect 2995 445 3285 475
rect 3315 445 3605 475
rect 3635 445 3925 475
rect 3955 445 4245 475
rect 4275 445 4565 475
rect 4595 445 4885 475
rect 4915 445 10640 475
rect -480 440 10640 445
rect -320 360 10640 400
rect -320 315 10960 320
rect -320 285 5365 315
rect 5395 285 5525 315
rect 5555 285 5685 315
rect 5715 285 6005 315
rect 6035 285 6165 315
rect 6195 285 6325 315
rect 6355 285 6485 315
rect 6515 285 6645 315
rect 6675 285 6805 315
rect 6835 285 6965 315
rect 6995 285 7285 315
rect 7315 285 7445 315
rect 7475 285 7605 315
rect 7635 285 7925 315
rect 7955 285 8085 315
rect 8115 285 8245 315
rect 8275 285 8565 315
rect 8595 285 8725 315
rect 8755 285 8885 315
rect 8915 285 9045 315
rect 9075 285 9205 315
rect 9235 285 9365 315
rect 9395 285 9525 315
rect 9555 285 9845 315
rect 9875 285 10005 315
rect 10035 285 10165 315
rect 10195 285 10925 315
rect 10955 285 10960 315
rect -320 280 10960 285
rect -720 235 11040 240
rect -720 205 -715 235
rect -685 205 -555 235
rect -525 205 -395 235
rect -365 205 10685 235
rect 10715 205 10845 235
rect 10875 205 11005 235
rect 11035 205 11040 235
rect -720 200 11040 205
rect -720 155 -360 160
rect -720 125 -715 155
rect -685 125 -555 155
rect -525 125 -395 155
rect -365 125 -360 155
rect -720 120 -360 125
rect -320 155 10800 160
rect -320 125 10 155
rect 190 125 330 155
rect 510 125 650 155
rect 830 125 970 155
rect 1150 125 1205 155
rect 1235 125 1290 155
rect 1470 125 1610 155
rect 1790 125 1930 155
rect 2110 125 2250 155
rect 2430 125 2570 155
rect 2750 125 2890 155
rect 3070 125 3210 155
rect 3390 125 3530 155
rect 3710 125 3765 155
rect 3795 125 3850 155
rect 4030 125 4170 155
rect 4350 125 4490 155
rect 4670 125 4810 155
rect 4990 125 5045 155
rect 5075 125 5290 155
rect 5470 125 5610 155
rect 5790 125 5930 155
rect 6110 125 6250 155
rect 6430 125 6570 155
rect 6750 125 6890 155
rect 7070 125 7210 155
rect 7390 125 7530 155
rect 7710 125 7850 155
rect 8030 125 8170 155
rect 8350 125 8490 155
rect 8670 125 8810 155
rect 8990 125 9130 155
rect 9310 125 9450 155
rect 9630 125 9770 155
rect 9950 125 10090 155
rect 10270 125 10765 155
rect 10795 125 10800 155
rect -320 120 10800 125
rect -720 75 10640 80
rect -720 45 -715 75
rect -685 45 -555 75
rect -525 45 -395 75
rect -365 45 -75 75
rect -45 45 2485 75
rect 2515 45 5045 75
rect 5075 45 5205 75
rect 5235 45 7765 75
rect 7795 45 10325 75
rect 10355 45 10640 75
rect -720 40 10640 45
rect -720 -5 10640 0
rect -720 -35 -715 -5
rect -685 -35 -555 -5
rect -525 -35 -395 -5
rect -365 -35 -75 -5
rect -45 -35 2485 -5
rect 2515 -35 5045 -5
rect 5075 -35 5205 -5
rect 5235 -35 7765 -5
rect 7795 -35 10325 -5
rect 10355 -35 10640 -5
rect -720 -40 10640 -35
rect -720 -120 10640 -80
<< via2 >>
rect -715 1005 -685 1035
rect -635 765 -605 795
rect -635 685 -605 715
rect -475 445 -445 475
rect 10925 285 10955 315
rect -715 205 -685 235
rect -555 205 -525 235
rect -395 205 -365 235
rect 10685 205 10715 235
rect 10845 205 10875 235
rect 11005 205 11035 235
rect -715 125 -685 155
rect -555 125 -525 155
rect -395 125 -365 155
rect 10765 125 10795 155
rect -715 45 -685 75
rect -555 45 -525 75
rect -395 45 -365 75
rect -715 -35 -685 -5
rect -555 -35 -525 -5
rect -395 -35 -365 -5
<< metal3 >>
rect -720 1035 -680 1040
rect -720 1005 -715 1035
rect -685 1005 -680 1035
rect -720 235 -680 1005
rect -720 205 -715 235
rect -685 205 -680 235
rect -720 155 -680 205
rect -720 125 -715 155
rect -685 125 -680 155
rect -720 75 -680 125
rect -720 45 -715 75
rect -685 45 -680 75
rect -720 -5 -680 45
rect -720 -35 -715 -5
rect -685 -35 -680 -5
rect -720 -120 -680 -35
rect -640 795 -600 1080
rect -640 765 -635 795
rect -605 765 -600 795
rect -640 715 -600 765
rect -640 685 -635 715
rect -605 685 -600 715
rect -640 -120 -600 685
rect -560 235 -520 1040
rect -560 205 -555 235
rect -525 205 -520 235
rect -560 155 -520 205
rect -560 125 -555 155
rect -525 125 -520 155
rect -560 75 -520 125
rect -560 45 -555 75
rect -525 45 -520 75
rect -560 -5 -520 45
rect -560 -35 -555 -5
rect -525 -35 -520 -5
rect -560 -120 -520 -35
rect -480 475 -440 1080
rect -480 445 -475 475
rect -445 445 -440 475
rect -480 -120 -440 445
rect -400 235 -360 1040
rect -400 205 -395 235
rect -365 205 -360 235
rect -400 155 -360 205
rect -400 125 -395 155
rect -365 125 -360 155
rect -400 75 -360 125
rect -400 45 -395 75
rect -365 45 -360 75
rect -400 -5 -360 45
rect -400 -35 -395 -5
rect -365 -35 -360 -5
rect -400 -120 -360 -35
rect 10680 235 10720 1040
rect 10680 205 10685 235
rect 10715 205 10720 235
rect 10680 -120 10720 205
rect 10760 155 10800 1080
rect 10760 125 10765 155
rect 10795 125 10800 155
rect 10760 -120 10800 125
rect 10840 235 10880 1040
rect 10840 205 10845 235
rect 10875 205 10880 235
rect 10840 -120 10880 205
rect 10920 315 10960 1080
rect 10920 285 10925 315
rect 10955 285 10960 315
rect 10920 -120 10960 285
rect 11000 235 11040 1080
rect 11000 205 11005 235
rect 11035 205 11040 235
rect 11000 -120 11040 205
<< labels >>
rlabel metal3 -640 1040 -600 1080 0 ii
port 1 nsew
rlabel metal3 -480 1040 -440 1080 0 vi
port 2 nsew
rlabel metal3 10760 1040 10800 1080 0 n
rlabel metal3 10920 1040 10960 1080 0 vo
port 3 nsew
rlabel metal3 11000 1040 11040 1080 0 vssa
port 4 nsew
<< end >>
