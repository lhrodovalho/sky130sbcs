* SPICE3 file created from vref5v0.ext - technology: sky130A

.subckt vref5v0 ii vi vo vssa
X0 a_16080_1320# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X1 a_6800_n760# n a_6160_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X2 a_19920_0# n a_19280_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X3 a_14800_0# n a_14160_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X4 vo n a_1680_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X5 a_5520_0# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X6 ii vo a_16080_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X7 a_12240_1320# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X8 a_5520_n2080# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X9 a_9360_0# n a_8720_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X10 a_4240_0# n a_3600_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X11 a_18640_n2080# vi a_18000_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X12 a_18640_n760# n n vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X13 a_7440_1320# vi a_6800_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X14 a_14160_n760# n a_13520_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X15 a_2960_1320# vi a_2320_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X16 a_2960_n2080# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X17 a_14800_n760# n a_14160_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X18 a_3600_1320# vi a_2960_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X19 a_16080_n2080# vi a_15440_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X20 vssa n a_4240_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X21 a_1040_n760# n a_400_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X22 a_16080_0# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X23 a_10960_0# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X24 vssa n a_19920_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X25 vssa n a_19920_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X26 vo vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X27 a_5520_n760# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X28 a_1680_0# n a_1040_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X29 ii vo a_2960_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X30 ii vo a_14800_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X31 a_16720_n2080# vi a_16080_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X32 vo vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X33 vo n a_17360_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X34 ii vo vo ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X35 a_9360_n760# n a_8720_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X36 a_8720_0# n a_8080_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X37 a_3600_0# n a_2960_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X38 ii vo vo ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X39 a_14160_n2080# vi a_13520_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X40 n n a_12240_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X41 a_1680_1320# vi a_1040_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X42 ii vo a_18640_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X43 vssa n a_9360_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X44 n n a_1680_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X45 a_13520_n760# n n vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X46 a_19920_1320# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X47 vssa n a_14800_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X48 a_14800_n2080# vi a_14160_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X49 a_17360_n760# n a_16720_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X50 a_19280_0# n a_18640_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X51 a_14160_0# n a_13520_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X52 a_6160_1320# vi a_5520_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X53 a_12240_n2080# vi a_11600_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X54 ii vo a_400_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X55 vssa n a_4240_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X56 n n a_17360_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X57 a_6800_1320# vi a_6160_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X58 a_2320_1320# vi a_1680_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X59 a_8080_n760# n vo vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X60 a_1680_n2080# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X61 a_8720_n760# n a_8080_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X62 a_6800_0# n a_6160_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X63 a_4240_n760# n a_3600_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X64 a_18640_1320# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X65 a_8080_n2080# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X66 ii vo a_13520_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X67 a_400_n760# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X68 a_15440_n2080# vi a_14800_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X69 a_18640_0# n vo vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X70 a_13520_0# n vo vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X71 a_14800_1320# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X72 a_16080_n760# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X73 a_1040_1320# vi a_400_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X74 a_4880_1320# vi a_4240_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X75 ii vi a_19920_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X76 ii vo a_8080_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X77 ii vo a_19920_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X78 a_17360_0# n a_16720_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X79 a_12240_0# n a_11600_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X80 a_12880_n2080# vi a_12240_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X81 a_16720_n760# n a_16080_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X82 a_5520_1320# vi a_4880_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X83 a_12240_n760# n a_11600_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X84 a_8080_0# n n vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X85 a_2960_0# n n vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X86 ii vo a_5520_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X87 vo n a_6800_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X88 a_19280_n2080# vi a_18640_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X89 a_2960_n760# n vo vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X90 a_9360_1320# vi a_8720_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X91 a_13520_n2080# vi a_12880_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X92 ii vo a_12240_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X93 vssa n a_9360_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X94 a_3600_n760# n a_2960_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X95 n vi a_9360_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X96 a_6800_n2080# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X97 a_13520_1320# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X98 a_10960_n2080# vi n ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X99 a_19920_n2080# vi a_19280_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X100 a_11600_0# n a_10960_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X101 a_4240_n2080# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X102 a_16720_0# n a_16080_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X103 a_400_0# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X104 vssa n a_14800_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7e+11p pd=2.9e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X105 a_400_n2080# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X106 a_10960_n760# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=7e+11p ps=2.9e+06u w=1e+06u l=2e+06u
X107 a_17360_n2080# vi a_16720_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X108 a_17360_1320# vo ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X109 n n a_6800_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X110 a_11600_n2080# vi a_10960_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X111 a_11600_n760# n a_10960_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X112 ii vo a_17360_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X113 a_1680_n760# n a_1040_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X114 a_19280_n760# n a_18640_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X115 a_6160_0# n a_5520_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X116 a_8080_1320# vi a_7440_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X117 a_18000_n2080# vi a_17360_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X118 a_19920_n760# n a_19280_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X119 a_8720_1320# vi a_8080_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X120 a_4240_1320# vi a_3600_1320# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X121 ii vo a_1680_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X122 ii vo a_6800_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X123 vo n a_12240_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X124 a_400_1320# vi ii ii sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.35294e+11p ps=2.44706e+06u w=1e+06u l=2e+06u
X125 a_6160_n760# n a_5520_n760# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X126 ii vo a_4240_n2080# ii sky130_fd_pr__pfet_g5v0d10v5 ad=6.35294e+11p pd=2.44706e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X127 a_1040_0# n a_400_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
C0 ii vo 23.34fF
C1 ii vi 21.01fF
C2 n vo 12.22fF
C3 vi vo 14.55fF
C4 n vssa 282.42fF
.ends
