* NGSPICE file created from sbcs5v0_.ext - technology: sky130A

.subckt sbcs5v0_ io vdda vssa x
X0 a_3920_3840# n a_3280_3840# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X1 a_3280_6120# p2 a_2720_6120# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X2 a_4560_0# y z vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X3 a_4560_6560# p0 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X4 a_3280_2720# p1 a_2720_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X5 a_1040_2280# p2 x vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X6 io p2 a_400_9960# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.66667e+11p pd=2.66667e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X7 p1 p2 a_3280_6120# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X8 p1 s a_1040_7680# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.22222e+11p pd=2.35556e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X9 a_3280_0# x vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X10 a_1040_3840# y a_400_3840# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X11 vssa n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X12 vdda p1 a_3280_2720# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X13 p0 p2 a_400_6120# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X14 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X15 n s p1 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X16 y y a_4560_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X17 a_1040_2280# p1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X18 a_1680_6560# p0 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X19 vdda p2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X20 vdda p1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X21 a_6160_7680# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X22 a_5200_6120# p0 a_4560_6560# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X23 a_1680_0# x z vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X24 a_6800_7680# n a_6160_7680# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X25 n s p1 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X26 vssa n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X27 a_6160_6560# p2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X28 p1 s n vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X29 a_6800_6560# p2 a_6160_6560# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X30 a_2320_6120# p0 a_1680_6560# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X31 vdda p0 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X32 n s p1 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7.42857e+11p pd=3.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X33 x x a_1680_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X34 a_8080_2280# p2 a_7440_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X35 a_3280_6560# p0 a_2720_6120# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X36 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X37 vssa n a_7440_3840# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X38 a_1040_7680# s p1 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.22222e+11p ps=2.35556e+06u w=1e+06u l=2e+06u
X39 vdda p1 a_400_10400# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X40 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X41 vdda p0 a_3280_6560# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X42 p2 p2 a_7440_6120# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X43 vssa n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X44 a_1680_10400# p1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X45 x p2 a_n160_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X46 a_8080_2280# p1 a_7440_2720# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X47 a_400_9960# p2 io vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.66667e+11p ps=2.66667e+06u w=1e+06u l=2e+06u
X48 vdda p0 a_400_6560# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X49 a_400_3840# y vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X50 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X51 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X52 a_400_6120# p2 a_n160_6120# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X53 a_6800_0# n a_6160_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X54 vdda p1 a_n160_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X55 a_7440_2280# p2 n vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X56 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X57 a_7440_3840# n p2 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X58 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X59 a_7440_6120# p2 a_6800_6120# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X60 a_7440_2720# p1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X61 a_4560_2280# p2 y vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X62 s n a_7440_7680# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X63 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X64 n n a_7440_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7.42857e+11p pd=3.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X65 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X66 a_4560_3840# n a_3920_3840# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X67 z x a_3280_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X68 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X69 vssa n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X70 a_4560_6120# p2 p1 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X71 p2 p2 a_7440_6560# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X72 p1 s n vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X73 a_4560_2720# p1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X74 x p2 a_1040_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X75 a_1680_9960# p2 io vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.66667e+11p ps=2.66667e+06u w=1e+06u l=2e+06u
X76 vdda p2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X77 a_400_10400# p1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X78 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X79 a_1680_3840# y a_1040_3840# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X80 vssa n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X81 a_400_6560# p0 a_n160_6120# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X82 a_400_0# x vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X83 a_5200_2280# p2 a_4560_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X84 a_1680_6120# p2 p0 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X85 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X86 vdda p2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X87 a_7440_0# n a_6800_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X88 vdda p1 a_1040_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X89 p1 n a_4560_3840# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.22222e+11p pd=2.35556e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X90 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X91 vdda p1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X92 a_6160_2280# p2 a_5600_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X93 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X94 a_5200_6120# p2 a_4560_6120# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X95 a_7440_7680# n a_6800_7680# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X96 a_2320_9960# p1 a_1680_10400# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X97 a_6160_0# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X98 a_6160_3840# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X99 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X100 n p2 a_6160_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X101 a_5200_2280# p1 a_4560_2720# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X102 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X103 a_2320_2280# p2 x vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X104 a_2320_9960# p2 a_1680_9960# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X105 vdda p2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X106 a_6160_6120# p2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X107 vdda p2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X108 p2 n a_6160_3840# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X109 p0 y a_1680_3840# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X110 vssa n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X111 a_7440_6560# p2 a_6800_6560# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X112 a_6160_2720# p1 a_5600_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X113 a_3280_2280# p2 a_2720_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X114 a_6800_6120# p2 a_6160_6120# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X115 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X116 a_2320_6120# p2 a_1680_6120# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X117 vdda p2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X118 p1 s n vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.22222e+11p pd=2.35556e+06u as=7.42857e+11p ps=3.2e+06u w=1e+06u l=2e+06u
X119 a_3280_3840# n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=8e+11p ps=3.6e+06u w=1e+06u l=2e+06u
X120 vdda p1 a_6160_2720# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X121 y p2 a_3280_2280# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X122 a_2320_2280# p1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=3.6e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X123 vdda s vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
X124 z x a_400_0# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X125 vdda p1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=6.9589e+11p pd=2.87123e+06u as=6.9589e+11p ps=2.87123e+06u w=1e+06u l=2e+06u
.ends

