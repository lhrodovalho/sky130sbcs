* 1.8 V CMOS only voltage reference testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0

.include "../mag/vref5v0.spice"
.include "../../sbcs5v0/mag/sbcs5v0.spice"

* supply voltages
vdda	vdda 0 3.3
vssa	vssa 0 0.0

* DUT
x0 io vdda vssa x sbcs5v0
vo io ii 0.0

x1 ii x ref vssa vref5v0

.option gmin=1e-12
.control
  dc vdda 10m 5.0 10m
  plot x ref
  plot i(vo)
  plot abs(deriv(ref)/ref) ylog
  
  dc temp -40 125 1
  meas dc r27 find ref at=27
  let refN = ref/r27
  plot refN
  
.endc

.end
