magic
tech sky130A
timestamp 1640957228
<< nwell >>
rect -200 480 10520 920
<< pmoslvt >>
rect 0 660 200 760
rect 320 660 520 760
rect 640 660 840 760
rect 960 660 1160 760
rect 1280 660 1480 760
rect 1600 660 1800 760
rect 1920 660 2120 760
rect 2240 660 2440 760
rect 2560 660 2760 760
rect 2880 660 3080 760
rect 3200 660 3400 760
rect 3520 660 3720 760
rect 3840 660 4040 760
rect 4160 660 4360 760
rect 4480 660 4680 760
rect 4800 660 5000 760
rect 5280 660 5480 760
rect 5600 660 5800 760
rect 5920 660 6120 760
rect 6240 660 6440 760
rect 6560 660 6760 760
rect 6880 660 7080 760
rect 7200 660 7400 760
rect 7520 660 7720 760
rect 7840 660 8040 760
rect 8160 660 8360 760
rect 8480 660 8680 760
rect 8800 660 9000 760
rect 9120 660 9320 760
rect 9440 660 9640 760
rect 9760 660 9960 760
rect 10080 660 10280 760
<< nmoslvt >>
rect 0 0 200 100
rect 320 0 520 100
rect 640 0 840 100
rect 960 0 1160 100
rect 1280 0 1480 100
rect 1600 0 1800 100
rect 1920 0 2120 100
rect 2240 0 2440 100
rect 2560 0 2760 100
rect 2880 0 3080 100
rect 3200 0 3400 100
rect 3520 0 3720 100
rect 3840 0 4040 100
rect 4160 0 4360 100
rect 4480 0 4680 100
rect 4800 0 5000 100
rect 5280 0 5480 100
rect 5600 0 5800 100
rect 5920 0 6120 100
rect 6240 0 6440 100
rect 6560 0 6760 100
rect 6880 0 7080 100
rect 7200 0 7400 100
rect 7520 0 7720 100
rect 7840 0 8040 100
rect 8160 0 8360 100
rect 8480 0 8680 100
rect 8800 0 9000 100
rect 9120 0 9320 100
rect 9440 0 9640 100
rect 9760 0 9960 100
rect 10080 0 10280 100
<< ndiff >>
rect -80 90 0 100
rect -80 10 -75 90
rect -45 10 0 90
rect -80 0 0 10
rect 200 90 320 100
rect 200 10 245 90
rect 275 10 320 90
rect 200 0 320 10
rect 520 90 640 100
rect 520 10 565 90
rect 595 10 640 90
rect 520 0 640 10
rect 840 90 960 100
rect 840 10 885 90
rect 915 10 960 90
rect 840 0 960 10
rect 1160 90 1280 100
rect 1160 10 1205 90
rect 1235 10 1280 90
rect 1160 0 1280 10
rect 1480 90 1600 100
rect 1480 10 1525 90
rect 1555 10 1600 90
rect 1480 0 1600 10
rect 1800 90 1920 100
rect 1800 10 1845 90
rect 1875 10 1920 90
rect 1800 0 1920 10
rect 2120 90 2240 100
rect 2120 10 2165 90
rect 2195 10 2240 90
rect 2120 0 2240 10
rect 2440 90 2560 100
rect 2440 10 2485 90
rect 2515 10 2560 90
rect 2440 0 2560 10
rect 2760 90 2880 100
rect 2760 10 2805 90
rect 2835 10 2880 90
rect 2760 0 2880 10
rect 3080 90 3200 100
rect 3080 10 3125 90
rect 3155 10 3200 90
rect 3080 0 3200 10
rect 3400 90 3520 100
rect 3400 10 3445 90
rect 3475 10 3520 90
rect 3400 0 3520 10
rect 3720 90 3840 100
rect 3720 10 3765 90
rect 3795 10 3840 90
rect 3720 0 3840 10
rect 4040 90 4160 100
rect 4040 10 4085 90
rect 4115 10 4160 90
rect 4040 0 4160 10
rect 4360 90 4480 100
rect 4360 10 4405 90
rect 4435 10 4480 90
rect 4360 0 4480 10
rect 4680 90 4800 100
rect 4680 10 4725 90
rect 4755 10 4800 90
rect 4680 0 4800 10
rect 5000 90 5080 100
rect 5000 10 5045 90
rect 5075 10 5080 90
rect 5000 0 5080 10
rect 5200 90 5280 100
rect 5200 10 5205 90
rect 5235 10 5280 90
rect 5200 0 5280 10
rect 5480 90 5600 100
rect 5480 10 5525 90
rect 5555 10 5600 90
rect 5480 0 5600 10
rect 5800 90 5920 100
rect 5800 10 5845 90
rect 5875 10 5920 90
rect 5800 0 5920 10
rect 6120 90 6240 100
rect 6120 10 6165 90
rect 6195 10 6240 90
rect 6120 0 6240 10
rect 6440 90 6560 100
rect 6440 10 6485 90
rect 6515 10 6560 90
rect 6440 0 6560 10
rect 6760 90 6880 100
rect 6760 10 6805 90
rect 6835 10 6880 90
rect 6760 0 6880 10
rect 7080 90 7200 100
rect 7080 10 7125 90
rect 7155 10 7200 90
rect 7080 0 7200 10
rect 7400 90 7520 100
rect 7400 10 7445 90
rect 7475 10 7520 90
rect 7400 0 7520 10
rect 7720 90 7840 100
rect 7720 10 7765 90
rect 7795 10 7840 90
rect 7720 0 7840 10
rect 8040 90 8160 100
rect 8040 10 8085 90
rect 8115 10 8160 90
rect 8040 0 8160 10
rect 8360 90 8480 100
rect 8360 10 8405 90
rect 8435 10 8480 90
rect 8360 0 8480 10
rect 8680 90 8800 100
rect 8680 10 8725 90
rect 8755 10 8800 90
rect 8680 0 8800 10
rect 9000 90 9120 100
rect 9000 10 9045 90
rect 9075 10 9120 90
rect 9000 0 9120 10
rect 9320 90 9440 100
rect 9320 10 9365 90
rect 9395 10 9440 90
rect 9320 0 9440 10
rect 9640 90 9760 100
rect 9640 10 9685 90
rect 9715 10 9760 90
rect 9640 0 9760 10
rect 9960 90 10080 100
rect 9960 10 10005 90
rect 10035 10 10080 90
rect 9960 0 10080 10
rect 10280 90 10360 100
rect 10280 10 10325 90
rect 10355 10 10360 90
rect 10280 0 10360 10
<< pdiff >>
rect -80 750 0 760
rect -80 670 -75 750
rect -45 670 0 750
rect -80 660 0 670
rect 200 750 320 760
rect 200 670 245 750
rect 275 670 320 750
rect 200 660 320 670
rect 520 750 640 760
rect 520 670 565 750
rect 595 670 640 750
rect 520 660 640 670
rect 840 750 960 760
rect 840 670 885 750
rect 915 670 960 750
rect 840 660 960 670
rect 1160 750 1280 760
rect 1160 670 1205 750
rect 1235 670 1280 750
rect 1160 660 1280 670
rect 1480 750 1600 760
rect 1480 670 1525 750
rect 1555 670 1600 750
rect 1480 660 1600 670
rect 1800 750 1920 760
rect 1800 670 1845 750
rect 1875 670 1920 750
rect 1800 660 1920 670
rect 2120 750 2240 760
rect 2120 670 2165 750
rect 2195 670 2240 750
rect 2120 660 2240 670
rect 2440 750 2560 760
rect 2440 670 2485 750
rect 2515 670 2560 750
rect 2440 660 2560 670
rect 2760 750 2880 760
rect 2760 670 2805 750
rect 2835 670 2880 750
rect 2760 660 2880 670
rect 3080 750 3200 760
rect 3080 670 3125 750
rect 3155 670 3200 750
rect 3080 660 3200 670
rect 3400 750 3520 760
rect 3400 670 3445 750
rect 3475 670 3520 750
rect 3400 660 3520 670
rect 3720 750 3840 760
rect 3720 670 3765 750
rect 3795 670 3840 750
rect 3720 660 3840 670
rect 4040 750 4160 760
rect 4040 670 4085 750
rect 4115 670 4160 750
rect 4040 660 4160 670
rect 4360 750 4480 760
rect 4360 670 4405 750
rect 4435 670 4480 750
rect 4360 660 4480 670
rect 4680 750 4800 760
rect 4680 670 4725 750
rect 4755 670 4800 750
rect 4680 660 4800 670
rect 5000 750 5080 760
rect 5000 670 5045 750
rect 5075 670 5080 750
rect 5000 660 5080 670
rect 5200 750 5280 760
rect 5200 670 5205 750
rect 5235 670 5280 750
rect 5200 660 5280 670
rect 5480 750 5600 760
rect 5480 670 5525 750
rect 5555 670 5600 750
rect 5480 660 5600 670
rect 5800 750 5920 760
rect 5800 670 5845 750
rect 5875 670 5920 750
rect 5800 660 5920 670
rect 6120 750 6240 760
rect 6120 670 6165 750
rect 6195 670 6240 750
rect 6120 660 6240 670
rect 6440 750 6560 760
rect 6440 670 6485 750
rect 6515 670 6560 750
rect 6440 660 6560 670
rect 6760 750 6880 760
rect 6760 670 6805 750
rect 6835 670 6880 750
rect 6760 660 6880 670
rect 7080 750 7200 760
rect 7080 670 7125 750
rect 7155 670 7200 750
rect 7080 660 7200 670
rect 7400 750 7520 760
rect 7400 670 7445 750
rect 7475 670 7520 750
rect 7400 660 7520 670
rect 7720 750 7840 760
rect 7720 670 7765 750
rect 7795 670 7840 750
rect 7720 660 7840 670
rect 8040 750 8160 760
rect 8040 670 8085 750
rect 8115 670 8160 750
rect 8040 660 8160 670
rect 8360 750 8480 760
rect 8360 670 8405 750
rect 8435 670 8480 750
rect 8360 660 8480 670
rect 8680 750 8800 760
rect 8680 670 8725 750
rect 8755 670 8800 750
rect 8680 660 8800 670
rect 9000 750 9120 760
rect 9000 670 9045 750
rect 9075 670 9120 750
rect 9000 660 9120 670
rect 9320 750 9440 760
rect 9320 670 9365 750
rect 9395 670 9440 750
rect 9320 660 9440 670
rect 9640 750 9760 760
rect 9640 670 9685 750
rect 9715 670 9760 750
rect 9640 660 9760 670
rect 9960 750 10080 760
rect 9960 670 10005 750
rect 10035 670 10080 750
rect 9960 660 10080 670
rect 10280 750 10360 760
rect 10280 670 10325 750
rect 10355 670 10360 750
rect 10280 660 10360 670
<< ndiffc >>
rect -75 10 -45 90
rect 245 10 275 90
rect 565 10 595 90
rect 885 10 915 90
rect 1205 10 1235 90
rect 1525 10 1555 90
rect 1845 10 1875 90
rect 2165 10 2195 90
rect 2485 10 2515 90
rect 2805 10 2835 90
rect 3125 10 3155 90
rect 3445 10 3475 90
rect 3765 10 3795 90
rect 4085 10 4115 90
rect 4405 10 4435 90
rect 4725 10 4755 90
rect 5045 10 5075 90
rect 5205 10 5235 90
rect 5525 10 5555 90
rect 5845 10 5875 90
rect 6165 10 6195 90
rect 6485 10 6515 90
rect 6805 10 6835 90
rect 7125 10 7155 90
rect 7445 10 7475 90
rect 7765 10 7795 90
rect 8085 10 8115 90
rect 8405 10 8435 90
rect 8725 10 8755 90
rect 9045 10 9075 90
rect 9365 10 9395 90
rect 9685 10 9715 90
rect 10005 10 10035 90
rect 10325 10 10355 90
<< pdiffc >>
rect -75 670 -45 750
rect 245 670 275 750
rect 565 670 595 750
rect 885 670 915 750
rect 1205 670 1235 750
rect 1525 670 1555 750
rect 1845 670 1875 750
rect 2165 670 2195 750
rect 2485 670 2515 750
rect 2805 670 2835 750
rect 3125 670 3155 750
rect 3445 670 3475 750
rect 3765 670 3795 750
rect 4085 670 4115 750
rect 4405 670 4435 750
rect 4725 670 4755 750
rect 5045 670 5075 750
rect 5205 670 5235 750
rect 5525 670 5555 750
rect 5845 670 5875 750
rect 6165 670 6195 750
rect 6485 670 6515 750
rect 6805 670 6835 750
rect 7125 670 7155 750
rect 7445 670 7475 750
rect 7765 670 7795 750
rect 8085 670 8115 750
rect 8405 670 8435 750
rect 8725 670 8755 750
rect 9045 670 9075 750
rect 9365 670 9395 750
rect 9685 670 9715 750
rect 10005 670 10035 750
rect 10325 670 10355 750
<< psubdiff >>
rect -320 1000 -40 1040
rect 240 1000 280 1040
rect 560 1000 600 1040
rect 880 1000 920 1040
rect 1200 1000 1240 1040
rect 1520 1000 1560 1040
rect 1840 1000 1880 1040
rect 2160 1000 2200 1040
rect 2480 1000 2520 1040
rect 2800 1000 2840 1040
rect 3120 1000 3160 1040
rect 3440 1000 3480 1040
rect 3760 1000 3800 1040
rect 4080 1000 4120 1040
rect 4400 1000 4440 1040
rect 4720 1000 4760 1040
rect 5040 1000 5240 1040
rect 5520 1000 5560 1040
rect 5840 1000 5880 1040
rect 6160 1000 6200 1040
rect 6480 1000 6520 1040
rect 6800 1000 6840 1040
rect 7120 1000 7160 1040
rect 7440 1000 7480 1040
rect 7760 1000 7800 1040
rect 8080 1000 8120 1040
rect 8400 1000 8440 1040
rect 8720 1000 8760 1040
rect 9040 1000 9080 1040
rect 9360 1000 9400 1040
rect 9680 1000 9720 1040
rect 10000 1000 10040 1040
rect 10320 1000 10600 1040
rect -320 960 -280 1000
rect 10560 960 10600 1000
rect -280 360 -40 400
rect 240 360 280 400
rect 560 360 600 400
rect 880 360 920 400
rect 1200 360 1240 400
rect 1520 360 1560 400
rect 1840 360 1880 400
rect 2160 360 2200 400
rect 2480 360 2520 400
rect 2800 360 2840 400
rect 3120 360 3160 400
rect 3440 360 3480 400
rect 3760 360 3800 400
rect 4080 360 4120 400
rect 4400 360 4440 400
rect 4720 360 4760 400
rect 5040 360 5240 400
rect 5520 360 5560 400
rect 5840 360 5880 400
rect 6160 360 6200 400
rect 6480 360 6520 400
rect 6800 360 6840 400
rect 7120 360 7160 400
rect 7440 360 7480 400
rect 7760 360 7800 400
rect 8080 360 8120 400
rect 8400 360 8440 400
rect 8720 360 8760 400
rect 9040 360 9080 400
rect 9360 360 9400 400
rect 9680 360 9720 400
rect 10000 360 10040 400
rect 10320 360 10560 400
rect -320 -80 -280 -40
rect -160 200 -40 240
rect 240 200 280 240
rect 560 200 600 240
rect 880 200 920 240
rect 1200 200 1240 240
rect 1520 200 1560 240
rect 1840 200 1880 240
rect 2160 200 2200 240
rect 2480 200 2520 240
rect 2800 200 2840 240
rect 3120 200 3160 240
rect 3440 200 3480 240
rect 3760 200 3800 240
rect 4080 200 4120 240
rect 4400 200 4440 240
rect 4720 200 4760 240
rect 5040 200 5240 240
rect 5520 200 5560 240
rect 5840 200 5880 240
rect 6160 200 6200 240
rect 6480 200 6520 240
rect 6800 200 6840 240
rect 7120 200 7160 240
rect 7440 200 7480 240
rect 7760 200 7800 240
rect 8080 200 8120 240
rect 8400 200 8440 240
rect 8720 200 8760 240
rect 9040 200 9080 240
rect 9360 200 9400 240
rect 9680 200 9720 240
rect 10000 200 10040 240
rect 10320 200 10480 240
rect -160 160 -120 200
rect 5120 160 5160 200
rect 10400 160 10440 200
rect -160 -80 -120 -40
rect 5120 -80 5160 -40
rect 10400 -80 10440 -40
rect 10560 -80 10600 -40
rect -320 -120 -40 -80
rect 240 -120 280 -80
rect 560 -120 600 -80
rect 880 -120 920 -80
rect 1200 -120 1240 -80
rect 1520 -120 1560 -80
rect 1840 -120 1880 -80
rect 2160 -120 2200 -80
rect 2480 -120 2520 -80
rect 2800 -120 2840 -80
rect 3120 -120 3160 -80
rect 3440 -120 3480 -80
rect 3760 -120 3800 -80
rect 4080 -120 4120 -80
rect 4400 -120 4440 -80
rect 4720 -120 4760 -80
rect 5040 -120 5240 -80
rect 5520 -120 5560 -80
rect 5840 -120 5880 -80
rect 6160 -120 6200 -80
rect 6480 -120 6520 -80
rect 6800 -120 6840 -80
rect 7120 -120 7160 -80
rect 7440 -120 7480 -80
rect 7760 -120 7800 -80
rect 8080 -120 8120 -80
rect 8400 -120 8440 -80
rect 8720 -120 8760 -80
rect 9040 -120 9080 -80
rect 9360 -120 9400 -80
rect 9680 -120 9720 -80
rect 10000 -120 10040 -80
rect 10320 -120 10600 -80
<< nsubdiff >>
rect -160 840 -40 880
rect 240 840 280 880
rect 560 840 600 880
rect 880 840 920 880
rect 1200 840 1240 880
rect 1520 840 1560 880
rect 1840 840 1880 880
rect 2160 840 2200 880
rect 2480 840 2520 880
rect 2800 840 2840 880
rect 3120 840 3160 880
rect 3440 840 3480 880
rect 3760 840 3800 880
rect 4080 840 4120 880
rect 4400 840 4440 880
rect 4720 840 4760 880
rect 5040 840 5240 880
rect 5520 840 5560 880
rect 5840 840 5880 880
rect 6160 840 6200 880
rect 6480 840 6520 880
rect 6800 840 6840 880
rect 7120 840 7160 880
rect 7440 840 7480 880
rect 7760 840 7800 880
rect 8080 840 8120 880
rect 8400 840 8440 880
rect 8720 840 8760 880
rect 9040 840 9080 880
rect 9360 840 9400 880
rect 9680 840 9720 880
rect 10000 840 10040 880
rect 10320 840 10480 880
rect -160 800 -120 840
rect 5120 800 5160 840
rect 10400 800 10440 840
rect -160 560 -120 600
rect 5120 560 5160 600
rect 10400 560 10440 600
rect -160 520 -40 560
rect 240 520 280 560
rect 560 520 600 560
rect 880 520 920 560
rect 1200 520 1240 560
rect 1520 520 1560 560
rect 1840 520 1880 560
rect 2160 520 2200 560
rect 2480 520 2520 560
rect 2800 520 2840 560
rect 3120 520 3160 560
rect 3440 520 3480 560
rect 3760 520 3800 560
rect 4080 520 4120 560
rect 4400 520 4440 560
rect 4720 520 4760 560
rect 5040 520 5240 560
rect 5520 520 5560 560
rect 5840 520 5880 560
rect 6160 520 6200 560
rect 6480 520 6520 560
rect 6800 520 6840 560
rect 7120 520 7160 560
rect 7440 520 7480 560
rect 7760 520 7800 560
rect 8080 520 8120 560
rect 8400 520 8440 560
rect 8720 520 8760 560
rect 9040 520 9080 560
rect 9360 520 9400 560
rect 9680 520 9720 560
rect 10000 520 10040 560
rect 10320 520 10480 560
<< psubdiffcont >>
rect -40 1000 240 1040
rect 280 1000 560 1040
rect 600 1000 880 1040
rect 920 1000 1200 1040
rect 1240 1000 1520 1040
rect 1560 1000 1840 1040
rect 1880 1000 2160 1040
rect 2200 1000 2480 1040
rect 2520 1000 2800 1040
rect 2840 1000 3120 1040
rect 3160 1000 3440 1040
rect 3480 1000 3760 1040
rect 3800 1000 4080 1040
rect 4120 1000 4400 1040
rect 4440 1000 4720 1040
rect 4760 1000 5040 1040
rect 5240 1000 5520 1040
rect 5560 1000 5840 1040
rect 5880 1000 6160 1040
rect 6200 1000 6480 1040
rect 6520 1000 6800 1040
rect 6840 1000 7120 1040
rect 7160 1000 7440 1040
rect 7480 1000 7760 1040
rect 7800 1000 8080 1040
rect 8120 1000 8400 1040
rect 8440 1000 8720 1040
rect 8760 1000 9040 1040
rect 9080 1000 9360 1040
rect 9400 1000 9680 1040
rect 9720 1000 10000 1040
rect 10040 1000 10320 1040
rect -320 -40 -280 960
rect -40 360 240 400
rect 280 360 560 400
rect 600 360 880 400
rect 920 360 1200 400
rect 1240 360 1520 400
rect 1560 360 1840 400
rect 1880 360 2160 400
rect 2200 360 2480 400
rect 2520 360 2800 400
rect 2840 360 3120 400
rect 3160 360 3440 400
rect 3480 360 3760 400
rect 3800 360 4080 400
rect 4120 360 4400 400
rect 4440 360 4720 400
rect 4760 360 5040 400
rect 5240 360 5520 400
rect 5560 360 5840 400
rect 5880 360 6160 400
rect 6200 360 6480 400
rect 6520 360 6800 400
rect 6840 360 7120 400
rect 7160 360 7440 400
rect 7480 360 7760 400
rect 7800 360 8080 400
rect 8120 360 8400 400
rect 8440 360 8720 400
rect 8760 360 9040 400
rect 9080 360 9360 400
rect 9400 360 9680 400
rect 9720 360 10000 400
rect 10040 360 10320 400
rect -40 200 240 240
rect 280 200 560 240
rect 600 200 880 240
rect 920 200 1200 240
rect 1240 200 1520 240
rect 1560 200 1840 240
rect 1880 200 2160 240
rect 2200 200 2480 240
rect 2520 200 2800 240
rect 2840 200 3120 240
rect 3160 200 3440 240
rect 3480 200 3760 240
rect 3800 200 4080 240
rect 4120 200 4400 240
rect 4440 200 4720 240
rect 4760 200 5040 240
rect 5240 200 5520 240
rect 5560 200 5840 240
rect 5880 200 6160 240
rect 6200 200 6480 240
rect 6520 200 6800 240
rect 6840 200 7120 240
rect 7160 200 7440 240
rect 7480 200 7760 240
rect 7800 200 8080 240
rect 8120 200 8400 240
rect 8440 200 8720 240
rect 8760 200 9040 240
rect 9080 200 9360 240
rect 9400 200 9680 240
rect 9720 200 10000 240
rect 10040 200 10320 240
rect -160 -40 -120 160
rect 5120 -40 5160 160
rect 10400 -40 10440 160
rect 10560 -40 10600 960
rect -40 -120 240 -80
rect 280 -120 560 -80
rect 600 -120 880 -80
rect 920 -120 1200 -80
rect 1240 -120 1520 -80
rect 1560 -120 1840 -80
rect 1880 -120 2160 -80
rect 2200 -120 2480 -80
rect 2520 -120 2800 -80
rect 2840 -120 3120 -80
rect 3160 -120 3440 -80
rect 3480 -120 3760 -80
rect 3800 -120 4080 -80
rect 4120 -120 4400 -80
rect 4440 -120 4720 -80
rect 4760 -120 5040 -80
rect 5240 -120 5520 -80
rect 5560 -120 5840 -80
rect 5880 -120 6160 -80
rect 6200 -120 6480 -80
rect 6520 -120 6800 -80
rect 6840 -120 7120 -80
rect 7160 -120 7440 -80
rect 7480 -120 7760 -80
rect 7800 -120 8080 -80
rect 8120 -120 8400 -80
rect 8440 -120 8720 -80
rect 8760 -120 9040 -80
rect 9080 -120 9360 -80
rect 9400 -120 9680 -80
rect 9720 -120 10000 -80
rect 10040 -120 10320 -80
<< nsubdiffcont >>
rect -40 840 240 880
rect 280 840 560 880
rect 600 840 880 880
rect 920 840 1200 880
rect 1240 840 1520 880
rect 1560 840 1840 880
rect 1880 840 2160 880
rect 2200 840 2480 880
rect 2520 840 2800 880
rect 2840 840 3120 880
rect 3160 840 3440 880
rect 3480 840 3760 880
rect 3800 840 4080 880
rect 4120 840 4400 880
rect 4440 840 4720 880
rect 4760 840 5040 880
rect 5240 840 5520 880
rect 5560 840 5840 880
rect 5880 840 6160 880
rect 6200 840 6480 880
rect 6520 840 6800 880
rect 6840 840 7120 880
rect 7160 840 7440 880
rect 7480 840 7760 880
rect 7800 840 8080 880
rect 8120 840 8400 880
rect 8440 840 8720 880
rect 8760 840 9040 880
rect 9080 840 9360 880
rect 9400 840 9680 880
rect 9720 840 10000 880
rect 10040 840 10320 880
rect -160 600 -120 800
rect 5120 600 5160 800
rect 10400 600 10440 800
rect -40 520 240 560
rect 280 520 560 560
rect 600 520 880 560
rect 920 520 1200 560
rect 1240 520 1520 560
rect 1560 520 1840 560
rect 1880 520 2160 560
rect 2200 520 2480 560
rect 2520 520 2800 560
rect 2840 520 3120 560
rect 3160 520 3440 560
rect 3480 520 3760 560
rect 3800 520 4080 560
rect 4120 520 4400 560
rect 4440 520 4720 560
rect 4760 520 5040 560
rect 5240 520 5520 560
rect 5560 520 5840 560
rect 5880 520 6160 560
rect 6200 520 6480 560
rect 6520 520 6800 560
rect 6840 520 7120 560
rect 7160 520 7440 560
rect 7480 520 7760 560
rect 7800 520 8080 560
rect 8120 520 8400 560
rect 8440 520 8720 560
rect 8760 520 9040 560
rect 9080 520 9360 560
rect 9400 520 9680 560
rect 9720 520 10000 560
rect 10040 520 10320 560
<< poly >>
rect 0 760 200 780
rect 320 760 520 780
rect 640 760 840 780
rect 960 760 1160 780
rect 1280 760 1480 780
rect 1600 760 1800 780
rect 1920 760 2120 780
rect 2240 760 2440 780
rect 2560 760 2760 780
rect 2880 760 3080 780
rect 3200 760 3400 780
rect 3520 760 3720 780
rect 3840 760 4040 780
rect 4160 760 4360 780
rect 4480 760 4680 780
rect 4800 760 5000 780
rect 0 635 200 660
rect 0 605 10 635
rect 190 605 200 635
rect 0 600 200 605
rect 320 635 520 660
rect 320 605 330 635
rect 510 605 520 635
rect 320 600 520 605
rect 640 635 840 660
rect 640 605 650 635
rect 830 605 840 635
rect 640 600 840 605
rect 960 635 1160 660
rect 960 605 970 635
rect 1150 605 1160 635
rect 960 600 1160 605
rect 1280 635 1480 660
rect 1280 605 1290 635
rect 1470 605 1480 635
rect 1280 600 1480 605
rect 1600 635 1800 660
rect 1600 605 1610 635
rect 1790 605 1800 635
rect 1600 600 1800 605
rect 1920 635 2120 660
rect 1920 605 1930 635
rect 2110 605 2120 635
rect 1920 600 2120 605
rect 2240 635 2440 660
rect 2240 605 2250 635
rect 2430 605 2440 635
rect 2240 600 2440 605
rect 2560 635 2760 660
rect 2560 605 2570 635
rect 2750 605 2760 635
rect 2560 600 2760 605
rect 2880 635 3080 660
rect 2880 605 2890 635
rect 3070 605 3080 635
rect 2880 600 3080 605
rect 3200 635 3400 660
rect 3200 605 3210 635
rect 3390 605 3400 635
rect 3200 600 3400 605
rect 3520 635 3720 660
rect 3520 605 3530 635
rect 3710 605 3720 635
rect 3520 600 3720 605
rect 3840 635 4040 660
rect 3840 605 3850 635
rect 4030 605 4040 635
rect 3840 600 4040 605
rect 4160 635 4360 660
rect 4160 605 4170 635
rect 4350 605 4360 635
rect 4160 600 4360 605
rect 4480 635 4680 660
rect 4480 605 4490 635
rect 4670 605 4680 635
rect 4480 600 4680 605
rect 4800 635 5000 660
rect 4800 605 4810 635
rect 4990 605 5000 635
rect 4800 600 5000 605
rect 5280 760 5480 780
rect 5600 760 5800 780
rect 5920 760 6120 780
rect 6240 760 6440 780
rect 6560 760 6760 780
rect 6880 760 7080 780
rect 7200 760 7400 780
rect 7520 760 7720 780
rect 7840 760 8040 780
rect 8160 760 8360 780
rect 8480 760 8680 780
rect 8800 760 9000 780
rect 9120 760 9320 780
rect 9440 760 9640 780
rect 9760 760 9960 780
rect 10080 760 10280 780
rect 5280 635 5480 660
rect 5280 605 5290 635
rect 5470 605 5480 635
rect 5280 600 5480 605
rect 5600 635 5800 660
rect 5600 605 5610 635
rect 5790 605 5800 635
rect 5600 600 5800 605
rect 5920 635 6120 660
rect 5920 605 5930 635
rect 6110 605 6120 635
rect 5920 600 6120 605
rect 6240 635 6440 660
rect 6240 605 6250 635
rect 6430 605 6440 635
rect 6240 600 6440 605
rect 6560 635 6760 660
rect 6560 605 6570 635
rect 6750 605 6760 635
rect 6560 600 6760 605
rect 6880 635 7080 660
rect 6880 605 6890 635
rect 7070 605 7080 635
rect 6880 600 7080 605
rect 7200 635 7400 660
rect 7200 605 7210 635
rect 7390 605 7400 635
rect 7200 600 7400 605
rect 7520 635 7720 660
rect 7520 605 7530 635
rect 7710 605 7720 635
rect 7520 600 7720 605
rect 7840 635 8040 660
rect 7840 605 7850 635
rect 8030 605 8040 635
rect 7840 600 8040 605
rect 8160 635 8360 660
rect 8160 605 8170 635
rect 8350 605 8360 635
rect 8160 600 8360 605
rect 8480 635 8680 660
rect 8480 605 8490 635
rect 8670 605 8680 635
rect 8480 600 8680 605
rect 8800 635 9000 660
rect 8800 605 8810 635
rect 8990 605 9000 635
rect 8800 600 9000 605
rect 9120 635 9320 660
rect 9120 605 9130 635
rect 9310 605 9320 635
rect 9120 600 9320 605
rect 9440 635 9640 660
rect 9440 605 9450 635
rect 9630 605 9640 635
rect 9440 600 9640 605
rect 9760 635 9960 660
rect 9760 605 9770 635
rect 9950 605 9960 635
rect 9760 600 9960 605
rect 10080 635 10280 660
rect 10080 605 10090 635
rect 10270 605 10280 635
rect 10080 600 10280 605
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 100 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 100 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 100 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 100 1160 125
rect 1280 155 1480 160
rect 1280 125 1290 155
rect 1470 125 1480 155
rect 1280 100 1480 125
rect 1600 155 1800 160
rect 1600 125 1610 155
rect 1790 125 1800 155
rect 1600 100 1800 125
rect 1920 155 2120 160
rect 1920 125 1930 155
rect 2110 125 2120 155
rect 1920 100 2120 125
rect 2240 155 2440 160
rect 2240 125 2250 155
rect 2430 125 2440 155
rect 2240 100 2440 125
rect 2560 155 2760 160
rect 2560 125 2570 155
rect 2750 125 2760 155
rect 2560 100 2760 125
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 100 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 100 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 100 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 100 4040 125
rect 4160 155 4360 160
rect 4160 125 4170 155
rect 4350 125 4360 155
rect 4160 100 4360 125
rect 4480 155 4680 160
rect 4480 125 4490 155
rect 4670 125 4680 155
rect 4480 100 4680 125
rect 4800 155 5000 160
rect 4800 125 4810 155
rect 4990 125 5000 155
rect 4800 100 5000 125
rect 0 -20 200 0
rect 320 -20 520 0
rect 640 -20 840 0
rect 960 -20 1160 0
rect 1280 -20 1480 0
rect 1600 -20 1800 0
rect 1920 -20 2120 0
rect 2240 -20 2440 0
rect 2560 -20 2760 0
rect 2880 -20 3080 0
rect 3200 -20 3400 0
rect 3520 -20 3720 0
rect 3840 -20 4040 0
rect 4160 -20 4360 0
rect 4480 -20 4680 0
rect 4800 -20 5000 0
rect 5280 155 5480 160
rect 5280 125 5290 155
rect 5470 125 5480 155
rect 5280 100 5480 125
rect 5600 155 5800 160
rect 5600 125 5610 155
rect 5790 125 5800 155
rect 5600 100 5800 125
rect 5920 155 6120 160
rect 5920 125 5930 155
rect 6110 125 6120 155
rect 5920 100 6120 125
rect 6240 155 6440 160
rect 6240 125 6250 155
rect 6430 125 6440 155
rect 6240 100 6440 125
rect 6560 155 6760 160
rect 6560 125 6570 155
rect 6750 125 6760 155
rect 6560 100 6760 125
rect 6880 155 7080 160
rect 6880 125 6890 155
rect 7070 125 7080 155
rect 6880 100 7080 125
rect 7200 155 7400 160
rect 7200 125 7210 155
rect 7390 125 7400 155
rect 7200 100 7400 125
rect 7520 155 7720 160
rect 7520 125 7530 155
rect 7710 125 7720 155
rect 7520 100 7720 125
rect 7840 155 8040 160
rect 7840 125 7850 155
rect 8030 125 8040 155
rect 7840 100 8040 125
rect 8160 155 8360 160
rect 8160 125 8170 155
rect 8350 125 8360 155
rect 8160 100 8360 125
rect 8480 155 8680 160
rect 8480 125 8490 155
rect 8670 125 8680 155
rect 8480 100 8680 125
rect 8800 155 9000 160
rect 8800 125 8810 155
rect 8990 125 9000 155
rect 8800 100 9000 125
rect 9120 155 9320 160
rect 9120 125 9130 155
rect 9310 125 9320 155
rect 9120 100 9320 125
rect 9440 155 9640 160
rect 9440 125 9450 155
rect 9630 125 9640 155
rect 9440 100 9640 125
rect 9760 155 9960 160
rect 9760 125 9770 155
rect 9950 125 9960 155
rect 9760 100 9960 125
rect 10080 155 10280 160
rect 10080 125 10090 155
rect 10270 125 10280 155
rect 10080 100 10280 125
rect 5280 -20 5480 0
rect 5600 -20 5800 0
rect 5920 -20 6120 0
rect 6240 -20 6440 0
rect 6560 -20 6760 0
rect 6880 -20 7080 0
rect 7200 -20 7400 0
rect 7520 -20 7720 0
rect 7840 -20 8040 0
rect 8160 -20 8360 0
rect 8480 -20 8680 0
rect 8800 -20 9000 0
rect 9120 -20 9320 0
rect 9440 -20 9640 0
rect 9760 -20 9960 0
rect 10080 -20 10280 0
<< polycont >>
rect 10 605 190 635
rect 330 605 510 635
rect 650 605 830 635
rect 970 605 1150 635
rect 1290 605 1470 635
rect 1610 605 1790 635
rect 1930 605 2110 635
rect 2250 605 2430 635
rect 2570 605 2750 635
rect 2890 605 3070 635
rect 3210 605 3390 635
rect 3530 605 3710 635
rect 3850 605 4030 635
rect 4170 605 4350 635
rect 4490 605 4670 635
rect 4810 605 4990 635
rect 5290 605 5470 635
rect 5610 605 5790 635
rect 5930 605 6110 635
rect 6250 605 6430 635
rect 6570 605 6750 635
rect 6890 605 7070 635
rect 7210 605 7390 635
rect 7530 605 7710 635
rect 7850 605 8030 635
rect 8170 605 8350 635
rect 8490 605 8670 635
rect 8810 605 8990 635
rect 9130 605 9310 635
rect 9450 605 9630 635
rect 9770 605 9950 635
rect 10090 605 10270 635
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect 1290 125 1470 155
rect 1610 125 1790 155
rect 1930 125 2110 155
rect 2250 125 2430 155
rect 2570 125 2750 155
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3850 125 4030 155
rect 4170 125 4350 155
rect 4490 125 4670 155
rect 4810 125 4990 155
rect 5290 125 5470 155
rect 5610 125 5790 155
rect 5930 125 6110 155
rect 6250 125 6430 155
rect 6570 125 6750 155
rect 6890 125 7070 155
rect 7210 125 7390 155
rect 7530 125 7710 155
rect 7850 125 8030 155
rect 8170 125 8350 155
rect 8490 125 8670 155
rect 8810 125 8990 155
rect 9130 125 9310 155
rect 9450 125 9630 155
rect 9770 125 9950 155
rect 10090 125 10270 155
<< locali >>
rect -320 1000 -40 1040
rect 240 1000 280 1040
rect 560 1000 600 1040
rect 880 1000 920 1040
rect 1200 1000 1240 1040
rect 1520 1000 1560 1040
rect 1840 1000 1880 1040
rect 2160 1000 2200 1040
rect 2480 1000 2520 1040
rect 2800 1000 2840 1040
rect 3120 1000 3160 1040
rect 3440 1000 3480 1040
rect 3760 1000 3800 1040
rect 4080 1000 4120 1040
rect 4400 1000 4440 1040
rect 4720 1000 4760 1040
rect 5040 1000 5240 1040
rect 5520 1000 5560 1040
rect 5840 1000 5880 1040
rect 6160 1000 6200 1040
rect 6480 1000 6520 1040
rect 6800 1000 6840 1040
rect 7120 1000 7160 1040
rect 7440 1000 7480 1040
rect 7760 1000 7800 1040
rect 8080 1000 8120 1040
rect 8400 1000 8440 1040
rect 8720 1000 8760 1040
rect 9040 1000 9080 1040
rect 9360 1000 9400 1040
rect 9680 1000 9720 1040
rect 10000 1000 10040 1040
rect 10320 1000 10600 1040
rect -320 960 -280 1000
rect 10560 960 10600 1000
rect -160 840 -40 880
rect 240 840 280 880
rect 560 840 600 880
rect 880 840 920 880
rect 1200 840 1240 880
rect 1520 840 1560 880
rect 1840 840 1880 880
rect 2160 840 2200 880
rect 2480 840 2520 880
rect 2800 840 2840 880
rect 3120 840 3160 880
rect 3440 840 3480 880
rect 3760 840 3800 880
rect 4080 840 4120 880
rect 4400 840 4440 880
rect 4720 840 4760 880
rect 5040 840 5240 880
rect 5520 840 5560 880
rect -160 800 -120 840
rect -160 560 -120 600
rect -80 750 -40 840
rect 5120 800 5160 840
rect -80 670 -75 750
rect -45 670 -40 750
rect -80 560 -40 670
rect 240 750 280 760
rect 240 670 245 750
rect 275 670 280 750
rect 240 660 280 670
rect 560 750 600 760
rect 560 670 565 750
rect 595 670 600 750
rect 560 660 600 670
rect 880 750 920 760
rect 880 670 885 750
rect 915 670 920 750
rect 880 660 920 670
rect 1200 750 1240 760
rect 1200 670 1205 750
rect 1235 670 1240 750
rect 1200 660 1240 670
rect 1520 750 1560 760
rect 1520 670 1525 750
rect 1555 670 1560 750
rect 1520 660 1560 670
rect 1840 750 1880 760
rect 1840 670 1845 750
rect 1875 670 1880 750
rect 1840 660 1880 670
rect 2160 750 2200 760
rect 2160 670 2165 750
rect 2195 670 2200 750
rect 2160 660 2200 670
rect 2480 750 2520 760
rect 2480 670 2485 750
rect 2515 670 2520 750
rect 2480 660 2520 670
rect 2800 750 2840 760
rect 2800 670 2805 750
rect 2835 670 2840 750
rect 2800 660 2840 670
rect 3120 750 3160 760
rect 3120 670 3125 750
rect 3155 670 3160 750
rect 3120 660 3160 670
rect 3440 750 3480 760
rect 3440 670 3445 750
rect 3475 670 3480 750
rect 3440 660 3480 670
rect 3760 750 3800 760
rect 3760 670 3765 750
rect 3795 670 3800 750
rect 3760 660 3800 670
rect 4080 750 4120 760
rect 4080 670 4085 750
rect 4115 670 4120 750
rect 4080 660 4120 670
rect 4400 750 4440 760
rect 4400 670 4405 750
rect 4435 670 4440 750
rect 4400 660 4440 670
rect 4720 750 4760 760
rect 4720 670 4725 750
rect 4755 670 4760 750
rect 4720 660 4760 670
rect 5040 750 5080 760
rect 5040 670 5045 750
rect 5075 670 5080 750
rect 5040 660 5080 670
rect 0 635 200 640
rect 0 605 10 635
rect 190 605 200 635
rect 0 600 200 605
rect 320 635 520 640
rect 320 605 330 635
rect 510 605 520 635
rect 320 600 520 605
rect 640 635 840 640
rect 640 605 650 635
rect 830 605 840 635
rect 640 600 840 605
rect 960 635 1160 640
rect 960 605 970 635
rect 1150 605 1160 635
rect 960 600 1160 605
rect 1280 635 1480 640
rect 1280 605 1290 635
rect 1470 605 1480 635
rect 1280 600 1480 605
rect 1600 635 1800 640
rect 1600 605 1610 635
rect 1790 605 1800 635
rect 1600 600 1800 605
rect 1920 635 2120 640
rect 1920 605 1930 635
rect 2110 605 2120 635
rect 1920 600 2120 605
rect 2240 635 2440 640
rect 2240 605 2250 635
rect 2430 605 2440 635
rect 2240 600 2440 605
rect 2560 635 2760 640
rect 2560 605 2570 635
rect 2750 605 2760 635
rect 2560 600 2760 605
rect 2880 635 3080 640
rect 2880 605 2890 635
rect 3070 605 3080 635
rect 2880 600 3080 605
rect 3200 635 3400 640
rect 3200 605 3210 635
rect 3390 605 3400 635
rect 3200 600 3400 605
rect 3520 635 3720 640
rect 3520 605 3530 635
rect 3710 605 3720 635
rect 3520 600 3720 605
rect 3840 635 4040 640
rect 3840 605 3850 635
rect 4030 605 4040 635
rect 3840 600 4040 605
rect 4160 635 4360 640
rect 4160 605 4170 635
rect 4350 605 4360 635
rect 4160 600 4360 605
rect 4480 635 4680 640
rect 4480 605 4490 635
rect 4670 605 4680 635
rect 4480 600 4680 605
rect 4800 635 5000 640
rect 4800 605 4810 635
rect 4990 605 5000 635
rect 4800 600 5000 605
rect 5120 560 5160 600
rect 5200 750 5240 840
rect 5200 670 5205 750
rect 5235 670 5240 750
rect 5200 560 5240 670
rect 5520 750 5560 760
rect 5520 670 5525 750
rect 5555 670 5560 750
rect 5520 660 5560 670
rect 5840 750 5880 880
rect 6160 840 6200 880
rect 5840 670 5845 750
rect 5875 670 5880 750
rect 5280 635 5480 640
rect 5280 605 5290 635
rect 5470 605 5480 635
rect 5280 600 5480 605
rect 5600 635 5800 640
rect 5600 605 5610 635
rect 5790 605 5800 635
rect 5600 600 5800 605
rect -160 520 -40 560
rect 240 520 280 560
rect 560 520 600 560
rect 880 520 920 560
rect 1200 520 1240 560
rect 1520 520 1560 560
rect 1840 520 1880 560
rect 2160 520 2200 560
rect 2480 520 2520 560
rect 2800 520 2840 560
rect 3120 520 3160 560
rect 3440 520 3480 560
rect 3760 520 3800 560
rect 4080 520 4120 560
rect 4400 520 4440 560
rect 4720 520 4760 560
rect 5040 520 5240 560
rect 5520 520 5560 560
rect 5840 520 5880 670
rect 6160 750 6200 760
rect 6160 670 6165 750
rect 6195 670 6200 750
rect 6160 660 6200 670
rect 6480 750 6520 880
rect 6800 840 6840 880
rect 6480 670 6485 750
rect 6515 670 6520 750
rect 5920 635 6120 640
rect 5920 605 5930 635
rect 6110 605 6120 635
rect 5920 600 6120 605
rect 6240 635 6440 640
rect 6240 605 6250 635
rect 6430 605 6440 635
rect 6240 600 6440 605
rect 6160 520 6200 560
rect 6480 520 6520 670
rect 6800 750 6840 760
rect 6800 670 6805 750
rect 6835 670 6840 750
rect 6800 660 6840 670
rect 7120 750 7160 880
rect 7440 840 7480 880
rect 7120 670 7125 750
rect 7155 670 7160 750
rect 6560 635 6760 640
rect 6560 605 6570 635
rect 6750 605 6760 635
rect 6560 600 6760 605
rect 6880 635 7080 640
rect 6880 605 6890 635
rect 7070 605 7080 635
rect 6880 600 7080 605
rect 6800 520 6840 560
rect 7120 520 7160 670
rect 7440 750 7480 760
rect 7440 670 7445 750
rect 7475 670 7480 750
rect 7440 660 7480 670
rect 7760 750 7800 880
rect 8080 840 8120 880
rect 7760 670 7765 750
rect 7795 670 7800 750
rect 7200 635 7400 640
rect 7200 605 7210 635
rect 7390 605 7400 635
rect 7200 600 7400 605
rect 7520 635 7720 640
rect 7520 605 7530 635
rect 7710 605 7720 635
rect 7520 600 7720 605
rect 7440 520 7480 560
rect 7760 520 7800 670
rect 8080 750 8120 760
rect 8080 670 8085 750
rect 8115 670 8120 750
rect 8080 660 8120 670
rect 8400 750 8440 880
rect 8720 840 8760 880
rect 8400 670 8405 750
rect 8435 670 8440 750
rect 7840 635 8040 640
rect 7840 605 7850 635
rect 8030 605 8040 635
rect 7840 600 8040 605
rect 8160 635 8360 640
rect 8160 605 8170 635
rect 8350 605 8360 635
rect 8160 600 8360 605
rect 8080 520 8120 560
rect 8400 520 8440 670
rect 8720 750 8760 760
rect 8720 670 8725 750
rect 8755 670 8760 750
rect 8720 660 8760 670
rect 9040 750 9080 880
rect 9360 840 9400 880
rect 9040 670 9045 750
rect 9075 670 9080 750
rect 8480 635 8680 640
rect 8480 605 8490 635
rect 8670 605 8680 635
rect 8480 600 8680 605
rect 8800 635 9000 640
rect 8800 605 8810 635
rect 8990 605 9000 635
rect 8800 600 9000 605
rect 8720 520 8760 560
rect 9040 520 9080 670
rect 9360 750 9400 760
rect 9360 670 9365 750
rect 9395 670 9400 750
rect 9360 660 9400 670
rect 9680 750 9720 880
rect 10000 840 10040 880
rect 10320 840 10480 880
rect 9680 670 9685 750
rect 9715 670 9720 750
rect 9120 635 9320 640
rect 9120 605 9130 635
rect 9310 605 9320 635
rect 9120 600 9320 605
rect 9440 635 9640 640
rect 9440 605 9450 635
rect 9630 605 9640 635
rect 9440 600 9640 605
rect 9360 520 9400 560
rect 9680 520 9720 670
rect 10000 750 10040 760
rect 10000 670 10005 750
rect 10035 670 10040 750
rect 10000 660 10040 670
rect 10320 750 10360 840
rect 10320 670 10325 750
rect 10355 670 10360 750
rect 9760 635 9960 640
rect 9760 605 9770 635
rect 9950 605 9960 635
rect 9760 600 9960 605
rect 10080 635 10280 640
rect 10080 605 10090 635
rect 10270 605 10280 635
rect 10080 600 10280 605
rect 10320 560 10360 670
rect 10400 800 10440 840
rect 10400 560 10440 600
rect 10000 520 10040 560
rect 10320 520 10480 560
rect -280 360 -40 400
rect 240 360 280 400
rect 560 360 600 400
rect 880 360 920 400
rect 1200 360 1240 400
rect 1520 360 1560 400
rect 1840 360 1880 400
rect 2160 360 2200 400
rect 2480 360 2520 400
rect 2800 360 2840 400
rect 3120 360 3160 400
rect 3440 360 3480 400
rect 3760 360 3800 400
rect 4080 360 4120 400
rect 4400 360 4440 400
rect 4720 360 4760 400
rect 5040 360 5240 400
rect 5520 360 5560 400
rect 5840 360 5880 400
rect 6160 360 6200 400
rect 6480 360 6520 400
rect 6800 360 6840 400
rect 7120 360 7160 400
rect 7440 360 7480 400
rect 7760 360 7800 400
rect 8080 360 8120 400
rect 8400 360 8440 400
rect 8720 360 8760 400
rect 9040 360 9080 400
rect 9360 360 9400 400
rect 9680 360 9720 400
rect 10000 360 10040 400
rect 10320 360 10560 400
rect -320 -80 -280 -40
rect -160 200 -40 240
rect 240 200 280 240
rect 560 200 600 240
rect 880 200 920 240
rect 1200 200 1240 240
rect 1520 200 1560 240
rect 1840 200 1880 240
rect 2160 200 2200 240
rect -160 160 -120 200
rect -160 -80 -120 -40
rect -80 90 -40 200
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 120 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 120 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 120 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 120 1160 125
rect 1280 155 1480 160
rect 1280 125 1290 155
rect 1470 125 1480 155
rect 1280 120 1480 125
rect 1600 155 1800 160
rect 1600 125 1610 155
rect 1790 125 1800 155
rect 1600 120 1800 125
rect 1920 155 2120 160
rect 1920 125 1930 155
rect 2110 125 2120 155
rect 1920 120 2120 125
rect 2240 155 2440 160
rect 2240 125 2250 155
rect 2430 125 2440 155
rect 2240 120 2440 125
rect -80 10 -75 90
rect -45 10 -40 90
rect -80 -80 -40 10
rect 240 90 280 100
rect 240 10 245 90
rect 275 10 280 90
rect 240 0 280 10
rect 560 90 600 100
rect 560 10 565 90
rect 595 10 600 90
rect 560 0 600 10
rect 880 90 920 100
rect 880 10 885 90
rect 915 10 920 90
rect 880 0 920 10
rect 1200 90 1240 100
rect 1200 10 1205 90
rect 1235 10 1240 90
rect 1200 0 1240 10
rect 1520 90 1560 100
rect 1520 10 1525 90
rect 1555 10 1560 90
rect 1520 0 1560 10
rect 1840 90 1880 100
rect 1840 10 1845 90
rect 1875 10 1880 90
rect 1840 0 1880 10
rect 2160 90 2200 100
rect 2160 10 2165 90
rect 2195 10 2200 90
rect 2160 0 2200 10
rect 2480 90 2520 240
rect 2800 200 2840 240
rect 3120 200 3160 240
rect 3440 200 3480 240
rect 3760 200 3800 240
rect 4080 200 4120 240
rect 4400 200 4440 240
rect 4720 200 4760 240
rect 5040 200 5240 240
rect 5520 200 5560 240
rect 5840 200 5880 240
rect 6160 200 6200 240
rect 6480 200 6520 240
rect 6800 200 6840 240
rect 7120 200 7160 240
rect 7440 200 7480 240
rect 2560 155 2760 160
rect 2560 125 2570 155
rect 2750 125 2760 155
rect 2560 120 2760 125
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 120 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 120 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 120 3720 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 120 4040 125
rect 4160 155 4360 160
rect 4160 125 4170 155
rect 4350 125 4360 155
rect 4160 120 4360 125
rect 4480 155 4680 160
rect 4480 125 4490 155
rect 4670 125 4680 155
rect 4480 120 4680 125
rect 4800 155 5000 160
rect 4800 125 4810 155
rect 4990 125 5000 155
rect 4800 120 5000 125
rect 2480 10 2485 90
rect 2515 10 2520 90
rect -320 -120 -40 -80
rect 240 -120 280 -80
rect 560 -120 600 -80
rect 880 -120 920 -80
rect 1200 -120 1240 -80
rect 1520 -120 1560 -80
rect 1840 -120 1880 -80
rect 2160 -120 2200 -80
rect 2480 -120 2520 10
rect 2800 90 2840 100
rect 2800 10 2805 90
rect 2835 10 2840 90
rect 2800 0 2840 10
rect 3120 90 3160 100
rect 3120 10 3125 90
rect 3155 10 3160 90
rect 3120 0 3160 10
rect 3440 90 3480 100
rect 3440 10 3445 90
rect 3475 10 3480 90
rect 3440 0 3480 10
rect 3760 90 3800 100
rect 3760 10 3765 90
rect 3795 10 3800 90
rect 3760 0 3800 10
rect 4080 90 4120 100
rect 4080 10 4085 90
rect 4115 10 4120 90
rect 4080 0 4120 10
rect 4400 90 4440 100
rect 4400 10 4405 90
rect 4435 10 4440 90
rect 4400 0 4440 10
rect 4720 90 4760 100
rect 4720 10 4725 90
rect 4755 10 4760 90
rect 4720 0 4760 10
rect 5040 90 5080 200
rect 5040 10 5045 90
rect 5075 10 5080 90
rect 5040 -80 5080 10
rect 5120 160 5160 200
rect 5120 -80 5160 -40
rect 5200 90 5240 200
rect 5280 155 5480 160
rect 5280 125 5290 155
rect 5470 125 5480 155
rect 5280 120 5480 125
rect 5600 155 5800 160
rect 5600 125 5610 155
rect 5790 125 5800 155
rect 5600 120 5800 125
rect 5920 155 6120 160
rect 5920 125 5930 155
rect 6110 125 6120 155
rect 5920 120 6120 125
rect 6240 155 6440 160
rect 6240 125 6250 155
rect 6430 125 6440 155
rect 6240 120 6440 125
rect 6560 155 6760 160
rect 6560 125 6570 155
rect 6750 125 6760 155
rect 6560 120 6760 125
rect 6880 155 7080 160
rect 6880 125 6890 155
rect 7070 125 7080 155
rect 6880 120 7080 125
rect 7200 155 7400 160
rect 7200 125 7210 155
rect 7390 125 7400 155
rect 7200 120 7400 125
rect 7520 155 7720 160
rect 7520 125 7530 155
rect 7710 125 7720 155
rect 7520 120 7720 125
rect 5200 10 5205 90
rect 5235 10 5240 90
rect 5200 -80 5240 10
rect 5520 90 5560 100
rect 5520 10 5525 90
rect 5555 10 5560 90
rect 5520 0 5560 10
rect 5840 90 5880 100
rect 5840 10 5845 90
rect 5875 10 5880 90
rect 5840 0 5880 10
rect 6160 90 6200 100
rect 6160 10 6165 90
rect 6195 10 6200 90
rect 6160 0 6200 10
rect 6480 90 6520 100
rect 6480 10 6485 90
rect 6515 10 6520 90
rect 6480 0 6520 10
rect 6800 90 6840 100
rect 6800 10 6805 90
rect 6835 10 6840 90
rect 6800 0 6840 10
rect 7120 90 7160 100
rect 7120 10 7125 90
rect 7155 10 7160 90
rect 7120 0 7160 10
rect 7440 90 7480 100
rect 7440 10 7445 90
rect 7475 10 7480 90
rect 7440 0 7480 10
rect 7760 90 7800 240
rect 8080 200 8120 240
rect 8400 200 8440 240
rect 8720 200 8760 240
rect 9040 200 9080 240
rect 9360 200 9400 240
rect 9680 200 9720 240
rect 10000 200 10040 240
rect 10320 200 10480 240
rect 7840 155 8040 160
rect 7840 125 7850 155
rect 8030 125 8040 155
rect 7840 120 8040 125
rect 8160 155 8360 160
rect 8160 125 8170 155
rect 8350 125 8360 155
rect 8160 120 8360 125
rect 8480 155 8680 160
rect 8480 125 8490 155
rect 8670 125 8680 155
rect 8480 120 8680 125
rect 8800 155 9000 160
rect 8800 125 8810 155
rect 8990 125 9000 155
rect 8800 120 9000 125
rect 9120 155 9320 160
rect 9120 125 9130 155
rect 9310 125 9320 155
rect 9120 120 9320 125
rect 9440 155 9640 160
rect 9440 125 9450 155
rect 9630 125 9640 155
rect 9440 120 9640 125
rect 9760 155 9960 160
rect 9760 125 9770 155
rect 9950 125 9960 155
rect 9760 120 9960 125
rect 10080 155 10280 160
rect 10080 125 10090 155
rect 10270 125 10280 155
rect 10080 120 10280 125
rect 7760 10 7765 90
rect 7795 10 7800 90
rect 2800 -120 2840 -80
rect 3120 -120 3160 -80
rect 3440 -120 3480 -80
rect 3760 -120 3800 -80
rect 4080 -120 4120 -80
rect 4400 -120 4440 -80
rect 4720 -120 4760 -80
rect 5040 -120 5240 -80
rect 5520 -120 5560 -80
rect 5840 -120 5880 -80
rect 6160 -120 6200 -80
rect 6480 -120 6520 -80
rect 6800 -120 6840 -80
rect 7120 -120 7160 -80
rect 7440 -120 7480 -80
rect 7760 -120 7800 10
rect 8080 90 8120 100
rect 8080 10 8085 90
rect 8115 10 8120 90
rect 8080 0 8120 10
rect 8400 90 8440 100
rect 8400 10 8405 90
rect 8435 10 8440 90
rect 8400 0 8440 10
rect 8720 90 8760 100
rect 8720 10 8725 90
rect 8755 10 8760 90
rect 8720 0 8760 10
rect 9040 90 9080 100
rect 9040 10 9045 90
rect 9075 10 9080 90
rect 9040 0 9080 10
rect 9360 90 9400 100
rect 9360 10 9365 90
rect 9395 10 9400 90
rect 9360 0 9400 10
rect 9680 90 9720 100
rect 9680 10 9685 90
rect 9715 10 9720 90
rect 9680 0 9720 10
rect 10000 90 10040 100
rect 10000 10 10005 90
rect 10035 10 10040 90
rect 10000 0 10040 10
rect 10320 90 10360 200
rect 10320 10 10325 90
rect 10355 10 10360 90
rect 10320 -80 10360 10
rect 10400 160 10440 200
rect 10400 -80 10440 -40
rect 10560 -80 10600 -40
rect 8080 -120 8120 -80
rect 8400 -120 8440 -80
rect 8720 -120 8760 -80
rect 9040 -120 9080 -80
rect 9360 -120 9400 -80
rect 9680 -120 9720 -80
rect 10000 -120 10040 -80
rect 10320 -120 10600 -80
<< viali >>
rect -75 670 -45 750
rect 245 670 275 750
rect 565 670 595 750
rect 885 670 915 750
rect 1205 670 1235 750
rect 1525 670 1555 750
rect 1845 670 1875 750
rect 2165 670 2195 750
rect 2485 670 2515 750
rect 2805 670 2835 750
rect 3125 670 3155 750
rect 3445 670 3475 750
rect 3765 670 3795 750
rect 4085 670 4115 750
rect 4405 670 4435 750
rect 4725 670 4755 750
rect 5045 670 5075 750
rect 10 605 190 635
rect 330 605 510 635
rect 650 605 830 635
rect 970 605 1150 635
rect 1290 605 1470 635
rect 1610 605 1790 635
rect 1930 605 2110 635
rect 2250 605 2430 635
rect 2570 605 2750 635
rect 2890 605 3070 635
rect 3210 605 3390 635
rect 3530 605 3710 635
rect 3850 605 4030 635
rect 4170 605 4350 635
rect 4490 605 4670 635
rect 4810 605 4990 635
rect 5205 670 5235 750
rect 5525 670 5555 750
rect 5845 670 5875 750
rect 5290 605 5470 635
rect 5610 605 5790 635
rect 6165 670 6195 750
rect 6485 670 6515 750
rect 5930 605 6110 635
rect 6250 605 6430 635
rect 6805 670 6835 750
rect 7125 670 7155 750
rect 6570 605 6750 635
rect 6890 605 7070 635
rect 7445 670 7475 750
rect 7765 670 7795 750
rect 7210 605 7390 635
rect 7530 605 7710 635
rect 8085 670 8115 750
rect 8405 670 8435 750
rect 7850 605 8030 635
rect 8170 605 8350 635
rect 8725 670 8755 750
rect 9045 670 9075 750
rect 8490 605 8670 635
rect 8810 605 8990 635
rect 9365 670 9395 750
rect 9685 670 9715 750
rect 9130 605 9310 635
rect 9450 605 9630 635
rect 10005 670 10035 750
rect 10325 670 10355 750
rect 9770 605 9950 635
rect 10090 605 10270 635
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect 1290 125 1470 155
rect 1610 125 1790 155
rect 1930 125 2110 155
rect 2250 125 2430 155
rect -75 10 -45 90
rect 245 10 275 90
rect 565 10 595 90
rect 885 10 915 90
rect 1205 10 1235 90
rect 1525 10 1555 90
rect 1845 10 1875 90
rect 2165 10 2195 90
rect 2570 125 2750 155
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3850 125 4030 155
rect 4170 125 4350 155
rect 4490 125 4670 155
rect 4810 125 4990 155
rect 2485 10 2515 90
rect 2805 10 2835 90
rect 3125 10 3155 90
rect 3445 10 3475 90
rect 3765 10 3795 90
rect 4085 10 4115 90
rect 4405 10 4435 90
rect 4725 10 4755 90
rect 5045 10 5075 90
rect 5290 125 5470 155
rect 5610 125 5790 155
rect 5930 125 6110 155
rect 6250 125 6430 155
rect 6570 125 6750 155
rect 6890 125 7070 155
rect 7210 125 7390 155
rect 7530 125 7710 155
rect 5205 10 5235 90
rect 5525 10 5555 90
rect 5845 10 5875 90
rect 6165 10 6195 90
rect 6485 10 6515 90
rect 6805 10 6835 90
rect 7125 10 7155 90
rect 7445 10 7475 90
rect 7850 125 8030 155
rect 8170 125 8350 155
rect 8490 125 8670 155
rect 8810 125 8990 155
rect 9130 125 9310 155
rect 9450 125 9630 155
rect 9770 125 9950 155
rect 10090 125 10270 155
rect 7765 10 7795 90
rect 8085 10 8115 90
rect 8405 10 8435 90
rect 8725 10 8755 90
rect 9045 10 9075 90
rect 9365 10 9395 90
rect 9685 10 9715 90
rect 10005 10 10035 90
rect 10325 10 10355 90
<< metal1 >>
rect -720 1035 -680 1040
rect -720 1005 -715 1035
rect -685 1005 -680 1035
rect -720 1000 -680 1005
rect -560 1035 -520 1040
rect -560 1005 -555 1035
rect -525 1005 -520 1035
rect -560 1000 -520 1005
rect -400 1035 -360 1040
rect -400 1005 -395 1035
rect -365 1005 -360 1035
rect -400 1000 -360 1005
rect 10640 1035 10680 1040
rect 10640 1005 10645 1035
rect 10675 1005 10680 1035
rect 10640 1000 10680 1005
rect 10800 1035 10840 1040
rect 10800 1005 10805 1035
rect 10835 1005 10840 1035
rect 10800 1000 10840 1005
rect 10960 1035 11000 1040
rect 10960 1005 10965 1035
rect 10995 1005 11000 1035
rect 10960 1000 11000 1005
rect -720 955 -680 960
rect -720 925 -715 955
rect -685 925 -680 955
rect -720 920 -680 925
rect -560 955 -520 960
rect -560 925 -555 955
rect -525 925 -520 955
rect -560 920 -520 925
rect -400 955 -360 960
rect -400 925 -395 955
rect -365 925 -360 955
rect -400 920 -360 925
rect 10640 955 10680 960
rect 10640 925 10645 955
rect 10675 925 10680 955
rect 10640 920 10680 925
rect 10800 955 10840 960
rect 10800 925 10805 955
rect 10835 925 10840 955
rect 10800 920 10840 925
rect 10960 955 11000 960
rect 10960 925 10965 955
rect 10995 925 11000 955
rect 10960 920 11000 925
rect -720 875 -680 880
rect -720 845 -715 875
rect -685 845 -680 875
rect -720 840 -680 845
rect -560 875 -520 880
rect -560 845 -555 875
rect -525 845 -520 875
rect -560 840 -520 845
rect -400 875 -360 880
rect -400 845 -395 875
rect -365 845 -360 875
rect -400 840 -360 845
rect 10640 875 10680 880
rect 10640 845 10645 875
rect 10675 845 10680 875
rect 10640 840 10680 845
rect 10800 875 10840 880
rect 10800 845 10805 875
rect 10835 845 10840 875
rect 10800 840 10840 845
rect 10960 875 11000 880
rect 10960 845 10965 875
rect 10995 845 11000 875
rect 10960 840 11000 845
rect -80 795 -40 800
rect -80 765 -75 795
rect -45 765 -40 795
rect -80 750 -40 765
rect 5200 795 5240 800
rect 5200 765 5205 795
rect 5235 765 5240 795
rect -80 670 -75 750
rect -45 670 -40 750
rect -80 660 -40 670
rect 240 750 280 760
rect 240 670 245 750
rect 275 670 280 750
rect 240 660 280 670
rect 560 750 600 760
rect 560 670 565 750
rect 595 670 600 750
rect 560 660 600 670
rect 880 750 920 760
rect 880 670 885 750
rect 915 670 920 750
rect 880 660 920 670
rect 1200 750 1240 760
rect 1200 670 1205 750
rect 1235 670 1240 750
rect 1200 660 1240 670
rect 1520 750 1560 760
rect 1520 670 1525 750
rect 1555 670 1560 750
rect 1520 660 1560 670
rect 1840 750 1880 760
rect 1840 670 1845 750
rect 1875 670 1880 750
rect 1840 660 1880 670
rect 2160 750 2200 760
rect 2160 670 2165 750
rect 2195 670 2200 750
rect 2160 660 2200 670
rect 2480 750 2520 760
rect 2480 670 2485 750
rect 2515 670 2520 750
rect 2480 660 2520 670
rect 2800 750 2840 760
rect 2800 670 2805 750
rect 2835 670 2840 750
rect 2800 660 2840 670
rect 3120 750 3160 760
rect 3120 670 3125 750
rect 3155 670 3160 750
rect 3120 660 3160 670
rect 3440 750 3480 760
rect 3440 670 3445 750
rect 3475 670 3480 750
rect 3440 660 3480 670
rect 3760 750 3800 760
rect 3760 670 3765 750
rect 3795 670 3800 750
rect 3760 660 3800 670
rect 4080 750 4120 760
rect 4080 670 4085 750
rect 4115 670 4120 750
rect 4080 660 4120 670
rect 4400 750 4440 760
rect 4400 670 4405 750
rect 4435 670 4440 750
rect 4400 660 4440 670
rect 4720 750 4760 760
rect 4720 670 4725 750
rect 4755 670 4760 750
rect 4720 660 4760 670
rect 5040 750 5080 760
rect 5040 670 5045 750
rect 5075 670 5080 750
rect -720 635 -680 640
rect -720 605 -715 635
rect -685 605 -680 635
rect -720 600 -680 605
rect -560 635 -520 640
rect -560 605 -555 635
rect -525 605 -520 635
rect -560 600 -520 605
rect -400 635 -360 640
rect -400 605 -395 635
rect -365 605 -360 635
rect -400 600 -360 605
rect 0 635 200 640
rect 0 605 10 635
rect 190 605 200 635
rect 0 600 200 605
rect 320 635 520 640
rect 320 605 330 635
rect 510 605 520 635
rect 320 600 520 605
rect 640 635 840 640
rect 640 605 650 635
rect 830 605 840 635
rect 640 600 840 605
rect 960 635 1160 640
rect 960 605 970 635
rect 1150 605 1160 635
rect 960 600 1160 605
rect 1280 635 1480 640
rect 1280 605 1290 635
rect 1470 605 1480 635
rect 1280 600 1480 605
rect 1600 635 1800 640
rect 1600 605 1610 635
rect 1790 605 1800 635
rect 1600 600 1800 605
rect 1920 635 2120 640
rect 1920 605 1930 635
rect 2110 605 2120 635
rect 1920 600 2120 605
rect 2240 635 2440 640
rect 2240 605 2250 635
rect 2430 605 2440 635
rect 2240 600 2440 605
rect 2560 635 2760 640
rect 2560 605 2570 635
rect 2750 605 2760 635
rect 2560 600 2760 605
rect 2880 635 3080 640
rect 2880 605 2890 635
rect 3070 605 3080 635
rect 2880 600 3080 605
rect 3200 635 3400 640
rect 3200 605 3210 635
rect 3390 605 3400 635
rect 3200 600 3400 605
rect 3520 635 3720 640
rect 3520 605 3530 635
rect 3710 605 3720 635
rect 3520 600 3720 605
rect 3840 635 4040 640
rect 3840 605 3850 635
rect 4030 605 4040 635
rect 3840 600 4040 605
rect 4160 635 4360 640
rect 4160 605 4170 635
rect 4350 605 4360 635
rect 4160 600 4360 605
rect 4480 635 4680 640
rect 4480 605 4490 635
rect 4670 605 4680 635
rect 4480 600 4680 605
rect 4800 635 5000 640
rect 4800 605 4810 635
rect 4990 605 5000 635
rect 4800 600 5000 605
rect -720 555 -680 560
rect -720 525 -715 555
rect -685 525 -680 555
rect -720 520 -680 525
rect -560 555 -520 560
rect -560 525 -555 555
rect -525 525 -520 555
rect -560 520 -520 525
rect -400 555 -360 560
rect -400 525 -395 555
rect -365 525 -360 555
rect -400 520 -360 525
rect -720 475 -680 480
rect -720 445 -715 475
rect -685 445 -680 475
rect -720 440 -680 445
rect -560 475 -520 480
rect -560 445 -555 475
rect -525 445 -520 475
rect -560 440 -520 445
rect 80 475 120 600
rect 80 445 85 475
rect 115 445 120 475
rect 80 440 120 445
rect 400 475 440 600
rect 400 445 405 475
rect 435 445 440 475
rect 400 440 440 445
rect 720 475 760 600
rect 720 445 725 475
rect 755 445 760 475
rect 720 440 760 445
rect 1040 475 1080 600
rect 1040 445 1045 475
rect 1075 445 1080 475
rect 1040 440 1080 445
rect 1360 475 1400 600
rect 1360 445 1365 475
rect 1395 445 1400 475
rect 1360 440 1400 445
rect 1680 475 1720 600
rect 1680 445 1685 475
rect 1715 445 1720 475
rect 1680 440 1720 445
rect 2000 475 2040 600
rect 2000 445 2005 475
rect 2035 445 2040 475
rect 2000 440 2040 445
rect 2320 475 2360 600
rect 2320 445 2325 475
rect 2355 445 2360 475
rect 2320 440 2360 445
rect 2640 475 2680 600
rect 2640 445 2645 475
rect 2675 445 2680 475
rect 2640 440 2680 445
rect 2960 475 3000 600
rect 2960 445 2965 475
rect 2995 445 3000 475
rect 2960 440 3000 445
rect 3280 475 3320 600
rect 3280 445 3285 475
rect 3315 445 3320 475
rect 3280 440 3320 445
rect 3600 475 3640 600
rect 3600 445 3605 475
rect 3635 445 3640 475
rect 3600 440 3640 445
rect 3920 475 3960 600
rect 3920 445 3925 475
rect 3955 445 3960 475
rect 3920 440 3960 445
rect 4240 475 4280 600
rect 4240 445 4245 475
rect 4275 445 4280 475
rect 4240 440 4280 445
rect 4560 475 4600 600
rect 4560 445 4565 475
rect 4595 445 4600 475
rect 4560 440 4600 445
rect 4880 475 4920 600
rect 4880 445 4885 475
rect 4915 445 4920 475
rect 4880 440 4920 445
rect -720 395 -680 400
rect -720 365 -715 395
rect -685 365 -680 395
rect -720 360 -680 365
rect -560 395 -520 400
rect -560 365 -555 395
rect -525 365 -520 395
rect -560 360 -520 365
rect -400 395 -360 400
rect -400 365 -395 395
rect -365 365 -360 395
rect -400 360 -360 365
rect -720 315 -680 320
rect -720 285 -715 315
rect -685 285 -680 315
rect -720 280 -680 285
rect -560 315 -520 320
rect -560 285 -555 315
rect -525 285 -520 315
rect -560 280 -520 285
rect -400 315 -360 320
rect -400 285 -395 315
rect -365 285 -360 315
rect -400 280 -360 285
rect -720 235 -680 240
rect -720 205 -715 235
rect -685 205 -680 235
rect -720 200 -680 205
rect -560 235 -520 240
rect -560 205 -555 235
rect -525 205 -520 235
rect -560 200 -520 205
rect -400 235 -360 240
rect -400 205 -395 235
rect -365 205 -360 235
rect -400 200 -360 205
rect -720 155 -680 160
rect -720 125 -715 155
rect -685 125 -680 155
rect -720 120 -680 125
rect -560 155 -520 160
rect -560 125 -555 155
rect -525 125 -520 155
rect -560 120 -520 125
rect -400 155 -360 160
rect -400 125 -395 155
rect -365 125 -360 155
rect -400 120 -360 125
rect 0 155 200 160
rect 0 125 10 155
rect 190 125 200 155
rect 0 120 200 125
rect 320 155 520 160
rect 320 125 330 155
rect 510 125 520 155
rect 320 120 520 125
rect 640 155 840 160
rect 640 125 650 155
rect 830 125 840 155
rect 640 120 840 125
rect 960 155 1160 160
rect 960 125 970 155
rect 1150 125 1160 155
rect 960 120 1160 125
rect 1200 155 1240 160
rect 1200 125 1205 155
rect 1235 125 1240 155
rect -80 90 -40 100
rect -720 75 -680 80
rect -720 45 -715 75
rect -685 45 -680 75
rect -720 40 -680 45
rect -560 75 -520 80
rect -560 45 -555 75
rect -525 45 -520 75
rect -560 40 -520 45
rect -400 75 -360 80
rect -400 45 -395 75
rect -365 45 -360 75
rect -400 40 -360 45
rect -80 10 -75 90
rect -45 10 -40 90
rect -720 -5 -680 0
rect -720 -35 -715 -5
rect -685 -35 -680 -5
rect -720 -40 -680 -35
rect -560 -5 -520 0
rect -560 -35 -555 -5
rect -525 -35 -520 -5
rect -560 -40 -520 -35
rect -400 -5 -360 0
rect -400 -35 -395 -5
rect -365 -35 -360 -5
rect -400 -40 -360 -35
rect -80 -5 -40 10
rect 240 90 280 100
rect 240 10 245 90
rect 275 10 280 90
rect 240 0 280 10
rect 560 90 600 100
rect 560 10 565 90
rect 595 10 600 90
rect 560 0 600 10
rect 880 90 920 100
rect 880 10 885 90
rect 915 10 920 90
rect 880 0 920 10
rect 1200 90 1240 125
rect 1280 155 1480 160
rect 1280 125 1290 155
rect 1470 125 1480 155
rect 1280 120 1480 125
rect 1600 155 1800 160
rect 1600 125 1610 155
rect 1790 125 1800 155
rect 1600 120 1800 125
rect 1920 155 2120 160
rect 1920 125 1930 155
rect 2110 125 2120 155
rect 1920 120 2120 125
rect 2240 155 2440 160
rect 2240 125 2250 155
rect 2430 125 2440 155
rect 2240 120 2440 125
rect 2560 155 2760 160
rect 2560 125 2570 155
rect 2750 125 2760 155
rect 2560 120 2760 125
rect 2880 155 3080 160
rect 2880 125 2890 155
rect 3070 125 3080 155
rect 2880 120 3080 125
rect 3200 155 3400 160
rect 3200 125 3210 155
rect 3390 125 3400 155
rect 3200 120 3400 125
rect 3520 155 3720 160
rect 3520 125 3530 155
rect 3710 125 3720 155
rect 3520 120 3720 125
rect 3760 155 3800 160
rect 3760 125 3765 155
rect 3795 125 3800 155
rect 1200 10 1205 90
rect 1235 10 1240 90
rect 1200 0 1240 10
rect 1520 90 1560 100
rect 1520 10 1525 90
rect 1555 10 1560 90
rect 1520 0 1560 10
rect 1840 90 1880 100
rect 1840 10 1845 90
rect 1875 10 1880 90
rect 1840 0 1880 10
rect 2160 90 2200 100
rect 2160 10 2165 90
rect 2195 10 2200 90
rect 2160 0 2200 10
rect 2480 90 2520 100
rect 2480 10 2485 90
rect 2515 10 2520 90
rect -80 -35 -75 -5
rect -45 -35 -40 -5
rect -80 -40 -40 -35
rect 2480 -5 2520 10
rect 2800 90 2840 100
rect 2800 10 2805 90
rect 2835 10 2840 90
rect 2800 0 2840 10
rect 3120 90 3160 100
rect 3120 10 3125 90
rect 3155 10 3160 90
rect 3120 0 3160 10
rect 3440 90 3480 100
rect 3440 10 3445 90
rect 3475 10 3480 90
rect 3440 0 3480 10
rect 3760 90 3800 125
rect 3840 155 4040 160
rect 3840 125 3850 155
rect 4030 125 4040 155
rect 3840 120 4040 125
rect 4160 155 4360 160
rect 4160 125 4170 155
rect 4350 125 4360 155
rect 4160 120 4360 125
rect 4480 155 4680 160
rect 4480 125 4490 155
rect 4670 125 4680 155
rect 4480 120 4680 125
rect 4800 155 5000 160
rect 4800 125 4810 155
rect 4990 125 5000 155
rect 4800 120 5000 125
rect 5040 155 5080 670
rect 5200 750 5240 765
rect 5840 795 5880 800
rect 5840 765 5845 795
rect 5875 765 5880 795
rect 5200 670 5205 750
rect 5235 670 5240 750
rect 5200 660 5240 670
rect 5520 750 5560 760
rect 5520 670 5525 750
rect 5555 670 5560 750
rect 5280 635 5480 640
rect 5280 605 5290 635
rect 5470 605 5480 635
rect 5280 600 5480 605
rect 5360 315 5400 600
rect 5360 285 5365 315
rect 5395 285 5400 315
rect 5360 280 5400 285
rect 5520 315 5560 670
rect 5840 750 5880 765
rect 6480 795 6520 800
rect 6480 765 6485 795
rect 6515 765 6520 795
rect 5840 670 5845 750
rect 5875 670 5880 750
rect 5840 660 5880 670
rect 6160 750 6200 760
rect 6160 670 6165 750
rect 6195 670 6200 750
rect 6160 660 6200 670
rect 6480 750 6520 765
rect 7120 795 7160 800
rect 7120 765 7125 795
rect 7155 765 7160 795
rect 6480 670 6485 750
rect 6515 670 6520 750
rect 6480 660 6520 670
rect 6800 750 6840 760
rect 6800 670 6805 750
rect 6835 670 6840 750
rect 6800 660 6840 670
rect 7120 750 7160 765
rect 7760 795 7800 800
rect 7760 765 7765 795
rect 7795 765 7800 795
rect 7120 670 7125 750
rect 7155 670 7160 750
rect 7120 660 7160 670
rect 7440 750 7480 760
rect 7440 670 7445 750
rect 7475 670 7480 750
rect 7440 660 7480 670
rect 7760 750 7800 765
rect 8400 795 8440 800
rect 8400 765 8405 795
rect 8435 765 8440 795
rect 7760 670 7765 750
rect 7795 670 7800 750
rect 7760 660 7800 670
rect 8080 750 8120 760
rect 8080 670 8085 750
rect 8115 670 8120 750
rect 8080 660 8120 670
rect 8400 750 8440 765
rect 9040 795 9080 800
rect 9040 765 9045 795
rect 9075 765 9080 795
rect 8400 670 8405 750
rect 8435 670 8440 750
rect 8400 660 8440 670
rect 8720 750 8760 760
rect 8720 670 8725 750
rect 8755 670 8760 750
rect 8720 660 8760 670
rect 9040 750 9080 765
rect 9680 795 9720 800
rect 9680 765 9685 795
rect 9715 765 9720 795
rect 9040 670 9045 750
rect 9075 670 9080 750
rect 9040 660 9080 670
rect 9360 750 9400 760
rect 9360 670 9365 750
rect 9395 670 9400 750
rect 9360 660 9400 670
rect 9680 750 9720 765
rect 10320 795 10360 800
rect 10320 765 10325 795
rect 10355 765 10360 795
rect 9680 670 9685 750
rect 9715 670 9720 750
rect 9680 660 9720 670
rect 10000 750 10040 760
rect 10000 670 10005 750
rect 10035 670 10040 750
rect 10000 660 10040 670
rect 10320 750 10360 765
rect 10640 795 10680 800
rect 10640 765 10645 795
rect 10675 765 10680 795
rect 10640 760 10680 765
rect 10800 795 10840 800
rect 10800 765 10805 795
rect 10835 765 10840 795
rect 10800 760 10840 765
rect 10960 795 11000 800
rect 10960 765 10965 795
rect 10995 765 11000 795
rect 10960 760 11000 765
rect 10320 670 10325 750
rect 10355 670 10360 750
rect 10640 715 10680 720
rect 10640 685 10645 715
rect 10675 685 10680 715
rect 10640 680 10680 685
rect 10800 715 10840 720
rect 10800 685 10805 715
rect 10835 685 10840 715
rect 10800 680 10840 685
rect 10960 715 11000 720
rect 10960 685 10965 715
rect 10995 685 11000 715
rect 10960 680 11000 685
rect 10320 660 10360 670
rect 5600 635 5800 640
rect 5600 605 5610 635
rect 5790 605 5800 635
rect 5600 600 5800 605
rect 5920 635 6120 640
rect 5920 605 5930 635
rect 6110 605 6120 635
rect 5920 600 6120 605
rect 6240 635 6440 640
rect 6240 605 6250 635
rect 6430 605 6440 635
rect 6240 600 6440 605
rect 6560 635 6760 640
rect 6560 605 6570 635
rect 6750 605 6760 635
rect 6560 600 6760 605
rect 6880 635 7080 640
rect 6880 605 6890 635
rect 7070 605 7080 635
rect 6880 600 7080 605
rect 7200 635 7400 640
rect 7200 605 7210 635
rect 7390 605 7400 635
rect 7200 600 7400 605
rect 7520 635 7720 640
rect 7520 605 7530 635
rect 7710 605 7720 635
rect 7520 600 7720 605
rect 7840 635 8040 640
rect 7840 605 7850 635
rect 8030 605 8040 635
rect 7840 600 8040 605
rect 8160 635 8360 640
rect 8160 605 8170 635
rect 8350 605 8360 635
rect 8160 600 8360 605
rect 8480 635 8680 640
rect 8480 605 8490 635
rect 8670 605 8680 635
rect 8480 600 8680 605
rect 8800 635 9000 640
rect 8800 605 8810 635
rect 8990 605 9000 635
rect 8800 600 9000 605
rect 9120 635 9320 640
rect 9120 605 9130 635
rect 9310 605 9320 635
rect 9120 600 9320 605
rect 9440 635 9640 640
rect 9440 605 9450 635
rect 9630 605 9640 635
rect 9440 600 9640 605
rect 9760 635 9960 640
rect 9760 605 9770 635
rect 9950 605 9960 635
rect 9760 600 9960 605
rect 10080 635 10280 640
rect 10080 605 10090 635
rect 10270 605 10280 635
rect 10080 600 10280 605
rect 10640 635 10680 640
rect 10640 605 10645 635
rect 10675 605 10680 635
rect 10640 600 10680 605
rect 10800 635 10840 640
rect 10800 605 10805 635
rect 10835 605 10840 635
rect 10800 600 10840 605
rect 10960 635 11000 640
rect 10960 605 10965 635
rect 10995 605 11000 635
rect 10960 600 11000 605
rect 5520 285 5525 315
rect 5555 285 5560 315
rect 5520 280 5560 285
rect 5680 315 5720 600
rect 5680 285 5685 315
rect 5715 285 5720 315
rect 5680 280 5720 285
rect 6000 315 6040 600
rect 6000 285 6005 315
rect 6035 285 6040 315
rect 6000 280 6040 285
rect 6160 315 6200 600
rect 6160 285 6165 315
rect 6195 285 6200 315
rect 6160 280 6200 285
rect 6320 315 6360 600
rect 6320 285 6325 315
rect 6355 285 6360 315
rect 6320 280 6360 285
rect 6480 315 6520 320
rect 6480 285 6485 315
rect 6515 285 6520 315
rect 5040 125 5045 155
rect 5075 125 5080 155
rect 5040 120 5080 125
rect 5280 155 5480 160
rect 5280 125 5290 155
rect 5470 125 5480 155
rect 5280 120 5480 125
rect 5600 155 5800 160
rect 5600 125 5610 155
rect 5790 125 5800 155
rect 5600 120 5800 125
rect 5920 155 6120 160
rect 5920 125 5930 155
rect 6110 125 6120 155
rect 5920 120 6120 125
rect 6240 155 6440 160
rect 6240 125 6250 155
rect 6430 125 6440 155
rect 6240 120 6440 125
rect 3760 10 3765 90
rect 3795 10 3800 90
rect 3760 0 3800 10
rect 4080 90 4120 100
rect 4080 10 4085 90
rect 4115 10 4120 90
rect 4080 0 4120 10
rect 4400 90 4440 100
rect 4400 10 4405 90
rect 4435 10 4440 90
rect 4400 0 4440 10
rect 4720 90 4760 100
rect 4720 10 4725 90
rect 4755 10 4760 90
rect 4720 0 4760 10
rect 5040 90 5080 100
rect 5040 10 5045 90
rect 5075 10 5080 90
rect 2480 -35 2485 -5
rect 2515 -35 2520 -5
rect 2480 -40 2520 -35
rect 5040 -5 5080 10
rect 5040 -35 5045 -5
rect 5075 -35 5080 -5
rect 5040 -40 5080 -35
rect 5200 90 5240 100
rect 5200 10 5205 90
rect 5235 10 5240 90
rect 5200 -5 5240 10
rect 5520 90 5560 100
rect 5520 10 5525 90
rect 5555 10 5560 90
rect 5520 0 5560 10
rect 5840 90 5880 100
rect 5840 10 5845 90
rect 5875 10 5880 90
rect 5840 0 5880 10
rect 6160 90 6200 100
rect 6160 10 6165 90
rect 6195 10 6200 90
rect 6160 0 6200 10
rect 6480 90 6520 285
rect 6640 315 6680 600
rect 6640 285 6645 315
rect 6675 285 6680 315
rect 6640 280 6680 285
rect 6800 315 6840 600
rect 6800 285 6805 315
rect 6835 285 6840 315
rect 6800 280 6840 285
rect 6960 315 7000 600
rect 6960 285 6965 315
rect 6995 285 7000 315
rect 6960 280 7000 285
rect 7280 315 7320 600
rect 7280 285 7285 315
rect 7315 285 7320 315
rect 7280 280 7320 285
rect 7440 315 7480 600
rect 7440 285 7445 315
rect 7475 285 7480 315
rect 7440 280 7480 285
rect 7600 315 7640 600
rect 7600 285 7605 315
rect 7635 285 7640 315
rect 7600 280 7640 285
rect 7920 315 7960 600
rect 7920 285 7925 315
rect 7955 285 7960 315
rect 7920 280 7960 285
rect 8080 315 8120 600
rect 8080 285 8085 315
rect 8115 285 8120 315
rect 8080 280 8120 285
rect 8240 315 8280 600
rect 8240 285 8245 315
rect 8275 285 8280 315
rect 8240 280 8280 285
rect 8560 315 8600 600
rect 8560 285 8565 315
rect 8595 285 8600 315
rect 8560 280 8600 285
rect 8720 315 8760 600
rect 8720 285 8725 315
rect 8755 285 8760 315
rect 8720 280 8760 285
rect 8880 315 8920 600
rect 8880 285 8885 315
rect 8915 285 8920 315
rect 8880 280 8920 285
rect 9040 315 9080 320
rect 9040 285 9045 315
rect 9075 285 9080 315
rect 6560 155 6760 160
rect 6560 125 6570 155
rect 6750 125 6760 155
rect 6560 120 6760 125
rect 6880 155 7080 160
rect 6880 125 6890 155
rect 7070 125 7080 155
rect 6880 120 7080 125
rect 7200 155 7400 160
rect 7200 125 7210 155
rect 7390 125 7400 155
rect 7200 120 7400 125
rect 7520 155 7720 160
rect 7520 125 7530 155
rect 7710 125 7720 155
rect 7520 120 7720 125
rect 7840 155 8040 160
rect 7840 125 7850 155
rect 8030 125 8040 155
rect 7840 120 8040 125
rect 8160 155 8360 160
rect 8160 125 8170 155
rect 8350 125 8360 155
rect 8160 120 8360 125
rect 8480 155 8680 160
rect 8480 125 8490 155
rect 8670 125 8680 155
rect 8480 120 8680 125
rect 8800 155 9000 160
rect 8800 125 8810 155
rect 8990 125 9000 155
rect 8800 120 9000 125
rect 6480 10 6485 90
rect 6515 10 6520 90
rect 6480 0 6520 10
rect 6800 90 6840 100
rect 6800 10 6805 90
rect 6835 10 6840 90
rect 6800 0 6840 10
rect 7120 90 7160 100
rect 7120 10 7125 90
rect 7155 10 7160 90
rect 7120 0 7160 10
rect 7440 90 7480 100
rect 7440 10 7445 90
rect 7475 10 7480 90
rect 7440 0 7480 10
rect 7760 90 7800 100
rect 7760 10 7765 90
rect 7795 10 7800 90
rect 5200 -35 5205 -5
rect 5235 -35 5240 -5
rect 5200 -40 5240 -35
rect 7760 -5 7800 10
rect 8080 90 8120 100
rect 8080 10 8085 90
rect 8115 10 8120 90
rect 8080 0 8120 10
rect 8400 90 8440 100
rect 8400 10 8405 90
rect 8435 10 8440 90
rect 8400 0 8440 10
rect 8720 90 8760 100
rect 8720 10 8725 90
rect 8755 10 8760 90
rect 8720 0 8760 10
rect 9040 90 9080 285
rect 9200 315 9240 600
rect 9200 285 9205 315
rect 9235 285 9240 315
rect 9200 280 9240 285
rect 9360 315 9400 600
rect 9360 285 9365 315
rect 9395 285 9400 315
rect 9360 280 9400 285
rect 9520 315 9560 600
rect 9520 285 9525 315
rect 9555 285 9560 315
rect 9520 280 9560 285
rect 9840 315 9880 600
rect 9840 285 9845 315
rect 9875 285 9880 315
rect 9840 280 9880 285
rect 10000 315 10040 600
rect 10000 285 10005 315
rect 10035 285 10040 315
rect 10000 280 10040 285
rect 10160 315 10200 600
rect 10640 555 10680 560
rect 10640 525 10645 555
rect 10675 525 10680 555
rect 10640 520 10680 525
rect 10800 555 10840 560
rect 10800 525 10805 555
rect 10835 525 10840 555
rect 10800 520 10840 525
rect 10960 555 11000 560
rect 10960 525 10965 555
rect 10995 525 11000 555
rect 10960 520 11000 525
rect 10640 475 10680 480
rect 10640 445 10645 475
rect 10675 445 10680 475
rect 10640 440 10680 445
rect 10800 475 10840 480
rect 10800 445 10805 475
rect 10835 445 10840 475
rect 10800 440 10840 445
rect 10960 475 11000 480
rect 10960 445 10965 475
rect 10995 445 11000 475
rect 10960 440 11000 445
rect 10640 395 10680 400
rect 10640 365 10645 395
rect 10675 365 10680 395
rect 10640 360 10680 365
rect 10800 395 10840 400
rect 10800 365 10805 395
rect 10835 365 10840 395
rect 10800 360 10840 365
rect 10960 395 11000 400
rect 10960 365 10965 395
rect 10995 365 11000 395
rect 10960 360 11000 365
rect 10160 285 10165 315
rect 10195 285 10200 315
rect 10160 280 10200 285
rect 10640 235 10680 240
rect 10640 205 10645 235
rect 10675 205 10680 235
rect 10640 200 10680 205
rect 10800 235 10840 240
rect 10800 205 10805 235
rect 10835 205 10840 235
rect 10800 200 10840 205
rect 10960 235 11000 240
rect 10960 205 10965 235
rect 10995 205 11000 235
rect 10960 200 11000 205
rect 9120 155 9320 160
rect 9120 125 9130 155
rect 9310 125 9320 155
rect 9120 120 9320 125
rect 9440 155 9640 160
rect 9440 125 9450 155
rect 9630 125 9640 155
rect 9440 120 9640 125
rect 9760 155 9960 160
rect 9760 125 9770 155
rect 9950 125 9960 155
rect 9760 120 9960 125
rect 10080 155 10280 160
rect 10080 125 10090 155
rect 10270 125 10280 155
rect 10080 120 10280 125
rect 10800 155 10840 160
rect 10800 125 10805 155
rect 10835 125 10840 155
rect 10800 120 10840 125
rect 10960 155 11000 160
rect 10960 125 10965 155
rect 10995 125 11000 155
rect 10960 120 11000 125
rect 9040 10 9045 90
rect 9075 10 9080 90
rect 9040 0 9080 10
rect 9360 90 9400 100
rect 9360 10 9365 90
rect 9395 10 9400 90
rect 9360 0 9400 10
rect 9680 90 9720 100
rect 9680 10 9685 90
rect 9715 10 9720 90
rect 9680 0 9720 10
rect 10000 90 10040 100
rect 10000 10 10005 90
rect 10035 10 10040 90
rect 10000 0 10040 10
rect 10320 90 10360 100
rect 10320 10 10325 90
rect 10355 10 10360 90
rect 10640 75 10680 80
rect 10640 45 10645 75
rect 10675 45 10680 75
rect 10640 40 10680 45
rect 10800 75 10840 80
rect 10800 45 10805 75
rect 10835 45 10840 75
rect 10800 40 10840 45
rect 10960 75 11000 80
rect 10960 45 10965 75
rect 10995 45 11000 75
rect 10960 40 11000 45
rect 7760 -35 7765 -5
rect 7795 -35 7800 -5
rect 7760 -40 7800 -35
rect 10320 -5 10360 10
rect 10320 -35 10325 -5
rect 10355 -35 10360 -5
rect 10320 -40 10360 -35
rect 10640 -5 10680 0
rect 10640 -35 10645 -5
rect 10675 -35 10680 -5
rect 10640 -40 10680 -35
rect 10800 -5 10840 0
rect 10800 -35 10805 -5
rect 10835 -35 10840 -5
rect 10800 -40 10840 -35
rect 10960 -5 11000 0
rect 10960 -35 10965 -5
rect 10995 -35 11000 -5
rect 10960 -40 11000 -35
rect -720 -85 -680 -80
rect -720 -115 -715 -85
rect -685 -115 -680 -85
rect -720 -120 -680 -115
rect -560 -85 -520 -80
rect -560 -115 -555 -85
rect -525 -115 -520 -85
rect -560 -120 -520 -115
rect -400 -85 -360 -80
rect -400 -115 -395 -85
rect -365 -115 -360 -85
rect -400 -120 -360 -115
rect 10640 -85 10680 -80
rect 10640 -115 10645 -85
rect 10675 -115 10680 -85
rect 10640 -120 10680 -115
rect 10800 -85 10840 -80
rect 10800 -115 10805 -85
rect 10835 -115 10840 -85
rect 10800 -120 10840 -115
rect 10960 -85 11000 -80
rect 10960 -115 10965 -85
rect 10995 -115 11000 -85
rect 10960 -120 11000 -115
<< via1 >>
rect -715 1005 -685 1035
rect -555 1005 -525 1035
rect -395 1005 -365 1035
rect 10645 1005 10675 1035
rect 10805 1005 10835 1035
rect 10965 1005 10995 1035
rect -715 925 -685 955
rect -555 925 -525 955
rect -395 925 -365 955
rect 10645 925 10675 955
rect 10805 925 10835 955
rect 10965 925 10995 955
rect -715 845 -685 875
rect -555 845 -525 875
rect -395 845 -365 875
rect 10645 845 10675 875
rect 10805 845 10835 875
rect 10965 845 10995 875
rect -75 765 -45 795
rect 5205 765 5235 795
rect -75 685 -45 715
rect -715 605 -685 635
rect -555 605 -525 635
rect -395 605 -365 635
rect -715 525 -685 555
rect -555 525 -525 555
rect -395 525 -365 555
rect -715 445 -685 475
rect -555 445 -525 475
rect 85 445 115 475
rect 405 445 435 475
rect 725 445 755 475
rect 1045 445 1075 475
rect 1365 445 1395 475
rect 1685 445 1715 475
rect 2005 445 2035 475
rect 2325 445 2355 475
rect 2645 445 2675 475
rect 2965 445 2995 475
rect 3285 445 3315 475
rect 3605 445 3635 475
rect 3925 445 3955 475
rect 4245 445 4275 475
rect 4565 445 4595 475
rect 4885 445 4915 475
rect -715 365 -685 395
rect -555 365 -525 395
rect -395 365 -365 395
rect -715 285 -685 315
rect -555 285 -525 315
rect -395 285 -365 315
rect -715 205 -685 235
rect -555 205 -525 235
rect -395 205 -365 235
rect -715 125 -685 155
rect -555 125 -525 155
rect -395 125 -365 155
rect 10 125 190 155
rect 330 125 510 155
rect 650 125 830 155
rect 970 125 1150 155
rect 1205 125 1235 155
rect -715 45 -685 75
rect -555 45 -525 75
rect -395 45 -365 75
rect -75 45 -45 75
rect -715 -35 -685 -5
rect -555 -35 -525 -5
rect -395 -35 -365 -5
rect 1290 125 1470 155
rect 1610 125 1790 155
rect 1930 125 2110 155
rect 2250 125 2430 155
rect 2570 125 2750 155
rect 2890 125 3070 155
rect 3210 125 3390 155
rect 3530 125 3710 155
rect 3765 125 3795 155
rect 2485 45 2515 75
rect -75 -35 -45 -5
rect 3850 125 4030 155
rect 4170 125 4350 155
rect 4490 125 4670 155
rect 4810 125 4990 155
rect 5845 765 5875 795
rect 5205 685 5235 715
rect 5365 285 5395 315
rect 6485 765 6515 795
rect 5845 685 5875 715
rect 7125 765 7155 795
rect 6485 685 6515 715
rect 7765 765 7795 795
rect 7125 685 7155 715
rect 8405 765 8435 795
rect 7765 685 7795 715
rect 9045 765 9075 795
rect 8405 685 8435 715
rect 9685 765 9715 795
rect 9045 685 9075 715
rect 10325 765 10355 795
rect 9685 685 9715 715
rect 10645 765 10675 795
rect 10805 765 10835 795
rect 10965 765 10995 795
rect 10325 685 10355 715
rect 10645 685 10675 715
rect 10805 685 10835 715
rect 10965 685 10995 715
rect 10645 605 10675 635
rect 10805 605 10835 635
rect 10965 605 10995 635
rect 5525 285 5555 315
rect 5685 285 5715 315
rect 6005 285 6035 315
rect 6165 285 6195 315
rect 6325 285 6355 315
rect 6485 285 6515 315
rect 5045 125 5075 155
rect 5290 125 5470 155
rect 5610 125 5790 155
rect 5930 125 6110 155
rect 6250 125 6430 155
rect 5045 45 5075 75
rect 2485 -35 2515 -5
rect 5045 -35 5075 -5
rect 5205 45 5235 75
rect 6645 285 6675 315
rect 6805 285 6835 315
rect 6965 285 6995 315
rect 7285 285 7315 315
rect 7445 285 7475 315
rect 7605 285 7635 315
rect 7925 285 7955 315
rect 8085 285 8115 315
rect 8245 285 8275 315
rect 8565 285 8595 315
rect 8725 285 8755 315
rect 8885 285 8915 315
rect 9045 285 9075 315
rect 6570 125 6750 155
rect 6890 125 7070 155
rect 7210 125 7390 155
rect 7530 125 7710 155
rect 7850 125 8030 155
rect 8170 125 8350 155
rect 8490 125 8670 155
rect 8810 125 8990 155
rect 7765 45 7795 75
rect 5205 -35 5235 -5
rect 9205 285 9235 315
rect 9365 285 9395 315
rect 9525 285 9555 315
rect 9845 285 9875 315
rect 10005 285 10035 315
rect 10645 525 10675 555
rect 10805 525 10835 555
rect 10965 525 10995 555
rect 10645 445 10675 475
rect 10805 445 10835 475
rect 10965 445 10995 475
rect 10645 365 10675 395
rect 10805 365 10835 395
rect 10965 365 10995 395
rect 10165 285 10195 315
rect 10645 205 10675 235
rect 10805 205 10835 235
rect 10965 205 10995 235
rect 9130 125 9310 155
rect 9450 125 9630 155
rect 9770 125 9950 155
rect 10090 125 10270 155
rect 10805 125 10835 155
rect 10965 125 10995 155
rect 10325 45 10355 75
rect 10645 45 10675 75
rect 10805 45 10835 75
rect 10965 45 10995 75
rect 7765 -35 7795 -5
rect 10325 -35 10355 -5
rect 10645 -35 10675 -5
rect 10805 -35 10835 -5
rect 10965 -35 10995 -5
rect -715 -115 -685 -85
rect -555 -115 -525 -85
rect -395 -115 -365 -85
rect 10645 -115 10675 -85
rect 10805 -115 10835 -85
rect 10965 -115 10995 -85
<< metal2 >>
rect -720 1035 11000 1040
rect -720 1005 -715 1035
rect -685 1005 -555 1035
rect -525 1005 -395 1035
rect -365 1005 -315 1035
rect -285 1005 -235 1035
rect -205 1005 -155 1035
rect -125 1005 -75 1035
rect -45 1005 5 1035
rect 35 1005 85 1035
rect 115 1005 165 1035
rect 195 1005 245 1035
rect 275 1005 325 1035
rect 355 1005 405 1035
rect 435 1005 485 1035
rect 515 1005 565 1035
rect 595 1005 645 1035
rect 675 1005 725 1035
rect 755 1005 805 1035
rect 835 1005 885 1035
rect 915 1005 965 1035
rect 995 1005 1045 1035
rect 1075 1005 1125 1035
rect 1155 1005 1205 1035
rect 1235 1005 1285 1035
rect 1315 1005 1365 1035
rect 1395 1005 1445 1035
rect 1475 1005 1525 1035
rect 1555 1005 1605 1035
rect 1635 1005 1685 1035
rect 1715 1005 1765 1035
rect 1795 1005 1845 1035
rect 1875 1005 1925 1035
rect 1955 1005 2005 1035
rect 2035 1005 2085 1035
rect 2115 1005 2165 1035
rect 2195 1005 2245 1035
rect 2275 1005 2325 1035
rect 2355 1005 2405 1035
rect 2435 1005 2485 1035
rect 2515 1005 2565 1035
rect 2595 1005 2645 1035
rect 2675 1005 2725 1035
rect 2755 1005 2805 1035
rect 2835 1005 2885 1035
rect 2915 1005 2965 1035
rect 2995 1005 3045 1035
rect 3075 1005 3125 1035
rect 3155 1005 3205 1035
rect 3235 1005 3285 1035
rect 3315 1005 3365 1035
rect 3395 1005 3445 1035
rect 3475 1005 3525 1035
rect 3555 1005 3605 1035
rect 3635 1005 3685 1035
rect 3715 1005 3765 1035
rect 3795 1005 3845 1035
rect 3875 1005 3925 1035
rect 3955 1005 4005 1035
rect 4035 1005 4085 1035
rect 4115 1005 4165 1035
rect 4195 1005 4245 1035
rect 4275 1005 4325 1035
rect 4355 1005 4405 1035
rect 4435 1005 4485 1035
rect 4515 1005 4565 1035
rect 4595 1005 4645 1035
rect 4675 1005 4725 1035
rect 4755 1005 4805 1035
rect 4835 1005 4885 1035
rect 4915 1005 4965 1035
rect 4995 1005 5045 1035
rect 5075 1005 5125 1035
rect 5155 1005 5205 1035
rect 5235 1005 5285 1035
rect 5315 1005 5365 1035
rect 5395 1005 5445 1035
rect 5475 1005 5525 1035
rect 5555 1005 5605 1035
rect 5635 1005 5685 1035
rect 5715 1005 5765 1035
rect 5795 1005 5845 1035
rect 5875 1005 5925 1035
rect 5955 1005 6005 1035
rect 6035 1005 6085 1035
rect 6115 1005 6165 1035
rect 6195 1005 6245 1035
rect 6275 1005 6325 1035
rect 6355 1005 6405 1035
rect 6435 1005 6485 1035
rect 6515 1005 6565 1035
rect 6595 1005 6645 1035
rect 6675 1005 6725 1035
rect 6755 1005 6805 1035
rect 6835 1005 6885 1035
rect 6915 1005 6965 1035
rect 6995 1005 7045 1035
rect 7075 1005 7125 1035
rect 7155 1005 7205 1035
rect 7235 1005 7285 1035
rect 7315 1005 7365 1035
rect 7395 1005 7445 1035
rect 7475 1005 7525 1035
rect 7555 1005 7605 1035
rect 7635 1005 7685 1035
rect 7715 1005 7765 1035
rect 7795 1005 7845 1035
rect 7875 1005 7925 1035
rect 7955 1005 8005 1035
rect 8035 1005 8085 1035
rect 8115 1005 8165 1035
rect 8195 1005 8245 1035
rect 8275 1005 8325 1035
rect 8355 1005 8405 1035
rect 8435 1005 8485 1035
rect 8515 1005 8565 1035
rect 8595 1005 8645 1035
rect 8675 1005 8725 1035
rect 8755 1005 8805 1035
rect 8835 1005 8885 1035
rect 8915 1005 8965 1035
rect 8995 1005 9045 1035
rect 9075 1005 9125 1035
rect 9155 1005 9205 1035
rect 9235 1005 9285 1035
rect 9315 1005 9365 1035
rect 9395 1005 9445 1035
rect 9475 1005 9525 1035
rect 9555 1005 9605 1035
rect 9635 1005 9685 1035
rect 9715 1005 9765 1035
rect 9795 1005 9845 1035
rect 9875 1005 9925 1035
rect 9955 1005 10005 1035
rect 10035 1005 10085 1035
rect 10115 1005 10165 1035
rect 10195 1005 10245 1035
rect 10275 1005 10325 1035
rect 10355 1005 10405 1035
rect 10435 1005 10485 1035
rect 10515 1005 10645 1035
rect 10675 1005 10805 1035
rect 10835 1005 10965 1035
rect 10995 1005 11000 1035
rect -720 1000 11000 1005
rect -720 955 11000 960
rect -720 925 -715 955
rect -685 925 -555 955
rect -525 925 -395 955
rect -365 925 -315 955
rect -285 925 -235 955
rect -205 925 -155 955
rect -125 925 -75 955
rect -45 925 5 955
rect 35 925 85 955
rect 115 925 165 955
rect 195 925 245 955
rect 275 925 325 955
rect 355 925 405 955
rect 435 925 485 955
rect 515 925 565 955
rect 595 925 645 955
rect 675 925 725 955
rect 755 925 805 955
rect 835 925 885 955
rect 915 925 965 955
rect 995 925 1045 955
rect 1075 925 1125 955
rect 1155 925 1205 955
rect 1235 925 1285 955
rect 1315 925 1365 955
rect 1395 925 1445 955
rect 1475 925 1525 955
rect 1555 925 1605 955
rect 1635 925 1685 955
rect 1715 925 1765 955
rect 1795 925 1845 955
rect 1875 925 1925 955
rect 1955 925 2005 955
rect 2035 925 2085 955
rect 2115 925 2165 955
rect 2195 925 2245 955
rect 2275 925 2325 955
rect 2355 925 2405 955
rect 2435 925 2485 955
rect 2515 925 2565 955
rect 2595 925 2645 955
rect 2675 925 2725 955
rect 2755 925 2805 955
rect 2835 925 2885 955
rect 2915 925 2965 955
rect 2995 925 3045 955
rect 3075 925 3125 955
rect 3155 925 3205 955
rect 3235 925 3285 955
rect 3315 925 3365 955
rect 3395 925 3445 955
rect 3475 925 3525 955
rect 3555 925 3605 955
rect 3635 925 3685 955
rect 3715 925 3765 955
rect 3795 925 3845 955
rect 3875 925 3925 955
rect 3955 925 4005 955
rect 4035 925 4085 955
rect 4115 925 4165 955
rect 4195 925 4245 955
rect 4275 925 4325 955
rect 4355 925 4405 955
rect 4435 925 4485 955
rect 4515 925 4565 955
rect 4595 925 4645 955
rect 4675 925 4725 955
rect 4755 925 4805 955
rect 4835 925 4885 955
rect 4915 925 4965 955
rect 4995 925 5045 955
rect 5075 925 5125 955
rect 5155 925 5205 955
rect 5235 925 5285 955
rect 5315 925 5365 955
rect 5395 925 5445 955
rect 5475 925 5525 955
rect 5555 925 5605 955
rect 5635 925 5685 955
rect 5715 925 5765 955
rect 5795 925 5845 955
rect 5875 925 5925 955
rect 5955 925 6005 955
rect 6035 925 6085 955
rect 6115 925 6165 955
rect 6195 925 6245 955
rect 6275 925 6325 955
rect 6355 925 6405 955
rect 6435 925 6485 955
rect 6515 925 6565 955
rect 6595 925 6645 955
rect 6675 925 6725 955
rect 6755 925 6805 955
rect 6835 925 6885 955
rect 6915 925 6965 955
rect 6995 925 7045 955
rect 7075 925 7125 955
rect 7155 925 7205 955
rect 7235 925 7285 955
rect 7315 925 7365 955
rect 7395 925 7445 955
rect 7475 925 7525 955
rect 7555 925 7605 955
rect 7635 925 7685 955
rect 7715 925 7765 955
rect 7795 925 7845 955
rect 7875 925 7925 955
rect 7955 925 8005 955
rect 8035 925 8085 955
rect 8115 925 8165 955
rect 8195 925 8245 955
rect 8275 925 8325 955
rect 8355 925 8405 955
rect 8435 925 8485 955
rect 8515 925 8565 955
rect 8595 925 8645 955
rect 8675 925 8725 955
rect 8755 925 8805 955
rect 8835 925 8885 955
rect 8915 925 8965 955
rect 8995 925 9045 955
rect 9075 925 9125 955
rect 9155 925 9205 955
rect 9235 925 9285 955
rect 9315 925 9365 955
rect 9395 925 9445 955
rect 9475 925 9525 955
rect 9555 925 9605 955
rect 9635 925 9685 955
rect 9715 925 9765 955
rect 9795 925 9845 955
rect 9875 925 9925 955
rect 9955 925 10005 955
rect 10035 925 10085 955
rect 10115 925 10165 955
rect 10195 925 10245 955
rect 10275 925 10325 955
rect 10355 925 10405 955
rect 10435 925 10485 955
rect 10515 925 10645 955
rect 10675 925 10805 955
rect 10835 925 10965 955
rect 10995 925 11000 955
rect -720 920 11000 925
rect -720 875 11000 880
rect -720 845 -715 875
rect -685 845 -555 875
rect -525 845 -395 875
rect -365 845 -315 875
rect -285 845 -235 875
rect -205 845 -155 875
rect -125 845 -75 875
rect -45 845 5 875
rect 35 845 85 875
rect 115 845 165 875
rect 195 845 245 875
rect 275 845 325 875
rect 355 845 405 875
rect 435 845 485 875
rect 515 845 565 875
rect 595 845 645 875
rect 675 845 725 875
rect 755 845 805 875
rect 835 845 885 875
rect 915 845 965 875
rect 995 845 1045 875
rect 1075 845 1125 875
rect 1155 845 1205 875
rect 1235 845 1285 875
rect 1315 845 1365 875
rect 1395 845 1445 875
rect 1475 845 1525 875
rect 1555 845 1605 875
rect 1635 845 1685 875
rect 1715 845 1765 875
rect 1795 845 1845 875
rect 1875 845 1925 875
rect 1955 845 2005 875
rect 2035 845 2085 875
rect 2115 845 2165 875
rect 2195 845 2245 875
rect 2275 845 2325 875
rect 2355 845 2405 875
rect 2435 845 2485 875
rect 2515 845 2565 875
rect 2595 845 2645 875
rect 2675 845 2725 875
rect 2755 845 2805 875
rect 2835 845 2885 875
rect 2915 845 2965 875
rect 2995 845 3045 875
rect 3075 845 3125 875
rect 3155 845 3205 875
rect 3235 845 3285 875
rect 3315 845 3365 875
rect 3395 845 3445 875
rect 3475 845 3525 875
rect 3555 845 3605 875
rect 3635 845 3685 875
rect 3715 845 3765 875
rect 3795 845 3845 875
rect 3875 845 3925 875
rect 3955 845 4005 875
rect 4035 845 4085 875
rect 4115 845 4165 875
rect 4195 845 4245 875
rect 4275 845 4325 875
rect 4355 845 4405 875
rect 4435 845 4485 875
rect 4515 845 4565 875
rect 4595 845 4645 875
rect 4675 845 4725 875
rect 4755 845 4805 875
rect 4835 845 4885 875
rect 4915 845 4965 875
rect 4995 845 5045 875
rect 5075 845 5125 875
rect 5155 845 5205 875
rect 5235 845 5285 875
rect 5315 845 5365 875
rect 5395 845 5445 875
rect 5475 845 5525 875
rect 5555 845 5605 875
rect 5635 845 5685 875
rect 5715 845 5765 875
rect 5795 845 5845 875
rect 5875 845 5925 875
rect 5955 845 6005 875
rect 6035 845 6085 875
rect 6115 845 6165 875
rect 6195 845 6245 875
rect 6275 845 6325 875
rect 6355 845 6405 875
rect 6435 845 6485 875
rect 6515 845 6565 875
rect 6595 845 6645 875
rect 6675 845 6725 875
rect 6755 845 6805 875
rect 6835 845 6885 875
rect 6915 845 6965 875
rect 6995 845 7045 875
rect 7075 845 7125 875
rect 7155 845 7205 875
rect 7235 845 7285 875
rect 7315 845 7365 875
rect 7395 845 7445 875
rect 7475 845 7525 875
rect 7555 845 7605 875
rect 7635 845 7685 875
rect 7715 845 7765 875
rect 7795 845 7845 875
rect 7875 845 7925 875
rect 7955 845 8005 875
rect 8035 845 8085 875
rect 8115 845 8165 875
rect 8195 845 8245 875
rect 8275 845 8325 875
rect 8355 845 8405 875
rect 8435 845 8485 875
rect 8515 845 8565 875
rect 8595 845 8645 875
rect 8675 845 8725 875
rect 8755 845 8805 875
rect 8835 845 8885 875
rect 8915 845 8965 875
rect 8995 845 9045 875
rect 9075 845 9125 875
rect 9155 845 9205 875
rect 9235 845 9285 875
rect 9315 845 9365 875
rect 9395 845 9445 875
rect 9475 845 9525 875
rect 9555 845 9605 875
rect 9635 845 9685 875
rect 9715 845 9765 875
rect 9795 845 9845 875
rect 9875 845 9925 875
rect 9955 845 10005 875
rect 10035 845 10085 875
rect 10115 845 10165 875
rect 10195 845 10245 875
rect 10275 845 10325 875
rect 10355 845 10405 875
rect 10435 845 10485 875
rect 10515 845 10645 875
rect 10675 845 10805 875
rect 10835 845 10965 875
rect 10995 845 11000 875
rect -720 840 11000 845
rect -640 795 10600 800
rect -640 765 -635 795
rect -605 765 -75 795
rect -45 765 5205 795
rect 5235 765 5845 795
rect 5875 765 6485 795
rect 6515 765 7125 795
rect 7155 765 7765 795
rect 7795 765 8405 795
rect 8435 765 9045 795
rect 9075 765 9685 795
rect 9715 765 10325 795
rect 10355 765 10600 795
rect -640 760 10600 765
rect 10640 795 11000 800
rect 10640 765 10645 795
rect 10675 765 10805 795
rect 10835 765 10965 795
rect 10995 765 11000 795
rect 10640 760 11000 765
rect -640 715 10600 720
rect -640 685 -635 715
rect -605 685 -75 715
rect -45 685 5205 715
rect 5235 685 5845 715
rect 5875 685 6485 715
rect 6515 685 7125 715
rect 7155 685 7765 715
rect 7795 685 8405 715
rect 8435 685 9045 715
rect 9075 685 9685 715
rect 9715 685 10325 715
rect 10355 685 10600 715
rect -640 680 10600 685
rect 10640 715 11000 720
rect 10640 685 10645 715
rect 10675 685 10805 715
rect 10835 685 10965 715
rect 10995 685 11000 715
rect 10640 680 11000 685
rect -720 635 11000 640
rect -720 605 -715 635
rect -685 605 -555 635
rect -525 605 -395 635
rect -365 605 -315 635
rect -285 605 -235 635
rect -205 605 -155 635
rect -125 605 -75 635
rect -45 605 5 635
rect 35 605 85 635
rect 115 605 165 635
rect 195 605 245 635
rect 275 605 325 635
rect 355 605 405 635
rect 435 605 485 635
rect 515 605 565 635
rect 595 605 645 635
rect 675 605 725 635
rect 755 605 805 635
rect 835 605 885 635
rect 915 605 965 635
rect 995 605 1045 635
rect 1075 605 1125 635
rect 1155 605 1205 635
rect 1235 605 1285 635
rect 1315 605 1365 635
rect 1395 605 1445 635
rect 1475 605 1525 635
rect 1555 605 1605 635
rect 1635 605 1685 635
rect 1715 605 1765 635
rect 1795 605 1845 635
rect 1875 605 1925 635
rect 1955 605 2005 635
rect 2035 605 2085 635
rect 2115 605 2165 635
rect 2195 605 2245 635
rect 2275 605 2325 635
rect 2355 605 2405 635
rect 2435 605 2485 635
rect 2515 605 2565 635
rect 2595 605 2645 635
rect 2675 605 2725 635
rect 2755 605 2805 635
rect 2835 605 2885 635
rect 2915 605 2965 635
rect 2995 605 3045 635
rect 3075 605 3125 635
rect 3155 605 3205 635
rect 3235 605 3285 635
rect 3315 605 3365 635
rect 3395 605 3445 635
rect 3475 605 3525 635
rect 3555 605 3605 635
rect 3635 605 3685 635
rect 3715 605 3765 635
rect 3795 605 3845 635
rect 3875 605 3925 635
rect 3955 605 4005 635
rect 4035 605 4085 635
rect 4115 605 4165 635
rect 4195 605 4245 635
rect 4275 605 4325 635
rect 4355 605 4405 635
rect 4435 605 4485 635
rect 4515 605 4565 635
rect 4595 605 4645 635
rect 4675 605 4725 635
rect 4755 605 4805 635
rect 4835 605 4885 635
rect 4915 605 4965 635
rect 4995 605 5045 635
rect 5075 605 5125 635
rect 5155 605 5205 635
rect 5235 605 5285 635
rect 5315 605 5365 635
rect 5395 605 5445 635
rect 5475 605 5525 635
rect 5555 605 5605 635
rect 5635 605 5685 635
rect 5715 605 5765 635
rect 5795 605 5845 635
rect 5875 605 5925 635
rect 5955 605 6005 635
rect 6035 605 6085 635
rect 6115 605 6165 635
rect 6195 605 6245 635
rect 6275 605 6325 635
rect 6355 605 6405 635
rect 6435 605 6485 635
rect 6515 605 6565 635
rect 6595 605 6645 635
rect 6675 605 6725 635
rect 6755 605 6805 635
rect 6835 605 6885 635
rect 6915 605 6965 635
rect 6995 605 7045 635
rect 7075 605 7125 635
rect 7155 605 7205 635
rect 7235 605 7285 635
rect 7315 605 7365 635
rect 7395 605 7445 635
rect 7475 605 7525 635
rect 7555 605 7605 635
rect 7635 605 7685 635
rect 7715 605 7765 635
rect 7795 605 7845 635
rect 7875 605 7925 635
rect 7955 605 8005 635
rect 8035 605 8085 635
rect 8115 605 8165 635
rect 8195 605 8245 635
rect 8275 605 8325 635
rect 8355 605 8405 635
rect 8435 605 8485 635
rect 8515 605 8565 635
rect 8595 605 8645 635
rect 8675 605 8725 635
rect 8755 605 8805 635
rect 8835 605 8885 635
rect 8915 605 8965 635
rect 8995 605 9045 635
rect 9075 605 9125 635
rect 9155 605 9205 635
rect 9235 605 9285 635
rect 9315 605 9365 635
rect 9395 605 9445 635
rect 9475 605 9525 635
rect 9555 605 9605 635
rect 9635 605 9685 635
rect 9715 605 9765 635
rect 9795 605 9845 635
rect 9875 605 9925 635
rect 9955 605 10005 635
rect 10035 605 10085 635
rect 10115 605 10165 635
rect 10195 605 10245 635
rect 10275 605 10325 635
rect 10355 605 10405 635
rect 10435 605 10485 635
rect 10515 605 10645 635
rect 10675 605 10805 635
rect 10835 605 10965 635
rect 10995 605 11000 635
rect -720 600 11000 605
rect -720 555 11000 560
rect -720 525 -715 555
rect -685 525 -555 555
rect -525 525 -395 555
rect -365 525 -315 555
rect -285 525 -235 555
rect -205 525 -155 555
rect -125 525 -75 555
rect -45 525 5 555
rect 35 525 85 555
rect 115 525 165 555
rect 195 525 245 555
rect 275 525 325 555
rect 355 525 405 555
rect 435 525 485 555
rect 515 525 565 555
rect 595 525 645 555
rect 675 525 725 555
rect 755 525 805 555
rect 835 525 885 555
rect 915 525 965 555
rect 995 525 1045 555
rect 1075 525 1125 555
rect 1155 525 1205 555
rect 1235 525 1285 555
rect 1315 525 1365 555
rect 1395 525 1445 555
rect 1475 525 1525 555
rect 1555 525 1605 555
rect 1635 525 1685 555
rect 1715 525 1765 555
rect 1795 525 1845 555
rect 1875 525 1925 555
rect 1955 525 2005 555
rect 2035 525 2085 555
rect 2115 525 2165 555
rect 2195 525 2245 555
rect 2275 525 2325 555
rect 2355 525 2405 555
rect 2435 525 2485 555
rect 2515 525 2565 555
rect 2595 525 2645 555
rect 2675 525 2725 555
rect 2755 525 2805 555
rect 2835 525 2885 555
rect 2915 525 2965 555
rect 2995 525 3045 555
rect 3075 525 3125 555
rect 3155 525 3205 555
rect 3235 525 3285 555
rect 3315 525 3365 555
rect 3395 525 3445 555
rect 3475 525 3525 555
rect 3555 525 3605 555
rect 3635 525 3685 555
rect 3715 525 3765 555
rect 3795 525 3845 555
rect 3875 525 3925 555
rect 3955 525 4005 555
rect 4035 525 4085 555
rect 4115 525 4165 555
rect 4195 525 4245 555
rect 4275 525 4325 555
rect 4355 525 4405 555
rect 4435 525 4485 555
rect 4515 525 4565 555
rect 4595 525 4645 555
rect 4675 525 4725 555
rect 4755 525 4805 555
rect 4835 525 4885 555
rect 4915 525 4965 555
rect 4995 525 5045 555
rect 5075 525 5125 555
rect 5155 525 5205 555
rect 5235 525 5285 555
rect 5315 525 5365 555
rect 5395 525 5445 555
rect 5475 525 5525 555
rect 5555 525 5605 555
rect 5635 525 5685 555
rect 5715 525 5765 555
rect 5795 525 5845 555
rect 5875 525 5925 555
rect 5955 525 6005 555
rect 6035 525 6085 555
rect 6115 525 6165 555
rect 6195 525 6245 555
rect 6275 525 6325 555
rect 6355 525 6405 555
rect 6435 525 6485 555
rect 6515 525 6565 555
rect 6595 525 6645 555
rect 6675 525 6725 555
rect 6755 525 6805 555
rect 6835 525 6885 555
rect 6915 525 6965 555
rect 6995 525 7045 555
rect 7075 525 7125 555
rect 7155 525 7205 555
rect 7235 525 7285 555
rect 7315 525 7365 555
rect 7395 525 7445 555
rect 7475 525 7525 555
rect 7555 525 7605 555
rect 7635 525 7685 555
rect 7715 525 7765 555
rect 7795 525 7845 555
rect 7875 525 7925 555
rect 7955 525 8005 555
rect 8035 525 8085 555
rect 8115 525 8165 555
rect 8195 525 8245 555
rect 8275 525 8325 555
rect 8355 525 8405 555
rect 8435 525 8485 555
rect 8515 525 8565 555
rect 8595 525 8645 555
rect 8675 525 8725 555
rect 8755 525 8805 555
rect 8835 525 8885 555
rect 8915 525 8965 555
rect 8995 525 9045 555
rect 9075 525 9125 555
rect 9155 525 9205 555
rect 9235 525 9285 555
rect 9315 525 9365 555
rect 9395 525 9445 555
rect 9475 525 9525 555
rect 9555 525 9605 555
rect 9635 525 9685 555
rect 9715 525 9765 555
rect 9795 525 9845 555
rect 9875 525 9925 555
rect 9955 525 10005 555
rect 10035 525 10085 555
rect 10115 525 10165 555
rect 10195 525 10245 555
rect 10275 525 10325 555
rect 10355 525 10405 555
rect 10435 525 10485 555
rect 10515 525 10645 555
rect 10675 525 10805 555
rect 10835 525 10965 555
rect 10995 525 11000 555
rect -720 520 11000 525
rect -720 475 -520 480
rect -720 445 -715 475
rect -685 445 -555 475
rect -525 445 -520 475
rect -720 440 -520 445
rect -480 475 10600 480
rect -480 445 -475 475
rect -445 445 85 475
rect 115 445 405 475
rect 435 445 725 475
rect 755 445 1045 475
rect 1075 445 1365 475
rect 1395 445 1685 475
rect 1715 445 2005 475
rect 2035 445 2325 475
rect 2355 445 2645 475
rect 2675 445 2965 475
rect 2995 445 3285 475
rect 3315 445 3605 475
rect 3635 445 3925 475
rect 3955 445 4245 475
rect 4275 445 4565 475
rect 4595 445 4885 475
rect 4915 445 10600 475
rect -480 440 10600 445
rect 10640 475 11000 480
rect 10640 445 10645 475
rect 10675 445 10805 475
rect 10835 445 10965 475
rect 10995 445 11000 475
rect 10640 440 11000 445
rect -720 395 11000 400
rect -720 365 -715 395
rect -685 365 -555 395
rect -525 365 -395 395
rect -365 365 -315 395
rect -285 365 -235 395
rect -205 365 -155 395
rect -125 365 -75 395
rect -45 365 5 395
rect 35 365 85 395
rect 115 365 165 395
rect 195 365 245 395
rect 275 365 325 395
rect 355 365 405 395
rect 435 365 485 395
rect 515 365 565 395
rect 595 365 645 395
rect 675 365 725 395
rect 755 365 805 395
rect 835 365 885 395
rect 915 365 965 395
rect 995 365 1045 395
rect 1075 365 1125 395
rect 1155 365 1205 395
rect 1235 365 1285 395
rect 1315 365 1365 395
rect 1395 365 1445 395
rect 1475 365 1525 395
rect 1555 365 1605 395
rect 1635 365 1685 395
rect 1715 365 1765 395
rect 1795 365 1845 395
rect 1875 365 1925 395
rect 1955 365 2005 395
rect 2035 365 2085 395
rect 2115 365 2165 395
rect 2195 365 2245 395
rect 2275 365 2325 395
rect 2355 365 2405 395
rect 2435 365 2485 395
rect 2515 365 2565 395
rect 2595 365 2645 395
rect 2675 365 2725 395
rect 2755 365 2805 395
rect 2835 365 2885 395
rect 2915 365 2965 395
rect 2995 365 3045 395
rect 3075 365 3125 395
rect 3155 365 3205 395
rect 3235 365 3285 395
rect 3315 365 3365 395
rect 3395 365 3445 395
rect 3475 365 3525 395
rect 3555 365 3605 395
rect 3635 365 3685 395
rect 3715 365 3765 395
rect 3795 365 3845 395
rect 3875 365 3925 395
rect 3955 365 4005 395
rect 4035 365 4085 395
rect 4115 365 4165 395
rect 4195 365 4245 395
rect 4275 365 4325 395
rect 4355 365 4405 395
rect 4435 365 4485 395
rect 4515 365 4565 395
rect 4595 365 4645 395
rect 4675 365 4725 395
rect 4755 365 4805 395
rect 4835 365 4885 395
rect 4915 365 4965 395
rect 4995 365 5045 395
rect 5075 365 5125 395
rect 5155 365 5205 395
rect 5235 365 5285 395
rect 5315 365 5365 395
rect 5395 365 5445 395
rect 5475 365 5525 395
rect 5555 365 5605 395
rect 5635 365 5685 395
rect 5715 365 5765 395
rect 5795 365 5845 395
rect 5875 365 5925 395
rect 5955 365 6005 395
rect 6035 365 6085 395
rect 6115 365 6165 395
rect 6195 365 6245 395
rect 6275 365 6325 395
rect 6355 365 6405 395
rect 6435 365 6485 395
rect 6515 365 6565 395
rect 6595 365 6645 395
rect 6675 365 6725 395
rect 6755 365 6805 395
rect 6835 365 6885 395
rect 6915 365 6965 395
rect 6995 365 7045 395
rect 7075 365 7125 395
rect 7155 365 7205 395
rect 7235 365 7285 395
rect 7315 365 7365 395
rect 7395 365 7445 395
rect 7475 365 7525 395
rect 7555 365 7605 395
rect 7635 365 7685 395
rect 7715 365 7765 395
rect 7795 365 7845 395
rect 7875 365 7925 395
rect 7955 365 8005 395
rect 8035 365 8085 395
rect 8115 365 8165 395
rect 8195 365 8245 395
rect 8275 365 8325 395
rect 8355 365 8405 395
rect 8435 365 8485 395
rect 8515 365 8565 395
rect 8595 365 8645 395
rect 8675 365 8725 395
rect 8755 365 8805 395
rect 8835 365 8885 395
rect 8915 365 8965 395
rect 8995 365 9045 395
rect 9075 365 9125 395
rect 9155 365 9205 395
rect 9235 365 9285 395
rect 9315 365 9365 395
rect 9395 365 9445 395
rect 9475 365 9525 395
rect 9555 365 9605 395
rect 9635 365 9685 395
rect 9715 365 9765 395
rect 9795 365 9845 395
rect 9875 365 9925 395
rect 9955 365 10005 395
rect 10035 365 10085 395
rect 10115 365 10165 395
rect 10195 365 10245 395
rect 10275 365 10325 395
rect 10355 365 10405 395
rect 10435 365 10485 395
rect 10515 365 10645 395
rect 10675 365 10805 395
rect 10835 365 10965 395
rect 10995 365 11000 395
rect -720 360 11000 365
rect -720 315 -360 320
rect -720 285 -715 315
rect -685 285 -555 315
rect -525 285 -395 315
rect -365 285 -360 315
rect -720 280 -360 285
rect -320 315 10920 320
rect -320 285 5365 315
rect 5395 285 5525 315
rect 5555 285 5685 315
rect 5715 285 6005 315
rect 6035 285 6165 315
rect 6195 285 6325 315
rect 6355 285 6485 315
rect 6515 285 6645 315
rect 6675 285 6805 315
rect 6835 285 6965 315
rect 6995 285 7285 315
rect 7315 285 7445 315
rect 7475 285 7605 315
rect 7635 285 7925 315
rect 7955 285 8085 315
rect 8115 285 8245 315
rect 8275 285 8565 315
rect 8595 285 8725 315
rect 8755 285 8885 315
rect 8915 285 9045 315
rect 9075 285 9205 315
rect 9235 285 9365 315
rect 9395 285 9525 315
rect 9555 285 9845 315
rect 9875 285 10005 315
rect 10035 285 10165 315
rect 10195 285 10885 315
rect 10915 285 10920 315
rect -320 280 10920 285
rect 10960 280 11000 320
rect -720 235 11000 240
rect -720 205 -715 235
rect -685 205 -555 235
rect -525 205 -395 235
rect -365 205 -315 235
rect -285 205 -235 235
rect -205 205 -155 235
rect -125 205 -75 235
rect -45 205 5 235
rect 35 205 85 235
rect 115 205 165 235
rect 195 205 245 235
rect 275 205 325 235
rect 355 205 405 235
rect 435 205 485 235
rect 515 205 565 235
rect 595 205 645 235
rect 675 205 725 235
rect 755 205 805 235
rect 835 205 885 235
rect 915 205 965 235
rect 995 205 1045 235
rect 1075 205 1125 235
rect 1155 205 1205 235
rect 1235 205 1285 235
rect 1315 205 1365 235
rect 1395 205 1445 235
rect 1475 205 1525 235
rect 1555 205 1605 235
rect 1635 205 1685 235
rect 1715 205 1765 235
rect 1795 205 1845 235
rect 1875 205 1925 235
rect 1955 205 2005 235
rect 2035 205 2085 235
rect 2115 205 2165 235
rect 2195 205 2245 235
rect 2275 205 2325 235
rect 2355 205 2405 235
rect 2435 205 2485 235
rect 2515 205 2565 235
rect 2595 205 2645 235
rect 2675 205 2725 235
rect 2755 205 2805 235
rect 2835 205 2885 235
rect 2915 205 2965 235
rect 2995 205 3045 235
rect 3075 205 3125 235
rect 3155 205 3205 235
rect 3235 205 3285 235
rect 3315 205 3365 235
rect 3395 205 3445 235
rect 3475 205 3525 235
rect 3555 205 3605 235
rect 3635 205 3685 235
rect 3715 205 3765 235
rect 3795 205 3845 235
rect 3875 205 3925 235
rect 3955 205 4005 235
rect 4035 205 4085 235
rect 4115 205 4165 235
rect 4195 205 4245 235
rect 4275 205 4325 235
rect 4355 205 4405 235
rect 4435 205 4485 235
rect 4515 205 4565 235
rect 4595 205 4645 235
rect 4675 205 4725 235
rect 4755 205 4805 235
rect 4835 205 4885 235
rect 4915 205 4965 235
rect 4995 205 5045 235
rect 5075 205 5125 235
rect 5155 205 5205 235
rect 5235 205 5285 235
rect 5315 205 5365 235
rect 5395 205 5445 235
rect 5475 205 5525 235
rect 5555 205 5605 235
rect 5635 205 5685 235
rect 5715 205 5765 235
rect 5795 205 5845 235
rect 5875 205 5925 235
rect 5955 205 6005 235
rect 6035 205 6085 235
rect 6115 205 6165 235
rect 6195 205 6245 235
rect 6275 205 6325 235
rect 6355 205 6405 235
rect 6435 205 6485 235
rect 6515 205 6565 235
rect 6595 205 6645 235
rect 6675 205 6725 235
rect 6755 205 6805 235
rect 6835 205 6885 235
rect 6915 205 6965 235
rect 6995 205 7045 235
rect 7075 205 7125 235
rect 7155 205 7205 235
rect 7235 205 7285 235
rect 7315 205 7365 235
rect 7395 205 7445 235
rect 7475 205 7525 235
rect 7555 205 7605 235
rect 7635 205 7685 235
rect 7715 205 7765 235
rect 7795 205 7845 235
rect 7875 205 7925 235
rect 7955 205 8005 235
rect 8035 205 8085 235
rect 8115 205 8165 235
rect 8195 205 8245 235
rect 8275 205 8325 235
rect 8355 205 8405 235
rect 8435 205 8485 235
rect 8515 205 8565 235
rect 8595 205 8645 235
rect 8675 205 8725 235
rect 8755 205 8805 235
rect 8835 205 8885 235
rect 8915 205 8965 235
rect 8995 205 9045 235
rect 9075 205 9125 235
rect 9155 205 9205 235
rect 9235 205 9285 235
rect 9315 205 9365 235
rect 9395 205 9445 235
rect 9475 205 9525 235
rect 9555 205 9605 235
rect 9635 205 9685 235
rect 9715 205 9765 235
rect 9795 205 9845 235
rect 9875 205 9925 235
rect 9955 205 10005 235
rect 10035 205 10085 235
rect 10115 205 10165 235
rect 10195 205 10245 235
rect 10275 205 10325 235
rect 10355 205 10405 235
rect 10435 205 10485 235
rect 10515 205 10645 235
rect 10675 205 10805 235
rect 10835 205 10965 235
rect 10995 205 11000 235
rect -720 200 11000 205
rect -720 155 -360 160
rect -720 125 -715 155
rect -685 125 -555 155
rect -525 125 -395 155
rect -365 125 -360 155
rect -720 120 -360 125
rect -320 155 10760 160
rect -320 125 10 155
rect 190 125 330 155
rect 510 125 650 155
rect 830 125 970 155
rect 1150 125 1205 155
rect 1235 125 1290 155
rect 1470 125 1610 155
rect 1790 125 1930 155
rect 2110 125 2250 155
rect 2430 125 2570 155
rect 2750 125 2890 155
rect 3070 125 3210 155
rect 3390 125 3530 155
rect 3710 125 3765 155
rect 3795 125 3850 155
rect 4030 125 4170 155
rect 4350 125 4490 155
rect 4670 125 4810 155
rect 4990 125 5045 155
rect 5075 125 5290 155
rect 5470 125 5610 155
rect 5790 125 5930 155
rect 6110 125 6250 155
rect 6430 125 6570 155
rect 6750 125 6890 155
rect 7070 125 7210 155
rect 7390 125 7530 155
rect 7710 125 7850 155
rect 8030 125 8170 155
rect 8350 125 8490 155
rect 8670 125 8810 155
rect 8990 125 9130 155
rect 9310 125 9450 155
rect 9630 125 9770 155
rect 9950 125 10090 155
rect 10270 125 10725 155
rect 10755 125 10760 155
rect -320 120 10760 125
rect 10800 155 11000 160
rect 10800 125 10805 155
rect 10835 125 10965 155
rect 10995 125 11000 155
rect 10800 120 11000 125
rect -720 75 11000 80
rect -720 45 -715 75
rect -685 45 -555 75
rect -525 45 -395 75
rect -365 45 -315 75
rect -285 45 -235 75
rect -205 45 -155 75
rect -125 45 -75 75
rect -45 45 5 75
rect 35 45 85 75
rect 115 45 165 75
rect 195 45 245 75
rect 275 45 325 75
rect 355 45 405 75
rect 435 45 485 75
rect 515 45 565 75
rect 595 45 645 75
rect 675 45 725 75
rect 755 45 805 75
rect 835 45 885 75
rect 915 45 965 75
rect 995 45 1045 75
rect 1075 45 1125 75
rect 1155 45 1205 75
rect 1235 45 1285 75
rect 1315 45 1365 75
rect 1395 45 1445 75
rect 1475 45 1525 75
rect 1555 45 1605 75
rect 1635 45 1685 75
rect 1715 45 1765 75
rect 1795 45 1845 75
rect 1875 45 1925 75
rect 1955 45 2005 75
rect 2035 45 2085 75
rect 2115 45 2165 75
rect 2195 45 2245 75
rect 2275 45 2325 75
rect 2355 45 2405 75
rect 2435 45 2485 75
rect 2515 45 2565 75
rect 2595 45 2645 75
rect 2675 45 2725 75
rect 2755 45 2805 75
rect 2835 45 2885 75
rect 2915 45 2965 75
rect 2995 45 3045 75
rect 3075 45 3125 75
rect 3155 45 3205 75
rect 3235 45 3285 75
rect 3315 45 3365 75
rect 3395 45 3445 75
rect 3475 45 3525 75
rect 3555 45 3605 75
rect 3635 45 3685 75
rect 3715 45 3765 75
rect 3795 45 3845 75
rect 3875 45 3925 75
rect 3955 45 4005 75
rect 4035 45 4085 75
rect 4115 45 4165 75
rect 4195 45 4245 75
rect 4275 45 4325 75
rect 4355 45 4405 75
rect 4435 45 4485 75
rect 4515 45 4565 75
rect 4595 45 4645 75
rect 4675 45 4725 75
rect 4755 45 4805 75
rect 4835 45 4885 75
rect 4915 45 4965 75
rect 4995 45 5045 75
rect 5075 45 5125 75
rect 5155 45 5205 75
rect 5235 45 5285 75
rect 5315 45 5365 75
rect 5395 45 5445 75
rect 5475 45 5525 75
rect 5555 45 5605 75
rect 5635 45 5685 75
rect 5715 45 5765 75
rect 5795 45 5845 75
rect 5875 45 5925 75
rect 5955 45 6005 75
rect 6035 45 6085 75
rect 6115 45 6165 75
rect 6195 45 6245 75
rect 6275 45 6325 75
rect 6355 45 6405 75
rect 6435 45 6485 75
rect 6515 45 6565 75
rect 6595 45 6645 75
rect 6675 45 6725 75
rect 6755 45 6805 75
rect 6835 45 6885 75
rect 6915 45 6965 75
rect 6995 45 7045 75
rect 7075 45 7125 75
rect 7155 45 7205 75
rect 7235 45 7285 75
rect 7315 45 7365 75
rect 7395 45 7445 75
rect 7475 45 7525 75
rect 7555 45 7605 75
rect 7635 45 7685 75
rect 7715 45 7765 75
rect 7795 45 7845 75
rect 7875 45 7925 75
rect 7955 45 8005 75
rect 8035 45 8085 75
rect 8115 45 8165 75
rect 8195 45 8245 75
rect 8275 45 8325 75
rect 8355 45 8405 75
rect 8435 45 8485 75
rect 8515 45 8565 75
rect 8595 45 8645 75
rect 8675 45 8725 75
rect 8755 45 8805 75
rect 8835 45 8885 75
rect 8915 45 8965 75
rect 8995 45 9045 75
rect 9075 45 9125 75
rect 9155 45 9205 75
rect 9235 45 9285 75
rect 9315 45 9365 75
rect 9395 45 9445 75
rect 9475 45 9525 75
rect 9555 45 9605 75
rect 9635 45 9685 75
rect 9715 45 9765 75
rect 9795 45 9845 75
rect 9875 45 9925 75
rect 9955 45 10005 75
rect 10035 45 10085 75
rect 10115 45 10165 75
rect 10195 45 10245 75
rect 10275 45 10325 75
rect 10355 45 10405 75
rect 10435 45 10485 75
rect 10515 45 10645 75
rect 10675 45 10805 75
rect 10835 45 10965 75
rect 10995 45 11000 75
rect -720 40 11000 45
rect -720 -5 11000 0
rect -720 -35 -715 -5
rect -685 -35 -555 -5
rect -525 -35 -395 -5
rect -365 -35 -315 -5
rect -285 -35 -235 -5
rect -205 -35 -155 -5
rect -125 -35 -75 -5
rect -45 -35 5 -5
rect 35 -35 85 -5
rect 115 -35 165 -5
rect 195 -35 245 -5
rect 275 -35 325 -5
rect 355 -35 405 -5
rect 435 -35 485 -5
rect 515 -35 565 -5
rect 595 -35 645 -5
rect 675 -35 725 -5
rect 755 -35 805 -5
rect 835 -35 885 -5
rect 915 -35 965 -5
rect 995 -35 1045 -5
rect 1075 -35 1125 -5
rect 1155 -35 1205 -5
rect 1235 -35 1285 -5
rect 1315 -35 1365 -5
rect 1395 -35 1445 -5
rect 1475 -35 1525 -5
rect 1555 -35 1605 -5
rect 1635 -35 1685 -5
rect 1715 -35 1765 -5
rect 1795 -35 1845 -5
rect 1875 -35 1925 -5
rect 1955 -35 2005 -5
rect 2035 -35 2085 -5
rect 2115 -35 2165 -5
rect 2195 -35 2245 -5
rect 2275 -35 2325 -5
rect 2355 -35 2405 -5
rect 2435 -35 2485 -5
rect 2515 -35 2565 -5
rect 2595 -35 2645 -5
rect 2675 -35 2725 -5
rect 2755 -35 2805 -5
rect 2835 -35 2885 -5
rect 2915 -35 2965 -5
rect 2995 -35 3045 -5
rect 3075 -35 3125 -5
rect 3155 -35 3205 -5
rect 3235 -35 3285 -5
rect 3315 -35 3365 -5
rect 3395 -35 3445 -5
rect 3475 -35 3525 -5
rect 3555 -35 3605 -5
rect 3635 -35 3685 -5
rect 3715 -35 3765 -5
rect 3795 -35 3845 -5
rect 3875 -35 3925 -5
rect 3955 -35 4005 -5
rect 4035 -35 4085 -5
rect 4115 -35 4165 -5
rect 4195 -35 4245 -5
rect 4275 -35 4325 -5
rect 4355 -35 4405 -5
rect 4435 -35 4485 -5
rect 4515 -35 4565 -5
rect 4595 -35 4645 -5
rect 4675 -35 4725 -5
rect 4755 -35 4805 -5
rect 4835 -35 4885 -5
rect 4915 -35 4965 -5
rect 4995 -35 5045 -5
rect 5075 -35 5125 -5
rect 5155 -35 5205 -5
rect 5235 -35 5285 -5
rect 5315 -35 5365 -5
rect 5395 -35 5445 -5
rect 5475 -35 5525 -5
rect 5555 -35 5605 -5
rect 5635 -35 5685 -5
rect 5715 -35 5765 -5
rect 5795 -35 5845 -5
rect 5875 -35 5925 -5
rect 5955 -35 6005 -5
rect 6035 -35 6085 -5
rect 6115 -35 6165 -5
rect 6195 -35 6245 -5
rect 6275 -35 6325 -5
rect 6355 -35 6405 -5
rect 6435 -35 6485 -5
rect 6515 -35 6565 -5
rect 6595 -35 6645 -5
rect 6675 -35 6725 -5
rect 6755 -35 6805 -5
rect 6835 -35 6885 -5
rect 6915 -35 6965 -5
rect 6995 -35 7045 -5
rect 7075 -35 7125 -5
rect 7155 -35 7205 -5
rect 7235 -35 7285 -5
rect 7315 -35 7365 -5
rect 7395 -35 7445 -5
rect 7475 -35 7525 -5
rect 7555 -35 7605 -5
rect 7635 -35 7685 -5
rect 7715 -35 7765 -5
rect 7795 -35 7845 -5
rect 7875 -35 7925 -5
rect 7955 -35 8005 -5
rect 8035 -35 8085 -5
rect 8115 -35 8165 -5
rect 8195 -35 8245 -5
rect 8275 -35 8325 -5
rect 8355 -35 8405 -5
rect 8435 -35 8485 -5
rect 8515 -35 8565 -5
rect 8595 -35 8645 -5
rect 8675 -35 8725 -5
rect 8755 -35 8805 -5
rect 8835 -35 8885 -5
rect 8915 -35 8965 -5
rect 8995 -35 9045 -5
rect 9075 -35 9125 -5
rect 9155 -35 9205 -5
rect 9235 -35 9285 -5
rect 9315 -35 9365 -5
rect 9395 -35 9445 -5
rect 9475 -35 9525 -5
rect 9555 -35 9605 -5
rect 9635 -35 9685 -5
rect 9715 -35 9765 -5
rect 9795 -35 9845 -5
rect 9875 -35 9925 -5
rect 9955 -35 10005 -5
rect 10035 -35 10085 -5
rect 10115 -35 10165 -5
rect 10195 -35 10245 -5
rect 10275 -35 10325 -5
rect 10355 -35 10405 -5
rect 10435 -35 10485 -5
rect 10515 -35 10645 -5
rect 10675 -35 10805 -5
rect 10835 -35 10965 -5
rect 10995 -35 11000 -5
rect -720 -40 11000 -35
rect -720 -85 11000 -80
rect -720 -115 -715 -85
rect -685 -115 -555 -85
rect -525 -115 -395 -85
rect -365 -115 -315 -85
rect -285 -115 -235 -85
rect -205 -115 -155 -85
rect -125 -115 -75 -85
rect -45 -115 5 -85
rect 35 -115 85 -85
rect 115 -115 165 -85
rect 195 -115 245 -85
rect 275 -115 325 -85
rect 355 -115 405 -85
rect 435 -115 485 -85
rect 515 -115 565 -85
rect 595 -115 645 -85
rect 675 -115 725 -85
rect 755 -115 805 -85
rect 835 -115 885 -85
rect 915 -115 965 -85
rect 995 -115 1045 -85
rect 1075 -115 1125 -85
rect 1155 -115 1205 -85
rect 1235 -115 1285 -85
rect 1315 -115 1365 -85
rect 1395 -115 1445 -85
rect 1475 -115 1525 -85
rect 1555 -115 1605 -85
rect 1635 -115 1685 -85
rect 1715 -115 1765 -85
rect 1795 -115 1845 -85
rect 1875 -115 1925 -85
rect 1955 -115 2005 -85
rect 2035 -115 2085 -85
rect 2115 -115 2165 -85
rect 2195 -115 2245 -85
rect 2275 -115 2325 -85
rect 2355 -115 2405 -85
rect 2435 -115 2485 -85
rect 2515 -115 2565 -85
rect 2595 -115 2645 -85
rect 2675 -115 2725 -85
rect 2755 -115 2805 -85
rect 2835 -115 2885 -85
rect 2915 -115 2965 -85
rect 2995 -115 3045 -85
rect 3075 -115 3125 -85
rect 3155 -115 3205 -85
rect 3235 -115 3285 -85
rect 3315 -115 3365 -85
rect 3395 -115 3445 -85
rect 3475 -115 3525 -85
rect 3555 -115 3605 -85
rect 3635 -115 3685 -85
rect 3715 -115 3765 -85
rect 3795 -115 3845 -85
rect 3875 -115 3925 -85
rect 3955 -115 4005 -85
rect 4035 -115 4085 -85
rect 4115 -115 4165 -85
rect 4195 -115 4245 -85
rect 4275 -115 4325 -85
rect 4355 -115 4405 -85
rect 4435 -115 4485 -85
rect 4515 -115 4565 -85
rect 4595 -115 4645 -85
rect 4675 -115 4725 -85
rect 4755 -115 4805 -85
rect 4835 -115 4885 -85
rect 4915 -115 4965 -85
rect 4995 -115 5045 -85
rect 5075 -115 5125 -85
rect 5155 -115 5205 -85
rect 5235 -115 5285 -85
rect 5315 -115 5365 -85
rect 5395 -115 5445 -85
rect 5475 -115 5525 -85
rect 5555 -115 5605 -85
rect 5635 -115 5685 -85
rect 5715 -115 5765 -85
rect 5795 -115 5845 -85
rect 5875 -115 5925 -85
rect 5955 -115 6005 -85
rect 6035 -115 6085 -85
rect 6115 -115 6165 -85
rect 6195 -115 6245 -85
rect 6275 -115 6325 -85
rect 6355 -115 6405 -85
rect 6435 -115 6485 -85
rect 6515 -115 6565 -85
rect 6595 -115 6645 -85
rect 6675 -115 6725 -85
rect 6755 -115 6805 -85
rect 6835 -115 6885 -85
rect 6915 -115 6965 -85
rect 6995 -115 7045 -85
rect 7075 -115 7125 -85
rect 7155 -115 7205 -85
rect 7235 -115 7285 -85
rect 7315 -115 7365 -85
rect 7395 -115 7445 -85
rect 7475 -115 7525 -85
rect 7555 -115 7605 -85
rect 7635 -115 7685 -85
rect 7715 -115 7765 -85
rect 7795 -115 7845 -85
rect 7875 -115 7925 -85
rect 7955 -115 8005 -85
rect 8035 -115 8085 -85
rect 8115 -115 8165 -85
rect 8195 -115 8245 -85
rect 8275 -115 8325 -85
rect 8355 -115 8405 -85
rect 8435 -115 8485 -85
rect 8515 -115 8565 -85
rect 8595 -115 8645 -85
rect 8675 -115 8725 -85
rect 8755 -115 8805 -85
rect 8835 -115 8885 -85
rect 8915 -115 8965 -85
rect 8995 -115 9045 -85
rect 9075 -115 9125 -85
rect 9155 -115 9205 -85
rect 9235 -115 9285 -85
rect 9315 -115 9365 -85
rect 9395 -115 9445 -85
rect 9475 -115 9525 -85
rect 9555 -115 9605 -85
rect 9635 -115 9685 -85
rect 9715 -115 9765 -85
rect 9795 -115 9845 -85
rect 9875 -115 9925 -85
rect 9955 -115 10005 -85
rect 10035 -115 10085 -85
rect 10115 -115 10165 -85
rect 10195 -115 10245 -85
rect 10275 -115 10325 -85
rect 10355 -115 10405 -85
rect 10435 -115 10485 -85
rect 10515 -115 10645 -85
rect 10675 -115 10805 -85
rect 10835 -115 10965 -85
rect 10995 -115 11000 -85
rect -720 -120 11000 -115
<< via2 >>
rect -715 1005 -685 1035
rect -555 1005 -525 1035
rect -395 1005 -365 1035
rect -315 1005 -285 1035
rect -235 1005 -205 1035
rect -155 1005 -125 1035
rect -75 1005 -45 1035
rect 5 1005 35 1035
rect 85 1005 115 1035
rect 165 1005 195 1035
rect 245 1005 275 1035
rect 325 1005 355 1035
rect 405 1005 435 1035
rect 485 1005 515 1035
rect 565 1005 595 1035
rect 645 1005 675 1035
rect 725 1005 755 1035
rect 805 1005 835 1035
rect 885 1005 915 1035
rect 965 1005 995 1035
rect 1045 1005 1075 1035
rect 1125 1005 1155 1035
rect 1205 1005 1235 1035
rect 1285 1005 1315 1035
rect 1365 1005 1395 1035
rect 1445 1005 1475 1035
rect 1525 1005 1555 1035
rect 1605 1005 1635 1035
rect 1685 1005 1715 1035
rect 1765 1005 1795 1035
rect 1845 1005 1875 1035
rect 1925 1005 1955 1035
rect 2005 1005 2035 1035
rect 2085 1005 2115 1035
rect 2165 1005 2195 1035
rect 2245 1005 2275 1035
rect 2325 1005 2355 1035
rect 2405 1005 2435 1035
rect 2485 1005 2515 1035
rect 2565 1005 2595 1035
rect 2645 1005 2675 1035
rect 2725 1005 2755 1035
rect 2805 1005 2835 1035
rect 2885 1005 2915 1035
rect 2965 1005 2995 1035
rect 3045 1005 3075 1035
rect 3125 1005 3155 1035
rect 3205 1005 3235 1035
rect 3285 1005 3315 1035
rect 3365 1005 3395 1035
rect 3445 1005 3475 1035
rect 3525 1005 3555 1035
rect 3605 1005 3635 1035
rect 3685 1005 3715 1035
rect 3765 1005 3795 1035
rect 3845 1005 3875 1035
rect 3925 1005 3955 1035
rect 4005 1005 4035 1035
rect 4085 1005 4115 1035
rect 4165 1005 4195 1035
rect 4245 1005 4275 1035
rect 4325 1005 4355 1035
rect 4405 1005 4435 1035
rect 4485 1005 4515 1035
rect 4565 1005 4595 1035
rect 4645 1005 4675 1035
rect 4725 1005 4755 1035
rect 4805 1005 4835 1035
rect 4885 1005 4915 1035
rect 4965 1005 4995 1035
rect 5045 1005 5075 1035
rect 5125 1005 5155 1035
rect 5205 1005 5235 1035
rect 5285 1005 5315 1035
rect 5365 1005 5395 1035
rect 5445 1005 5475 1035
rect 5525 1005 5555 1035
rect 5605 1005 5635 1035
rect 5685 1005 5715 1035
rect 5765 1005 5795 1035
rect 5845 1005 5875 1035
rect 5925 1005 5955 1035
rect 6005 1005 6035 1035
rect 6085 1005 6115 1035
rect 6165 1005 6195 1035
rect 6245 1005 6275 1035
rect 6325 1005 6355 1035
rect 6405 1005 6435 1035
rect 6485 1005 6515 1035
rect 6565 1005 6595 1035
rect 6645 1005 6675 1035
rect 6725 1005 6755 1035
rect 6805 1005 6835 1035
rect 6885 1005 6915 1035
rect 6965 1005 6995 1035
rect 7045 1005 7075 1035
rect 7125 1005 7155 1035
rect 7205 1005 7235 1035
rect 7285 1005 7315 1035
rect 7365 1005 7395 1035
rect 7445 1005 7475 1035
rect 7525 1005 7555 1035
rect 7605 1005 7635 1035
rect 7685 1005 7715 1035
rect 7765 1005 7795 1035
rect 7845 1005 7875 1035
rect 7925 1005 7955 1035
rect 8005 1005 8035 1035
rect 8085 1005 8115 1035
rect 8165 1005 8195 1035
rect 8245 1005 8275 1035
rect 8325 1005 8355 1035
rect 8405 1005 8435 1035
rect 8485 1005 8515 1035
rect 8565 1005 8595 1035
rect 8645 1005 8675 1035
rect 8725 1005 8755 1035
rect 8805 1005 8835 1035
rect 8885 1005 8915 1035
rect 8965 1005 8995 1035
rect 9045 1005 9075 1035
rect 9125 1005 9155 1035
rect 9205 1005 9235 1035
rect 9285 1005 9315 1035
rect 9365 1005 9395 1035
rect 9445 1005 9475 1035
rect 9525 1005 9555 1035
rect 9605 1005 9635 1035
rect 9685 1005 9715 1035
rect 9765 1005 9795 1035
rect 9845 1005 9875 1035
rect 9925 1005 9955 1035
rect 10005 1005 10035 1035
rect 10085 1005 10115 1035
rect 10165 1005 10195 1035
rect 10245 1005 10275 1035
rect 10325 1005 10355 1035
rect 10405 1005 10435 1035
rect 10485 1005 10515 1035
rect 10645 1005 10675 1035
rect 10805 1005 10835 1035
rect 10965 1005 10995 1035
rect -715 925 -685 955
rect -555 925 -525 955
rect -395 925 -365 955
rect -315 925 -285 955
rect -235 925 -205 955
rect -155 925 -125 955
rect -75 925 -45 955
rect 5 925 35 955
rect 85 925 115 955
rect 165 925 195 955
rect 245 925 275 955
rect 325 925 355 955
rect 405 925 435 955
rect 485 925 515 955
rect 565 925 595 955
rect 645 925 675 955
rect 725 925 755 955
rect 805 925 835 955
rect 885 925 915 955
rect 965 925 995 955
rect 1045 925 1075 955
rect 1125 925 1155 955
rect 1205 925 1235 955
rect 1285 925 1315 955
rect 1365 925 1395 955
rect 1445 925 1475 955
rect 1525 925 1555 955
rect 1605 925 1635 955
rect 1685 925 1715 955
rect 1765 925 1795 955
rect 1845 925 1875 955
rect 1925 925 1955 955
rect 2005 925 2035 955
rect 2085 925 2115 955
rect 2165 925 2195 955
rect 2245 925 2275 955
rect 2325 925 2355 955
rect 2405 925 2435 955
rect 2485 925 2515 955
rect 2565 925 2595 955
rect 2645 925 2675 955
rect 2725 925 2755 955
rect 2805 925 2835 955
rect 2885 925 2915 955
rect 2965 925 2995 955
rect 3045 925 3075 955
rect 3125 925 3155 955
rect 3205 925 3235 955
rect 3285 925 3315 955
rect 3365 925 3395 955
rect 3445 925 3475 955
rect 3525 925 3555 955
rect 3605 925 3635 955
rect 3685 925 3715 955
rect 3765 925 3795 955
rect 3845 925 3875 955
rect 3925 925 3955 955
rect 4005 925 4035 955
rect 4085 925 4115 955
rect 4165 925 4195 955
rect 4245 925 4275 955
rect 4325 925 4355 955
rect 4405 925 4435 955
rect 4485 925 4515 955
rect 4565 925 4595 955
rect 4645 925 4675 955
rect 4725 925 4755 955
rect 4805 925 4835 955
rect 4885 925 4915 955
rect 4965 925 4995 955
rect 5045 925 5075 955
rect 5125 925 5155 955
rect 5205 925 5235 955
rect 5285 925 5315 955
rect 5365 925 5395 955
rect 5445 925 5475 955
rect 5525 925 5555 955
rect 5605 925 5635 955
rect 5685 925 5715 955
rect 5765 925 5795 955
rect 5845 925 5875 955
rect 5925 925 5955 955
rect 6005 925 6035 955
rect 6085 925 6115 955
rect 6165 925 6195 955
rect 6245 925 6275 955
rect 6325 925 6355 955
rect 6405 925 6435 955
rect 6485 925 6515 955
rect 6565 925 6595 955
rect 6645 925 6675 955
rect 6725 925 6755 955
rect 6805 925 6835 955
rect 6885 925 6915 955
rect 6965 925 6995 955
rect 7045 925 7075 955
rect 7125 925 7155 955
rect 7205 925 7235 955
rect 7285 925 7315 955
rect 7365 925 7395 955
rect 7445 925 7475 955
rect 7525 925 7555 955
rect 7605 925 7635 955
rect 7685 925 7715 955
rect 7765 925 7795 955
rect 7845 925 7875 955
rect 7925 925 7955 955
rect 8005 925 8035 955
rect 8085 925 8115 955
rect 8165 925 8195 955
rect 8245 925 8275 955
rect 8325 925 8355 955
rect 8405 925 8435 955
rect 8485 925 8515 955
rect 8565 925 8595 955
rect 8645 925 8675 955
rect 8725 925 8755 955
rect 8805 925 8835 955
rect 8885 925 8915 955
rect 8965 925 8995 955
rect 9045 925 9075 955
rect 9125 925 9155 955
rect 9205 925 9235 955
rect 9285 925 9315 955
rect 9365 925 9395 955
rect 9445 925 9475 955
rect 9525 925 9555 955
rect 9605 925 9635 955
rect 9685 925 9715 955
rect 9765 925 9795 955
rect 9845 925 9875 955
rect 9925 925 9955 955
rect 10005 925 10035 955
rect 10085 925 10115 955
rect 10165 925 10195 955
rect 10245 925 10275 955
rect 10325 925 10355 955
rect 10405 925 10435 955
rect 10485 925 10515 955
rect 10645 925 10675 955
rect 10805 925 10835 955
rect 10965 925 10995 955
rect -715 845 -685 875
rect -555 845 -525 875
rect -395 845 -365 875
rect -315 845 -285 875
rect -235 845 -205 875
rect -155 845 -125 875
rect -75 845 -45 875
rect 5 845 35 875
rect 85 845 115 875
rect 165 845 195 875
rect 245 845 275 875
rect 325 845 355 875
rect 405 845 435 875
rect 485 845 515 875
rect 565 845 595 875
rect 645 845 675 875
rect 725 845 755 875
rect 805 845 835 875
rect 885 845 915 875
rect 965 845 995 875
rect 1045 845 1075 875
rect 1125 845 1155 875
rect 1205 845 1235 875
rect 1285 845 1315 875
rect 1365 845 1395 875
rect 1445 845 1475 875
rect 1525 845 1555 875
rect 1605 845 1635 875
rect 1685 845 1715 875
rect 1765 845 1795 875
rect 1845 845 1875 875
rect 1925 845 1955 875
rect 2005 845 2035 875
rect 2085 845 2115 875
rect 2165 845 2195 875
rect 2245 845 2275 875
rect 2325 845 2355 875
rect 2405 845 2435 875
rect 2485 845 2515 875
rect 2565 845 2595 875
rect 2645 845 2675 875
rect 2725 845 2755 875
rect 2805 845 2835 875
rect 2885 845 2915 875
rect 2965 845 2995 875
rect 3045 845 3075 875
rect 3125 845 3155 875
rect 3205 845 3235 875
rect 3285 845 3315 875
rect 3365 845 3395 875
rect 3445 845 3475 875
rect 3525 845 3555 875
rect 3605 845 3635 875
rect 3685 845 3715 875
rect 3765 845 3795 875
rect 3845 845 3875 875
rect 3925 845 3955 875
rect 4005 845 4035 875
rect 4085 845 4115 875
rect 4165 845 4195 875
rect 4245 845 4275 875
rect 4325 845 4355 875
rect 4405 845 4435 875
rect 4485 845 4515 875
rect 4565 845 4595 875
rect 4645 845 4675 875
rect 4725 845 4755 875
rect 4805 845 4835 875
rect 4885 845 4915 875
rect 4965 845 4995 875
rect 5045 845 5075 875
rect 5125 845 5155 875
rect 5205 845 5235 875
rect 5285 845 5315 875
rect 5365 845 5395 875
rect 5445 845 5475 875
rect 5525 845 5555 875
rect 5605 845 5635 875
rect 5685 845 5715 875
rect 5765 845 5795 875
rect 5845 845 5875 875
rect 5925 845 5955 875
rect 6005 845 6035 875
rect 6085 845 6115 875
rect 6165 845 6195 875
rect 6245 845 6275 875
rect 6325 845 6355 875
rect 6405 845 6435 875
rect 6485 845 6515 875
rect 6565 845 6595 875
rect 6645 845 6675 875
rect 6725 845 6755 875
rect 6805 845 6835 875
rect 6885 845 6915 875
rect 6965 845 6995 875
rect 7045 845 7075 875
rect 7125 845 7155 875
rect 7205 845 7235 875
rect 7285 845 7315 875
rect 7365 845 7395 875
rect 7445 845 7475 875
rect 7525 845 7555 875
rect 7605 845 7635 875
rect 7685 845 7715 875
rect 7765 845 7795 875
rect 7845 845 7875 875
rect 7925 845 7955 875
rect 8005 845 8035 875
rect 8085 845 8115 875
rect 8165 845 8195 875
rect 8245 845 8275 875
rect 8325 845 8355 875
rect 8405 845 8435 875
rect 8485 845 8515 875
rect 8565 845 8595 875
rect 8645 845 8675 875
rect 8725 845 8755 875
rect 8805 845 8835 875
rect 8885 845 8915 875
rect 8965 845 8995 875
rect 9045 845 9075 875
rect 9125 845 9155 875
rect 9205 845 9235 875
rect 9285 845 9315 875
rect 9365 845 9395 875
rect 9445 845 9475 875
rect 9525 845 9555 875
rect 9605 845 9635 875
rect 9685 845 9715 875
rect 9765 845 9795 875
rect 9845 845 9875 875
rect 9925 845 9955 875
rect 10005 845 10035 875
rect 10085 845 10115 875
rect 10165 845 10195 875
rect 10245 845 10275 875
rect 10325 845 10355 875
rect 10405 845 10435 875
rect 10485 845 10515 875
rect 10645 845 10675 875
rect 10805 845 10835 875
rect 10965 845 10995 875
rect -635 765 -605 795
rect 10645 765 10675 795
rect 10805 765 10835 795
rect 10965 765 10995 795
rect -635 685 -605 715
rect 10645 685 10675 715
rect 10805 685 10835 715
rect 10965 685 10995 715
rect -715 605 -685 635
rect -555 605 -525 635
rect -395 605 -365 635
rect -315 605 -285 635
rect -235 605 -205 635
rect -155 605 -125 635
rect -75 605 -45 635
rect 5 605 35 635
rect 85 605 115 635
rect 165 605 195 635
rect 245 605 275 635
rect 325 605 355 635
rect 405 605 435 635
rect 485 605 515 635
rect 565 605 595 635
rect 645 605 675 635
rect 725 605 755 635
rect 805 605 835 635
rect 885 605 915 635
rect 965 605 995 635
rect 1045 605 1075 635
rect 1125 605 1155 635
rect 1205 605 1235 635
rect 1285 605 1315 635
rect 1365 605 1395 635
rect 1445 605 1475 635
rect 1525 605 1555 635
rect 1605 605 1635 635
rect 1685 605 1715 635
rect 1765 605 1795 635
rect 1845 605 1875 635
rect 1925 605 1955 635
rect 2005 605 2035 635
rect 2085 605 2115 635
rect 2165 605 2195 635
rect 2245 605 2275 635
rect 2325 605 2355 635
rect 2405 605 2435 635
rect 2485 605 2515 635
rect 2565 605 2595 635
rect 2645 605 2675 635
rect 2725 605 2755 635
rect 2805 605 2835 635
rect 2885 605 2915 635
rect 2965 605 2995 635
rect 3045 605 3075 635
rect 3125 605 3155 635
rect 3205 605 3235 635
rect 3285 605 3315 635
rect 3365 605 3395 635
rect 3445 605 3475 635
rect 3525 605 3555 635
rect 3605 605 3635 635
rect 3685 605 3715 635
rect 3765 605 3795 635
rect 3845 605 3875 635
rect 3925 605 3955 635
rect 4005 605 4035 635
rect 4085 605 4115 635
rect 4165 605 4195 635
rect 4245 605 4275 635
rect 4325 605 4355 635
rect 4405 605 4435 635
rect 4485 605 4515 635
rect 4565 605 4595 635
rect 4645 605 4675 635
rect 4725 605 4755 635
rect 4805 605 4835 635
rect 4885 605 4915 635
rect 4965 605 4995 635
rect 5045 605 5075 635
rect 5125 605 5155 635
rect 5205 605 5235 635
rect 5285 605 5315 635
rect 5365 605 5395 635
rect 5445 605 5475 635
rect 5525 605 5555 635
rect 5605 605 5635 635
rect 5685 605 5715 635
rect 5765 605 5795 635
rect 5845 605 5875 635
rect 5925 605 5955 635
rect 6005 605 6035 635
rect 6085 605 6115 635
rect 6165 605 6195 635
rect 6245 605 6275 635
rect 6325 605 6355 635
rect 6405 605 6435 635
rect 6485 605 6515 635
rect 6565 605 6595 635
rect 6645 605 6675 635
rect 6725 605 6755 635
rect 6805 605 6835 635
rect 6885 605 6915 635
rect 6965 605 6995 635
rect 7045 605 7075 635
rect 7125 605 7155 635
rect 7205 605 7235 635
rect 7285 605 7315 635
rect 7365 605 7395 635
rect 7445 605 7475 635
rect 7525 605 7555 635
rect 7605 605 7635 635
rect 7685 605 7715 635
rect 7765 605 7795 635
rect 7845 605 7875 635
rect 7925 605 7955 635
rect 8005 605 8035 635
rect 8085 605 8115 635
rect 8165 605 8195 635
rect 8245 605 8275 635
rect 8325 605 8355 635
rect 8405 605 8435 635
rect 8485 605 8515 635
rect 8565 605 8595 635
rect 8645 605 8675 635
rect 8725 605 8755 635
rect 8805 605 8835 635
rect 8885 605 8915 635
rect 8965 605 8995 635
rect 9045 605 9075 635
rect 9125 605 9155 635
rect 9205 605 9235 635
rect 9285 605 9315 635
rect 9365 605 9395 635
rect 9445 605 9475 635
rect 9525 605 9555 635
rect 9605 605 9635 635
rect 9685 605 9715 635
rect 9765 605 9795 635
rect 9845 605 9875 635
rect 9925 605 9955 635
rect 10005 605 10035 635
rect 10085 605 10115 635
rect 10165 605 10195 635
rect 10245 605 10275 635
rect 10325 605 10355 635
rect 10405 605 10435 635
rect 10485 605 10515 635
rect 10645 605 10675 635
rect 10805 605 10835 635
rect 10965 605 10995 635
rect -715 525 -685 555
rect -555 525 -525 555
rect -395 525 -365 555
rect -315 525 -285 555
rect -235 525 -205 555
rect -155 525 -125 555
rect -75 525 -45 555
rect 5 525 35 555
rect 85 525 115 555
rect 165 525 195 555
rect 245 525 275 555
rect 325 525 355 555
rect 405 525 435 555
rect 485 525 515 555
rect 565 525 595 555
rect 645 525 675 555
rect 725 525 755 555
rect 805 525 835 555
rect 885 525 915 555
rect 965 525 995 555
rect 1045 525 1075 555
rect 1125 525 1155 555
rect 1205 525 1235 555
rect 1285 525 1315 555
rect 1365 525 1395 555
rect 1445 525 1475 555
rect 1525 525 1555 555
rect 1605 525 1635 555
rect 1685 525 1715 555
rect 1765 525 1795 555
rect 1845 525 1875 555
rect 1925 525 1955 555
rect 2005 525 2035 555
rect 2085 525 2115 555
rect 2165 525 2195 555
rect 2245 525 2275 555
rect 2325 525 2355 555
rect 2405 525 2435 555
rect 2485 525 2515 555
rect 2565 525 2595 555
rect 2645 525 2675 555
rect 2725 525 2755 555
rect 2805 525 2835 555
rect 2885 525 2915 555
rect 2965 525 2995 555
rect 3045 525 3075 555
rect 3125 525 3155 555
rect 3205 525 3235 555
rect 3285 525 3315 555
rect 3365 525 3395 555
rect 3445 525 3475 555
rect 3525 525 3555 555
rect 3605 525 3635 555
rect 3685 525 3715 555
rect 3765 525 3795 555
rect 3845 525 3875 555
rect 3925 525 3955 555
rect 4005 525 4035 555
rect 4085 525 4115 555
rect 4165 525 4195 555
rect 4245 525 4275 555
rect 4325 525 4355 555
rect 4405 525 4435 555
rect 4485 525 4515 555
rect 4565 525 4595 555
rect 4645 525 4675 555
rect 4725 525 4755 555
rect 4805 525 4835 555
rect 4885 525 4915 555
rect 4965 525 4995 555
rect 5045 525 5075 555
rect 5125 525 5155 555
rect 5205 525 5235 555
rect 5285 525 5315 555
rect 5365 525 5395 555
rect 5445 525 5475 555
rect 5525 525 5555 555
rect 5605 525 5635 555
rect 5685 525 5715 555
rect 5765 525 5795 555
rect 5845 525 5875 555
rect 5925 525 5955 555
rect 6005 525 6035 555
rect 6085 525 6115 555
rect 6165 525 6195 555
rect 6245 525 6275 555
rect 6325 525 6355 555
rect 6405 525 6435 555
rect 6485 525 6515 555
rect 6565 525 6595 555
rect 6645 525 6675 555
rect 6725 525 6755 555
rect 6805 525 6835 555
rect 6885 525 6915 555
rect 6965 525 6995 555
rect 7045 525 7075 555
rect 7125 525 7155 555
rect 7205 525 7235 555
rect 7285 525 7315 555
rect 7365 525 7395 555
rect 7445 525 7475 555
rect 7525 525 7555 555
rect 7605 525 7635 555
rect 7685 525 7715 555
rect 7765 525 7795 555
rect 7845 525 7875 555
rect 7925 525 7955 555
rect 8005 525 8035 555
rect 8085 525 8115 555
rect 8165 525 8195 555
rect 8245 525 8275 555
rect 8325 525 8355 555
rect 8405 525 8435 555
rect 8485 525 8515 555
rect 8565 525 8595 555
rect 8645 525 8675 555
rect 8725 525 8755 555
rect 8805 525 8835 555
rect 8885 525 8915 555
rect 8965 525 8995 555
rect 9045 525 9075 555
rect 9125 525 9155 555
rect 9205 525 9235 555
rect 9285 525 9315 555
rect 9365 525 9395 555
rect 9445 525 9475 555
rect 9525 525 9555 555
rect 9605 525 9635 555
rect 9685 525 9715 555
rect 9765 525 9795 555
rect 9845 525 9875 555
rect 9925 525 9955 555
rect 10005 525 10035 555
rect 10085 525 10115 555
rect 10165 525 10195 555
rect 10245 525 10275 555
rect 10325 525 10355 555
rect 10405 525 10435 555
rect 10485 525 10515 555
rect 10645 525 10675 555
rect 10805 525 10835 555
rect 10965 525 10995 555
rect -715 445 -685 475
rect -555 445 -525 475
rect -475 445 -445 475
rect 10645 445 10675 475
rect 10805 445 10835 475
rect 10965 445 10995 475
rect -715 365 -685 395
rect -555 365 -525 395
rect -395 365 -365 395
rect -315 365 -285 395
rect -235 365 -205 395
rect -155 365 -125 395
rect -75 365 -45 395
rect 5 365 35 395
rect 85 365 115 395
rect 165 365 195 395
rect 245 365 275 395
rect 325 365 355 395
rect 405 365 435 395
rect 485 365 515 395
rect 565 365 595 395
rect 645 365 675 395
rect 725 365 755 395
rect 805 365 835 395
rect 885 365 915 395
rect 965 365 995 395
rect 1045 365 1075 395
rect 1125 365 1155 395
rect 1205 365 1235 395
rect 1285 365 1315 395
rect 1365 365 1395 395
rect 1445 365 1475 395
rect 1525 365 1555 395
rect 1605 365 1635 395
rect 1685 365 1715 395
rect 1765 365 1795 395
rect 1845 365 1875 395
rect 1925 365 1955 395
rect 2005 365 2035 395
rect 2085 365 2115 395
rect 2165 365 2195 395
rect 2245 365 2275 395
rect 2325 365 2355 395
rect 2405 365 2435 395
rect 2485 365 2515 395
rect 2565 365 2595 395
rect 2645 365 2675 395
rect 2725 365 2755 395
rect 2805 365 2835 395
rect 2885 365 2915 395
rect 2965 365 2995 395
rect 3045 365 3075 395
rect 3125 365 3155 395
rect 3205 365 3235 395
rect 3285 365 3315 395
rect 3365 365 3395 395
rect 3445 365 3475 395
rect 3525 365 3555 395
rect 3605 365 3635 395
rect 3685 365 3715 395
rect 3765 365 3795 395
rect 3845 365 3875 395
rect 3925 365 3955 395
rect 4005 365 4035 395
rect 4085 365 4115 395
rect 4165 365 4195 395
rect 4245 365 4275 395
rect 4325 365 4355 395
rect 4405 365 4435 395
rect 4485 365 4515 395
rect 4565 365 4595 395
rect 4645 365 4675 395
rect 4725 365 4755 395
rect 4805 365 4835 395
rect 4885 365 4915 395
rect 4965 365 4995 395
rect 5045 365 5075 395
rect 5125 365 5155 395
rect 5205 365 5235 395
rect 5285 365 5315 395
rect 5365 365 5395 395
rect 5445 365 5475 395
rect 5525 365 5555 395
rect 5605 365 5635 395
rect 5685 365 5715 395
rect 5765 365 5795 395
rect 5845 365 5875 395
rect 5925 365 5955 395
rect 6005 365 6035 395
rect 6085 365 6115 395
rect 6165 365 6195 395
rect 6245 365 6275 395
rect 6325 365 6355 395
rect 6405 365 6435 395
rect 6485 365 6515 395
rect 6565 365 6595 395
rect 6645 365 6675 395
rect 6725 365 6755 395
rect 6805 365 6835 395
rect 6885 365 6915 395
rect 6965 365 6995 395
rect 7045 365 7075 395
rect 7125 365 7155 395
rect 7205 365 7235 395
rect 7285 365 7315 395
rect 7365 365 7395 395
rect 7445 365 7475 395
rect 7525 365 7555 395
rect 7605 365 7635 395
rect 7685 365 7715 395
rect 7765 365 7795 395
rect 7845 365 7875 395
rect 7925 365 7955 395
rect 8005 365 8035 395
rect 8085 365 8115 395
rect 8165 365 8195 395
rect 8245 365 8275 395
rect 8325 365 8355 395
rect 8405 365 8435 395
rect 8485 365 8515 395
rect 8565 365 8595 395
rect 8645 365 8675 395
rect 8725 365 8755 395
rect 8805 365 8835 395
rect 8885 365 8915 395
rect 8965 365 8995 395
rect 9045 365 9075 395
rect 9125 365 9155 395
rect 9205 365 9235 395
rect 9285 365 9315 395
rect 9365 365 9395 395
rect 9445 365 9475 395
rect 9525 365 9555 395
rect 9605 365 9635 395
rect 9685 365 9715 395
rect 9765 365 9795 395
rect 9845 365 9875 395
rect 9925 365 9955 395
rect 10005 365 10035 395
rect 10085 365 10115 395
rect 10165 365 10195 395
rect 10245 365 10275 395
rect 10325 365 10355 395
rect 10405 365 10435 395
rect 10485 365 10515 395
rect 10645 365 10675 395
rect 10805 365 10835 395
rect 10965 365 10995 395
rect -715 285 -685 315
rect -555 285 -525 315
rect -395 285 -365 315
rect 10885 285 10915 315
rect -715 205 -685 235
rect -555 205 -525 235
rect -395 205 -365 235
rect -315 205 -285 235
rect -235 205 -205 235
rect -155 205 -125 235
rect -75 205 -45 235
rect 5 205 35 235
rect 85 205 115 235
rect 165 205 195 235
rect 245 205 275 235
rect 325 205 355 235
rect 405 205 435 235
rect 485 205 515 235
rect 565 205 595 235
rect 645 205 675 235
rect 725 205 755 235
rect 805 205 835 235
rect 885 205 915 235
rect 965 205 995 235
rect 1045 205 1075 235
rect 1125 205 1155 235
rect 1205 205 1235 235
rect 1285 205 1315 235
rect 1365 205 1395 235
rect 1445 205 1475 235
rect 1525 205 1555 235
rect 1605 205 1635 235
rect 1685 205 1715 235
rect 1765 205 1795 235
rect 1845 205 1875 235
rect 1925 205 1955 235
rect 2005 205 2035 235
rect 2085 205 2115 235
rect 2165 205 2195 235
rect 2245 205 2275 235
rect 2325 205 2355 235
rect 2405 205 2435 235
rect 2485 205 2515 235
rect 2565 205 2595 235
rect 2645 205 2675 235
rect 2725 205 2755 235
rect 2805 205 2835 235
rect 2885 205 2915 235
rect 2965 205 2995 235
rect 3045 205 3075 235
rect 3125 205 3155 235
rect 3205 205 3235 235
rect 3285 205 3315 235
rect 3365 205 3395 235
rect 3445 205 3475 235
rect 3525 205 3555 235
rect 3605 205 3635 235
rect 3685 205 3715 235
rect 3765 205 3795 235
rect 3845 205 3875 235
rect 3925 205 3955 235
rect 4005 205 4035 235
rect 4085 205 4115 235
rect 4165 205 4195 235
rect 4245 205 4275 235
rect 4325 205 4355 235
rect 4405 205 4435 235
rect 4485 205 4515 235
rect 4565 205 4595 235
rect 4645 205 4675 235
rect 4725 205 4755 235
rect 4805 205 4835 235
rect 4885 205 4915 235
rect 4965 205 4995 235
rect 5045 205 5075 235
rect 5125 205 5155 235
rect 5205 205 5235 235
rect 5285 205 5315 235
rect 5365 205 5395 235
rect 5445 205 5475 235
rect 5525 205 5555 235
rect 5605 205 5635 235
rect 5685 205 5715 235
rect 5765 205 5795 235
rect 5845 205 5875 235
rect 5925 205 5955 235
rect 6005 205 6035 235
rect 6085 205 6115 235
rect 6165 205 6195 235
rect 6245 205 6275 235
rect 6325 205 6355 235
rect 6405 205 6435 235
rect 6485 205 6515 235
rect 6565 205 6595 235
rect 6645 205 6675 235
rect 6725 205 6755 235
rect 6805 205 6835 235
rect 6885 205 6915 235
rect 6965 205 6995 235
rect 7045 205 7075 235
rect 7125 205 7155 235
rect 7205 205 7235 235
rect 7285 205 7315 235
rect 7365 205 7395 235
rect 7445 205 7475 235
rect 7525 205 7555 235
rect 7605 205 7635 235
rect 7685 205 7715 235
rect 7765 205 7795 235
rect 7845 205 7875 235
rect 7925 205 7955 235
rect 8005 205 8035 235
rect 8085 205 8115 235
rect 8165 205 8195 235
rect 8245 205 8275 235
rect 8325 205 8355 235
rect 8405 205 8435 235
rect 8485 205 8515 235
rect 8565 205 8595 235
rect 8645 205 8675 235
rect 8725 205 8755 235
rect 8805 205 8835 235
rect 8885 205 8915 235
rect 8965 205 8995 235
rect 9045 205 9075 235
rect 9125 205 9155 235
rect 9205 205 9235 235
rect 9285 205 9315 235
rect 9365 205 9395 235
rect 9445 205 9475 235
rect 9525 205 9555 235
rect 9605 205 9635 235
rect 9685 205 9715 235
rect 9765 205 9795 235
rect 9845 205 9875 235
rect 9925 205 9955 235
rect 10005 205 10035 235
rect 10085 205 10115 235
rect 10165 205 10195 235
rect 10245 205 10275 235
rect 10325 205 10355 235
rect 10405 205 10435 235
rect 10485 205 10515 235
rect 10645 205 10675 235
rect 10805 205 10835 235
rect 10965 205 10995 235
rect -715 125 -685 155
rect -555 125 -525 155
rect -395 125 -365 155
rect 10725 125 10755 155
rect 10805 125 10835 155
rect 10965 125 10995 155
rect -715 45 -685 75
rect -555 45 -525 75
rect -395 45 -365 75
rect -315 45 -285 75
rect -235 45 -205 75
rect -155 45 -125 75
rect -75 45 -45 75
rect 5 45 35 75
rect 85 45 115 75
rect 165 45 195 75
rect 245 45 275 75
rect 325 45 355 75
rect 405 45 435 75
rect 485 45 515 75
rect 565 45 595 75
rect 645 45 675 75
rect 725 45 755 75
rect 805 45 835 75
rect 885 45 915 75
rect 965 45 995 75
rect 1045 45 1075 75
rect 1125 45 1155 75
rect 1205 45 1235 75
rect 1285 45 1315 75
rect 1365 45 1395 75
rect 1445 45 1475 75
rect 1525 45 1555 75
rect 1605 45 1635 75
rect 1685 45 1715 75
rect 1765 45 1795 75
rect 1845 45 1875 75
rect 1925 45 1955 75
rect 2005 45 2035 75
rect 2085 45 2115 75
rect 2165 45 2195 75
rect 2245 45 2275 75
rect 2325 45 2355 75
rect 2405 45 2435 75
rect 2485 45 2515 75
rect 2565 45 2595 75
rect 2645 45 2675 75
rect 2725 45 2755 75
rect 2805 45 2835 75
rect 2885 45 2915 75
rect 2965 45 2995 75
rect 3045 45 3075 75
rect 3125 45 3155 75
rect 3205 45 3235 75
rect 3285 45 3315 75
rect 3365 45 3395 75
rect 3445 45 3475 75
rect 3525 45 3555 75
rect 3605 45 3635 75
rect 3685 45 3715 75
rect 3765 45 3795 75
rect 3845 45 3875 75
rect 3925 45 3955 75
rect 4005 45 4035 75
rect 4085 45 4115 75
rect 4165 45 4195 75
rect 4245 45 4275 75
rect 4325 45 4355 75
rect 4405 45 4435 75
rect 4485 45 4515 75
rect 4565 45 4595 75
rect 4645 45 4675 75
rect 4725 45 4755 75
rect 4805 45 4835 75
rect 4885 45 4915 75
rect 4965 45 4995 75
rect 5045 45 5075 75
rect 5125 45 5155 75
rect 5205 45 5235 75
rect 5285 45 5315 75
rect 5365 45 5395 75
rect 5445 45 5475 75
rect 5525 45 5555 75
rect 5605 45 5635 75
rect 5685 45 5715 75
rect 5765 45 5795 75
rect 5845 45 5875 75
rect 5925 45 5955 75
rect 6005 45 6035 75
rect 6085 45 6115 75
rect 6165 45 6195 75
rect 6245 45 6275 75
rect 6325 45 6355 75
rect 6405 45 6435 75
rect 6485 45 6515 75
rect 6565 45 6595 75
rect 6645 45 6675 75
rect 6725 45 6755 75
rect 6805 45 6835 75
rect 6885 45 6915 75
rect 6965 45 6995 75
rect 7045 45 7075 75
rect 7125 45 7155 75
rect 7205 45 7235 75
rect 7285 45 7315 75
rect 7365 45 7395 75
rect 7445 45 7475 75
rect 7525 45 7555 75
rect 7605 45 7635 75
rect 7685 45 7715 75
rect 7765 45 7795 75
rect 7845 45 7875 75
rect 7925 45 7955 75
rect 8005 45 8035 75
rect 8085 45 8115 75
rect 8165 45 8195 75
rect 8245 45 8275 75
rect 8325 45 8355 75
rect 8405 45 8435 75
rect 8485 45 8515 75
rect 8565 45 8595 75
rect 8645 45 8675 75
rect 8725 45 8755 75
rect 8805 45 8835 75
rect 8885 45 8915 75
rect 8965 45 8995 75
rect 9045 45 9075 75
rect 9125 45 9155 75
rect 9205 45 9235 75
rect 9285 45 9315 75
rect 9365 45 9395 75
rect 9445 45 9475 75
rect 9525 45 9555 75
rect 9605 45 9635 75
rect 9685 45 9715 75
rect 9765 45 9795 75
rect 9845 45 9875 75
rect 9925 45 9955 75
rect 10005 45 10035 75
rect 10085 45 10115 75
rect 10165 45 10195 75
rect 10245 45 10275 75
rect 10325 45 10355 75
rect 10405 45 10435 75
rect 10485 45 10515 75
rect 10645 45 10675 75
rect 10805 45 10835 75
rect 10965 45 10995 75
rect -715 -35 -685 -5
rect -555 -35 -525 -5
rect -395 -35 -365 -5
rect -315 -35 -285 -5
rect -235 -35 -205 -5
rect -155 -35 -125 -5
rect -75 -35 -45 -5
rect 5 -35 35 -5
rect 85 -35 115 -5
rect 165 -35 195 -5
rect 245 -35 275 -5
rect 325 -35 355 -5
rect 405 -35 435 -5
rect 485 -35 515 -5
rect 565 -35 595 -5
rect 645 -35 675 -5
rect 725 -35 755 -5
rect 805 -35 835 -5
rect 885 -35 915 -5
rect 965 -35 995 -5
rect 1045 -35 1075 -5
rect 1125 -35 1155 -5
rect 1205 -35 1235 -5
rect 1285 -35 1315 -5
rect 1365 -35 1395 -5
rect 1445 -35 1475 -5
rect 1525 -35 1555 -5
rect 1605 -35 1635 -5
rect 1685 -35 1715 -5
rect 1765 -35 1795 -5
rect 1845 -35 1875 -5
rect 1925 -35 1955 -5
rect 2005 -35 2035 -5
rect 2085 -35 2115 -5
rect 2165 -35 2195 -5
rect 2245 -35 2275 -5
rect 2325 -35 2355 -5
rect 2405 -35 2435 -5
rect 2485 -35 2515 -5
rect 2565 -35 2595 -5
rect 2645 -35 2675 -5
rect 2725 -35 2755 -5
rect 2805 -35 2835 -5
rect 2885 -35 2915 -5
rect 2965 -35 2995 -5
rect 3045 -35 3075 -5
rect 3125 -35 3155 -5
rect 3205 -35 3235 -5
rect 3285 -35 3315 -5
rect 3365 -35 3395 -5
rect 3445 -35 3475 -5
rect 3525 -35 3555 -5
rect 3605 -35 3635 -5
rect 3685 -35 3715 -5
rect 3765 -35 3795 -5
rect 3845 -35 3875 -5
rect 3925 -35 3955 -5
rect 4005 -35 4035 -5
rect 4085 -35 4115 -5
rect 4165 -35 4195 -5
rect 4245 -35 4275 -5
rect 4325 -35 4355 -5
rect 4405 -35 4435 -5
rect 4485 -35 4515 -5
rect 4565 -35 4595 -5
rect 4645 -35 4675 -5
rect 4725 -35 4755 -5
rect 4805 -35 4835 -5
rect 4885 -35 4915 -5
rect 4965 -35 4995 -5
rect 5045 -35 5075 -5
rect 5125 -35 5155 -5
rect 5205 -35 5235 -5
rect 5285 -35 5315 -5
rect 5365 -35 5395 -5
rect 5445 -35 5475 -5
rect 5525 -35 5555 -5
rect 5605 -35 5635 -5
rect 5685 -35 5715 -5
rect 5765 -35 5795 -5
rect 5845 -35 5875 -5
rect 5925 -35 5955 -5
rect 6005 -35 6035 -5
rect 6085 -35 6115 -5
rect 6165 -35 6195 -5
rect 6245 -35 6275 -5
rect 6325 -35 6355 -5
rect 6405 -35 6435 -5
rect 6485 -35 6515 -5
rect 6565 -35 6595 -5
rect 6645 -35 6675 -5
rect 6725 -35 6755 -5
rect 6805 -35 6835 -5
rect 6885 -35 6915 -5
rect 6965 -35 6995 -5
rect 7045 -35 7075 -5
rect 7125 -35 7155 -5
rect 7205 -35 7235 -5
rect 7285 -35 7315 -5
rect 7365 -35 7395 -5
rect 7445 -35 7475 -5
rect 7525 -35 7555 -5
rect 7605 -35 7635 -5
rect 7685 -35 7715 -5
rect 7765 -35 7795 -5
rect 7845 -35 7875 -5
rect 7925 -35 7955 -5
rect 8005 -35 8035 -5
rect 8085 -35 8115 -5
rect 8165 -35 8195 -5
rect 8245 -35 8275 -5
rect 8325 -35 8355 -5
rect 8405 -35 8435 -5
rect 8485 -35 8515 -5
rect 8565 -35 8595 -5
rect 8645 -35 8675 -5
rect 8725 -35 8755 -5
rect 8805 -35 8835 -5
rect 8885 -35 8915 -5
rect 8965 -35 8995 -5
rect 9045 -35 9075 -5
rect 9125 -35 9155 -5
rect 9205 -35 9235 -5
rect 9285 -35 9315 -5
rect 9365 -35 9395 -5
rect 9445 -35 9475 -5
rect 9525 -35 9555 -5
rect 9605 -35 9635 -5
rect 9685 -35 9715 -5
rect 9765 -35 9795 -5
rect 9845 -35 9875 -5
rect 9925 -35 9955 -5
rect 10005 -35 10035 -5
rect 10085 -35 10115 -5
rect 10165 -35 10195 -5
rect 10245 -35 10275 -5
rect 10325 -35 10355 -5
rect 10405 -35 10435 -5
rect 10485 -35 10515 -5
rect 10645 -35 10675 -5
rect 10805 -35 10835 -5
rect 10965 -35 10995 -5
rect -715 -115 -685 -85
rect -555 -115 -525 -85
rect -395 -115 -365 -85
rect -315 -115 -285 -85
rect -235 -115 -205 -85
rect -155 -115 -125 -85
rect -75 -115 -45 -85
rect 5 -115 35 -85
rect 85 -115 115 -85
rect 165 -115 195 -85
rect 245 -115 275 -85
rect 325 -115 355 -85
rect 405 -115 435 -85
rect 485 -115 515 -85
rect 565 -115 595 -85
rect 645 -115 675 -85
rect 725 -115 755 -85
rect 805 -115 835 -85
rect 885 -115 915 -85
rect 965 -115 995 -85
rect 1045 -115 1075 -85
rect 1125 -115 1155 -85
rect 1205 -115 1235 -85
rect 1285 -115 1315 -85
rect 1365 -115 1395 -85
rect 1445 -115 1475 -85
rect 1525 -115 1555 -85
rect 1605 -115 1635 -85
rect 1685 -115 1715 -85
rect 1765 -115 1795 -85
rect 1845 -115 1875 -85
rect 1925 -115 1955 -85
rect 2005 -115 2035 -85
rect 2085 -115 2115 -85
rect 2165 -115 2195 -85
rect 2245 -115 2275 -85
rect 2325 -115 2355 -85
rect 2405 -115 2435 -85
rect 2485 -115 2515 -85
rect 2565 -115 2595 -85
rect 2645 -115 2675 -85
rect 2725 -115 2755 -85
rect 2805 -115 2835 -85
rect 2885 -115 2915 -85
rect 2965 -115 2995 -85
rect 3045 -115 3075 -85
rect 3125 -115 3155 -85
rect 3205 -115 3235 -85
rect 3285 -115 3315 -85
rect 3365 -115 3395 -85
rect 3445 -115 3475 -85
rect 3525 -115 3555 -85
rect 3605 -115 3635 -85
rect 3685 -115 3715 -85
rect 3765 -115 3795 -85
rect 3845 -115 3875 -85
rect 3925 -115 3955 -85
rect 4005 -115 4035 -85
rect 4085 -115 4115 -85
rect 4165 -115 4195 -85
rect 4245 -115 4275 -85
rect 4325 -115 4355 -85
rect 4405 -115 4435 -85
rect 4485 -115 4515 -85
rect 4565 -115 4595 -85
rect 4645 -115 4675 -85
rect 4725 -115 4755 -85
rect 4805 -115 4835 -85
rect 4885 -115 4915 -85
rect 4965 -115 4995 -85
rect 5045 -115 5075 -85
rect 5125 -115 5155 -85
rect 5205 -115 5235 -85
rect 5285 -115 5315 -85
rect 5365 -115 5395 -85
rect 5445 -115 5475 -85
rect 5525 -115 5555 -85
rect 5605 -115 5635 -85
rect 5685 -115 5715 -85
rect 5765 -115 5795 -85
rect 5845 -115 5875 -85
rect 5925 -115 5955 -85
rect 6005 -115 6035 -85
rect 6085 -115 6115 -85
rect 6165 -115 6195 -85
rect 6245 -115 6275 -85
rect 6325 -115 6355 -85
rect 6405 -115 6435 -85
rect 6485 -115 6515 -85
rect 6565 -115 6595 -85
rect 6645 -115 6675 -85
rect 6725 -115 6755 -85
rect 6805 -115 6835 -85
rect 6885 -115 6915 -85
rect 6965 -115 6995 -85
rect 7045 -115 7075 -85
rect 7125 -115 7155 -85
rect 7205 -115 7235 -85
rect 7285 -115 7315 -85
rect 7365 -115 7395 -85
rect 7445 -115 7475 -85
rect 7525 -115 7555 -85
rect 7605 -115 7635 -85
rect 7685 -115 7715 -85
rect 7765 -115 7795 -85
rect 7845 -115 7875 -85
rect 7925 -115 7955 -85
rect 8005 -115 8035 -85
rect 8085 -115 8115 -85
rect 8165 -115 8195 -85
rect 8245 -115 8275 -85
rect 8325 -115 8355 -85
rect 8405 -115 8435 -85
rect 8485 -115 8515 -85
rect 8565 -115 8595 -85
rect 8645 -115 8675 -85
rect 8725 -115 8755 -85
rect 8805 -115 8835 -85
rect 8885 -115 8915 -85
rect 8965 -115 8995 -85
rect 9045 -115 9075 -85
rect 9125 -115 9155 -85
rect 9205 -115 9235 -85
rect 9285 -115 9315 -85
rect 9365 -115 9395 -85
rect 9445 -115 9475 -85
rect 9525 -115 9555 -85
rect 9605 -115 9635 -85
rect 9685 -115 9715 -85
rect 9765 -115 9795 -85
rect 9845 -115 9875 -85
rect 9925 -115 9955 -85
rect 10005 -115 10035 -85
rect 10085 -115 10115 -85
rect 10165 -115 10195 -85
rect 10245 -115 10275 -85
rect 10325 -115 10355 -85
rect 10405 -115 10435 -85
rect 10485 -115 10515 -85
rect 10645 -115 10675 -85
rect 10805 -115 10835 -85
rect 10965 -115 10995 -85
<< metal3 >>
rect -720 1036 -680 1040
rect -720 1004 -716 1036
rect -684 1004 -680 1036
rect -720 956 -680 1004
rect -720 924 -716 956
rect -684 924 -680 956
rect -720 876 -680 924
rect -720 844 -716 876
rect -684 844 -680 876
rect -720 796 -680 844
rect -720 764 -716 796
rect -684 764 -680 796
rect -720 716 -680 764
rect -720 684 -716 716
rect -684 684 -680 716
rect -720 636 -680 684
rect -720 604 -716 636
rect -684 604 -680 636
rect -720 556 -680 604
rect -720 524 -716 556
rect -684 524 -680 556
rect -720 476 -680 524
rect -720 444 -716 476
rect -684 444 -680 476
rect -720 396 -680 444
rect -720 364 -716 396
rect -684 364 -680 396
rect -720 316 -680 364
rect -720 284 -716 316
rect -684 284 -680 316
rect -720 236 -680 284
rect -720 204 -716 236
rect -684 204 -680 236
rect -720 156 -680 204
rect -720 124 -716 156
rect -684 124 -680 156
rect -720 76 -680 124
rect -720 44 -716 76
rect -684 44 -680 76
rect -720 -4 -680 44
rect -720 -36 -716 -4
rect -684 -36 -680 -4
rect -720 -84 -680 -36
rect -720 -116 -716 -84
rect -684 -116 -680 -84
rect -720 -120 -680 -116
rect -640 795 -600 1080
rect -640 765 -635 795
rect -605 765 -600 795
rect -640 715 -600 765
rect -640 685 -635 715
rect -605 685 -600 715
rect -640 -120 -600 685
rect -560 1036 -520 1040
rect -560 1004 -556 1036
rect -524 1004 -520 1036
rect -560 956 -520 1004
rect -560 924 -556 956
rect -524 924 -520 956
rect -560 876 -520 924
rect -560 844 -556 876
rect -524 844 -520 876
rect -560 796 -520 844
rect -560 764 -556 796
rect -524 764 -520 796
rect -560 716 -520 764
rect -560 684 -556 716
rect -524 684 -520 716
rect -560 636 -520 684
rect -560 604 -556 636
rect -524 604 -520 636
rect -560 556 -520 604
rect -560 524 -556 556
rect -524 524 -520 556
rect -560 476 -520 524
rect -560 444 -556 476
rect -524 444 -520 476
rect -560 396 -520 444
rect -560 364 -556 396
rect -524 364 -520 396
rect -560 316 -520 364
rect -560 284 -556 316
rect -524 284 -520 316
rect -560 236 -520 284
rect -560 204 -556 236
rect -524 204 -520 236
rect -560 156 -520 204
rect -560 124 -556 156
rect -524 124 -520 156
rect -560 76 -520 124
rect -560 44 -556 76
rect -524 44 -520 76
rect -560 -4 -520 44
rect -560 -36 -556 -4
rect -524 -36 -520 -4
rect -560 -84 -520 -36
rect -560 -116 -556 -84
rect -524 -116 -520 -84
rect -560 -120 -520 -116
rect -480 475 -440 1080
rect -480 445 -475 475
rect -445 445 -440 475
rect -480 -120 -440 445
rect -400 1036 -360 1040
rect -400 1004 -396 1036
rect -364 1004 -360 1036
rect -400 956 -360 1004
rect -400 924 -396 956
rect -364 924 -360 956
rect -400 876 -360 924
rect -400 844 -396 876
rect -364 844 -360 876
rect -400 796 -360 844
rect -400 764 -396 796
rect -364 764 -360 796
rect -400 716 -360 764
rect -400 684 -396 716
rect -364 684 -360 716
rect -400 636 -360 684
rect -400 604 -396 636
rect -364 604 -360 636
rect -400 556 -360 604
rect -400 524 -396 556
rect -364 524 -360 556
rect -400 476 -360 524
rect -400 444 -396 476
rect -364 444 -360 476
rect -400 396 -360 444
rect -400 364 -396 396
rect -364 364 -360 396
rect -400 316 -360 364
rect -400 284 -396 316
rect -364 284 -360 316
rect -400 236 -360 284
rect -400 204 -396 236
rect -364 204 -360 236
rect -400 156 -360 204
rect -400 124 -396 156
rect -364 124 -360 156
rect -400 76 -360 124
rect -400 44 -396 76
rect -364 44 -360 76
rect -400 -4 -360 44
rect -400 -36 -396 -4
rect -364 -36 -360 -4
rect -400 -84 -360 -36
rect -400 -116 -396 -84
rect -364 -116 -360 -84
rect -400 -120 -360 -116
rect -320 1036 -280 1040
rect -320 1004 -316 1036
rect -284 1004 -280 1036
rect -320 956 -280 1004
rect -320 924 -316 956
rect -284 924 -280 956
rect -320 876 -280 924
rect -320 844 -316 876
rect -284 844 -280 876
rect -320 796 -280 844
rect -320 764 -316 796
rect -284 764 -280 796
rect -320 716 -280 764
rect -320 684 -316 716
rect -284 684 -280 716
rect -320 636 -280 684
rect -320 604 -316 636
rect -284 604 -280 636
rect -320 556 -280 604
rect -320 524 -316 556
rect -284 524 -280 556
rect -320 476 -280 524
rect -320 444 -316 476
rect -284 444 -280 476
rect -320 396 -280 444
rect -320 364 -316 396
rect -284 364 -280 396
rect -320 316 -280 364
rect -320 284 -316 316
rect -284 284 -280 316
rect -320 236 -280 284
rect -320 204 -316 236
rect -284 204 -280 236
rect -320 156 -280 204
rect -320 124 -316 156
rect -284 124 -280 156
rect -320 76 -280 124
rect -320 44 -316 76
rect -284 44 -280 76
rect -320 -4 -280 44
rect -320 -36 -316 -4
rect -284 -36 -280 -4
rect -320 -84 -280 -36
rect -320 -116 -316 -84
rect -284 -116 -280 -84
rect -320 -120 -280 -116
rect -240 1036 -200 1040
rect -240 1004 -236 1036
rect -204 1004 -200 1036
rect -240 956 -200 1004
rect -240 924 -236 956
rect -204 924 -200 956
rect -240 876 -200 924
rect -240 844 -236 876
rect -204 844 -200 876
rect -240 796 -200 844
rect -240 764 -236 796
rect -204 764 -200 796
rect -240 716 -200 764
rect -240 684 -236 716
rect -204 684 -200 716
rect -240 636 -200 684
rect -240 604 -236 636
rect -204 604 -200 636
rect -240 556 -200 604
rect -240 524 -236 556
rect -204 524 -200 556
rect -240 476 -200 524
rect -240 444 -236 476
rect -204 444 -200 476
rect -240 396 -200 444
rect -240 364 -236 396
rect -204 364 -200 396
rect -240 316 -200 364
rect -240 284 -236 316
rect -204 284 -200 316
rect -240 236 -200 284
rect -240 204 -236 236
rect -204 204 -200 236
rect -240 156 -200 204
rect -240 124 -236 156
rect -204 124 -200 156
rect -240 76 -200 124
rect -240 44 -236 76
rect -204 44 -200 76
rect -240 -4 -200 44
rect -240 -36 -236 -4
rect -204 -36 -200 -4
rect -240 -84 -200 -36
rect -240 -116 -236 -84
rect -204 -116 -200 -84
rect -240 -120 -200 -116
rect -160 1036 -120 1040
rect -160 1004 -156 1036
rect -124 1004 -120 1036
rect -160 956 -120 1004
rect -160 924 -156 956
rect -124 924 -120 956
rect -160 876 -120 924
rect -160 844 -156 876
rect -124 844 -120 876
rect -160 796 -120 844
rect -160 764 -156 796
rect -124 764 -120 796
rect -160 716 -120 764
rect -160 684 -156 716
rect -124 684 -120 716
rect -160 636 -120 684
rect -160 604 -156 636
rect -124 604 -120 636
rect -160 556 -120 604
rect -160 524 -156 556
rect -124 524 -120 556
rect -160 476 -120 524
rect -160 444 -156 476
rect -124 444 -120 476
rect -160 396 -120 444
rect -160 364 -156 396
rect -124 364 -120 396
rect -160 316 -120 364
rect -160 284 -156 316
rect -124 284 -120 316
rect -160 236 -120 284
rect -160 204 -156 236
rect -124 204 -120 236
rect -160 156 -120 204
rect -160 124 -156 156
rect -124 124 -120 156
rect -160 76 -120 124
rect -160 44 -156 76
rect -124 44 -120 76
rect -160 -4 -120 44
rect -160 -36 -156 -4
rect -124 -36 -120 -4
rect -160 -84 -120 -36
rect -160 -116 -156 -84
rect -124 -116 -120 -84
rect -160 -120 -120 -116
rect -80 1036 -40 1040
rect -80 1004 -76 1036
rect -44 1004 -40 1036
rect -80 956 -40 1004
rect -80 924 -76 956
rect -44 924 -40 956
rect -80 876 -40 924
rect -80 844 -76 876
rect -44 844 -40 876
rect -80 796 -40 844
rect -80 764 -76 796
rect -44 764 -40 796
rect -80 716 -40 764
rect -80 684 -76 716
rect -44 684 -40 716
rect -80 636 -40 684
rect -80 604 -76 636
rect -44 604 -40 636
rect -80 556 -40 604
rect -80 524 -76 556
rect -44 524 -40 556
rect -80 476 -40 524
rect -80 444 -76 476
rect -44 444 -40 476
rect -80 396 -40 444
rect -80 364 -76 396
rect -44 364 -40 396
rect -80 316 -40 364
rect -80 284 -76 316
rect -44 284 -40 316
rect -80 236 -40 284
rect -80 204 -76 236
rect -44 204 -40 236
rect -80 156 -40 204
rect -80 124 -76 156
rect -44 124 -40 156
rect -80 76 -40 124
rect -80 44 -76 76
rect -44 44 -40 76
rect -80 -4 -40 44
rect -80 -36 -76 -4
rect -44 -36 -40 -4
rect -80 -84 -40 -36
rect -80 -116 -76 -84
rect -44 -116 -40 -84
rect -80 -120 -40 -116
rect 0 1036 40 1040
rect 0 1004 4 1036
rect 36 1004 40 1036
rect 0 956 40 1004
rect 0 924 4 956
rect 36 924 40 956
rect 0 876 40 924
rect 0 844 4 876
rect 36 844 40 876
rect 0 796 40 844
rect 0 764 4 796
rect 36 764 40 796
rect 0 716 40 764
rect 0 684 4 716
rect 36 684 40 716
rect 0 636 40 684
rect 0 604 4 636
rect 36 604 40 636
rect 0 556 40 604
rect 0 524 4 556
rect 36 524 40 556
rect 0 476 40 524
rect 0 444 4 476
rect 36 444 40 476
rect 0 396 40 444
rect 0 364 4 396
rect 36 364 40 396
rect 0 316 40 364
rect 0 284 4 316
rect 36 284 40 316
rect 0 236 40 284
rect 0 204 4 236
rect 36 204 40 236
rect 0 156 40 204
rect 0 124 4 156
rect 36 124 40 156
rect 0 76 40 124
rect 0 44 4 76
rect 36 44 40 76
rect 0 -4 40 44
rect 0 -36 4 -4
rect 36 -36 40 -4
rect 0 -84 40 -36
rect 0 -116 4 -84
rect 36 -116 40 -84
rect 0 -120 40 -116
rect 80 1036 120 1040
rect 80 1004 84 1036
rect 116 1004 120 1036
rect 80 956 120 1004
rect 80 924 84 956
rect 116 924 120 956
rect 80 876 120 924
rect 80 844 84 876
rect 116 844 120 876
rect 80 796 120 844
rect 80 764 84 796
rect 116 764 120 796
rect 80 716 120 764
rect 80 684 84 716
rect 116 684 120 716
rect 80 636 120 684
rect 80 604 84 636
rect 116 604 120 636
rect 80 556 120 604
rect 80 524 84 556
rect 116 524 120 556
rect 80 476 120 524
rect 80 444 84 476
rect 116 444 120 476
rect 80 396 120 444
rect 80 364 84 396
rect 116 364 120 396
rect 80 316 120 364
rect 80 284 84 316
rect 116 284 120 316
rect 80 236 120 284
rect 80 204 84 236
rect 116 204 120 236
rect 80 156 120 204
rect 80 124 84 156
rect 116 124 120 156
rect 80 76 120 124
rect 80 44 84 76
rect 116 44 120 76
rect 80 -4 120 44
rect 80 -36 84 -4
rect 116 -36 120 -4
rect 80 -84 120 -36
rect 80 -116 84 -84
rect 116 -116 120 -84
rect 80 -120 120 -116
rect 160 1036 200 1040
rect 160 1004 164 1036
rect 196 1004 200 1036
rect 160 956 200 1004
rect 160 924 164 956
rect 196 924 200 956
rect 160 876 200 924
rect 160 844 164 876
rect 196 844 200 876
rect 160 796 200 844
rect 160 764 164 796
rect 196 764 200 796
rect 160 716 200 764
rect 160 684 164 716
rect 196 684 200 716
rect 160 636 200 684
rect 160 604 164 636
rect 196 604 200 636
rect 160 556 200 604
rect 160 524 164 556
rect 196 524 200 556
rect 160 476 200 524
rect 160 444 164 476
rect 196 444 200 476
rect 160 396 200 444
rect 160 364 164 396
rect 196 364 200 396
rect 160 316 200 364
rect 160 284 164 316
rect 196 284 200 316
rect 160 236 200 284
rect 160 204 164 236
rect 196 204 200 236
rect 160 156 200 204
rect 160 124 164 156
rect 196 124 200 156
rect 160 76 200 124
rect 160 44 164 76
rect 196 44 200 76
rect 160 -4 200 44
rect 160 -36 164 -4
rect 196 -36 200 -4
rect 160 -84 200 -36
rect 160 -116 164 -84
rect 196 -116 200 -84
rect 160 -120 200 -116
rect 240 1036 280 1040
rect 240 1004 244 1036
rect 276 1004 280 1036
rect 240 956 280 1004
rect 240 924 244 956
rect 276 924 280 956
rect 240 876 280 924
rect 240 844 244 876
rect 276 844 280 876
rect 240 796 280 844
rect 240 764 244 796
rect 276 764 280 796
rect 240 716 280 764
rect 240 684 244 716
rect 276 684 280 716
rect 240 636 280 684
rect 240 604 244 636
rect 276 604 280 636
rect 240 556 280 604
rect 240 524 244 556
rect 276 524 280 556
rect 240 476 280 524
rect 240 444 244 476
rect 276 444 280 476
rect 240 396 280 444
rect 240 364 244 396
rect 276 364 280 396
rect 240 316 280 364
rect 240 284 244 316
rect 276 284 280 316
rect 240 236 280 284
rect 240 204 244 236
rect 276 204 280 236
rect 240 156 280 204
rect 240 124 244 156
rect 276 124 280 156
rect 240 76 280 124
rect 240 44 244 76
rect 276 44 280 76
rect 240 -4 280 44
rect 240 -36 244 -4
rect 276 -36 280 -4
rect 240 -84 280 -36
rect 240 -116 244 -84
rect 276 -116 280 -84
rect 240 -120 280 -116
rect 320 1036 360 1040
rect 320 1004 324 1036
rect 356 1004 360 1036
rect 320 956 360 1004
rect 320 924 324 956
rect 356 924 360 956
rect 320 876 360 924
rect 320 844 324 876
rect 356 844 360 876
rect 320 796 360 844
rect 320 764 324 796
rect 356 764 360 796
rect 320 716 360 764
rect 320 684 324 716
rect 356 684 360 716
rect 320 636 360 684
rect 320 604 324 636
rect 356 604 360 636
rect 320 556 360 604
rect 320 524 324 556
rect 356 524 360 556
rect 320 476 360 524
rect 320 444 324 476
rect 356 444 360 476
rect 320 396 360 444
rect 320 364 324 396
rect 356 364 360 396
rect 320 316 360 364
rect 320 284 324 316
rect 356 284 360 316
rect 320 236 360 284
rect 320 204 324 236
rect 356 204 360 236
rect 320 156 360 204
rect 320 124 324 156
rect 356 124 360 156
rect 320 76 360 124
rect 320 44 324 76
rect 356 44 360 76
rect 320 -4 360 44
rect 320 -36 324 -4
rect 356 -36 360 -4
rect 320 -84 360 -36
rect 320 -116 324 -84
rect 356 -116 360 -84
rect 320 -120 360 -116
rect 400 1036 440 1040
rect 400 1004 404 1036
rect 436 1004 440 1036
rect 400 956 440 1004
rect 400 924 404 956
rect 436 924 440 956
rect 400 876 440 924
rect 400 844 404 876
rect 436 844 440 876
rect 400 796 440 844
rect 400 764 404 796
rect 436 764 440 796
rect 400 716 440 764
rect 400 684 404 716
rect 436 684 440 716
rect 400 636 440 684
rect 400 604 404 636
rect 436 604 440 636
rect 400 556 440 604
rect 400 524 404 556
rect 436 524 440 556
rect 400 476 440 524
rect 400 444 404 476
rect 436 444 440 476
rect 400 396 440 444
rect 400 364 404 396
rect 436 364 440 396
rect 400 316 440 364
rect 400 284 404 316
rect 436 284 440 316
rect 400 236 440 284
rect 400 204 404 236
rect 436 204 440 236
rect 400 156 440 204
rect 400 124 404 156
rect 436 124 440 156
rect 400 76 440 124
rect 400 44 404 76
rect 436 44 440 76
rect 400 -4 440 44
rect 400 -36 404 -4
rect 436 -36 440 -4
rect 400 -84 440 -36
rect 400 -116 404 -84
rect 436 -116 440 -84
rect 400 -120 440 -116
rect 480 1036 520 1040
rect 480 1004 484 1036
rect 516 1004 520 1036
rect 480 956 520 1004
rect 480 924 484 956
rect 516 924 520 956
rect 480 876 520 924
rect 480 844 484 876
rect 516 844 520 876
rect 480 796 520 844
rect 480 764 484 796
rect 516 764 520 796
rect 480 716 520 764
rect 480 684 484 716
rect 516 684 520 716
rect 480 636 520 684
rect 480 604 484 636
rect 516 604 520 636
rect 480 556 520 604
rect 480 524 484 556
rect 516 524 520 556
rect 480 476 520 524
rect 480 444 484 476
rect 516 444 520 476
rect 480 396 520 444
rect 480 364 484 396
rect 516 364 520 396
rect 480 316 520 364
rect 480 284 484 316
rect 516 284 520 316
rect 480 236 520 284
rect 480 204 484 236
rect 516 204 520 236
rect 480 156 520 204
rect 480 124 484 156
rect 516 124 520 156
rect 480 76 520 124
rect 480 44 484 76
rect 516 44 520 76
rect 480 -4 520 44
rect 480 -36 484 -4
rect 516 -36 520 -4
rect 480 -84 520 -36
rect 480 -116 484 -84
rect 516 -116 520 -84
rect 480 -120 520 -116
rect 560 1036 600 1040
rect 560 1004 564 1036
rect 596 1004 600 1036
rect 560 956 600 1004
rect 560 924 564 956
rect 596 924 600 956
rect 560 876 600 924
rect 560 844 564 876
rect 596 844 600 876
rect 560 796 600 844
rect 560 764 564 796
rect 596 764 600 796
rect 560 716 600 764
rect 560 684 564 716
rect 596 684 600 716
rect 560 636 600 684
rect 560 604 564 636
rect 596 604 600 636
rect 560 556 600 604
rect 560 524 564 556
rect 596 524 600 556
rect 560 476 600 524
rect 560 444 564 476
rect 596 444 600 476
rect 560 396 600 444
rect 560 364 564 396
rect 596 364 600 396
rect 560 316 600 364
rect 560 284 564 316
rect 596 284 600 316
rect 560 236 600 284
rect 560 204 564 236
rect 596 204 600 236
rect 560 156 600 204
rect 560 124 564 156
rect 596 124 600 156
rect 560 76 600 124
rect 560 44 564 76
rect 596 44 600 76
rect 560 -4 600 44
rect 560 -36 564 -4
rect 596 -36 600 -4
rect 560 -84 600 -36
rect 560 -116 564 -84
rect 596 -116 600 -84
rect 560 -120 600 -116
rect 640 1036 680 1040
rect 640 1004 644 1036
rect 676 1004 680 1036
rect 640 956 680 1004
rect 640 924 644 956
rect 676 924 680 956
rect 640 876 680 924
rect 640 844 644 876
rect 676 844 680 876
rect 640 796 680 844
rect 640 764 644 796
rect 676 764 680 796
rect 640 716 680 764
rect 640 684 644 716
rect 676 684 680 716
rect 640 636 680 684
rect 640 604 644 636
rect 676 604 680 636
rect 640 556 680 604
rect 640 524 644 556
rect 676 524 680 556
rect 640 476 680 524
rect 640 444 644 476
rect 676 444 680 476
rect 640 396 680 444
rect 640 364 644 396
rect 676 364 680 396
rect 640 316 680 364
rect 640 284 644 316
rect 676 284 680 316
rect 640 236 680 284
rect 640 204 644 236
rect 676 204 680 236
rect 640 156 680 204
rect 640 124 644 156
rect 676 124 680 156
rect 640 76 680 124
rect 640 44 644 76
rect 676 44 680 76
rect 640 -4 680 44
rect 640 -36 644 -4
rect 676 -36 680 -4
rect 640 -84 680 -36
rect 640 -116 644 -84
rect 676 -116 680 -84
rect 640 -120 680 -116
rect 720 1036 760 1040
rect 720 1004 724 1036
rect 756 1004 760 1036
rect 720 956 760 1004
rect 720 924 724 956
rect 756 924 760 956
rect 720 876 760 924
rect 720 844 724 876
rect 756 844 760 876
rect 720 796 760 844
rect 720 764 724 796
rect 756 764 760 796
rect 720 716 760 764
rect 720 684 724 716
rect 756 684 760 716
rect 720 636 760 684
rect 720 604 724 636
rect 756 604 760 636
rect 720 556 760 604
rect 720 524 724 556
rect 756 524 760 556
rect 720 476 760 524
rect 720 444 724 476
rect 756 444 760 476
rect 720 396 760 444
rect 720 364 724 396
rect 756 364 760 396
rect 720 316 760 364
rect 720 284 724 316
rect 756 284 760 316
rect 720 236 760 284
rect 720 204 724 236
rect 756 204 760 236
rect 720 156 760 204
rect 720 124 724 156
rect 756 124 760 156
rect 720 76 760 124
rect 720 44 724 76
rect 756 44 760 76
rect 720 -4 760 44
rect 720 -36 724 -4
rect 756 -36 760 -4
rect 720 -84 760 -36
rect 720 -116 724 -84
rect 756 -116 760 -84
rect 720 -120 760 -116
rect 800 1036 840 1040
rect 800 1004 804 1036
rect 836 1004 840 1036
rect 800 956 840 1004
rect 800 924 804 956
rect 836 924 840 956
rect 800 876 840 924
rect 800 844 804 876
rect 836 844 840 876
rect 800 796 840 844
rect 800 764 804 796
rect 836 764 840 796
rect 800 716 840 764
rect 800 684 804 716
rect 836 684 840 716
rect 800 636 840 684
rect 800 604 804 636
rect 836 604 840 636
rect 800 556 840 604
rect 800 524 804 556
rect 836 524 840 556
rect 800 476 840 524
rect 800 444 804 476
rect 836 444 840 476
rect 800 396 840 444
rect 800 364 804 396
rect 836 364 840 396
rect 800 316 840 364
rect 800 284 804 316
rect 836 284 840 316
rect 800 236 840 284
rect 800 204 804 236
rect 836 204 840 236
rect 800 156 840 204
rect 800 124 804 156
rect 836 124 840 156
rect 800 76 840 124
rect 800 44 804 76
rect 836 44 840 76
rect 800 -4 840 44
rect 800 -36 804 -4
rect 836 -36 840 -4
rect 800 -84 840 -36
rect 800 -116 804 -84
rect 836 -116 840 -84
rect 800 -120 840 -116
rect 880 1036 920 1040
rect 880 1004 884 1036
rect 916 1004 920 1036
rect 880 956 920 1004
rect 880 924 884 956
rect 916 924 920 956
rect 880 876 920 924
rect 880 844 884 876
rect 916 844 920 876
rect 880 796 920 844
rect 880 764 884 796
rect 916 764 920 796
rect 880 716 920 764
rect 880 684 884 716
rect 916 684 920 716
rect 880 636 920 684
rect 880 604 884 636
rect 916 604 920 636
rect 880 556 920 604
rect 880 524 884 556
rect 916 524 920 556
rect 880 476 920 524
rect 880 444 884 476
rect 916 444 920 476
rect 880 396 920 444
rect 880 364 884 396
rect 916 364 920 396
rect 880 316 920 364
rect 880 284 884 316
rect 916 284 920 316
rect 880 236 920 284
rect 880 204 884 236
rect 916 204 920 236
rect 880 156 920 204
rect 880 124 884 156
rect 916 124 920 156
rect 880 76 920 124
rect 880 44 884 76
rect 916 44 920 76
rect 880 -4 920 44
rect 880 -36 884 -4
rect 916 -36 920 -4
rect 880 -84 920 -36
rect 880 -116 884 -84
rect 916 -116 920 -84
rect 880 -120 920 -116
rect 960 1036 1000 1040
rect 960 1004 964 1036
rect 996 1004 1000 1036
rect 960 956 1000 1004
rect 960 924 964 956
rect 996 924 1000 956
rect 960 876 1000 924
rect 960 844 964 876
rect 996 844 1000 876
rect 960 796 1000 844
rect 960 764 964 796
rect 996 764 1000 796
rect 960 716 1000 764
rect 960 684 964 716
rect 996 684 1000 716
rect 960 636 1000 684
rect 960 604 964 636
rect 996 604 1000 636
rect 960 556 1000 604
rect 960 524 964 556
rect 996 524 1000 556
rect 960 476 1000 524
rect 960 444 964 476
rect 996 444 1000 476
rect 960 396 1000 444
rect 960 364 964 396
rect 996 364 1000 396
rect 960 316 1000 364
rect 960 284 964 316
rect 996 284 1000 316
rect 960 236 1000 284
rect 960 204 964 236
rect 996 204 1000 236
rect 960 156 1000 204
rect 960 124 964 156
rect 996 124 1000 156
rect 960 76 1000 124
rect 960 44 964 76
rect 996 44 1000 76
rect 960 -4 1000 44
rect 960 -36 964 -4
rect 996 -36 1000 -4
rect 960 -84 1000 -36
rect 960 -116 964 -84
rect 996 -116 1000 -84
rect 960 -120 1000 -116
rect 1040 1036 1080 1040
rect 1040 1004 1044 1036
rect 1076 1004 1080 1036
rect 1040 956 1080 1004
rect 1040 924 1044 956
rect 1076 924 1080 956
rect 1040 876 1080 924
rect 1040 844 1044 876
rect 1076 844 1080 876
rect 1040 796 1080 844
rect 1040 764 1044 796
rect 1076 764 1080 796
rect 1040 716 1080 764
rect 1040 684 1044 716
rect 1076 684 1080 716
rect 1040 636 1080 684
rect 1040 604 1044 636
rect 1076 604 1080 636
rect 1040 556 1080 604
rect 1040 524 1044 556
rect 1076 524 1080 556
rect 1040 476 1080 524
rect 1040 444 1044 476
rect 1076 444 1080 476
rect 1040 396 1080 444
rect 1040 364 1044 396
rect 1076 364 1080 396
rect 1040 316 1080 364
rect 1040 284 1044 316
rect 1076 284 1080 316
rect 1040 236 1080 284
rect 1040 204 1044 236
rect 1076 204 1080 236
rect 1040 156 1080 204
rect 1040 124 1044 156
rect 1076 124 1080 156
rect 1040 76 1080 124
rect 1040 44 1044 76
rect 1076 44 1080 76
rect 1040 -4 1080 44
rect 1040 -36 1044 -4
rect 1076 -36 1080 -4
rect 1040 -84 1080 -36
rect 1040 -116 1044 -84
rect 1076 -116 1080 -84
rect 1040 -120 1080 -116
rect 1120 1036 1160 1040
rect 1120 1004 1124 1036
rect 1156 1004 1160 1036
rect 1120 956 1160 1004
rect 1120 924 1124 956
rect 1156 924 1160 956
rect 1120 876 1160 924
rect 1120 844 1124 876
rect 1156 844 1160 876
rect 1120 796 1160 844
rect 1120 764 1124 796
rect 1156 764 1160 796
rect 1120 716 1160 764
rect 1120 684 1124 716
rect 1156 684 1160 716
rect 1120 636 1160 684
rect 1120 604 1124 636
rect 1156 604 1160 636
rect 1120 556 1160 604
rect 1120 524 1124 556
rect 1156 524 1160 556
rect 1120 476 1160 524
rect 1120 444 1124 476
rect 1156 444 1160 476
rect 1120 396 1160 444
rect 1120 364 1124 396
rect 1156 364 1160 396
rect 1120 316 1160 364
rect 1120 284 1124 316
rect 1156 284 1160 316
rect 1120 236 1160 284
rect 1120 204 1124 236
rect 1156 204 1160 236
rect 1120 156 1160 204
rect 1120 124 1124 156
rect 1156 124 1160 156
rect 1120 76 1160 124
rect 1120 44 1124 76
rect 1156 44 1160 76
rect 1120 -4 1160 44
rect 1120 -36 1124 -4
rect 1156 -36 1160 -4
rect 1120 -84 1160 -36
rect 1120 -116 1124 -84
rect 1156 -116 1160 -84
rect 1120 -120 1160 -116
rect 1200 1036 1240 1040
rect 1200 1004 1204 1036
rect 1236 1004 1240 1036
rect 1200 956 1240 1004
rect 1200 924 1204 956
rect 1236 924 1240 956
rect 1200 876 1240 924
rect 1200 844 1204 876
rect 1236 844 1240 876
rect 1200 796 1240 844
rect 1200 764 1204 796
rect 1236 764 1240 796
rect 1200 716 1240 764
rect 1200 684 1204 716
rect 1236 684 1240 716
rect 1200 636 1240 684
rect 1200 604 1204 636
rect 1236 604 1240 636
rect 1200 556 1240 604
rect 1200 524 1204 556
rect 1236 524 1240 556
rect 1200 476 1240 524
rect 1200 444 1204 476
rect 1236 444 1240 476
rect 1200 396 1240 444
rect 1200 364 1204 396
rect 1236 364 1240 396
rect 1200 316 1240 364
rect 1200 284 1204 316
rect 1236 284 1240 316
rect 1200 236 1240 284
rect 1200 204 1204 236
rect 1236 204 1240 236
rect 1200 156 1240 204
rect 1200 124 1204 156
rect 1236 124 1240 156
rect 1200 76 1240 124
rect 1200 44 1204 76
rect 1236 44 1240 76
rect 1200 -4 1240 44
rect 1200 -36 1204 -4
rect 1236 -36 1240 -4
rect 1200 -84 1240 -36
rect 1200 -116 1204 -84
rect 1236 -116 1240 -84
rect 1200 -120 1240 -116
rect 1280 1036 1320 1040
rect 1280 1004 1284 1036
rect 1316 1004 1320 1036
rect 1280 956 1320 1004
rect 1280 924 1284 956
rect 1316 924 1320 956
rect 1280 876 1320 924
rect 1280 844 1284 876
rect 1316 844 1320 876
rect 1280 796 1320 844
rect 1280 764 1284 796
rect 1316 764 1320 796
rect 1280 716 1320 764
rect 1280 684 1284 716
rect 1316 684 1320 716
rect 1280 636 1320 684
rect 1280 604 1284 636
rect 1316 604 1320 636
rect 1280 556 1320 604
rect 1280 524 1284 556
rect 1316 524 1320 556
rect 1280 476 1320 524
rect 1280 444 1284 476
rect 1316 444 1320 476
rect 1280 396 1320 444
rect 1280 364 1284 396
rect 1316 364 1320 396
rect 1280 316 1320 364
rect 1280 284 1284 316
rect 1316 284 1320 316
rect 1280 236 1320 284
rect 1280 204 1284 236
rect 1316 204 1320 236
rect 1280 156 1320 204
rect 1280 124 1284 156
rect 1316 124 1320 156
rect 1280 76 1320 124
rect 1280 44 1284 76
rect 1316 44 1320 76
rect 1280 -4 1320 44
rect 1280 -36 1284 -4
rect 1316 -36 1320 -4
rect 1280 -84 1320 -36
rect 1280 -116 1284 -84
rect 1316 -116 1320 -84
rect 1280 -120 1320 -116
rect 1360 1036 1400 1040
rect 1360 1004 1364 1036
rect 1396 1004 1400 1036
rect 1360 956 1400 1004
rect 1360 924 1364 956
rect 1396 924 1400 956
rect 1360 876 1400 924
rect 1360 844 1364 876
rect 1396 844 1400 876
rect 1360 796 1400 844
rect 1360 764 1364 796
rect 1396 764 1400 796
rect 1360 716 1400 764
rect 1360 684 1364 716
rect 1396 684 1400 716
rect 1360 636 1400 684
rect 1360 604 1364 636
rect 1396 604 1400 636
rect 1360 556 1400 604
rect 1360 524 1364 556
rect 1396 524 1400 556
rect 1360 476 1400 524
rect 1360 444 1364 476
rect 1396 444 1400 476
rect 1360 396 1400 444
rect 1360 364 1364 396
rect 1396 364 1400 396
rect 1360 316 1400 364
rect 1360 284 1364 316
rect 1396 284 1400 316
rect 1360 236 1400 284
rect 1360 204 1364 236
rect 1396 204 1400 236
rect 1360 156 1400 204
rect 1360 124 1364 156
rect 1396 124 1400 156
rect 1360 76 1400 124
rect 1360 44 1364 76
rect 1396 44 1400 76
rect 1360 -4 1400 44
rect 1360 -36 1364 -4
rect 1396 -36 1400 -4
rect 1360 -84 1400 -36
rect 1360 -116 1364 -84
rect 1396 -116 1400 -84
rect 1360 -120 1400 -116
rect 1440 1036 1480 1040
rect 1440 1004 1444 1036
rect 1476 1004 1480 1036
rect 1440 956 1480 1004
rect 1440 924 1444 956
rect 1476 924 1480 956
rect 1440 876 1480 924
rect 1440 844 1444 876
rect 1476 844 1480 876
rect 1440 796 1480 844
rect 1440 764 1444 796
rect 1476 764 1480 796
rect 1440 716 1480 764
rect 1440 684 1444 716
rect 1476 684 1480 716
rect 1440 636 1480 684
rect 1440 604 1444 636
rect 1476 604 1480 636
rect 1440 556 1480 604
rect 1440 524 1444 556
rect 1476 524 1480 556
rect 1440 476 1480 524
rect 1440 444 1444 476
rect 1476 444 1480 476
rect 1440 396 1480 444
rect 1440 364 1444 396
rect 1476 364 1480 396
rect 1440 316 1480 364
rect 1440 284 1444 316
rect 1476 284 1480 316
rect 1440 236 1480 284
rect 1440 204 1444 236
rect 1476 204 1480 236
rect 1440 156 1480 204
rect 1440 124 1444 156
rect 1476 124 1480 156
rect 1440 76 1480 124
rect 1440 44 1444 76
rect 1476 44 1480 76
rect 1440 -4 1480 44
rect 1440 -36 1444 -4
rect 1476 -36 1480 -4
rect 1440 -84 1480 -36
rect 1440 -116 1444 -84
rect 1476 -116 1480 -84
rect 1440 -120 1480 -116
rect 1520 1036 1560 1040
rect 1520 1004 1524 1036
rect 1556 1004 1560 1036
rect 1520 956 1560 1004
rect 1520 924 1524 956
rect 1556 924 1560 956
rect 1520 876 1560 924
rect 1520 844 1524 876
rect 1556 844 1560 876
rect 1520 796 1560 844
rect 1520 764 1524 796
rect 1556 764 1560 796
rect 1520 716 1560 764
rect 1520 684 1524 716
rect 1556 684 1560 716
rect 1520 636 1560 684
rect 1520 604 1524 636
rect 1556 604 1560 636
rect 1520 556 1560 604
rect 1520 524 1524 556
rect 1556 524 1560 556
rect 1520 476 1560 524
rect 1520 444 1524 476
rect 1556 444 1560 476
rect 1520 396 1560 444
rect 1520 364 1524 396
rect 1556 364 1560 396
rect 1520 316 1560 364
rect 1520 284 1524 316
rect 1556 284 1560 316
rect 1520 236 1560 284
rect 1520 204 1524 236
rect 1556 204 1560 236
rect 1520 156 1560 204
rect 1520 124 1524 156
rect 1556 124 1560 156
rect 1520 76 1560 124
rect 1520 44 1524 76
rect 1556 44 1560 76
rect 1520 -4 1560 44
rect 1520 -36 1524 -4
rect 1556 -36 1560 -4
rect 1520 -84 1560 -36
rect 1520 -116 1524 -84
rect 1556 -116 1560 -84
rect 1520 -120 1560 -116
rect 1600 1036 1640 1040
rect 1600 1004 1604 1036
rect 1636 1004 1640 1036
rect 1600 956 1640 1004
rect 1600 924 1604 956
rect 1636 924 1640 956
rect 1600 876 1640 924
rect 1600 844 1604 876
rect 1636 844 1640 876
rect 1600 796 1640 844
rect 1600 764 1604 796
rect 1636 764 1640 796
rect 1600 716 1640 764
rect 1600 684 1604 716
rect 1636 684 1640 716
rect 1600 636 1640 684
rect 1600 604 1604 636
rect 1636 604 1640 636
rect 1600 556 1640 604
rect 1600 524 1604 556
rect 1636 524 1640 556
rect 1600 476 1640 524
rect 1600 444 1604 476
rect 1636 444 1640 476
rect 1600 396 1640 444
rect 1600 364 1604 396
rect 1636 364 1640 396
rect 1600 316 1640 364
rect 1600 284 1604 316
rect 1636 284 1640 316
rect 1600 236 1640 284
rect 1600 204 1604 236
rect 1636 204 1640 236
rect 1600 156 1640 204
rect 1600 124 1604 156
rect 1636 124 1640 156
rect 1600 76 1640 124
rect 1600 44 1604 76
rect 1636 44 1640 76
rect 1600 -4 1640 44
rect 1600 -36 1604 -4
rect 1636 -36 1640 -4
rect 1600 -84 1640 -36
rect 1600 -116 1604 -84
rect 1636 -116 1640 -84
rect 1600 -120 1640 -116
rect 1680 1036 1720 1040
rect 1680 1004 1684 1036
rect 1716 1004 1720 1036
rect 1680 956 1720 1004
rect 1680 924 1684 956
rect 1716 924 1720 956
rect 1680 876 1720 924
rect 1680 844 1684 876
rect 1716 844 1720 876
rect 1680 796 1720 844
rect 1680 764 1684 796
rect 1716 764 1720 796
rect 1680 716 1720 764
rect 1680 684 1684 716
rect 1716 684 1720 716
rect 1680 636 1720 684
rect 1680 604 1684 636
rect 1716 604 1720 636
rect 1680 556 1720 604
rect 1680 524 1684 556
rect 1716 524 1720 556
rect 1680 476 1720 524
rect 1680 444 1684 476
rect 1716 444 1720 476
rect 1680 396 1720 444
rect 1680 364 1684 396
rect 1716 364 1720 396
rect 1680 316 1720 364
rect 1680 284 1684 316
rect 1716 284 1720 316
rect 1680 236 1720 284
rect 1680 204 1684 236
rect 1716 204 1720 236
rect 1680 156 1720 204
rect 1680 124 1684 156
rect 1716 124 1720 156
rect 1680 76 1720 124
rect 1680 44 1684 76
rect 1716 44 1720 76
rect 1680 -4 1720 44
rect 1680 -36 1684 -4
rect 1716 -36 1720 -4
rect 1680 -84 1720 -36
rect 1680 -116 1684 -84
rect 1716 -116 1720 -84
rect 1680 -120 1720 -116
rect 1760 1036 1800 1040
rect 1760 1004 1764 1036
rect 1796 1004 1800 1036
rect 1760 956 1800 1004
rect 1760 924 1764 956
rect 1796 924 1800 956
rect 1760 876 1800 924
rect 1760 844 1764 876
rect 1796 844 1800 876
rect 1760 796 1800 844
rect 1760 764 1764 796
rect 1796 764 1800 796
rect 1760 716 1800 764
rect 1760 684 1764 716
rect 1796 684 1800 716
rect 1760 636 1800 684
rect 1760 604 1764 636
rect 1796 604 1800 636
rect 1760 556 1800 604
rect 1760 524 1764 556
rect 1796 524 1800 556
rect 1760 476 1800 524
rect 1760 444 1764 476
rect 1796 444 1800 476
rect 1760 396 1800 444
rect 1760 364 1764 396
rect 1796 364 1800 396
rect 1760 316 1800 364
rect 1760 284 1764 316
rect 1796 284 1800 316
rect 1760 236 1800 284
rect 1760 204 1764 236
rect 1796 204 1800 236
rect 1760 156 1800 204
rect 1760 124 1764 156
rect 1796 124 1800 156
rect 1760 76 1800 124
rect 1760 44 1764 76
rect 1796 44 1800 76
rect 1760 -4 1800 44
rect 1760 -36 1764 -4
rect 1796 -36 1800 -4
rect 1760 -84 1800 -36
rect 1760 -116 1764 -84
rect 1796 -116 1800 -84
rect 1760 -120 1800 -116
rect 1840 1036 1880 1040
rect 1840 1004 1844 1036
rect 1876 1004 1880 1036
rect 1840 956 1880 1004
rect 1840 924 1844 956
rect 1876 924 1880 956
rect 1840 876 1880 924
rect 1840 844 1844 876
rect 1876 844 1880 876
rect 1840 796 1880 844
rect 1840 764 1844 796
rect 1876 764 1880 796
rect 1840 716 1880 764
rect 1840 684 1844 716
rect 1876 684 1880 716
rect 1840 636 1880 684
rect 1840 604 1844 636
rect 1876 604 1880 636
rect 1840 556 1880 604
rect 1840 524 1844 556
rect 1876 524 1880 556
rect 1840 476 1880 524
rect 1840 444 1844 476
rect 1876 444 1880 476
rect 1840 396 1880 444
rect 1840 364 1844 396
rect 1876 364 1880 396
rect 1840 316 1880 364
rect 1840 284 1844 316
rect 1876 284 1880 316
rect 1840 236 1880 284
rect 1840 204 1844 236
rect 1876 204 1880 236
rect 1840 156 1880 204
rect 1840 124 1844 156
rect 1876 124 1880 156
rect 1840 76 1880 124
rect 1840 44 1844 76
rect 1876 44 1880 76
rect 1840 -4 1880 44
rect 1840 -36 1844 -4
rect 1876 -36 1880 -4
rect 1840 -84 1880 -36
rect 1840 -116 1844 -84
rect 1876 -116 1880 -84
rect 1840 -120 1880 -116
rect 1920 1036 1960 1040
rect 1920 1004 1924 1036
rect 1956 1004 1960 1036
rect 1920 956 1960 1004
rect 1920 924 1924 956
rect 1956 924 1960 956
rect 1920 876 1960 924
rect 1920 844 1924 876
rect 1956 844 1960 876
rect 1920 796 1960 844
rect 1920 764 1924 796
rect 1956 764 1960 796
rect 1920 716 1960 764
rect 1920 684 1924 716
rect 1956 684 1960 716
rect 1920 636 1960 684
rect 1920 604 1924 636
rect 1956 604 1960 636
rect 1920 556 1960 604
rect 1920 524 1924 556
rect 1956 524 1960 556
rect 1920 476 1960 524
rect 1920 444 1924 476
rect 1956 444 1960 476
rect 1920 396 1960 444
rect 1920 364 1924 396
rect 1956 364 1960 396
rect 1920 316 1960 364
rect 1920 284 1924 316
rect 1956 284 1960 316
rect 1920 236 1960 284
rect 1920 204 1924 236
rect 1956 204 1960 236
rect 1920 156 1960 204
rect 1920 124 1924 156
rect 1956 124 1960 156
rect 1920 76 1960 124
rect 1920 44 1924 76
rect 1956 44 1960 76
rect 1920 -4 1960 44
rect 1920 -36 1924 -4
rect 1956 -36 1960 -4
rect 1920 -84 1960 -36
rect 1920 -116 1924 -84
rect 1956 -116 1960 -84
rect 1920 -120 1960 -116
rect 2000 1036 2040 1040
rect 2000 1004 2004 1036
rect 2036 1004 2040 1036
rect 2000 956 2040 1004
rect 2000 924 2004 956
rect 2036 924 2040 956
rect 2000 876 2040 924
rect 2000 844 2004 876
rect 2036 844 2040 876
rect 2000 796 2040 844
rect 2000 764 2004 796
rect 2036 764 2040 796
rect 2000 716 2040 764
rect 2000 684 2004 716
rect 2036 684 2040 716
rect 2000 636 2040 684
rect 2000 604 2004 636
rect 2036 604 2040 636
rect 2000 556 2040 604
rect 2000 524 2004 556
rect 2036 524 2040 556
rect 2000 476 2040 524
rect 2000 444 2004 476
rect 2036 444 2040 476
rect 2000 396 2040 444
rect 2000 364 2004 396
rect 2036 364 2040 396
rect 2000 316 2040 364
rect 2000 284 2004 316
rect 2036 284 2040 316
rect 2000 236 2040 284
rect 2000 204 2004 236
rect 2036 204 2040 236
rect 2000 156 2040 204
rect 2000 124 2004 156
rect 2036 124 2040 156
rect 2000 76 2040 124
rect 2000 44 2004 76
rect 2036 44 2040 76
rect 2000 -4 2040 44
rect 2000 -36 2004 -4
rect 2036 -36 2040 -4
rect 2000 -84 2040 -36
rect 2000 -116 2004 -84
rect 2036 -116 2040 -84
rect 2000 -120 2040 -116
rect 2080 1036 2120 1040
rect 2080 1004 2084 1036
rect 2116 1004 2120 1036
rect 2080 956 2120 1004
rect 2080 924 2084 956
rect 2116 924 2120 956
rect 2080 876 2120 924
rect 2080 844 2084 876
rect 2116 844 2120 876
rect 2080 796 2120 844
rect 2080 764 2084 796
rect 2116 764 2120 796
rect 2080 716 2120 764
rect 2080 684 2084 716
rect 2116 684 2120 716
rect 2080 636 2120 684
rect 2080 604 2084 636
rect 2116 604 2120 636
rect 2080 556 2120 604
rect 2080 524 2084 556
rect 2116 524 2120 556
rect 2080 476 2120 524
rect 2080 444 2084 476
rect 2116 444 2120 476
rect 2080 396 2120 444
rect 2080 364 2084 396
rect 2116 364 2120 396
rect 2080 316 2120 364
rect 2080 284 2084 316
rect 2116 284 2120 316
rect 2080 236 2120 284
rect 2080 204 2084 236
rect 2116 204 2120 236
rect 2080 156 2120 204
rect 2080 124 2084 156
rect 2116 124 2120 156
rect 2080 76 2120 124
rect 2080 44 2084 76
rect 2116 44 2120 76
rect 2080 -4 2120 44
rect 2080 -36 2084 -4
rect 2116 -36 2120 -4
rect 2080 -84 2120 -36
rect 2080 -116 2084 -84
rect 2116 -116 2120 -84
rect 2080 -120 2120 -116
rect 2160 1036 2200 1040
rect 2160 1004 2164 1036
rect 2196 1004 2200 1036
rect 2160 956 2200 1004
rect 2160 924 2164 956
rect 2196 924 2200 956
rect 2160 876 2200 924
rect 2160 844 2164 876
rect 2196 844 2200 876
rect 2160 796 2200 844
rect 2160 764 2164 796
rect 2196 764 2200 796
rect 2160 716 2200 764
rect 2160 684 2164 716
rect 2196 684 2200 716
rect 2160 636 2200 684
rect 2160 604 2164 636
rect 2196 604 2200 636
rect 2160 556 2200 604
rect 2160 524 2164 556
rect 2196 524 2200 556
rect 2160 476 2200 524
rect 2160 444 2164 476
rect 2196 444 2200 476
rect 2160 396 2200 444
rect 2160 364 2164 396
rect 2196 364 2200 396
rect 2160 316 2200 364
rect 2160 284 2164 316
rect 2196 284 2200 316
rect 2160 236 2200 284
rect 2160 204 2164 236
rect 2196 204 2200 236
rect 2160 156 2200 204
rect 2160 124 2164 156
rect 2196 124 2200 156
rect 2160 76 2200 124
rect 2160 44 2164 76
rect 2196 44 2200 76
rect 2160 -4 2200 44
rect 2160 -36 2164 -4
rect 2196 -36 2200 -4
rect 2160 -84 2200 -36
rect 2160 -116 2164 -84
rect 2196 -116 2200 -84
rect 2160 -120 2200 -116
rect 2240 1036 2280 1040
rect 2240 1004 2244 1036
rect 2276 1004 2280 1036
rect 2240 956 2280 1004
rect 2240 924 2244 956
rect 2276 924 2280 956
rect 2240 876 2280 924
rect 2240 844 2244 876
rect 2276 844 2280 876
rect 2240 796 2280 844
rect 2240 764 2244 796
rect 2276 764 2280 796
rect 2240 716 2280 764
rect 2240 684 2244 716
rect 2276 684 2280 716
rect 2240 636 2280 684
rect 2240 604 2244 636
rect 2276 604 2280 636
rect 2240 556 2280 604
rect 2240 524 2244 556
rect 2276 524 2280 556
rect 2240 476 2280 524
rect 2240 444 2244 476
rect 2276 444 2280 476
rect 2240 396 2280 444
rect 2240 364 2244 396
rect 2276 364 2280 396
rect 2240 316 2280 364
rect 2240 284 2244 316
rect 2276 284 2280 316
rect 2240 236 2280 284
rect 2240 204 2244 236
rect 2276 204 2280 236
rect 2240 156 2280 204
rect 2240 124 2244 156
rect 2276 124 2280 156
rect 2240 76 2280 124
rect 2240 44 2244 76
rect 2276 44 2280 76
rect 2240 -4 2280 44
rect 2240 -36 2244 -4
rect 2276 -36 2280 -4
rect 2240 -84 2280 -36
rect 2240 -116 2244 -84
rect 2276 -116 2280 -84
rect 2240 -120 2280 -116
rect 2320 1036 2360 1040
rect 2320 1004 2324 1036
rect 2356 1004 2360 1036
rect 2320 956 2360 1004
rect 2320 924 2324 956
rect 2356 924 2360 956
rect 2320 876 2360 924
rect 2320 844 2324 876
rect 2356 844 2360 876
rect 2320 796 2360 844
rect 2320 764 2324 796
rect 2356 764 2360 796
rect 2320 716 2360 764
rect 2320 684 2324 716
rect 2356 684 2360 716
rect 2320 636 2360 684
rect 2320 604 2324 636
rect 2356 604 2360 636
rect 2320 556 2360 604
rect 2320 524 2324 556
rect 2356 524 2360 556
rect 2320 476 2360 524
rect 2320 444 2324 476
rect 2356 444 2360 476
rect 2320 396 2360 444
rect 2320 364 2324 396
rect 2356 364 2360 396
rect 2320 316 2360 364
rect 2320 284 2324 316
rect 2356 284 2360 316
rect 2320 236 2360 284
rect 2320 204 2324 236
rect 2356 204 2360 236
rect 2320 156 2360 204
rect 2320 124 2324 156
rect 2356 124 2360 156
rect 2320 76 2360 124
rect 2320 44 2324 76
rect 2356 44 2360 76
rect 2320 -4 2360 44
rect 2320 -36 2324 -4
rect 2356 -36 2360 -4
rect 2320 -84 2360 -36
rect 2320 -116 2324 -84
rect 2356 -116 2360 -84
rect 2320 -120 2360 -116
rect 2400 1036 2440 1040
rect 2400 1004 2404 1036
rect 2436 1004 2440 1036
rect 2400 956 2440 1004
rect 2400 924 2404 956
rect 2436 924 2440 956
rect 2400 876 2440 924
rect 2400 844 2404 876
rect 2436 844 2440 876
rect 2400 796 2440 844
rect 2400 764 2404 796
rect 2436 764 2440 796
rect 2400 716 2440 764
rect 2400 684 2404 716
rect 2436 684 2440 716
rect 2400 636 2440 684
rect 2400 604 2404 636
rect 2436 604 2440 636
rect 2400 556 2440 604
rect 2400 524 2404 556
rect 2436 524 2440 556
rect 2400 476 2440 524
rect 2400 444 2404 476
rect 2436 444 2440 476
rect 2400 396 2440 444
rect 2400 364 2404 396
rect 2436 364 2440 396
rect 2400 316 2440 364
rect 2400 284 2404 316
rect 2436 284 2440 316
rect 2400 236 2440 284
rect 2400 204 2404 236
rect 2436 204 2440 236
rect 2400 156 2440 204
rect 2400 124 2404 156
rect 2436 124 2440 156
rect 2400 76 2440 124
rect 2400 44 2404 76
rect 2436 44 2440 76
rect 2400 -4 2440 44
rect 2400 -36 2404 -4
rect 2436 -36 2440 -4
rect 2400 -84 2440 -36
rect 2400 -116 2404 -84
rect 2436 -116 2440 -84
rect 2400 -120 2440 -116
rect 2480 1036 2520 1040
rect 2480 1004 2484 1036
rect 2516 1004 2520 1036
rect 2480 956 2520 1004
rect 2480 924 2484 956
rect 2516 924 2520 956
rect 2480 876 2520 924
rect 2480 844 2484 876
rect 2516 844 2520 876
rect 2480 796 2520 844
rect 2480 764 2484 796
rect 2516 764 2520 796
rect 2480 716 2520 764
rect 2480 684 2484 716
rect 2516 684 2520 716
rect 2480 636 2520 684
rect 2480 604 2484 636
rect 2516 604 2520 636
rect 2480 556 2520 604
rect 2480 524 2484 556
rect 2516 524 2520 556
rect 2480 476 2520 524
rect 2480 444 2484 476
rect 2516 444 2520 476
rect 2480 396 2520 444
rect 2480 364 2484 396
rect 2516 364 2520 396
rect 2480 316 2520 364
rect 2480 284 2484 316
rect 2516 284 2520 316
rect 2480 236 2520 284
rect 2480 204 2484 236
rect 2516 204 2520 236
rect 2480 156 2520 204
rect 2480 124 2484 156
rect 2516 124 2520 156
rect 2480 76 2520 124
rect 2480 44 2484 76
rect 2516 44 2520 76
rect 2480 -4 2520 44
rect 2480 -36 2484 -4
rect 2516 -36 2520 -4
rect 2480 -84 2520 -36
rect 2480 -116 2484 -84
rect 2516 -116 2520 -84
rect 2480 -120 2520 -116
rect 2560 1036 2600 1040
rect 2560 1004 2564 1036
rect 2596 1004 2600 1036
rect 2560 956 2600 1004
rect 2560 924 2564 956
rect 2596 924 2600 956
rect 2560 876 2600 924
rect 2560 844 2564 876
rect 2596 844 2600 876
rect 2560 796 2600 844
rect 2560 764 2564 796
rect 2596 764 2600 796
rect 2560 716 2600 764
rect 2560 684 2564 716
rect 2596 684 2600 716
rect 2560 636 2600 684
rect 2560 604 2564 636
rect 2596 604 2600 636
rect 2560 556 2600 604
rect 2560 524 2564 556
rect 2596 524 2600 556
rect 2560 476 2600 524
rect 2560 444 2564 476
rect 2596 444 2600 476
rect 2560 396 2600 444
rect 2560 364 2564 396
rect 2596 364 2600 396
rect 2560 316 2600 364
rect 2560 284 2564 316
rect 2596 284 2600 316
rect 2560 236 2600 284
rect 2560 204 2564 236
rect 2596 204 2600 236
rect 2560 156 2600 204
rect 2560 124 2564 156
rect 2596 124 2600 156
rect 2560 76 2600 124
rect 2560 44 2564 76
rect 2596 44 2600 76
rect 2560 -4 2600 44
rect 2560 -36 2564 -4
rect 2596 -36 2600 -4
rect 2560 -84 2600 -36
rect 2560 -116 2564 -84
rect 2596 -116 2600 -84
rect 2560 -120 2600 -116
rect 2640 1036 2680 1040
rect 2640 1004 2644 1036
rect 2676 1004 2680 1036
rect 2640 956 2680 1004
rect 2640 924 2644 956
rect 2676 924 2680 956
rect 2640 876 2680 924
rect 2640 844 2644 876
rect 2676 844 2680 876
rect 2640 796 2680 844
rect 2640 764 2644 796
rect 2676 764 2680 796
rect 2640 716 2680 764
rect 2640 684 2644 716
rect 2676 684 2680 716
rect 2640 636 2680 684
rect 2640 604 2644 636
rect 2676 604 2680 636
rect 2640 556 2680 604
rect 2640 524 2644 556
rect 2676 524 2680 556
rect 2640 476 2680 524
rect 2640 444 2644 476
rect 2676 444 2680 476
rect 2640 396 2680 444
rect 2640 364 2644 396
rect 2676 364 2680 396
rect 2640 316 2680 364
rect 2640 284 2644 316
rect 2676 284 2680 316
rect 2640 236 2680 284
rect 2640 204 2644 236
rect 2676 204 2680 236
rect 2640 156 2680 204
rect 2640 124 2644 156
rect 2676 124 2680 156
rect 2640 76 2680 124
rect 2640 44 2644 76
rect 2676 44 2680 76
rect 2640 -4 2680 44
rect 2640 -36 2644 -4
rect 2676 -36 2680 -4
rect 2640 -84 2680 -36
rect 2640 -116 2644 -84
rect 2676 -116 2680 -84
rect 2640 -120 2680 -116
rect 2720 1036 2760 1040
rect 2720 1004 2724 1036
rect 2756 1004 2760 1036
rect 2720 956 2760 1004
rect 2720 924 2724 956
rect 2756 924 2760 956
rect 2720 876 2760 924
rect 2720 844 2724 876
rect 2756 844 2760 876
rect 2720 796 2760 844
rect 2720 764 2724 796
rect 2756 764 2760 796
rect 2720 716 2760 764
rect 2720 684 2724 716
rect 2756 684 2760 716
rect 2720 636 2760 684
rect 2720 604 2724 636
rect 2756 604 2760 636
rect 2720 556 2760 604
rect 2720 524 2724 556
rect 2756 524 2760 556
rect 2720 476 2760 524
rect 2720 444 2724 476
rect 2756 444 2760 476
rect 2720 396 2760 444
rect 2720 364 2724 396
rect 2756 364 2760 396
rect 2720 316 2760 364
rect 2720 284 2724 316
rect 2756 284 2760 316
rect 2720 236 2760 284
rect 2720 204 2724 236
rect 2756 204 2760 236
rect 2720 156 2760 204
rect 2720 124 2724 156
rect 2756 124 2760 156
rect 2720 76 2760 124
rect 2720 44 2724 76
rect 2756 44 2760 76
rect 2720 -4 2760 44
rect 2720 -36 2724 -4
rect 2756 -36 2760 -4
rect 2720 -84 2760 -36
rect 2720 -116 2724 -84
rect 2756 -116 2760 -84
rect 2720 -120 2760 -116
rect 2800 1036 2840 1040
rect 2800 1004 2804 1036
rect 2836 1004 2840 1036
rect 2800 956 2840 1004
rect 2800 924 2804 956
rect 2836 924 2840 956
rect 2800 876 2840 924
rect 2800 844 2804 876
rect 2836 844 2840 876
rect 2800 796 2840 844
rect 2800 764 2804 796
rect 2836 764 2840 796
rect 2800 716 2840 764
rect 2800 684 2804 716
rect 2836 684 2840 716
rect 2800 636 2840 684
rect 2800 604 2804 636
rect 2836 604 2840 636
rect 2800 556 2840 604
rect 2800 524 2804 556
rect 2836 524 2840 556
rect 2800 476 2840 524
rect 2800 444 2804 476
rect 2836 444 2840 476
rect 2800 396 2840 444
rect 2800 364 2804 396
rect 2836 364 2840 396
rect 2800 316 2840 364
rect 2800 284 2804 316
rect 2836 284 2840 316
rect 2800 236 2840 284
rect 2800 204 2804 236
rect 2836 204 2840 236
rect 2800 156 2840 204
rect 2800 124 2804 156
rect 2836 124 2840 156
rect 2800 76 2840 124
rect 2800 44 2804 76
rect 2836 44 2840 76
rect 2800 -4 2840 44
rect 2800 -36 2804 -4
rect 2836 -36 2840 -4
rect 2800 -84 2840 -36
rect 2800 -116 2804 -84
rect 2836 -116 2840 -84
rect 2800 -120 2840 -116
rect 2880 1036 2920 1040
rect 2880 1004 2884 1036
rect 2916 1004 2920 1036
rect 2880 956 2920 1004
rect 2880 924 2884 956
rect 2916 924 2920 956
rect 2880 876 2920 924
rect 2880 844 2884 876
rect 2916 844 2920 876
rect 2880 796 2920 844
rect 2880 764 2884 796
rect 2916 764 2920 796
rect 2880 716 2920 764
rect 2880 684 2884 716
rect 2916 684 2920 716
rect 2880 636 2920 684
rect 2880 604 2884 636
rect 2916 604 2920 636
rect 2880 556 2920 604
rect 2880 524 2884 556
rect 2916 524 2920 556
rect 2880 476 2920 524
rect 2880 444 2884 476
rect 2916 444 2920 476
rect 2880 396 2920 444
rect 2880 364 2884 396
rect 2916 364 2920 396
rect 2880 316 2920 364
rect 2880 284 2884 316
rect 2916 284 2920 316
rect 2880 236 2920 284
rect 2880 204 2884 236
rect 2916 204 2920 236
rect 2880 156 2920 204
rect 2880 124 2884 156
rect 2916 124 2920 156
rect 2880 76 2920 124
rect 2880 44 2884 76
rect 2916 44 2920 76
rect 2880 -4 2920 44
rect 2880 -36 2884 -4
rect 2916 -36 2920 -4
rect 2880 -84 2920 -36
rect 2880 -116 2884 -84
rect 2916 -116 2920 -84
rect 2880 -120 2920 -116
rect 2960 1036 3000 1040
rect 2960 1004 2964 1036
rect 2996 1004 3000 1036
rect 2960 956 3000 1004
rect 2960 924 2964 956
rect 2996 924 3000 956
rect 2960 876 3000 924
rect 2960 844 2964 876
rect 2996 844 3000 876
rect 2960 796 3000 844
rect 2960 764 2964 796
rect 2996 764 3000 796
rect 2960 716 3000 764
rect 2960 684 2964 716
rect 2996 684 3000 716
rect 2960 636 3000 684
rect 2960 604 2964 636
rect 2996 604 3000 636
rect 2960 556 3000 604
rect 2960 524 2964 556
rect 2996 524 3000 556
rect 2960 476 3000 524
rect 2960 444 2964 476
rect 2996 444 3000 476
rect 2960 396 3000 444
rect 2960 364 2964 396
rect 2996 364 3000 396
rect 2960 316 3000 364
rect 2960 284 2964 316
rect 2996 284 3000 316
rect 2960 236 3000 284
rect 2960 204 2964 236
rect 2996 204 3000 236
rect 2960 156 3000 204
rect 2960 124 2964 156
rect 2996 124 3000 156
rect 2960 76 3000 124
rect 2960 44 2964 76
rect 2996 44 3000 76
rect 2960 -4 3000 44
rect 2960 -36 2964 -4
rect 2996 -36 3000 -4
rect 2960 -84 3000 -36
rect 2960 -116 2964 -84
rect 2996 -116 3000 -84
rect 2960 -120 3000 -116
rect 3040 1036 3080 1040
rect 3040 1004 3044 1036
rect 3076 1004 3080 1036
rect 3040 956 3080 1004
rect 3040 924 3044 956
rect 3076 924 3080 956
rect 3040 876 3080 924
rect 3040 844 3044 876
rect 3076 844 3080 876
rect 3040 796 3080 844
rect 3040 764 3044 796
rect 3076 764 3080 796
rect 3040 716 3080 764
rect 3040 684 3044 716
rect 3076 684 3080 716
rect 3040 636 3080 684
rect 3040 604 3044 636
rect 3076 604 3080 636
rect 3040 556 3080 604
rect 3040 524 3044 556
rect 3076 524 3080 556
rect 3040 476 3080 524
rect 3040 444 3044 476
rect 3076 444 3080 476
rect 3040 396 3080 444
rect 3040 364 3044 396
rect 3076 364 3080 396
rect 3040 316 3080 364
rect 3040 284 3044 316
rect 3076 284 3080 316
rect 3040 236 3080 284
rect 3040 204 3044 236
rect 3076 204 3080 236
rect 3040 156 3080 204
rect 3040 124 3044 156
rect 3076 124 3080 156
rect 3040 76 3080 124
rect 3040 44 3044 76
rect 3076 44 3080 76
rect 3040 -4 3080 44
rect 3040 -36 3044 -4
rect 3076 -36 3080 -4
rect 3040 -84 3080 -36
rect 3040 -116 3044 -84
rect 3076 -116 3080 -84
rect 3040 -120 3080 -116
rect 3120 1036 3160 1040
rect 3120 1004 3124 1036
rect 3156 1004 3160 1036
rect 3120 956 3160 1004
rect 3120 924 3124 956
rect 3156 924 3160 956
rect 3120 876 3160 924
rect 3120 844 3124 876
rect 3156 844 3160 876
rect 3120 796 3160 844
rect 3120 764 3124 796
rect 3156 764 3160 796
rect 3120 716 3160 764
rect 3120 684 3124 716
rect 3156 684 3160 716
rect 3120 636 3160 684
rect 3120 604 3124 636
rect 3156 604 3160 636
rect 3120 556 3160 604
rect 3120 524 3124 556
rect 3156 524 3160 556
rect 3120 476 3160 524
rect 3120 444 3124 476
rect 3156 444 3160 476
rect 3120 396 3160 444
rect 3120 364 3124 396
rect 3156 364 3160 396
rect 3120 316 3160 364
rect 3120 284 3124 316
rect 3156 284 3160 316
rect 3120 236 3160 284
rect 3120 204 3124 236
rect 3156 204 3160 236
rect 3120 156 3160 204
rect 3120 124 3124 156
rect 3156 124 3160 156
rect 3120 76 3160 124
rect 3120 44 3124 76
rect 3156 44 3160 76
rect 3120 -4 3160 44
rect 3120 -36 3124 -4
rect 3156 -36 3160 -4
rect 3120 -84 3160 -36
rect 3120 -116 3124 -84
rect 3156 -116 3160 -84
rect 3120 -120 3160 -116
rect 3200 1036 3240 1040
rect 3200 1004 3204 1036
rect 3236 1004 3240 1036
rect 3200 956 3240 1004
rect 3200 924 3204 956
rect 3236 924 3240 956
rect 3200 876 3240 924
rect 3200 844 3204 876
rect 3236 844 3240 876
rect 3200 796 3240 844
rect 3200 764 3204 796
rect 3236 764 3240 796
rect 3200 716 3240 764
rect 3200 684 3204 716
rect 3236 684 3240 716
rect 3200 636 3240 684
rect 3200 604 3204 636
rect 3236 604 3240 636
rect 3200 556 3240 604
rect 3200 524 3204 556
rect 3236 524 3240 556
rect 3200 476 3240 524
rect 3200 444 3204 476
rect 3236 444 3240 476
rect 3200 396 3240 444
rect 3200 364 3204 396
rect 3236 364 3240 396
rect 3200 316 3240 364
rect 3200 284 3204 316
rect 3236 284 3240 316
rect 3200 236 3240 284
rect 3200 204 3204 236
rect 3236 204 3240 236
rect 3200 156 3240 204
rect 3200 124 3204 156
rect 3236 124 3240 156
rect 3200 76 3240 124
rect 3200 44 3204 76
rect 3236 44 3240 76
rect 3200 -4 3240 44
rect 3200 -36 3204 -4
rect 3236 -36 3240 -4
rect 3200 -84 3240 -36
rect 3200 -116 3204 -84
rect 3236 -116 3240 -84
rect 3200 -120 3240 -116
rect 3280 1036 3320 1040
rect 3280 1004 3284 1036
rect 3316 1004 3320 1036
rect 3280 956 3320 1004
rect 3280 924 3284 956
rect 3316 924 3320 956
rect 3280 876 3320 924
rect 3280 844 3284 876
rect 3316 844 3320 876
rect 3280 796 3320 844
rect 3280 764 3284 796
rect 3316 764 3320 796
rect 3280 716 3320 764
rect 3280 684 3284 716
rect 3316 684 3320 716
rect 3280 636 3320 684
rect 3280 604 3284 636
rect 3316 604 3320 636
rect 3280 556 3320 604
rect 3280 524 3284 556
rect 3316 524 3320 556
rect 3280 476 3320 524
rect 3280 444 3284 476
rect 3316 444 3320 476
rect 3280 396 3320 444
rect 3280 364 3284 396
rect 3316 364 3320 396
rect 3280 316 3320 364
rect 3280 284 3284 316
rect 3316 284 3320 316
rect 3280 236 3320 284
rect 3280 204 3284 236
rect 3316 204 3320 236
rect 3280 156 3320 204
rect 3280 124 3284 156
rect 3316 124 3320 156
rect 3280 76 3320 124
rect 3280 44 3284 76
rect 3316 44 3320 76
rect 3280 -4 3320 44
rect 3280 -36 3284 -4
rect 3316 -36 3320 -4
rect 3280 -84 3320 -36
rect 3280 -116 3284 -84
rect 3316 -116 3320 -84
rect 3280 -120 3320 -116
rect 3360 1036 3400 1040
rect 3360 1004 3364 1036
rect 3396 1004 3400 1036
rect 3360 956 3400 1004
rect 3360 924 3364 956
rect 3396 924 3400 956
rect 3360 876 3400 924
rect 3360 844 3364 876
rect 3396 844 3400 876
rect 3360 796 3400 844
rect 3360 764 3364 796
rect 3396 764 3400 796
rect 3360 716 3400 764
rect 3360 684 3364 716
rect 3396 684 3400 716
rect 3360 636 3400 684
rect 3360 604 3364 636
rect 3396 604 3400 636
rect 3360 556 3400 604
rect 3360 524 3364 556
rect 3396 524 3400 556
rect 3360 476 3400 524
rect 3360 444 3364 476
rect 3396 444 3400 476
rect 3360 396 3400 444
rect 3360 364 3364 396
rect 3396 364 3400 396
rect 3360 316 3400 364
rect 3360 284 3364 316
rect 3396 284 3400 316
rect 3360 236 3400 284
rect 3360 204 3364 236
rect 3396 204 3400 236
rect 3360 156 3400 204
rect 3360 124 3364 156
rect 3396 124 3400 156
rect 3360 76 3400 124
rect 3360 44 3364 76
rect 3396 44 3400 76
rect 3360 -4 3400 44
rect 3360 -36 3364 -4
rect 3396 -36 3400 -4
rect 3360 -84 3400 -36
rect 3360 -116 3364 -84
rect 3396 -116 3400 -84
rect 3360 -120 3400 -116
rect 3440 1036 3480 1040
rect 3440 1004 3444 1036
rect 3476 1004 3480 1036
rect 3440 956 3480 1004
rect 3440 924 3444 956
rect 3476 924 3480 956
rect 3440 876 3480 924
rect 3440 844 3444 876
rect 3476 844 3480 876
rect 3440 796 3480 844
rect 3440 764 3444 796
rect 3476 764 3480 796
rect 3440 716 3480 764
rect 3440 684 3444 716
rect 3476 684 3480 716
rect 3440 636 3480 684
rect 3440 604 3444 636
rect 3476 604 3480 636
rect 3440 556 3480 604
rect 3440 524 3444 556
rect 3476 524 3480 556
rect 3440 476 3480 524
rect 3440 444 3444 476
rect 3476 444 3480 476
rect 3440 396 3480 444
rect 3440 364 3444 396
rect 3476 364 3480 396
rect 3440 316 3480 364
rect 3440 284 3444 316
rect 3476 284 3480 316
rect 3440 236 3480 284
rect 3440 204 3444 236
rect 3476 204 3480 236
rect 3440 156 3480 204
rect 3440 124 3444 156
rect 3476 124 3480 156
rect 3440 76 3480 124
rect 3440 44 3444 76
rect 3476 44 3480 76
rect 3440 -4 3480 44
rect 3440 -36 3444 -4
rect 3476 -36 3480 -4
rect 3440 -84 3480 -36
rect 3440 -116 3444 -84
rect 3476 -116 3480 -84
rect 3440 -120 3480 -116
rect 3520 1036 3560 1040
rect 3520 1004 3524 1036
rect 3556 1004 3560 1036
rect 3520 956 3560 1004
rect 3520 924 3524 956
rect 3556 924 3560 956
rect 3520 876 3560 924
rect 3520 844 3524 876
rect 3556 844 3560 876
rect 3520 796 3560 844
rect 3520 764 3524 796
rect 3556 764 3560 796
rect 3520 716 3560 764
rect 3520 684 3524 716
rect 3556 684 3560 716
rect 3520 636 3560 684
rect 3520 604 3524 636
rect 3556 604 3560 636
rect 3520 556 3560 604
rect 3520 524 3524 556
rect 3556 524 3560 556
rect 3520 476 3560 524
rect 3520 444 3524 476
rect 3556 444 3560 476
rect 3520 396 3560 444
rect 3520 364 3524 396
rect 3556 364 3560 396
rect 3520 316 3560 364
rect 3520 284 3524 316
rect 3556 284 3560 316
rect 3520 236 3560 284
rect 3520 204 3524 236
rect 3556 204 3560 236
rect 3520 156 3560 204
rect 3520 124 3524 156
rect 3556 124 3560 156
rect 3520 76 3560 124
rect 3520 44 3524 76
rect 3556 44 3560 76
rect 3520 -4 3560 44
rect 3520 -36 3524 -4
rect 3556 -36 3560 -4
rect 3520 -84 3560 -36
rect 3520 -116 3524 -84
rect 3556 -116 3560 -84
rect 3520 -120 3560 -116
rect 3600 1036 3640 1040
rect 3600 1004 3604 1036
rect 3636 1004 3640 1036
rect 3600 956 3640 1004
rect 3600 924 3604 956
rect 3636 924 3640 956
rect 3600 876 3640 924
rect 3600 844 3604 876
rect 3636 844 3640 876
rect 3600 796 3640 844
rect 3600 764 3604 796
rect 3636 764 3640 796
rect 3600 716 3640 764
rect 3600 684 3604 716
rect 3636 684 3640 716
rect 3600 636 3640 684
rect 3600 604 3604 636
rect 3636 604 3640 636
rect 3600 556 3640 604
rect 3600 524 3604 556
rect 3636 524 3640 556
rect 3600 476 3640 524
rect 3600 444 3604 476
rect 3636 444 3640 476
rect 3600 396 3640 444
rect 3600 364 3604 396
rect 3636 364 3640 396
rect 3600 316 3640 364
rect 3600 284 3604 316
rect 3636 284 3640 316
rect 3600 236 3640 284
rect 3600 204 3604 236
rect 3636 204 3640 236
rect 3600 156 3640 204
rect 3600 124 3604 156
rect 3636 124 3640 156
rect 3600 76 3640 124
rect 3600 44 3604 76
rect 3636 44 3640 76
rect 3600 -4 3640 44
rect 3600 -36 3604 -4
rect 3636 -36 3640 -4
rect 3600 -84 3640 -36
rect 3600 -116 3604 -84
rect 3636 -116 3640 -84
rect 3600 -120 3640 -116
rect 3680 1036 3720 1040
rect 3680 1004 3684 1036
rect 3716 1004 3720 1036
rect 3680 956 3720 1004
rect 3680 924 3684 956
rect 3716 924 3720 956
rect 3680 876 3720 924
rect 3680 844 3684 876
rect 3716 844 3720 876
rect 3680 796 3720 844
rect 3680 764 3684 796
rect 3716 764 3720 796
rect 3680 716 3720 764
rect 3680 684 3684 716
rect 3716 684 3720 716
rect 3680 636 3720 684
rect 3680 604 3684 636
rect 3716 604 3720 636
rect 3680 556 3720 604
rect 3680 524 3684 556
rect 3716 524 3720 556
rect 3680 476 3720 524
rect 3680 444 3684 476
rect 3716 444 3720 476
rect 3680 396 3720 444
rect 3680 364 3684 396
rect 3716 364 3720 396
rect 3680 316 3720 364
rect 3680 284 3684 316
rect 3716 284 3720 316
rect 3680 236 3720 284
rect 3680 204 3684 236
rect 3716 204 3720 236
rect 3680 156 3720 204
rect 3680 124 3684 156
rect 3716 124 3720 156
rect 3680 76 3720 124
rect 3680 44 3684 76
rect 3716 44 3720 76
rect 3680 -4 3720 44
rect 3680 -36 3684 -4
rect 3716 -36 3720 -4
rect 3680 -84 3720 -36
rect 3680 -116 3684 -84
rect 3716 -116 3720 -84
rect 3680 -120 3720 -116
rect 3760 1036 3800 1040
rect 3760 1004 3764 1036
rect 3796 1004 3800 1036
rect 3760 956 3800 1004
rect 3760 924 3764 956
rect 3796 924 3800 956
rect 3760 876 3800 924
rect 3760 844 3764 876
rect 3796 844 3800 876
rect 3760 796 3800 844
rect 3760 764 3764 796
rect 3796 764 3800 796
rect 3760 716 3800 764
rect 3760 684 3764 716
rect 3796 684 3800 716
rect 3760 636 3800 684
rect 3760 604 3764 636
rect 3796 604 3800 636
rect 3760 556 3800 604
rect 3760 524 3764 556
rect 3796 524 3800 556
rect 3760 476 3800 524
rect 3760 444 3764 476
rect 3796 444 3800 476
rect 3760 396 3800 444
rect 3760 364 3764 396
rect 3796 364 3800 396
rect 3760 316 3800 364
rect 3760 284 3764 316
rect 3796 284 3800 316
rect 3760 236 3800 284
rect 3760 204 3764 236
rect 3796 204 3800 236
rect 3760 156 3800 204
rect 3760 124 3764 156
rect 3796 124 3800 156
rect 3760 76 3800 124
rect 3760 44 3764 76
rect 3796 44 3800 76
rect 3760 -4 3800 44
rect 3760 -36 3764 -4
rect 3796 -36 3800 -4
rect 3760 -84 3800 -36
rect 3760 -116 3764 -84
rect 3796 -116 3800 -84
rect 3760 -120 3800 -116
rect 3840 1036 3880 1040
rect 3840 1004 3844 1036
rect 3876 1004 3880 1036
rect 3840 956 3880 1004
rect 3840 924 3844 956
rect 3876 924 3880 956
rect 3840 876 3880 924
rect 3840 844 3844 876
rect 3876 844 3880 876
rect 3840 796 3880 844
rect 3840 764 3844 796
rect 3876 764 3880 796
rect 3840 716 3880 764
rect 3840 684 3844 716
rect 3876 684 3880 716
rect 3840 636 3880 684
rect 3840 604 3844 636
rect 3876 604 3880 636
rect 3840 556 3880 604
rect 3840 524 3844 556
rect 3876 524 3880 556
rect 3840 476 3880 524
rect 3840 444 3844 476
rect 3876 444 3880 476
rect 3840 396 3880 444
rect 3840 364 3844 396
rect 3876 364 3880 396
rect 3840 316 3880 364
rect 3840 284 3844 316
rect 3876 284 3880 316
rect 3840 236 3880 284
rect 3840 204 3844 236
rect 3876 204 3880 236
rect 3840 156 3880 204
rect 3840 124 3844 156
rect 3876 124 3880 156
rect 3840 76 3880 124
rect 3840 44 3844 76
rect 3876 44 3880 76
rect 3840 -4 3880 44
rect 3840 -36 3844 -4
rect 3876 -36 3880 -4
rect 3840 -84 3880 -36
rect 3840 -116 3844 -84
rect 3876 -116 3880 -84
rect 3840 -120 3880 -116
rect 3920 1036 3960 1040
rect 3920 1004 3924 1036
rect 3956 1004 3960 1036
rect 3920 956 3960 1004
rect 3920 924 3924 956
rect 3956 924 3960 956
rect 3920 876 3960 924
rect 3920 844 3924 876
rect 3956 844 3960 876
rect 3920 796 3960 844
rect 3920 764 3924 796
rect 3956 764 3960 796
rect 3920 716 3960 764
rect 3920 684 3924 716
rect 3956 684 3960 716
rect 3920 636 3960 684
rect 3920 604 3924 636
rect 3956 604 3960 636
rect 3920 556 3960 604
rect 3920 524 3924 556
rect 3956 524 3960 556
rect 3920 476 3960 524
rect 3920 444 3924 476
rect 3956 444 3960 476
rect 3920 396 3960 444
rect 3920 364 3924 396
rect 3956 364 3960 396
rect 3920 316 3960 364
rect 3920 284 3924 316
rect 3956 284 3960 316
rect 3920 236 3960 284
rect 3920 204 3924 236
rect 3956 204 3960 236
rect 3920 156 3960 204
rect 3920 124 3924 156
rect 3956 124 3960 156
rect 3920 76 3960 124
rect 3920 44 3924 76
rect 3956 44 3960 76
rect 3920 -4 3960 44
rect 3920 -36 3924 -4
rect 3956 -36 3960 -4
rect 3920 -84 3960 -36
rect 3920 -116 3924 -84
rect 3956 -116 3960 -84
rect 3920 -120 3960 -116
rect 4000 1036 4040 1040
rect 4000 1004 4004 1036
rect 4036 1004 4040 1036
rect 4000 956 4040 1004
rect 4000 924 4004 956
rect 4036 924 4040 956
rect 4000 876 4040 924
rect 4000 844 4004 876
rect 4036 844 4040 876
rect 4000 796 4040 844
rect 4000 764 4004 796
rect 4036 764 4040 796
rect 4000 716 4040 764
rect 4000 684 4004 716
rect 4036 684 4040 716
rect 4000 636 4040 684
rect 4000 604 4004 636
rect 4036 604 4040 636
rect 4000 556 4040 604
rect 4000 524 4004 556
rect 4036 524 4040 556
rect 4000 476 4040 524
rect 4000 444 4004 476
rect 4036 444 4040 476
rect 4000 396 4040 444
rect 4000 364 4004 396
rect 4036 364 4040 396
rect 4000 316 4040 364
rect 4000 284 4004 316
rect 4036 284 4040 316
rect 4000 236 4040 284
rect 4000 204 4004 236
rect 4036 204 4040 236
rect 4000 156 4040 204
rect 4000 124 4004 156
rect 4036 124 4040 156
rect 4000 76 4040 124
rect 4000 44 4004 76
rect 4036 44 4040 76
rect 4000 -4 4040 44
rect 4000 -36 4004 -4
rect 4036 -36 4040 -4
rect 4000 -84 4040 -36
rect 4000 -116 4004 -84
rect 4036 -116 4040 -84
rect 4000 -120 4040 -116
rect 4080 1036 4120 1040
rect 4080 1004 4084 1036
rect 4116 1004 4120 1036
rect 4080 956 4120 1004
rect 4080 924 4084 956
rect 4116 924 4120 956
rect 4080 876 4120 924
rect 4080 844 4084 876
rect 4116 844 4120 876
rect 4080 796 4120 844
rect 4080 764 4084 796
rect 4116 764 4120 796
rect 4080 716 4120 764
rect 4080 684 4084 716
rect 4116 684 4120 716
rect 4080 636 4120 684
rect 4080 604 4084 636
rect 4116 604 4120 636
rect 4080 556 4120 604
rect 4080 524 4084 556
rect 4116 524 4120 556
rect 4080 476 4120 524
rect 4080 444 4084 476
rect 4116 444 4120 476
rect 4080 396 4120 444
rect 4080 364 4084 396
rect 4116 364 4120 396
rect 4080 316 4120 364
rect 4080 284 4084 316
rect 4116 284 4120 316
rect 4080 236 4120 284
rect 4080 204 4084 236
rect 4116 204 4120 236
rect 4080 156 4120 204
rect 4080 124 4084 156
rect 4116 124 4120 156
rect 4080 76 4120 124
rect 4080 44 4084 76
rect 4116 44 4120 76
rect 4080 -4 4120 44
rect 4080 -36 4084 -4
rect 4116 -36 4120 -4
rect 4080 -84 4120 -36
rect 4080 -116 4084 -84
rect 4116 -116 4120 -84
rect 4080 -120 4120 -116
rect 4160 1036 4200 1040
rect 4160 1004 4164 1036
rect 4196 1004 4200 1036
rect 4160 956 4200 1004
rect 4160 924 4164 956
rect 4196 924 4200 956
rect 4160 876 4200 924
rect 4160 844 4164 876
rect 4196 844 4200 876
rect 4160 796 4200 844
rect 4160 764 4164 796
rect 4196 764 4200 796
rect 4160 716 4200 764
rect 4160 684 4164 716
rect 4196 684 4200 716
rect 4160 636 4200 684
rect 4160 604 4164 636
rect 4196 604 4200 636
rect 4160 556 4200 604
rect 4160 524 4164 556
rect 4196 524 4200 556
rect 4160 476 4200 524
rect 4160 444 4164 476
rect 4196 444 4200 476
rect 4160 396 4200 444
rect 4160 364 4164 396
rect 4196 364 4200 396
rect 4160 316 4200 364
rect 4160 284 4164 316
rect 4196 284 4200 316
rect 4160 236 4200 284
rect 4160 204 4164 236
rect 4196 204 4200 236
rect 4160 156 4200 204
rect 4160 124 4164 156
rect 4196 124 4200 156
rect 4160 76 4200 124
rect 4160 44 4164 76
rect 4196 44 4200 76
rect 4160 -4 4200 44
rect 4160 -36 4164 -4
rect 4196 -36 4200 -4
rect 4160 -84 4200 -36
rect 4160 -116 4164 -84
rect 4196 -116 4200 -84
rect 4160 -120 4200 -116
rect 4240 1036 4280 1040
rect 4240 1004 4244 1036
rect 4276 1004 4280 1036
rect 4240 956 4280 1004
rect 4240 924 4244 956
rect 4276 924 4280 956
rect 4240 876 4280 924
rect 4240 844 4244 876
rect 4276 844 4280 876
rect 4240 796 4280 844
rect 4240 764 4244 796
rect 4276 764 4280 796
rect 4240 716 4280 764
rect 4240 684 4244 716
rect 4276 684 4280 716
rect 4240 636 4280 684
rect 4240 604 4244 636
rect 4276 604 4280 636
rect 4240 556 4280 604
rect 4240 524 4244 556
rect 4276 524 4280 556
rect 4240 476 4280 524
rect 4240 444 4244 476
rect 4276 444 4280 476
rect 4240 396 4280 444
rect 4240 364 4244 396
rect 4276 364 4280 396
rect 4240 316 4280 364
rect 4240 284 4244 316
rect 4276 284 4280 316
rect 4240 236 4280 284
rect 4240 204 4244 236
rect 4276 204 4280 236
rect 4240 156 4280 204
rect 4240 124 4244 156
rect 4276 124 4280 156
rect 4240 76 4280 124
rect 4240 44 4244 76
rect 4276 44 4280 76
rect 4240 -4 4280 44
rect 4240 -36 4244 -4
rect 4276 -36 4280 -4
rect 4240 -84 4280 -36
rect 4240 -116 4244 -84
rect 4276 -116 4280 -84
rect 4240 -120 4280 -116
rect 4320 1036 4360 1040
rect 4320 1004 4324 1036
rect 4356 1004 4360 1036
rect 4320 956 4360 1004
rect 4320 924 4324 956
rect 4356 924 4360 956
rect 4320 876 4360 924
rect 4320 844 4324 876
rect 4356 844 4360 876
rect 4320 796 4360 844
rect 4320 764 4324 796
rect 4356 764 4360 796
rect 4320 716 4360 764
rect 4320 684 4324 716
rect 4356 684 4360 716
rect 4320 636 4360 684
rect 4320 604 4324 636
rect 4356 604 4360 636
rect 4320 556 4360 604
rect 4320 524 4324 556
rect 4356 524 4360 556
rect 4320 476 4360 524
rect 4320 444 4324 476
rect 4356 444 4360 476
rect 4320 396 4360 444
rect 4320 364 4324 396
rect 4356 364 4360 396
rect 4320 316 4360 364
rect 4320 284 4324 316
rect 4356 284 4360 316
rect 4320 236 4360 284
rect 4320 204 4324 236
rect 4356 204 4360 236
rect 4320 156 4360 204
rect 4320 124 4324 156
rect 4356 124 4360 156
rect 4320 76 4360 124
rect 4320 44 4324 76
rect 4356 44 4360 76
rect 4320 -4 4360 44
rect 4320 -36 4324 -4
rect 4356 -36 4360 -4
rect 4320 -84 4360 -36
rect 4320 -116 4324 -84
rect 4356 -116 4360 -84
rect 4320 -120 4360 -116
rect 4400 1036 4440 1040
rect 4400 1004 4404 1036
rect 4436 1004 4440 1036
rect 4400 956 4440 1004
rect 4400 924 4404 956
rect 4436 924 4440 956
rect 4400 876 4440 924
rect 4400 844 4404 876
rect 4436 844 4440 876
rect 4400 796 4440 844
rect 4400 764 4404 796
rect 4436 764 4440 796
rect 4400 716 4440 764
rect 4400 684 4404 716
rect 4436 684 4440 716
rect 4400 636 4440 684
rect 4400 604 4404 636
rect 4436 604 4440 636
rect 4400 556 4440 604
rect 4400 524 4404 556
rect 4436 524 4440 556
rect 4400 476 4440 524
rect 4400 444 4404 476
rect 4436 444 4440 476
rect 4400 396 4440 444
rect 4400 364 4404 396
rect 4436 364 4440 396
rect 4400 316 4440 364
rect 4400 284 4404 316
rect 4436 284 4440 316
rect 4400 236 4440 284
rect 4400 204 4404 236
rect 4436 204 4440 236
rect 4400 156 4440 204
rect 4400 124 4404 156
rect 4436 124 4440 156
rect 4400 76 4440 124
rect 4400 44 4404 76
rect 4436 44 4440 76
rect 4400 -4 4440 44
rect 4400 -36 4404 -4
rect 4436 -36 4440 -4
rect 4400 -84 4440 -36
rect 4400 -116 4404 -84
rect 4436 -116 4440 -84
rect 4400 -120 4440 -116
rect 4480 1036 4520 1040
rect 4480 1004 4484 1036
rect 4516 1004 4520 1036
rect 4480 956 4520 1004
rect 4480 924 4484 956
rect 4516 924 4520 956
rect 4480 876 4520 924
rect 4480 844 4484 876
rect 4516 844 4520 876
rect 4480 796 4520 844
rect 4480 764 4484 796
rect 4516 764 4520 796
rect 4480 716 4520 764
rect 4480 684 4484 716
rect 4516 684 4520 716
rect 4480 636 4520 684
rect 4480 604 4484 636
rect 4516 604 4520 636
rect 4480 556 4520 604
rect 4480 524 4484 556
rect 4516 524 4520 556
rect 4480 476 4520 524
rect 4480 444 4484 476
rect 4516 444 4520 476
rect 4480 396 4520 444
rect 4480 364 4484 396
rect 4516 364 4520 396
rect 4480 316 4520 364
rect 4480 284 4484 316
rect 4516 284 4520 316
rect 4480 236 4520 284
rect 4480 204 4484 236
rect 4516 204 4520 236
rect 4480 156 4520 204
rect 4480 124 4484 156
rect 4516 124 4520 156
rect 4480 76 4520 124
rect 4480 44 4484 76
rect 4516 44 4520 76
rect 4480 -4 4520 44
rect 4480 -36 4484 -4
rect 4516 -36 4520 -4
rect 4480 -84 4520 -36
rect 4480 -116 4484 -84
rect 4516 -116 4520 -84
rect 4480 -120 4520 -116
rect 4560 1036 4600 1040
rect 4560 1004 4564 1036
rect 4596 1004 4600 1036
rect 4560 956 4600 1004
rect 4560 924 4564 956
rect 4596 924 4600 956
rect 4560 876 4600 924
rect 4560 844 4564 876
rect 4596 844 4600 876
rect 4560 796 4600 844
rect 4560 764 4564 796
rect 4596 764 4600 796
rect 4560 716 4600 764
rect 4560 684 4564 716
rect 4596 684 4600 716
rect 4560 636 4600 684
rect 4560 604 4564 636
rect 4596 604 4600 636
rect 4560 556 4600 604
rect 4560 524 4564 556
rect 4596 524 4600 556
rect 4560 476 4600 524
rect 4560 444 4564 476
rect 4596 444 4600 476
rect 4560 396 4600 444
rect 4560 364 4564 396
rect 4596 364 4600 396
rect 4560 316 4600 364
rect 4560 284 4564 316
rect 4596 284 4600 316
rect 4560 236 4600 284
rect 4560 204 4564 236
rect 4596 204 4600 236
rect 4560 156 4600 204
rect 4560 124 4564 156
rect 4596 124 4600 156
rect 4560 76 4600 124
rect 4560 44 4564 76
rect 4596 44 4600 76
rect 4560 -4 4600 44
rect 4560 -36 4564 -4
rect 4596 -36 4600 -4
rect 4560 -84 4600 -36
rect 4560 -116 4564 -84
rect 4596 -116 4600 -84
rect 4560 -120 4600 -116
rect 4640 1036 4680 1040
rect 4640 1004 4644 1036
rect 4676 1004 4680 1036
rect 4640 956 4680 1004
rect 4640 924 4644 956
rect 4676 924 4680 956
rect 4640 876 4680 924
rect 4640 844 4644 876
rect 4676 844 4680 876
rect 4640 796 4680 844
rect 4640 764 4644 796
rect 4676 764 4680 796
rect 4640 716 4680 764
rect 4640 684 4644 716
rect 4676 684 4680 716
rect 4640 636 4680 684
rect 4640 604 4644 636
rect 4676 604 4680 636
rect 4640 556 4680 604
rect 4640 524 4644 556
rect 4676 524 4680 556
rect 4640 476 4680 524
rect 4640 444 4644 476
rect 4676 444 4680 476
rect 4640 396 4680 444
rect 4640 364 4644 396
rect 4676 364 4680 396
rect 4640 316 4680 364
rect 4640 284 4644 316
rect 4676 284 4680 316
rect 4640 236 4680 284
rect 4640 204 4644 236
rect 4676 204 4680 236
rect 4640 156 4680 204
rect 4640 124 4644 156
rect 4676 124 4680 156
rect 4640 76 4680 124
rect 4640 44 4644 76
rect 4676 44 4680 76
rect 4640 -4 4680 44
rect 4640 -36 4644 -4
rect 4676 -36 4680 -4
rect 4640 -84 4680 -36
rect 4640 -116 4644 -84
rect 4676 -116 4680 -84
rect 4640 -120 4680 -116
rect 4720 1036 4760 1040
rect 4720 1004 4724 1036
rect 4756 1004 4760 1036
rect 4720 956 4760 1004
rect 4720 924 4724 956
rect 4756 924 4760 956
rect 4720 876 4760 924
rect 4720 844 4724 876
rect 4756 844 4760 876
rect 4720 796 4760 844
rect 4720 764 4724 796
rect 4756 764 4760 796
rect 4720 716 4760 764
rect 4720 684 4724 716
rect 4756 684 4760 716
rect 4720 636 4760 684
rect 4720 604 4724 636
rect 4756 604 4760 636
rect 4720 556 4760 604
rect 4720 524 4724 556
rect 4756 524 4760 556
rect 4720 476 4760 524
rect 4720 444 4724 476
rect 4756 444 4760 476
rect 4720 396 4760 444
rect 4720 364 4724 396
rect 4756 364 4760 396
rect 4720 316 4760 364
rect 4720 284 4724 316
rect 4756 284 4760 316
rect 4720 236 4760 284
rect 4720 204 4724 236
rect 4756 204 4760 236
rect 4720 156 4760 204
rect 4720 124 4724 156
rect 4756 124 4760 156
rect 4720 76 4760 124
rect 4720 44 4724 76
rect 4756 44 4760 76
rect 4720 -4 4760 44
rect 4720 -36 4724 -4
rect 4756 -36 4760 -4
rect 4720 -84 4760 -36
rect 4720 -116 4724 -84
rect 4756 -116 4760 -84
rect 4720 -120 4760 -116
rect 4800 1036 4840 1040
rect 4800 1004 4804 1036
rect 4836 1004 4840 1036
rect 4800 956 4840 1004
rect 4800 924 4804 956
rect 4836 924 4840 956
rect 4800 876 4840 924
rect 4800 844 4804 876
rect 4836 844 4840 876
rect 4800 796 4840 844
rect 4800 764 4804 796
rect 4836 764 4840 796
rect 4800 716 4840 764
rect 4800 684 4804 716
rect 4836 684 4840 716
rect 4800 636 4840 684
rect 4800 604 4804 636
rect 4836 604 4840 636
rect 4800 556 4840 604
rect 4800 524 4804 556
rect 4836 524 4840 556
rect 4800 476 4840 524
rect 4800 444 4804 476
rect 4836 444 4840 476
rect 4800 396 4840 444
rect 4800 364 4804 396
rect 4836 364 4840 396
rect 4800 316 4840 364
rect 4800 284 4804 316
rect 4836 284 4840 316
rect 4800 236 4840 284
rect 4800 204 4804 236
rect 4836 204 4840 236
rect 4800 156 4840 204
rect 4800 124 4804 156
rect 4836 124 4840 156
rect 4800 76 4840 124
rect 4800 44 4804 76
rect 4836 44 4840 76
rect 4800 -4 4840 44
rect 4800 -36 4804 -4
rect 4836 -36 4840 -4
rect 4800 -84 4840 -36
rect 4800 -116 4804 -84
rect 4836 -116 4840 -84
rect 4800 -120 4840 -116
rect 4880 1036 4920 1040
rect 4880 1004 4884 1036
rect 4916 1004 4920 1036
rect 4880 956 4920 1004
rect 4880 924 4884 956
rect 4916 924 4920 956
rect 4880 876 4920 924
rect 4880 844 4884 876
rect 4916 844 4920 876
rect 4880 796 4920 844
rect 4880 764 4884 796
rect 4916 764 4920 796
rect 4880 716 4920 764
rect 4880 684 4884 716
rect 4916 684 4920 716
rect 4880 636 4920 684
rect 4880 604 4884 636
rect 4916 604 4920 636
rect 4880 556 4920 604
rect 4880 524 4884 556
rect 4916 524 4920 556
rect 4880 476 4920 524
rect 4880 444 4884 476
rect 4916 444 4920 476
rect 4880 396 4920 444
rect 4880 364 4884 396
rect 4916 364 4920 396
rect 4880 316 4920 364
rect 4880 284 4884 316
rect 4916 284 4920 316
rect 4880 236 4920 284
rect 4880 204 4884 236
rect 4916 204 4920 236
rect 4880 156 4920 204
rect 4880 124 4884 156
rect 4916 124 4920 156
rect 4880 76 4920 124
rect 4880 44 4884 76
rect 4916 44 4920 76
rect 4880 -4 4920 44
rect 4880 -36 4884 -4
rect 4916 -36 4920 -4
rect 4880 -84 4920 -36
rect 4880 -116 4884 -84
rect 4916 -116 4920 -84
rect 4880 -120 4920 -116
rect 4960 1036 5000 1040
rect 4960 1004 4964 1036
rect 4996 1004 5000 1036
rect 4960 956 5000 1004
rect 4960 924 4964 956
rect 4996 924 5000 956
rect 4960 876 5000 924
rect 4960 844 4964 876
rect 4996 844 5000 876
rect 4960 796 5000 844
rect 4960 764 4964 796
rect 4996 764 5000 796
rect 4960 716 5000 764
rect 4960 684 4964 716
rect 4996 684 5000 716
rect 4960 636 5000 684
rect 4960 604 4964 636
rect 4996 604 5000 636
rect 4960 556 5000 604
rect 4960 524 4964 556
rect 4996 524 5000 556
rect 4960 476 5000 524
rect 4960 444 4964 476
rect 4996 444 5000 476
rect 4960 396 5000 444
rect 4960 364 4964 396
rect 4996 364 5000 396
rect 4960 316 5000 364
rect 4960 284 4964 316
rect 4996 284 5000 316
rect 4960 236 5000 284
rect 4960 204 4964 236
rect 4996 204 5000 236
rect 4960 156 5000 204
rect 4960 124 4964 156
rect 4996 124 5000 156
rect 4960 76 5000 124
rect 4960 44 4964 76
rect 4996 44 5000 76
rect 4960 -4 5000 44
rect 4960 -36 4964 -4
rect 4996 -36 5000 -4
rect 4960 -84 5000 -36
rect 4960 -116 4964 -84
rect 4996 -116 5000 -84
rect 4960 -120 5000 -116
rect 5040 1036 5080 1040
rect 5040 1004 5044 1036
rect 5076 1004 5080 1036
rect 5040 956 5080 1004
rect 5040 924 5044 956
rect 5076 924 5080 956
rect 5040 876 5080 924
rect 5040 844 5044 876
rect 5076 844 5080 876
rect 5040 796 5080 844
rect 5040 764 5044 796
rect 5076 764 5080 796
rect 5040 716 5080 764
rect 5040 684 5044 716
rect 5076 684 5080 716
rect 5040 636 5080 684
rect 5040 604 5044 636
rect 5076 604 5080 636
rect 5040 556 5080 604
rect 5040 524 5044 556
rect 5076 524 5080 556
rect 5040 476 5080 524
rect 5040 444 5044 476
rect 5076 444 5080 476
rect 5040 396 5080 444
rect 5040 364 5044 396
rect 5076 364 5080 396
rect 5040 316 5080 364
rect 5040 284 5044 316
rect 5076 284 5080 316
rect 5040 236 5080 284
rect 5040 204 5044 236
rect 5076 204 5080 236
rect 5040 156 5080 204
rect 5040 124 5044 156
rect 5076 124 5080 156
rect 5040 76 5080 124
rect 5040 44 5044 76
rect 5076 44 5080 76
rect 5040 -4 5080 44
rect 5040 -36 5044 -4
rect 5076 -36 5080 -4
rect 5040 -84 5080 -36
rect 5040 -116 5044 -84
rect 5076 -116 5080 -84
rect 5040 -120 5080 -116
rect 5120 1036 5160 1040
rect 5120 1004 5124 1036
rect 5156 1004 5160 1036
rect 5120 956 5160 1004
rect 5120 924 5124 956
rect 5156 924 5160 956
rect 5120 876 5160 924
rect 5120 844 5124 876
rect 5156 844 5160 876
rect 5120 796 5160 844
rect 5120 764 5124 796
rect 5156 764 5160 796
rect 5120 716 5160 764
rect 5120 684 5124 716
rect 5156 684 5160 716
rect 5120 636 5160 684
rect 5120 604 5124 636
rect 5156 604 5160 636
rect 5120 556 5160 604
rect 5120 524 5124 556
rect 5156 524 5160 556
rect 5120 476 5160 524
rect 5120 444 5124 476
rect 5156 444 5160 476
rect 5120 396 5160 444
rect 5120 364 5124 396
rect 5156 364 5160 396
rect 5120 316 5160 364
rect 5120 284 5124 316
rect 5156 284 5160 316
rect 5120 236 5160 284
rect 5120 204 5124 236
rect 5156 204 5160 236
rect 5120 156 5160 204
rect 5120 124 5124 156
rect 5156 124 5160 156
rect 5120 76 5160 124
rect 5120 44 5124 76
rect 5156 44 5160 76
rect 5120 -4 5160 44
rect 5120 -36 5124 -4
rect 5156 -36 5160 -4
rect 5120 -84 5160 -36
rect 5120 -116 5124 -84
rect 5156 -116 5160 -84
rect 5120 -120 5160 -116
rect 5200 1036 5240 1040
rect 5200 1004 5204 1036
rect 5236 1004 5240 1036
rect 5200 956 5240 1004
rect 5200 924 5204 956
rect 5236 924 5240 956
rect 5200 876 5240 924
rect 5200 844 5204 876
rect 5236 844 5240 876
rect 5200 796 5240 844
rect 5200 764 5204 796
rect 5236 764 5240 796
rect 5200 716 5240 764
rect 5200 684 5204 716
rect 5236 684 5240 716
rect 5200 636 5240 684
rect 5200 604 5204 636
rect 5236 604 5240 636
rect 5200 556 5240 604
rect 5200 524 5204 556
rect 5236 524 5240 556
rect 5200 476 5240 524
rect 5200 444 5204 476
rect 5236 444 5240 476
rect 5200 396 5240 444
rect 5200 364 5204 396
rect 5236 364 5240 396
rect 5200 316 5240 364
rect 5200 284 5204 316
rect 5236 284 5240 316
rect 5200 236 5240 284
rect 5200 204 5204 236
rect 5236 204 5240 236
rect 5200 156 5240 204
rect 5200 124 5204 156
rect 5236 124 5240 156
rect 5200 76 5240 124
rect 5200 44 5204 76
rect 5236 44 5240 76
rect 5200 -4 5240 44
rect 5200 -36 5204 -4
rect 5236 -36 5240 -4
rect 5200 -84 5240 -36
rect 5200 -116 5204 -84
rect 5236 -116 5240 -84
rect 5200 -120 5240 -116
rect 5280 1036 5320 1040
rect 5280 1004 5284 1036
rect 5316 1004 5320 1036
rect 5280 956 5320 1004
rect 5280 924 5284 956
rect 5316 924 5320 956
rect 5280 876 5320 924
rect 5280 844 5284 876
rect 5316 844 5320 876
rect 5280 796 5320 844
rect 5280 764 5284 796
rect 5316 764 5320 796
rect 5280 716 5320 764
rect 5280 684 5284 716
rect 5316 684 5320 716
rect 5280 636 5320 684
rect 5280 604 5284 636
rect 5316 604 5320 636
rect 5280 556 5320 604
rect 5280 524 5284 556
rect 5316 524 5320 556
rect 5280 476 5320 524
rect 5280 444 5284 476
rect 5316 444 5320 476
rect 5280 396 5320 444
rect 5280 364 5284 396
rect 5316 364 5320 396
rect 5280 316 5320 364
rect 5280 284 5284 316
rect 5316 284 5320 316
rect 5280 236 5320 284
rect 5280 204 5284 236
rect 5316 204 5320 236
rect 5280 156 5320 204
rect 5280 124 5284 156
rect 5316 124 5320 156
rect 5280 76 5320 124
rect 5280 44 5284 76
rect 5316 44 5320 76
rect 5280 -4 5320 44
rect 5280 -36 5284 -4
rect 5316 -36 5320 -4
rect 5280 -84 5320 -36
rect 5280 -116 5284 -84
rect 5316 -116 5320 -84
rect 5280 -120 5320 -116
rect 5360 1036 5400 1040
rect 5360 1004 5364 1036
rect 5396 1004 5400 1036
rect 5360 956 5400 1004
rect 5360 924 5364 956
rect 5396 924 5400 956
rect 5360 876 5400 924
rect 5360 844 5364 876
rect 5396 844 5400 876
rect 5360 796 5400 844
rect 5360 764 5364 796
rect 5396 764 5400 796
rect 5360 716 5400 764
rect 5360 684 5364 716
rect 5396 684 5400 716
rect 5360 636 5400 684
rect 5360 604 5364 636
rect 5396 604 5400 636
rect 5360 556 5400 604
rect 5360 524 5364 556
rect 5396 524 5400 556
rect 5360 476 5400 524
rect 5360 444 5364 476
rect 5396 444 5400 476
rect 5360 396 5400 444
rect 5360 364 5364 396
rect 5396 364 5400 396
rect 5360 316 5400 364
rect 5360 284 5364 316
rect 5396 284 5400 316
rect 5360 236 5400 284
rect 5360 204 5364 236
rect 5396 204 5400 236
rect 5360 156 5400 204
rect 5360 124 5364 156
rect 5396 124 5400 156
rect 5360 76 5400 124
rect 5360 44 5364 76
rect 5396 44 5400 76
rect 5360 -4 5400 44
rect 5360 -36 5364 -4
rect 5396 -36 5400 -4
rect 5360 -84 5400 -36
rect 5360 -116 5364 -84
rect 5396 -116 5400 -84
rect 5360 -120 5400 -116
rect 5440 1036 5480 1040
rect 5440 1004 5444 1036
rect 5476 1004 5480 1036
rect 5440 956 5480 1004
rect 5440 924 5444 956
rect 5476 924 5480 956
rect 5440 876 5480 924
rect 5440 844 5444 876
rect 5476 844 5480 876
rect 5440 796 5480 844
rect 5440 764 5444 796
rect 5476 764 5480 796
rect 5440 716 5480 764
rect 5440 684 5444 716
rect 5476 684 5480 716
rect 5440 636 5480 684
rect 5440 604 5444 636
rect 5476 604 5480 636
rect 5440 556 5480 604
rect 5440 524 5444 556
rect 5476 524 5480 556
rect 5440 476 5480 524
rect 5440 444 5444 476
rect 5476 444 5480 476
rect 5440 396 5480 444
rect 5440 364 5444 396
rect 5476 364 5480 396
rect 5440 316 5480 364
rect 5440 284 5444 316
rect 5476 284 5480 316
rect 5440 236 5480 284
rect 5440 204 5444 236
rect 5476 204 5480 236
rect 5440 156 5480 204
rect 5440 124 5444 156
rect 5476 124 5480 156
rect 5440 76 5480 124
rect 5440 44 5444 76
rect 5476 44 5480 76
rect 5440 -4 5480 44
rect 5440 -36 5444 -4
rect 5476 -36 5480 -4
rect 5440 -84 5480 -36
rect 5440 -116 5444 -84
rect 5476 -116 5480 -84
rect 5440 -120 5480 -116
rect 5520 1036 5560 1040
rect 5520 1004 5524 1036
rect 5556 1004 5560 1036
rect 5520 956 5560 1004
rect 5520 924 5524 956
rect 5556 924 5560 956
rect 5520 876 5560 924
rect 5520 844 5524 876
rect 5556 844 5560 876
rect 5520 796 5560 844
rect 5520 764 5524 796
rect 5556 764 5560 796
rect 5520 716 5560 764
rect 5520 684 5524 716
rect 5556 684 5560 716
rect 5520 636 5560 684
rect 5520 604 5524 636
rect 5556 604 5560 636
rect 5520 556 5560 604
rect 5520 524 5524 556
rect 5556 524 5560 556
rect 5520 476 5560 524
rect 5520 444 5524 476
rect 5556 444 5560 476
rect 5520 396 5560 444
rect 5520 364 5524 396
rect 5556 364 5560 396
rect 5520 316 5560 364
rect 5520 284 5524 316
rect 5556 284 5560 316
rect 5520 236 5560 284
rect 5520 204 5524 236
rect 5556 204 5560 236
rect 5520 156 5560 204
rect 5520 124 5524 156
rect 5556 124 5560 156
rect 5520 76 5560 124
rect 5520 44 5524 76
rect 5556 44 5560 76
rect 5520 -4 5560 44
rect 5520 -36 5524 -4
rect 5556 -36 5560 -4
rect 5520 -84 5560 -36
rect 5520 -116 5524 -84
rect 5556 -116 5560 -84
rect 5520 -120 5560 -116
rect 5600 1036 5640 1040
rect 5600 1004 5604 1036
rect 5636 1004 5640 1036
rect 5600 956 5640 1004
rect 5600 924 5604 956
rect 5636 924 5640 956
rect 5600 876 5640 924
rect 5600 844 5604 876
rect 5636 844 5640 876
rect 5600 796 5640 844
rect 5600 764 5604 796
rect 5636 764 5640 796
rect 5600 716 5640 764
rect 5600 684 5604 716
rect 5636 684 5640 716
rect 5600 636 5640 684
rect 5600 604 5604 636
rect 5636 604 5640 636
rect 5600 556 5640 604
rect 5600 524 5604 556
rect 5636 524 5640 556
rect 5600 476 5640 524
rect 5600 444 5604 476
rect 5636 444 5640 476
rect 5600 396 5640 444
rect 5600 364 5604 396
rect 5636 364 5640 396
rect 5600 316 5640 364
rect 5600 284 5604 316
rect 5636 284 5640 316
rect 5600 236 5640 284
rect 5600 204 5604 236
rect 5636 204 5640 236
rect 5600 156 5640 204
rect 5600 124 5604 156
rect 5636 124 5640 156
rect 5600 76 5640 124
rect 5600 44 5604 76
rect 5636 44 5640 76
rect 5600 -4 5640 44
rect 5600 -36 5604 -4
rect 5636 -36 5640 -4
rect 5600 -84 5640 -36
rect 5600 -116 5604 -84
rect 5636 -116 5640 -84
rect 5600 -120 5640 -116
rect 5680 1036 5720 1040
rect 5680 1004 5684 1036
rect 5716 1004 5720 1036
rect 5680 956 5720 1004
rect 5680 924 5684 956
rect 5716 924 5720 956
rect 5680 876 5720 924
rect 5680 844 5684 876
rect 5716 844 5720 876
rect 5680 796 5720 844
rect 5680 764 5684 796
rect 5716 764 5720 796
rect 5680 716 5720 764
rect 5680 684 5684 716
rect 5716 684 5720 716
rect 5680 636 5720 684
rect 5680 604 5684 636
rect 5716 604 5720 636
rect 5680 556 5720 604
rect 5680 524 5684 556
rect 5716 524 5720 556
rect 5680 476 5720 524
rect 5680 444 5684 476
rect 5716 444 5720 476
rect 5680 396 5720 444
rect 5680 364 5684 396
rect 5716 364 5720 396
rect 5680 316 5720 364
rect 5680 284 5684 316
rect 5716 284 5720 316
rect 5680 236 5720 284
rect 5680 204 5684 236
rect 5716 204 5720 236
rect 5680 156 5720 204
rect 5680 124 5684 156
rect 5716 124 5720 156
rect 5680 76 5720 124
rect 5680 44 5684 76
rect 5716 44 5720 76
rect 5680 -4 5720 44
rect 5680 -36 5684 -4
rect 5716 -36 5720 -4
rect 5680 -84 5720 -36
rect 5680 -116 5684 -84
rect 5716 -116 5720 -84
rect 5680 -120 5720 -116
rect 5760 1036 5800 1040
rect 5760 1004 5764 1036
rect 5796 1004 5800 1036
rect 5760 956 5800 1004
rect 5760 924 5764 956
rect 5796 924 5800 956
rect 5760 876 5800 924
rect 5760 844 5764 876
rect 5796 844 5800 876
rect 5760 796 5800 844
rect 5760 764 5764 796
rect 5796 764 5800 796
rect 5760 716 5800 764
rect 5760 684 5764 716
rect 5796 684 5800 716
rect 5760 636 5800 684
rect 5760 604 5764 636
rect 5796 604 5800 636
rect 5760 556 5800 604
rect 5760 524 5764 556
rect 5796 524 5800 556
rect 5760 476 5800 524
rect 5760 444 5764 476
rect 5796 444 5800 476
rect 5760 396 5800 444
rect 5760 364 5764 396
rect 5796 364 5800 396
rect 5760 316 5800 364
rect 5760 284 5764 316
rect 5796 284 5800 316
rect 5760 236 5800 284
rect 5760 204 5764 236
rect 5796 204 5800 236
rect 5760 156 5800 204
rect 5760 124 5764 156
rect 5796 124 5800 156
rect 5760 76 5800 124
rect 5760 44 5764 76
rect 5796 44 5800 76
rect 5760 -4 5800 44
rect 5760 -36 5764 -4
rect 5796 -36 5800 -4
rect 5760 -84 5800 -36
rect 5760 -116 5764 -84
rect 5796 -116 5800 -84
rect 5760 -120 5800 -116
rect 5840 1036 5880 1040
rect 5840 1004 5844 1036
rect 5876 1004 5880 1036
rect 5840 956 5880 1004
rect 5840 924 5844 956
rect 5876 924 5880 956
rect 5840 876 5880 924
rect 5840 844 5844 876
rect 5876 844 5880 876
rect 5840 796 5880 844
rect 5840 764 5844 796
rect 5876 764 5880 796
rect 5840 716 5880 764
rect 5840 684 5844 716
rect 5876 684 5880 716
rect 5840 636 5880 684
rect 5840 604 5844 636
rect 5876 604 5880 636
rect 5840 556 5880 604
rect 5840 524 5844 556
rect 5876 524 5880 556
rect 5840 476 5880 524
rect 5840 444 5844 476
rect 5876 444 5880 476
rect 5840 396 5880 444
rect 5840 364 5844 396
rect 5876 364 5880 396
rect 5840 316 5880 364
rect 5840 284 5844 316
rect 5876 284 5880 316
rect 5840 236 5880 284
rect 5840 204 5844 236
rect 5876 204 5880 236
rect 5840 156 5880 204
rect 5840 124 5844 156
rect 5876 124 5880 156
rect 5840 76 5880 124
rect 5840 44 5844 76
rect 5876 44 5880 76
rect 5840 -4 5880 44
rect 5840 -36 5844 -4
rect 5876 -36 5880 -4
rect 5840 -84 5880 -36
rect 5840 -116 5844 -84
rect 5876 -116 5880 -84
rect 5840 -120 5880 -116
rect 5920 1036 5960 1040
rect 5920 1004 5924 1036
rect 5956 1004 5960 1036
rect 5920 956 5960 1004
rect 5920 924 5924 956
rect 5956 924 5960 956
rect 5920 876 5960 924
rect 5920 844 5924 876
rect 5956 844 5960 876
rect 5920 796 5960 844
rect 5920 764 5924 796
rect 5956 764 5960 796
rect 5920 716 5960 764
rect 5920 684 5924 716
rect 5956 684 5960 716
rect 5920 636 5960 684
rect 5920 604 5924 636
rect 5956 604 5960 636
rect 5920 556 5960 604
rect 5920 524 5924 556
rect 5956 524 5960 556
rect 5920 476 5960 524
rect 5920 444 5924 476
rect 5956 444 5960 476
rect 5920 396 5960 444
rect 5920 364 5924 396
rect 5956 364 5960 396
rect 5920 316 5960 364
rect 5920 284 5924 316
rect 5956 284 5960 316
rect 5920 236 5960 284
rect 5920 204 5924 236
rect 5956 204 5960 236
rect 5920 156 5960 204
rect 5920 124 5924 156
rect 5956 124 5960 156
rect 5920 76 5960 124
rect 5920 44 5924 76
rect 5956 44 5960 76
rect 5920 -4 5960 44
rect 5920 -36 5924 -4
rect 5956 -36 5960 -4
rect 5920 -84 5960 -36
rect 5920 -116 5924 -84
rect 5956 -116 5960 -84
rect 5920 -120 5960 -116
rect 6000 1036 6040 1040
rect 6000 1004 6004 1036
rect 6036 1004 6040 1036
rect 6000 956 6040 1004
rect 6000 924 6004 956
rect 6036 924 6040 956
rect 6000 876 6040 924
rect 6000 844 6004 876
rect 6036 844 6040 876
rect 6000 796 6040 844
rect 6000 764 6004 796
rect 6036 764 6040 796
rect 6000 716 6040 764
rect 6000 684 6004 716
rect 6036 684 6040 716
rect 6000 636 6040 684
rect 6000 604 6004 636
rect 6036 604 6040 636
rect 6000 556 6040 604
rect 6000 524 6004 556
rect 6036 524 6040 556
rect 6000 476 6040 524
rect 6000 444 6004 476
rect 6036 444 6040 476
rect 6000 396 6040 444
rect 6000 364 6004 396
rect 6036 364 6040 396
rect 6000 316 6040 364
rect 6000 284 6004 316
rect 6036 284 6040 316
rect 6000 236 6040 284
rect 6000 204 6004 236
rect 6036 204 6040 236
rect 6000 156 6040 204
rect 6000 124 6004 156
rect 6036 124 6040 156
rect 6000 76 6040 124
rect 6000 44 6004 76
rect 6036 44 6040 76
rect 6000 -4 6040 44
rect 6000 -36 6004 -4
rect 6036 -36 6040 -4
rect 6000 -84 6040 -36
rect 6000 -116 6004 -84
rect 6036 -116 6040 -84
rect 6000 -120 6040 -116
rect 6080 1036 6120 1040
rect 6080 1004 6084 1036
rect 6116 1004 6120 1036
rect 6080 956 6120 1004
rect 6080 924 6084 956
rect 6116 924 6120 956
rect 6080 876 6120 924
rect 6080 844 6084 876
rect 6116 844 6120 876
rect 6080 796 6120 844
rect 6080 764 6084 796
rect 6116 764 6120 796
rect 6080 716 6120 764
rect 6080 684 6084 716
rect 6116 684 6120 716
rect 6080 636 6120 684
rect 6080 604 6084 636
rect 6116 604 6120 636
rect 6080 556 6120 604
rect 6080 524 6084 556
rect 6116 524 6120 556
rect 6080 476 6120 524
rect 6080 444 6084 476
rect 6116 444 6120 476
rect 6080 396 6120 444
rect 6080 364 6084 396
rect 6116 364 6120 396
rect 6080 316 6120 364
rect 6080 284 6084 316
rect 6116 284 6120 316
rect 6080 236 6120 284
rect 6080 204 6084 236
rect 6116 204 6120 236
rect 6080 156 6120 204
rect 6080 124 6084 156
rect 6116 124 6120 156
rect 6080 76 6120 124
rect 6080 44 6084 76
rect 6116 44 6120 76
rect 6080 -4 6120 44
rect 6080 -36 6084 -4
rect 6116 -36 6120 -4
rect 6080 -84 6120 -36
rect 6080 -116 6084 -84
rect 6116 -116 6120 -84
rect 6080 -120 6120 -116
rect 6160 1036 6200 1040
rect 6160 1004 6164 1036
rect 6196 1004 6200 1036
rect 6160 956 6200 1004
rect 6160 924 6164 956
rect 6196 924 6200 956
rect 6160 876 6200 924
rect 6160 844 6164 876
rect 6196 844 6200 876
rect 6160 796 6200 844
rect 6160 764 6164 796
rect 6196 764 6200 796
rect 6160 716 6200 764
rect 6160 684 6164 716
rect 6196 684 6200 716
rect 6160 636 6200 684
rect 6160 604 6164 636
rect 6196 604 6200 636
rect 6160 556 6200 604
rect 6160 524 6164 556
rect 6196 524 6200 556
rect 6160 476 6200 524
rect 6160 444 6164 476
rect 6196 444 6200 476
rect 6160 396 6200 444
rect 6160 364 6164 396
rect 6196 364 6200 396
rect 6160 316 6200 364
rect 6160 284 6164 316
rect 6196 284 6200 316
rect 6160 236 6200 284
rect 6160 204 6164 236
rect 6196 204 6200 236
rect 6160 156 6200 204
rect 6160 124 6164 156
rect 6196 124 6200 156
rect 6160 76 6200 124
rect 6160 44 6164 76
rect 6196 44 6200 76
rect 6160 -4 6200 44
rect 6160 -36 6164 -4
rect 6196 -36 6200 -4
rect 6160 -84 6200 -36
rect 6160 -116 6164 -84
rect 6196 -116 6200 -84
rect 6160 -120 6200 -116
rect 6240 1036 6280 1040
rect 6240 1004 6244 1036
rect 6276 1004 6280 1036
rect 6240 956 6280 1004
rect 6240 924 6244 956
rect 6276 924 6280 956
rect 6240 876 6280 924
rect 6240 844 6244 876
rect 6276 844 6280 876
rect 6240 796 6280 844
rect 6240 764 6244 796
rect 6276 764 6280 796
rect 6240 716 6280 764
rect 6240 684 6244 716
rect 6276 684 6280 716
rect 6240 636 6280 684
rect 6240 604 6244 636
rect 6276 604 6280 636
rect 6240 556 6280 604
rect 6240 524 6244 556
rect 6276 524 6280 556
rect 6240 476 6280 524
rect 6240 444 6244 476
rect 6276 444 6280 476
rect 6240 396 6280 444
rect 6240 364 6244 396
rect 6276 364 6280 396
rect 6240 316 6280 364
rect 6240 284 6244 316
rect 6276 284 6280 316
rect 6240 236 6280 284
rect 6240 204 6244 236
rect 6276 204 6280 236
rect 6240 156 6280 204
rect 6240 124 6244 156
rect 6276 124 6280 156
rect 6240 76 6280 124
rect 6240 44 6244 76
rect 6276 44 6280 76
rect 6240 -4 6280 44
rect 6240 -36 6244 -4
rect 6276 -36 6280 -4
rect 6240 -84 6280 -36
rect 6240 -116 6244 -84
rect 6276 -116 6280 -84
rect 6240 -120 6280 -116
rect 6320 1036 6360 1040
rect 6320 1004 6324 1036
rect 6356 1004 6360 1036
rect 6320 956 6360 1004
rect 6320 924 6324 956
rect 6356 924 6360 956
rect 6320 876 6360 924
rect 6320 844 6324 876
rect 6356 844 6360 876
rect 6320 796 6360 844
rect 6320 764 6324 796
rect 6356 764 6360 796
rect 6320 716 6360 764
rect 6320 684 6324 716
rect 6356 684 6360 716
rect 6320 636 6360 684
rect 6320 604 6324 636
rect 6356 604 6360 636
rect 6320 556 6360 604
rect 6320 524 6324 556
rect 6356 524 6360 556
rect 6320 476 6360 524
rect 6320 444 6324 476
rect 6356 444 6360 476
rect 6320 396 6360 444
rect 6320 364 6324 396
rect 6356 364 6360 396
rect 6320 316 6360 364
rect 6320 284 6324 316
rect 6356 284 6360 316
rect 6320 236 6360 284
rect 6320 204 6324 236
rect 6356 204 6360 236
rect 6320 156 6360 204
rect 6320 124 6324 156
rect 6356 124 6360 156
rect 6320 76 6360 124
rect 6320 44 6324 76
rect 6356 44 6360 76
rect 6320 -4 6360 44
rect 6320 -36 6324 -4
rect 6356 -36 6360 -4
rect 6320 -84 6360 -36
rect 6320 -116 6324 -84
rect 6356 -116 6360 -84
rect 6320 -120 6360 -116
rect 6400 1036 6440 1040
rect 6400 1004 6404 1036
rect 6436 1004 6440 1036
rect 6400 956 6440 1004
rect 6400 924 6404 956
rect 6436 924 6440 956
rect 6400 876 6440 924
rect 6400 844 6404 876
rect 6436 844 6440 876
rect 6400 796 6440 844
rect 6400 764 6404 796
rect 6436 764 6440 796
rect 6400 716 6440 764
rect 6400 684 6404 716
rect 6436 684 6440 716
rect 6400 636 6440 684
rect 6400 604 6404 636
rect 6436 604 6440 636
rect 6400 556 6440 604
rect 6400 524 6404 556
rect 6436 524 6440 556
rect 6400 476 6440 524
rect 6400 444 6404 476
rect 6436 444 6440 476
rect 6400 396 6440 444
rect 6400 364 6404 396
rect 6436 364 6440 396
rect 6400 316 6440 364
rect 6400 284 6404 316
rect 6436 284 6440 316
rect 6400 236 6440 284
rect 6400 204 6404 236
rect 6436 204 6440 236
rect 6400 156 6440 204
rect 6400 124 6404 156
rect 6436 124 6440 156
rect 6400 76 6440 124
rect 6400 44 6404 76
rect 6436 44 6440 76
rect 6400 -4 6440 44
rect 6400 -36 6404 -4
rect 6436 -36 6440 -4
rect 6400 -84 6440 -36
rect 6400 -116 6404 -84
rect 6436 -116 6440 -84
rect 6400 -120 6440 -116
rect 6480 1036 6520 1040
rect 6480 1004 6484 1036
rect 6516 1004 6520 1036
rect 6480 956 6520 1004
rect 6480 924 6484 956
rect 6516 924 6520 956
rect 6480 876 6520 924
rect 6480 844 6484 876
rect 6516 844 6520 876
rect 6480 796 6520 844
rect 6480 764 6484 796
rect 6516 764 6520 796
rect 6480 716 6520 764
rect 6480 684 6484 716
rect 6516 684 6520 716
rect 6480 636 6520 684
rect 6480 604 6484 636
rect 6516 604 6520 636
rect 6480 556 6520 604
rect 6480 524 6484 556
rect 6516 524 6520 556
rect 6480 476 6520 524
rect 6480 444 6484 476
rect 6516 444 6520 476
rect 6480 396 6520 444
rect 6480 364 6484 396
rect 6516 364 6520 396
rect 6480 316 6520 364
rect 6480 284 6484 316
rect 6516 284 6520 316
rect 6480 236 6520 284
rect 6480 204 6484 236
rect 6516 204 6520 236
rect 6480 156 6520 204
rect 6480 124 6484 156
rect 6516 124 6520 156
rect 6480 76 6520 124
rect 6480 44 6484 76
rect 6516 44 6520 76
rect 6480 -4 6520 44
rect 6480 -36 6484 -4
rect 6516 -36 6520 -4
rect 6480 -84 6520 -36
rect 6480 -116 6484 -84
rect 6516 -116 6520 -84
rect 6480 -120 6520 -116
rect 6560 1036 6600 1040
rect 6560 1004 6564 1036
rect 6596 1004 6600 1036
rect 6560 956 6600 1004
rect 6560 924 6564 956
rect 6596 924 6600 956
rect 6560 876 6600 924
rect 6560 844 6564 876
rect 6596 844 6600 876
rect 6560 796 6600 844
rect 6560 764 6564 796
rect 6596 764 6600 796
rect 6560 716 6600 764
rect 6560 684 6564 716
rect 6596 684 6600 716
rect 6560 636 6600 684
rect 6560 604 6564 636
rect 6596 604 6600 636
rect 6560 556 6600 604
rect 6560 524 6564 556
rect 6596 524 6600 556
rect 6560 476 6600 524
rect 6560 444 6564 476
rect 6596 444 6600 476
rect 6560 396 6600 444
rect 6560 364 6564 396
rect 6596 364 6600 396
rect 6560 316 6600 364
rect 6560 284 6564 316
rect 6596 284 6600 316
rect 6560 236 6600 284
rect 6560 204 6564 236
rect 6596 204 6600 236
rect 6560 156 6600 204
rect 6560 124 6564 156
rect 6596 124 6600 156
rect 6560 76 6600 124
rect 6560 44 6564 76
rect 6596 44 6600 76
rect 6560 -4 6600 44
rect 6560 -36 6564 -4
rect 6596 -36 6600 -4
rect 6560 -84 6600 -36
rect 6560 -116 6564 -84
rect 6596 -116 6600 -84
rect 6560 -120 6600 -116
rect 6640 1036 6680 1040
rect 6640 1004 6644 1036
rect 6676 1004 6680 1036
rect 6640 956 6680 1004
rect 6640 924 6644 956
rect 6676 924 6680 956
rect 6640 876 6680 924
rect 6640 844 6644 876
rect 6676 844 6680 876
rect 6640 796 6680 844
rect 6640 764 6644 796
rect 6676 764 6680 796
rect 6640 716 6680 764
rect 6640 684 6644 716
rect 6676 684 6680 716
rect 6640 636 6680 684
rect 6640 604 6644 636
rect 6676 604 6680 636
rect 6640 556 6680 604
rect 6640 524 6644 556
rect 6676 524 6680 556
rect 6640 476 6680 524
rect 6640 444 6644 476
rect 6676 444 6680 476
rect 6640 396 6680 444
rect 6640 364 6644 396
rect 6676 364 6680 396
rect 6640 316 6680 364
rect 6640 284 6644 316
rect 6676 284 6680 316
rect 6640 236 6680 284
rect 6640 204 6644 236
rect 6676 204 6680 236
rect 6640 156 6680 204
rect 6640 124 6644 156
rect 6676 124 6680 156
rect 6640 76 6680 124
rect 6640 44 6644 76
rect 6676 44 6680 76
rect 6640 -4 6680 44
rect 6640 -36 6644 -4
rect 6676 -36 6680 -4
rect 6640 -84 6680 -36
rect 6640 -116 6644 -84
rect 6676 -116 6680 -84
rect 6640 -120 6680 -116
rect 6720 1036 6760 1040
rect 6720 1004 6724 1036
rect 6756 1004 6760 1036
rect 6720 956 6760 1004
rect 6720 924 6724 956
rect 6756 924 6760 956
rect 6720 876 6760 924
rect 6720 844 6724 876
rect 6756 844 6760 876
rect 6720 796 6760 844
rect 6720 764 6724 796
rect 6756 764 6760 796
rect 6720 716 6760 764
rect 6720 684 6724 716
rect 6756 684 6760 716
rect 6720 636 6760 684
rect 6720 604 6724 636
rect 6756 604 6760 636
rect 6720 556 6760 604
rect 6720 524 6724 556
rect 6756 524 6760 556
rect 6720 476 6760 524
rect 6720 444 6724 476
rect 6756 444 6760 476
rect 6720 396 6760 444
rect 6720 364 6724 396
rect 6756 364 6760 396
rect 6720 316 6760 364
rect 6720 284 6724 316
rect 6756 284 6760 316
rect 6720 236 6760 284
rect 6720 204 6724 236
rect 6756 204 6760 236
rect 6720 156 6760 204
rect 6720 124 6724 156
rect 6756 124 6760 156
rect 6720 76 6760 124
rect 6720 44 6724 76
rect 6756 44 6760 76
rect 6720 -4 6760 44
rect 6720 -36 6724 -4
rect 6756 -36 6760 -4
rect 6720 -84 6760 -36
rect 6720 -116 6724 -84
rect 6756 -116 6760 -84
rect 6720 -120 6760 -116
rect 6800 1036 6840 1040
rect 6800 1004 6804 1036
rect 6836 1004 6840 1036
rect 6800 956 6840 1004
rect 6800 924 6804 956
rect 6836 924 6840 956
rect 6800 876 6840 924
rect 6800 844 6804 876
rect 6836 844 6840 876
rect 6800 796 6840 844
rect 6800 764 6804 796
rect 6836 764 6840 796
rect 6800 716 6840 764
rect 6800 684 6804 716
rect 6836 684 6840 716
rect 6800 636 6840 684
rect 6800 604 6804 636
rect 6836 604 6840 636
rect 6800 556 6840 604
rect 6800 524 6804 556
rect 6836 524 6840 556
rect 6800 476 6840 524
rect 6800 444 6804 476
rect 6836 444 6840 476
rect 6800 396 6840 444
rect 6800 364 6804 396
rect 6836 364 6840 396
rect 6800 316 6840 364
rect 6800 284 6804 316
rect 6836 284 6840 316
rect 6800 236 6840 284
rect 6800 204 6804 236
rect 6836 204 6840 236
rect 6800 156 6840 204
rect 6800 124 6804 156
rect 6836 124 6840 156
rect 6800 76 6840 124
rect 6800 44 6804 76
rect 6836 44 6840 76
rect 6800 -4 6840 44
rect 6800 -36 6804 -4
rect 6836 -36 6840 -4
rect 6800 -84 6840 -36
rect 6800 -116 6804 -84
rect 6836 -116 6840 -84
rect 6800 -120 6840 -116
rect 6880 1036 6920 1040
rect 6880 1004 6884 1036
rect 6916 1004 6920 1036
rect 6880 956 6920 1004
rect 6880 924 6884 956
rect 6916 924 6920 956
rect 6880 876 6920 924
rect 6880 844 6884 876
rect 6916 844 6920 876
rect 6880 796 6920 844
rect 6880 764 6884 796
rect 6916 764 6920 796
rect 6880 716 6920 764
rect 6880 684 6884 716
rect 6916 684 6920 716
rect 6880 636 6920 684
rect 6880 604 6884 636
rect 6916 604 6920 636
rect 6880 556 6920 604
rect 6880 524 6884 556
rect 6916 524 6920 556
rect 6880 476 6920 524
rect 6880 444 6884 476
rect 6916 444 6920 476
rect 6880 396 6920 444
rect 6880 364 6884 396
rect 6916 364 6920 396
rect 6880 316 6920 364
rect 6880 284 6884 316
rect 6916 284 6920 316
rect 6880 236 6920 284
rect 6880 204 6884 236
rect 6916 204 6920 236
rect 6880 156 6920 204
rect 6880 124 6884 156
rect 6916 124 6920 156
rect 6880 76 6920 124
rect 6880 44 6884 76
rect 6916 44 6920 76
rect 6880 -4 6920 44
rect 6880 -36 6884 -4
rect 6916 -36 6920 -4
rect 6880 -84 6920 -36
rect 6880 -116 6884 -84
rect 6916 -116 6920 -84
rect 6880 -120 6920 -116
rect 6960 1036 7000 1040
rect 6960 1004 6964 1036
rect 6996 1004 7000 1036
rect 6960 956 7000 1004
rect 6960 924 6964 956
rect 6996 924 7000 956
rect 6960 876 7000 924
rect 6960 844 6964 876
rect 6996 844 7000 876
rect 6960 796 7000 844
rect 6960 764 6964 796
rect 6996 764 7000 796
rect 6960 716 7000 764
rect 6960 684 6964 716
rect 6996 684 7000 716
rect 6960 636 7000 684
rect 6960 604 6964 636
rect 6996 604 7000 636
rect 6960 556 7000 604
rect 6960 524 6964 556
rect 6996 524 7000 556
rect 6960 476 7000 524
rect 6960 444 6964 476
rect 6996 444 7000 476
rect 6960 396 7000 444
rect 6960 364 6964 396
rect 6996 364 7000 396
rect 6960 316 7000 364
rect 6960 284 6964 316
rect 6996 284 7000 316
rect 6960 236 7000 284
rect 6960 204 6964 236
rect 6996 204 7000 236
rect 6960 156 7000 204
rect 6960 124 6964 156
rect 6996 124 7000 156
rect 6960 76 7000 124
rect 6960 44 6964 76
rect 6996 44 7000 76
rect 6960 -4 7000 44
rect 6960 -36 6964 -4
rect 6996 -36 7000 -4
rect 6960 -84 7000 -36
rect 6960 -116 6964 -84
rect 6996 -116 7000 -84
rect 6960 -120 7000 -116
rect 7040 1036 7080 1040
rect 7040 1004 7044 1036
rect 7076 1004 7080 1036
rect 7040 956 7080 1004
rect 7040 924 7044 956
rect 7076 924 7080 956
rect 7040 876 7080 924
rect 7040 844 7044 876
rect 7076 844 7080 876
rect 7040 796 7080 844
rect 7040 764 7044 796
rect 7076 764 7080 796
rect 7040 716 7080 764
rect 7040 684 7044 716
rect 7076 684 7080 716
rect 7040 636 7080 684
rect 7040 604 7044 636
rect 7076 604 7080 636
rect 7040 556 7080 604
rect 7040 524 7044 556
rect 7076 524 7080 556
rect 7040 476 7080 524
rect 7040 444 7044 476
rect 7076 444 7080 476
rect 7040 396 7080 444
rect 7040 364 7044 396
rect 7076 364 7080 396
rect 7040 316 7080 364
rect 7040 284 7044 316
rect 7076 284 7080 316
rect 7040 236 7080 284
rect 7040 204 7044 236
rect 7076 204 7080 236
rect 7040 156 7080 204
rect 7040 124 7044 156
rect 7076 124 7080 156
rect 7040 76 7080 124
rect 7040 44 7044 76
rect 7076 44 7080 76
rect 7040 -4 7080 44
rect 7040 -36 7044 -4
rect 7076 -36 7080 -4
rect 7040 -84 7080 -36
rect 7040 -116 7044 -84
rect 7076 -116 7080 -84
rect 7040 -120 7080 -116
rect 7120 1036 7160 1040
rect 7120 1004 7124 1036
rect 7156 1004 7160 1036
rect 7120 956 7160 1004
rect 7120 924 7124 956
rect 7156 924 7160 956
rect 7120 876 7160 924
rect 7120 844 7124 876
rect 7156 844 7160 876
rect 7120 796 7160 844
rect 7120 764 7124 796
rect 7156 764 7160 796
rect 7120 716 7160 764
rect 7120 684 7124 716
rect 7156 684 7160 716
rect 7120 636 7160 684
rect 7120 604 7124 636
rect 7156 604 7160 636
rect 7120 556 7160 604
rect 7120 524 7124 556
rect 7156 524 7160 556
rect 7120 476 7160 524
rect 7120 444 7124 476
rect 7156 444 7160 476
rect 7120 396 7160 444
rect 7120 364 7124 396
rect 7156 364 7160 396
rect 7120 316 7160 364
rect 7120 284 7124 316
rect 7156 284 7160 316
rect 7120 236 7160 284
rect 7120 204 7124 236
rect 7156 204 7160 236
rect 7120 156 7160 204
rect 7120 124 7124 156
rect 7156 124 7160 156
rect 7120 76 7160 124
rect 7120 44 7124 76
rect 7156 44 7160 76
rect 7120 -4 7160 44
rect 7120 -36 7124 -4
rect 7156 -36 7160 -4
rect 7120 -84 7160 -36
rect 7120 -116 7124 -84
rect 7156 -116 7160 -84
rect 7120 -120 7160 -116
rect 7200 1036 7240 1040
rect 7200 1004 7204 1036
rect 7236 1004 7240 1036
rect 7200 956 7240 1004
rect 7200 924 7204 956
rect 7236 924 7240 956
rect 7200 876 7240 924
rect 7200 844 7204 876
rect 7236 844 7240 876
rect 7200 796 7240 844
rect 7200 764 7204 796
rect 7236 764 7240 796
rect 7200 716 7240 764
rect 7200 684 7204 716
rect 7236 684 7240 716
rect 7200 636 7240 684
rect 7200 604 7204 636
rect 7236 604 7240 636
rect 7200 556 7240 604
rect 7200 524 7204 556
rect 7236 524 7240 556
rect 7200 476 7240 524
rect 7200 444 7204 476
rect 7236 444 7240 476
rect 7200 396 7240 444
rect 7200 364 7204 396
rect 7236 364 7240 396
rect 7200 316 7240 364
rect 7200 284 7204 316
rect 7236 284 7240 316
rect 7200 236 7240 284
rect 7200 204 7204 236
rect 7236 204 7240 236
rect 7200 156 7240 204
rect 7200 124 7204 156
rect 7236 124 7240 156
rect 7200 76 7240 124
rect 7200 44 7204 76
rect 7236 44 7240 76
rect 7200 -4 7240 44
rect 7200 -36 7204 -4
rect 7236 -36 7240 -4
rect 7200 -84 7240 -36
rect 7200 -116 7204 -84
rect 7236 -116 7240 -84
rect 7200 -120 7240 -116
rect 7280 1036 7320 1040
rect 7280 1004 7284 1036
rect 7316 1004 7320 1036
rect 7280 956 7320 1004
rect 7280 924 7284 956
rect 7316 924 7320 956
rect 7280 876 7320 924
rect 7280 844 7284 876
rect 7316 844 7320 876
rect 7280 796 7320 844
rect 7280 764 7284 796
rect 7316 764 7320 796
rect 7280 716 7320 764
rect 7280 684 7284 716
rect 7316 684 7320 716
rect 7280 636 7320 684
rect 7280 604 7284 636
rect 7316 604 7320 636
rect 7280 556 7320 604
rect 7280 524 7284 556
rect 7316 524 7320 556
rect 7280 476 7320 524
rect 7280 444 7284 476
rect 7316 444 7320 476
rect 7280 396 7320 444
rect 7280 364 7284 396
rect 7316 364 7320 396
rect 7280 316 7320 364
rect 7280 284 7284 316
rect 7316 284 7320 316
rect 7280 236 7320 284
rect 7280 204 7284 236
rect 7316 204 7320 236
rect 7280 156 7320 204
rect 7280 124 7284 156
rect 7316 124 7320 156
rect 7280 76 7320 124
rect 7280 44 7284 76
rect 7316 44 7320 76
rect 7280 -4 7320 44
rect 7280 -36 7284 -4
rect 7316 -36 7320 -4
rect 7280 -84 7320 -36
rect 7280 -116 7284 -84
rect 7316 -116 7320 -84
rect 7280 -120 7320 -116
rect 7360 1036 7400 1040
rect 7360 1004 7364 1036
rect 7396 1004 7400 1036
rect 7360 956 7400 1004
rect 7360 924 7364 956
rect 7396 924 7400 956
rect 7360 876 7400 924
rect 7360 844 7364 876
rect 7396 844 7400 876
rect 7360 796 7400 844
rect 7360 764 7364 796
rect 7396 764 7400 796
rect 7360 716 7400 764
rect 7360 684 7364 716
rect 7396 684 7400 716
rect 7360 636 7400 684
rect 7360 604 7364 636
rect 7396 604 7400 636
rect 7360 556 7400 604
rect 7360 524 7364 556
rect 7396 524 7400 556
rect 7360 476 7400 524
rect 7360 444 7364 476
rect 7396 444 7400 476
rect 7360 396 7400 444
rect 7360 364 7364 396
rect 7396 364 7400 396
rect 7360 316 7400 364
rect 7360 284 7364 316
rect 7396 284 7400 316
rect 7360 236 7400 284
rect 7360 204 7364 236
rect 7396 204 7400 236
rect 7360 156 7400 204
rect 7360 124 7364 156
rect 7396 124 7400 156
rect 7360 76 7400 124
rect 7360 44 7364 76
rect 7396 44 7400 76
rect 7360 -4 7400 44
rect 7360 -36 7364 -4
rect 7396 -36 7400 -4
rect 7360 -84 7400 -36
rect 7360 -116 7364 -84
rect 7396 -116 7400 -84
rect 7360 -120 7400 -116
rect 7440 1036 7480 1040
rect 7440 1004 7444 1036
rect 7476 1004 7480 1036
rect 7440 956 7480 1004
rect 7440 924 7444 956
rect 7476 924 7480 956
rect 7440 876 7480 924
rect 7440 844 7444 876
rect 7476 844 7480 876
rect 7440 796 7480 844
rect 7440 764 7444 796
rect 7476 764 7480 796
rect 7440 716 7480 764
rect 7440 684 7444 716
rect 7476 684 7480 716
rect 7440 636 7480 684
rect 7440 604 7444 636
rect 7476 604 7480 636
rect 7440 556 7480 604
rect 7440 524 7444 556
rect 7476 524 7480 556
rect 7440 476 7480 524
rect 7440 444 7444 476
rect 7476 444 7480 476
rect 7440 396 7480 444
rect 7440 364 7444 396
rect 7476 364 7480 396
rect 7440 316 7480 364
rect 7440 284 7444 316
rect 7476 284 7480 316
rect 7440 236 7480 284
rect 7440 204 7444 236
rect 7476 204 7480 236
rect 7440 156 7480 204
rect 7440 124 7444 156
rect 7476 124 7480 156
rect 7440 76 7480 124
rect 7440 44 7444 76
rect 7476 44 7480 76
rect 7440 -4 7480 44
rect 7440 -36 7444 -4
rect 7476 -36 7480 -4
rect 7440 -84 7480 -36
rect 7440 -116 7444 -84
rect 7476 -116 7480 -84
rect 7440 -120 7480 -116
rect 7520 1036 7560 1040
rect 7520 1004 7524 1036
rect 7556 1004 7560 1036
rect 7520 956 7560 1004
rect 7520 924 7524 956
rect 7556 924 7560 956
rect 7520 876 7560 924
rect 7520 844 7524 876
rect 7556 844 7560 876
rect 7520 796 7560 844
rect 7520 764 7524 796
rect 7556 764 7560 796
rect 7520 716 7560 764
rect 7520 684 7524 716
rect 7556 684 7560 716
rect 7520 636 7560 684
rect 7520 604 7524 636
rect 7556 604 7560 636
rect 7520 556 7560 604
rect 7520 524 7524 556
rect 7556 524 7560 556
rect 7520 476 7560 524
rect 7520 444 7524 476
rect 7556 444 7560 476
rect 7520 396 7560 444
rect 7520 364 7524 396
rect 7556 364 7560 396
rect 7520 316 7560 364
rect 7520 284 7524 316
rect 7556 284 7560 316
rect 7520 236 7560 284
rect 7520 204 7524 236
rect 7556 204 7560 236
rect 7520 156 7560 204
rect 7520 124 7524 156
rect 7556 124 7560 156
rect 7520 76 7560 124
rect 7520 44 7524 76
rect 7556 44 7560 76
rect 7520 -4 7560 44
rect 7520 -36 7524 -4
rect 7556 -36 7560 -4
rect 7520 -84 7560 -36
rect 7520 -116 7524 -84
rect 7556 -116 7560 -84
rect 7520 -120 7560 -116
rect 7600 1036 7640 1040
rect 7600 1004 7604 1036
rect 7636 1004 7640 1036
rect 7600 956 7640 1004
rect 7600 924 7604 956
rect 7636 924 7640 956
rect 7600 876 7640 924
rect 7600 844 7604 876
rect 7636 844 7640 876
rect 7600 796 7640 844
rect 7600 764 7604 796
rect 7636 764 7640 796
rect 7600 716 7640 764
rect 7600 684 7604 716
rect 7636 684 7640 716
rect 7600 636 7640 684
rect 7600 604 7604 636
rect 7636 604 7640 636
rect 7600 556 7640 604
rect 7600 524 7604 556
rect 7636 524 7640 556
rect 7600 476 7640 524
rect 7600 444 7604 476
rect 7636 444 7640 476
rect 7600 396 7640 444
rect 7600 364 7604 396
rect 7636 364 7640 396
rect 7600 316 7640 364
rect 7600 284 7604 316
rect 7636 284 7640 316
rect 7600 236 7640 284
rect 7600 204 7604 236
rect 7636 204 7640 236
rect 7600 156 7640 204
rect 7600 124 7604 156
rect 7636 124 7640 156
rect 7600 76 7640 124
rect 7600 44 7604 76
rect 7636 44 7640 76
rect 7600 -4 7640 44
rect 7600 -36 7604 -4
rect 7636 -36 7640 -4
rect 7600 -84 7640 -36
rect 7600 -116 7604 -84
rect 7636 -116 7640 -84
rect 7600 -120 7640 -116
rect 7680 1036 7720 1040
rect 7680 1004 7684 1036
rect 7716 1004 7720 1036
rect 7680 956 7720 1004
rect 7680 924 7684 956
rect 7716 924 7720 956
rect 7680 876 7720 924
rect 7680 844 7684 876
rect 7716 844 7720 876
rect 7680 796 7720 844
rect 7680 764 7684 796
rect 7716 764 7720 796
rect 7680 716 7720 764
rect 7680 684 7684 716
rect 7716 684 7720 716
rect 7680 636 7720 684
rect 7680 604 7684 636
rect 7716 604 7720 636
rect 7680 556 7720 604
rect 7680 524 7684 556
rect 7716 524 7720 556
rect 7680 476 7720 524
rect 7680 444 7684 476
rect 7716 444 7720 476
rect 7680 396 7720 444
rect 7680 364 7684 396
rect 7716 364 7720 396
rect 7680 316 7720 364
rect 7680 284 7684 316
rect 7716 284 7720 316
rect 7680 236 7720 284
rect 7680 204 7684 236
rect 7716 204 7720 236
rect 7680 156 7720 204
rect 7680 124 7684 156
rect 7716 124 7720 156
rect 7680 76 7720 124
rect 7680 44 7684 76
rect 7716 44 7720 76
rect 7680 -4 7720 44
rect 7680 -36 7684 -4
rect 7716 -36 7720 -4
rect 7680 -84 7720 -36
rect 7680 -116 7684 -84
rect 7716 -116 7720 -84
rect 7680 -120 7720 -116
rect 7760 1036 7800 1040
rect 7760 1004 7764 1036
rect 7796 1004 7800 1036
rect 7760 956 7800 1004
rect 7760 924 7764 956
rect 7796 924 7800 956
rect 7760 876 7800 924
rect 7760 844 7764 876
rect 7796 844 7800 876
rect 7760 796 7800 844
rect 7760 764 7764 796
rect 7796 764 7800 796
rect 7760 716 7800 764
rect 7760 684 7764 716
rect 7796 684 7800 716
rect 7760 636 7800 684
rect 7760 604 7764 636
rect 7796 604 7800 636
rect 7760 556 7800 604
rect 7760 524 7764 556
rect 7796 524 7800 556
rect 7760 476 7800 524
rect 7760 444 7764 476
rect 7796 444 7800 476
rect 7760 396 7800 444
rect 7760 364 7764 396
rect 7796 364 7800 396
rect 7760 316 7800 364
rect 7760 284 7764 316
rect 7796 284 7800 316
rect 7760 236 7800 284
rect 7760 204 7764 236
rect 7796 204 7800 236
rect 7760 156 7800 204
rect 7760 124 7764 156
rect 7796 124 7800 156
rect 7760 76 7800 124
rect 7760 44 7764 76
rect 7796 44 7800 76
rect 7760 -4 7800 44
rect 7760 -36 7764 -4
rect 7796 -36 7800 -4
rect 7760 -84 7800 -36
rect 7760 -116 7764 -84
rect 7796 -116 7800 -84
rect 7760 -120 7800 -116
rect 7840 1036 7880 1040
rect 7840 1004 7844 1036
rect 7876 1004 7880 1036
rect 7840 956 7880 1004
rect 7840 924 7844 956
rect 7876 924 7880 956
rect 7840 876 7880 924
rect 7840 844 7844 876
rect 7876 844 7880 876
rect 7840 796 7880 844
rect 7840 764 7844 796
rect 7876 764 7880 796
rect 7840 716 7880 764
rect 7840 684 7844 716
rect 7876 684 7880 716
rect 7840 636 7880 684
rect 7840 604 7844 636
rect 7876 604 7880 636
rect 7840 556 7880 604
rect 7840 524 7844 556
rect 7876 524 7880 556
rect 7840 476 7880 524
rect 7840 444 7844 476
rect 7876 444 7880 476
rect 7840 396 7880 444
rect 7840 364 7844 396
rect 7876 364 7880 396
rect 7840 316 7880 364
rect 7840 284 7844 316
rect 7876 284 7880 316
rect 7840 236 7880 284
rect 7840 204 7844 236
rect 7876 204 7880 236
rect 7840 156 7880 204
rect 7840 124 7844 156
rect 7876 124 7880 156
rect 7840 76 7880 124
rect 7840 44 7844 76
rect 7876 44 7880 76
rect 7840 -4 7880 44
rect 7840 -36 7844 -4
rect 7876 -36 7880 -4
rect 7840 -84 7880 -36
rect 7840 -116 7844 -84
rect 7876 -116 7880 -84
rect 7840 -120 7880 -116
rect 7920 1036 7960 1040
rect 7920 1004 7924 1036
rect 7956 1004 7960 1036
rect 7920 956 7960 1004
rect 7920 924 7924 956
rect 7956 924 7960 956
rect 7920 876 7960 924
rect 7920 844 7924 876
rect 7956 844 7960 876
rect 7920 796 7960 844
rect 7920 764 7924 796
rect 7956 764 7960 796
rect 7920 716 7960 764
rect 7920 684 7924 716
rect 7956 684 7960 716
rect 7920 636 7960 684
rect 7920 604 7924 636
rect 7956 604 7960 636
rect 7920 556 7960 604
rect 7920 524 7924 556
rect 7956 524 7960 556
rect 7920 476 7960 524
rect 7920 444 7924 476
rect 7956 444 7960 476
rect 7920 396 7960 444
rect 7920 364 7924 396
rect 7956 364 7960 396
rect 7920 316 7960 364
rect 7920 284 7924 316
rect 7956 284 7960 316
rect 7920 236 7960 284
rect 7920 204 7924 236
rect 7956 204 7960 236
rect 7920 156 7960 204
rect 7920 124 7924 156
rect 7956 124 7960 156
rect 7920 76 7960 124
rect 7920 44 7924 76
rect 7956 44 7960 76
rect 7920 -4 7960 44
rect 7920 -36 7924 -4
rect 7956 -36 7960 -4
rect 7920 -84 7960 -36
rect 7920 -116 7924 -84
rect 7956 -116 7960 -84
rect 7920 -120 7960 -116
rect 8000 1036 8040 1040
rect 8000 1004 8004 1036
rect 8036 1004 8040 1036
rect 8000 956 8040 1004
rect 8000 924 8004 956
rect 8036 924 8040 956
rect 8000 876 8040 924
rect 8000 844 8004 876
rect 8036 844 8040 876
rect 8000 796 8040 844
rect 8000 764 8004 796
rect 8036 764 8040 796
rect 8000 716 8040 764
rect 8000 684 8004 716
rect 8036 684 8040 716
rect 8000 636 8040 684
rect 8000 604 8004 636
rect 8036 604 8040 636
rect 8000 556 8040 604
rect 8000 524 8004 556
rect 8036 524 8040 556
rect 8000 476 8040 524
rect 8000 444 8004 476
rect 8036 444 8040 476
rect 8000 396 8040 444
rect 8000 364 8004 396
rect 8036 364 8040 396
rect 8000 316 8040 364
rect 8000 284 8004 316
rect 8036 284 8040 316
rect 8000 236 8040 284
rect 8000 204 8004 236
rect 8036 204 8040 236
rect 8000 156 8040 204
rect 8000 124 8004 156
rect 8036 124 8040 156
rect 8000 76 8040 124
rect 8000 44 8004 76
rect 8036 44 8040 76
rect 8000 -4 8040 44
rect 8000 -36 8004 -4
rect 8036 -36 8040 -4
rect 8000 -84 8040 -36
rect 8000 -116 8004 -84
rect 8036 -116 8040 -84
rect 8000 -120 8040 -116
rect 8080 1036 8120 1040
rect 8080 1004 8084 1036
rect 8116 1004 8120 1036
rect 8080 956 8120 1004
rect 8080 924 8084 956
rect 8116 924 8120 956
rect 8080 876 8120 924
rect 8080 844 8084 876
rect 8116 844 8120 876
rect 8080 796 8120 844
rect 8080 764 8084 796
rect 8116 764 8120 796
rect 8080 716 8120 764
rect 8080 684 8084 716
rect 8116 684 8120 716
rect 8080 636 8120 684
rect 8080 604 8084 636
rect 8116 604 8120 636
rect 8080 556 8120 604
rect 8080 524 8084 556
rect 8116 524 8120 556
rect 8080 476 8120 524
rect 8080 444 8084 476
rect 8116 444 8120 476
rect 8080 396 8120 444
rect 8080 364 8084 396
rect 8116 364 8120 396
rect 8080 316 8120 364
rect 8080 284 8084 316
rect 8116 284 8120 316
rect 8080 236 8120 284
rect 8080 204 8084 236
rect 8116 204 8120 236
rect 8080 156 8120 204
rect 8080 124 8084 156
rect 8116 124 8120 156
rect 8080 76 8120 124
rect 8080 44 8084 76
rect 8116 44 8120 76
rect 8080 -4 8120 44
rect 8080 -36 8084 -4
rect 8116 -36 8120 -4
rect 8080 -84 8120 -36
rect 8080 -116 8084 -84
rect 8116 -116 8120 -84
rect 8080 -120 8120 -116
rect 8160 1036 8200 1040
rect 8160 1004 8164 1036
rect 8196 1004 8200 1036
rect 8160 956 8200 1004
rect 8160 924 8164 956
rect 8196 924 8200 956
rect 8160 876 8200 924
rect 8160 844 8164 876
rect 8196 844 8200 876
rect 8160 796 8200 844
rect 8160 764 8164 796
rect 8196 764 8200 796
rect 8160 716 8200 764
rect 8160 684 8164 716
rect 8196 684 8200 716
rect 8160 636 8200 684
rect 8160 604 8164 636
rect 8196 604 8200 636
rect 8160 556 8200 604
rect 8160 524 8164 556
rect 8196 524 8200 556
rect 8160 476 8200 524
rect 8160 444 8164 476
rect 8196 444 8200 476
rect 8160 396 8200 444
rect 8160 364 8164 396
rect 8196 364 8200 396
rect 8160 316 8200 364
rect 8160 284 8164 316
rect 8196 284 8200 316
rect 8160 236 8200 284
rect 8160 204 8164 236
rect 8196 204 8200 236
rect 8160 156 8200 204
rect 8160 124 8164 156
rect 8196 124 8200 156
rect 8160 76 8200 124
rect 8160 44 8164 76
rect 8196 44 8200 76
rect 8160 -4 8200 44
rect 8160 -36 8164 -4
rect 8196 -36 8200 -4
rect 8160 -84 8200 -36
rect 8160 -116 8164 -84
rect 8196 -116 8200 -84
rect 8160 -120 8200 -116
rect 8240 1036 8280 1040
rect 8240 1004 8244 1036
rect 8276 1004 8280 1036
rect 8240 956 8280 1004
rect 8240 924 8244 956
rect 8276 924 8280 956
rect 8240 876 8280 924
rect 8240 844 8244 876
rect 8276 844 8280 876
rect 8240 796 8280 844
rect 8240 764 8244 796
rect 8276 764 8280 796
rect 8240 716 8280 764
rect 8240 684 8244 716
rect 8276 684 8280 716
rect 8240 636 8280 684
rect 8240 604 8244 636
rect 8276 604 8280 636
rect 8240 556 8280 604
rect 8240 524 8244 556
rect 8276 524 8280 556
rect 8240 476 8280 524
rect 8240 444 8244 476
rect 8276 444 8280 476
rect 8240 396 8280 444
rect 8240 364 8244 396
rect 8276 364 8280 396
rect 8240 316 8280 364
rect 8240 284 8244 316
rect 8276 284 8280 316
rect 8240 236 8280 284
rect 8240 204 8244 236
rect 8276 204 8280 236
rect 8240 156 8280 204
rect 8240 124 8244 156
rect 8276 124 8280 156
rect 8240 76 8280 124
rect 8240 44 8244 76
rect 8276 44 8280 76
rect 8240 -4 8280 44
rect 8240 -36 8244 -4
rect 8276 -36 8280 -4
rect 8240 -84 8280 -36
rect 8240 -116 8244 -84
rect 8276 -116 8280 -84
rect 8240 -120 8280 -116
rect 8320 1036 8360 1040
rect 8320 1004 8324 1036
rect 8356 1004 8360 1036
rect 8320 956 8360 1004
rect 8320 924 8324 956
rect 8356 924 8360 956
rect 8320 876 8360 924
rect 8320 844 8324 876
rect 8356 844 8360 876
rect 8320 796 8360 844
rect 8320 764 8324 796
rect 8356 764 8360 796
rect 8320 716 8360 764
rect 8320 684 8324 716
rect 8356 684 8360 716
rect 8320 636 8360 684
rect 8320 604 8324 636
rect 8356 604 8360 636
rect 8320 556 8360 604
rect 8320 524 8324 556
rect 8356 524 8360 556
rect 8320 476 8360 524
rect 8320 444 8324 476
rect 8356 444 8360 476
rect 8320 396 8360 444
rect 8320 364 8324 396
rect 8356 364 8360 396
rect 8320 316 8360 364
rect 8320 284 8324 316
rect 8356 284 8360 316
rect 8320 236 8360 284
rect 8320 204 8324 236
rect 8356 204 8360 236
rect 8320 156 8360 204
rect 8320 124 8324 156
rect 8356 124 8360 156
rect 8320 76 8360 124
rect 8320 44 8324 76
rect 8356 44 8360 76
rect 8320 -4 8360 44
rect 8320 -36 8324 -4
rect 8356 -36 8360 -4
rect 8320 -84 8360 -36
rect 8320 -116 8324 -84
rect 8356 -116 8360 -84
rect 8320 -120 8360 -116
rect 8400 1036 8440 1040
rect 8400 1004 8404 1036
rect 8436 1004 8440 1036
rect 8400 956 8440 1004
rect 8400 924 8404 956
rect 8436 924 8440 956
rect 8400 876 8440 924
rect 8400 844 8404 876
rect 8436 844 8440 876
rect 8400 796 8440 844
rect 8400 764 8404 796
rect 8436 764 8440 796
rect 8400 716 8440 764
rect 8400 684 8404 716
rect 8436 684 8440 716
rect 8400 636 8440 684
rect 8400 604 8404 636
rect 8436 604 8440 636
rect 8400 556 8440 604
rect 8400 524 8404 556
rect 8436 524 8440 556
rect 8400 476 8440 524
rect 8400 444 8404 476
rect 8436 444 8440 476
rect 8400 396 8440 444
rect 8400 364 8404 396
rect 8436 364 8440 396
rect 8400 316 8440 364
rect 8400 284 8404 316
rect 8436 284 8440 316
rect 8400 236 8440 284
rect 8400 204 8404 236
rect 8436 204 8440 236
rect 8400 156 8440 204
rect 8400 124 8404 156
rect 8436 124 8440 156
rect 8400 76 8440 124
rect 8400 44 8404 76
rect 8436 44 8440 76
rect 8400 -4 8440 44
rect 8400 -36 8404 -4
rect 8436 -36 8440 -4
rect 8400 -84 8440 -36
rect 8400 -116 8404 -84
rect 8436 -116 8440 -84
rect 8400 -120 8440 -116
rect 8480 1036 8520 1040
rect 8480 1004 8484 1036
rect 8516 1004 8520 1036
rect 8480 956 8520 1004
rect 8480 924 8484 956
rect 8516 924 8520 956
rect 8480 876 8520 924
rect 8480 844 8484 876
rect 8516 844 8520 876
rect 8480 796 8520 844
rect 8480 764 8484 796
rect 8516 764 8520 796
rect 8480 716 8520 764
rect 8480 684 8484 716
rect 8516 684 8520 716
rect 8480 636 8520 684
rect 8480 604 8484 636
rect 8516 604 8520 636
rect 8480 556 8520 604
rect 8480 524 8484 556
rect 8516 524 8520 556
rect 8480 476 8520 524
rect 8480 444 8484 476
rect 8516 444 8520 476
rect 8480 396 8520 444
rect 8480 364 8484 396
rect 8516 364 8520 396
rect 8480 316 8520 364
rect 8480 284 8484 316
rect 8516 284 8520 316
rect 8480 236 8520 284
rect 8480 204 8484 236
rect 8516 204 8520 236
rect 8480 156 8520 204
rect 8480 124 8484 156
rect 8516 124 8520 156
rect 8480 76 8520 124
rect 8480 44 8484 76
rect 8516 44 8520 76
rect 8480 -4 8520 44
rect 8480 -36 8484 -4
rect 8516 -36 8520 -4
rect 8480 -84 8520 -36
rect 8480 -116 8484 -84
rect 8516 -116 8520 -84
rect 8480 -120 8520 -116
rect 8560 1036 8600 1040
rect 8560 1004 8564 1036
rect 8596 1004 8600 1036
rect 8560 956 8600 1004
rect 8560 924 8564 956
rect 8596 924 8600 956
rect 8560 876 8600 924
rect 8560 844 8564 876
rect 8596 844 8600 876
rect 8560 796 8600 844
rect 8560 764 8564 796
rect 8596 764 8600 796
rect 8560 716 8600 764
rect 8560 684 8564 716
rect 8596 684 8600 716
rect 8560 636 8600 684
rect 8560 604 8564 636
rect 8596 604 8600 636
rect 8560 556 8600 604
rect 8560 524 8564 556
rect 8596 524 8600 556
rect 8560 476 8600 524
rect 8560 444 8564 476
rect 8596 444 8600 476
rect 8560 396 8600 444
rect 8560 364 8564 396
rect 8596 364 8600 396
rect 8560 316 8600 364
rect 8560 284 8564 316
rect 8596 284 8600 316
rect 8560 236 8600 284
rect 8560 204 8564 236
rect 8596 204 8600 236
rect 8560 156 8600 204
rect 8560 124 8564 156
rect 8596 124 8600 156
rect 8560 76 8600 124
rect 8560 44 8564 76
rect 8596 44 8600 76
rect 8560 -4 8600 44
rect 8560 -36 8564 -4
rect 8596 -36 8600 -4
rect 8560 -84 8600 -36
rect 8560 -116 8564 -84
rect 8596 -116 8600 -84
rect 8560 -120 8600 -116
rect 8640 1036 8680 1040
rect 8640 1004 8644 1036
rect 8676 1004 8680 1036
rect 8640 956 8680 1004
rect 8640 924 8644 956
rect 8676 924 8680 956
rect 8640 876 8680 924
rect 8640 844 8644 876
rect 8676 844 8680 876
rect 8640 796 8680 844
rect 8640 764 8644 796
rect 8676 764 8680 796
rect 8640 716 8680 764
rect 8640 684 8644 716
rect 8676 684 8680 716
rect 8640 636 8680 684
rect 8640 604 8644 636
rect 8676 604 8680 636
rect 8640 556 8680 604
rect 8640 524 8644 556
rect 8676 524 8680 556
rect 8640 476 8680 524
rect 8640 444 8644 476
rect 8676 444 8680 476
rect 8640 396 8680 444
rect 8640 364 8644 396
rect 8676 364 8680 396
rect 8640 316 8680 364
rect 8640 284 8644 316
rect 8676 284 8680 316
rect 8640 236 8680 284
rect 8640 204 8644 236
rect 8676 204 8680 236
rect 8640 156 8680 204
rect 8640 124 8644 156
rect 8676 124 8680 156
rect 8640 76 8680 124
rect 8640 44 8644 76
rect 8676 44 8680 76
rect 8640 -4 8680 44
rect 8640 -36 8644 -4
rect 8676 -36 8680 -4
rect 8640 -84 8680 -36
rect 8640 -116 8644 -84
rect 8676 -116 8680 -84
rect 8640 -120 8680 -116
rect 8720 1036 8760 1040
rect 8720 1004 8724 1036
rect 8756 1004 8760 1036
rect 8720 956 8760 1004
rect 8720 924 8724 956
rect 8756 924 8760 956
rect 8720 876 8760 924
rect 8720 844 8724 876
rect 8756 844 8760 876
rect 8720 796 8760 844
rect 8720 764 8724 796
rect 8756 764 8760 796
rect 8720 716 8760 764
rect 8720 684 8724 716
rect 8756 684 8760 716
rect 8720 636 8760 684
rect 8720 604 8724 636
rect 8756 604 8760 636
rect 8720 556 8760 604
rect 8720 524 8724 556
rect 8756 524 8760 556
rect 8720 476 8760 524
rect 8720 444 8724 476
rect 8756 444 8760 476
rect 8720 396 8760 444
rect 8720 364 8724 396
rect 8756 364 8760 396
rect 8720 316 8760 364
rect 8720 284 8724 316
rect 8756 284 8760 316
rect 8720 236 8760 284
rect 8720 204 8724 236
rect 8756 204 8760 236
rect 8720 156 8760 204
rect 8720 124 8724 156
rect 8756 124 8760 156
rect 8720 76 8760 124
rect 8720 44 8724 76
rect 8756 44 8760 76
rect 8720 -4 8760 44
rect 8720 -36 8724 -4
rect 8756 -36 8760 -4
rect 8720 -84 8760 -36
rect 8720 -116 8724 -84
rect 8756 -116 8760 -84
rect 8720 -120 8760 -116
rect 8800 1036 8840 1040
rect 8800 1004 8804 1036
rect 8836 1004 8840 1036
rect 8800 956 8840 1004
rect 8800 924 8804 956
rect 8836 924 8840 956
rect 8800 876 8840 924
rect 8800 844 8804 876
rect 8836 844 8840 876
rect 8800 796 8840 844
rect 8800 764 8804 796
rect 8836 764 8840 796
rect 8800 716 8840 764
rect 8800 684 8804 716
rect 8836 684 8840 716
rect 8800 636 8840 684
rect 8800 604 8804 636
rect 8836 604 8840 636
rect 8800 556 8840 604
rect 8800 524 8804 556
rect 8836 524 8840 556
rect 8800 476 8840 524
rect 8800 444 8804 476
rect 8836 444 8840 476
rect 8800 396 8840 444
rect 8800 364 8804 396
rect 8836 364 8840 396
rect 8800 316 8840 364
rect 8800 284 8804 316
rect 8836 284 8840 316
rect 8800 236 8840 284
rect 8800 204 8804 236
rect 8836 204 8840 236
rect 8800 156 8840 204
rect 8800 124 8804 156
rect 8836 124 8840 156
rect 8800 76 8840 124
rect 8800 44 8804 76
rect 8836 44 8840 76
rect 8800 -4 8840 44
rect 8800 -36 8804 -4
rect 8836 -36 8840 -4
rect 8800 -84 8840 -36
rect 8800 -116 8804 -84
rect 8836 -116 8840 -84
rect 8800 -120 8840 -116
rect 8880 1036 8920 1040
rect 8880 1004 8884 1036
rect 8916 1004 8920 1036
rect 8880 956 8920 1004
rect 8880 924 8884 956
rect 8916 924 8920 956
rect 8880 876 8920 924
rect 8880 844 8884 876
rect 8916 844 8920 876
rect 8880 796 8920 844
rect 8880 764 8884 796
rect 8916 764 8920 796
rect 8880 716 8920 764
rect 8880 684 8884 716
rect 8916 684 8920 716
rect 8880 636 8920 684
rect 8880 604 8884 636
rect 8916 604 8920 636
rect 8880 556 8920 604
rect 8880 524 8884 556
rect 8916 524 8920 556
rect 8880 476 8920 524
rect 8880 444 8884 476
rect 8916 444 8920 476
rect 8880 396 8920 444
rect 8880 364 8884 396
rect 8916 364 8920 396
rect 8880 316 8920 364
rect 8880 284 8884 316
rect 8916 284 8920 316
rect 8880 236 8920 284
rect 8880 204 8884 236
rect 8916 204 8920 236
rect 8880 156 8920 204
rect 8880 124 8884 156
rect 8916 124 8920 156
rect 8880 76 8920 124
rect 8880 44 8884 76
rect 8916 44 8920 76
rect 8880 -4 8920 44
rect 8880 -36 8884 -4
rect 8916 -36 8920 -4
rect 8880 -84 8920 -36
rect 8880 -116 8884 -84
rect 8916 -116 8920 -84
rect 8880 -120 8920 -116
rect 8960 1036 9000 1040
rect 8960 1004 8964 1036
rect 8996 1004 9000 1036
rect 8960 956 9000 1004
rect 8960 924 8964 956
rect 8996 924 9000 956
rect 8960 876 9000 924
rect 8960 844 8964 876
rect 8996 844 9000 876
rect 8960 796 9000 844
rect 8960 764 8964 796
rect 8996 764 9000 796
rect 8960 716 9000 764
rect 8960 684 8964 716
rect 8996 684 9000 716
rect 8960 636 9000 684
rect 8960 604 8964 636
rect 8996 604 9000 636
rect 8960 556 9000 604
rect 8960 524 8964 556
rect 8996 524 9000 556
rect 8960 476 9000 524
rect 8960 444 8964 476
rect 8996 444 9000 476
rect 8960 396 9000 444
rect 8960 364 8964 396
rect 8996 364 9000 396
rect 8960 316 9000 364
rect 8960 284 8964 316
rect 8996 284 9000 316
rect 8960 236 9000 284
rect 8960 204 8964 236
rect 8996 204 9000 236
rect 8960 156 9000 204
rect 8960 124 8964 156
rect 8996 124 9000 156
rect 8960 76 9000 124
rect 8960 44 8964 76
rect 8996 44 9000 76
rect 8960 -4 9000 44
rect 8960 -36 8964 -4
rect 8996 -36 9000 -4
rect 8960 -84 9000 -36
rect 8960 -116 8964 -84
rect 8996 -116 9000 -84
rect 8960 -120 9000 -116
rect 9040 1036 9080 1040
rect 9040 1004 9044 1036
rect 9076 1004 9080 1036
rect 9040 956 9080 1004
rect 9040 924 9044 956
rect 9076 924 9080 956
rect 9040 876 9080 924
rect 9040 844 9044 876
rect 9076 844 9080 876
rect 9040 796 9080 844
rect 9040 764 9044 796
rect 9076 764 9080 796
rect 9040 716 9080 764
rect 9040 684 9044 716
rect 9076 684 9080 716
rect 9040 636 9080 684
rect 9040 604 9044 636
rect 9076 604 9080 636
rect 9040 556 9080 604
rect 9040 524 9044 556
rect 9076 524 9080 556
rect 9040 476 9080 524
rect 9040 444 9044 476
rect 9076 444 9080 476
rect 9040 396 9080 444
rect 9040 364 9044 396
rect 9076 364 9080 396
rect 9040 316 9080 364
rect 9040 284 9044 316
rect 9076 284 9080 316
rect 9040 236 9080 284
rect 9040 204 9044 236
rect 9076 204 9080 236
rect 9040 156 9080 204
rect 9040 124 9044 156
rect 9076 124 9080 156
rect 9040 76 9080 124
rect 9040 44 9044 76
rect 9076 44 9080 76
rect 9040 -4 9080 44
rect 9040 -36 9044 -4
rect 9076 -36 9080 -4
rect 9040 -84 9080 -36
rect 9040 -116 9044 -84
rect 9076 -116 9080 -84
rect 9040 -120 9080 -116
rect 9120 1036 9160 1040
rect 9120 1004 9124 1036
rect 9156 1004 9160 1036
rect 9120 956 9160 1004
rect 9120 924 9124 956
rect 9156 924 9160 956
rect 9120 876 9160 924
rect 9120 844 9124 876
rect 9156 844 9160 876
rect 9120 796 9160 844
rect 9120 764 9124 796
rect 9156 764 9160 796
rect 9120 716 9160 764
rect 9120 684 9124 716
rect 9156 684 9160 716
rect 9120 636 9160 684
rect 9120 604 9124 636
rect 9156 604 9160 636
rect 9120 556 9160 604
rect 9120 524 9124 556
rect 9156 524 9160 556
rect 9120 476 9160 524
rect 9120 444 9124 476
rect 9156 444 9160 476
rect 9120 396 9160 444
rect 9120 364 9124 396
rect 9156 364 9160 396
rect 9120 316 9160 364
rect 9120 284 9124 316
rect 9156 284 9160 316
rect 9120 236 9160 284
rect 9120 204 9124 236
rect 9156 204 9160 236
rect 9120 156 9160 204
rect 9120 124 9124 156
rect 9156 124 9160 156
rect 9120 76 9160 124
rect 9120 44 9124 76
rect 9156 44 9160 76
rect 9120 -4 9160 44
rect 9120 -36 9124 -4
rect 9156 -36 9160 -4
rect 9120 -84 9160 -36
rect 9120 -116 9124 -84
rect 9156 -116 9160 -84
rect 9120 -120 9160 -116
rect 9200 1036 9240 1040
rect 9200 1004 9204 1036
rect 9236 1004 9240 1036
rect 9200 956 9240 1004
rect 9200 924 9204 956
rect 9236 924 9240 956
rect 9200 876 9240 924
rect 9200 844 9204 876
rect 9236 844 9240 876
rect 9200 796 9240 844
rect 9200 764 9204 796
rect 9236 764 9240 796
rect 9200 716 9240 764
rect 9200 684 9204 716
rect 9236 684 9240 716
rect 9200 636 9240 684
rect 9200 604 9204 636
rect 9236 604 9240 636
rect 9200 556 9240 604
rect 9200 524 9204 556
rect 9236 524 9240 556
rect 9200 476 9240 524
rect 9200 444 9204 476
rect 9236 444 9240 476
rect 9200 396 9240 444
rect 9200 364 9204 396
rect 9236 364 9240 396
rect 9200 316 9240 364
rect 9200 284 9204 316
rect 9236 284 9240 316
rect 9200 236 9240 284
rect 9200 204 9204 236
rect 9236 204 9240 236
rect 9200 156 9240 204
rect 9200 124 9204 156
rect 9236 124 9240 156
rect 9200 76 9240 124
rect 9200 44 9204 76
rect 9236 44 9240 76
rect 9200 -4 9240 44
rect 9200 -36 9204 -4
rect 9236 -36 9240 -4
rect 9200 -84 9240 -36
rect 9200 -116 9204 -84
rect 9236 -116 9240 -84
rect 9200 -120 9240 -116
rect 9280 1036 9320 1040
rect 9280 1004 9284 1036
rect 9316 1004 9320 1036
rect 9280 956 9320 1004
rect 9280 924 9284 956
rect 9316 924 9320 956
rect 9280 876 9320 924
rect 9280 844 9284 876
rect 9316 844 9320 876
rect 9280 796 9320 844
rect 9280 764 9284 796
rect 9316 764 9320 796
rect 9280 716 9320 764
rect 9280 684 9284 716
rect 9316 684 9320 716
rect 9280 636 9320 684
rect 9280 604 9284 636
rect 9316 604 9320 636
rect 9280 556 9320 604
rect 9280 524 9284 556
rect 9316 524 9320 556
rect 9280 476 9320 524
rect 9280 444 9284 476
rect 9316 444 9320 476
rect 9280 396 9320 444
rect 9280 364 9284 396
rect 9316 364 9320 396
rect 9280 316 9320 364
rect 9280 284 9284 316
rect 9316 284 9320 316
rect 9280 236 9320 284
rect 9280 204 9284 236
rect 9316 204 9320 236
rect 9280 156 9320 204
rect 9280 124 9284 156
rect 9316 124 9320 156
rect 9280 76 9320 124
rect 9280 44 9284 76
rect 9316 44 9320 76
rect 9280 -4 9320 44
rect 9280 -36 9284 -4
rect 9316 -36 9320 -4
rect 9280 -84 9320 -36
rect 9280 -116 9284 -84
rect 9316 -116 9320 -84
rect 9280 -120 9320 -116
rect 9360 1036 9400 1040
rect 9360 1004 9364 1036
rect 9396 1004 9400 1036
rect 9360 956 9400 1004
rect 9360 924 9364 956
rect 9396 924 9400 956
rect 9360 876 9400 924
rect 9360 844 9364 876
rect 9396 844 9400 876
rect 9360 796 9400 844
rect 9360 764 9364 796
rect 9396 764 9400 796
rect 9360 716 9400 764
rect 9360 684 9364 716
rect 9396 684 9400 716
rect 9360 636 9400 684
rect 9360 604 9364 636
rect 9396 604 9400 636
rect 9360 556 9400 604
rect 9360 524 9364 556
rect 9396 524 9400 556
rect 9360 476 9400 524
rect 9360 444 9364 476
rect 9396 444 9400 476
rect 9360 396 9400 444
rect 9360 364 9364 396
rect 9396 364 9400 396
rect 9360 316 9400 364
rect 9360 284 9364 316
rect 9396 284 9400 316
rect 9360 236 9400 284
rect 9360 204 9364 236
rect 9396 204 9400 236
rect 9360 156 9400 204
rect 9360 124 9364 156
rect 9396 124 9400 156
rect 9360 76 9400 124
rect 9360 44 9364 76
rect 9396 44 9400 76
rect 9360 -4 9400 44
rect 9360 -36 9364 -4
rect 9396 -36 9400 -4
rect 9360 -84 9400 -36
rect 9360 -116 9364 -84
rect 9396 -116 9400 -84
rect 9360 -120 9400 -116
rect 9440 1036 9480 1040
rect 9440 1004 9444 1036
rect 9476 1004 9480 1036
rect 9440 956 9480 1004
rect 9440 924 9444 956
rect 9476 924 9480 956
rect 9440 876 9480 924
rect 9440 844 9444 876
rect 9476 844 9480 876
rect 9440 796 9480 844
rect 9440 764 9444 796
rect 9476 764 9480 796
rect 9440 716 9480 764
rect 9440 684 9444 716
rect 9476 684 9480 716
rect 9440 636 9480 684
rect 9440 604 9444 636
rect 9476 604 9480 636
rect 9440 556 9480 604
rect 9440 524 9444 556
rect 9476 524 9480 556
rect 9440 476 9480 524
rect 9440 444 9444 476
rect 9476 444 9480 476
rect 9440 396 9480 444
rect 9440 364 9444 396
rect 9476 364 9480 396
rect 9440 316 9480 364
rect 9440 284 9444 316
rect 9476 284 9480 316
rect 9440 236 9480 284
rect 9440 204 9444 236
rect 9476 204 9480 236
rect 9440 156 9480 204
rect 9440 124 9444 156
rect 9476 124 9480 156
rect 9440 76 9480 124
rect 9440 44 9444 76
rect 9476 44 9480 76
rect 9440 -4 9480 44
rect 9440 -36 9444 -4
rect 9476 -36 9480 -4
rect 9440 -84 9480 -36
rect 9440 -116 9444 -84
rect 9476 -116 9480 -84
rect 9440 -120 9480 -116
rect 9520 1036 9560 1040
rect 9520 1004 9524 1036
rect 9556 1004 9560 1036
rect 9520 956 9560 1004
rect 9520 924 9524 956
rect 9556 924 9560 956
rect 9520 876 9560 924
rect 9520 844 9524 876
rect 9556 844 9560 876
rect 9520 796 9560 844
rect 9520 764 9524 796
rect 9556 764 9560 796
rect 9520 716 9560 764
rect 9520 684 9524 716
rect 9556 684 9560 716
rect 9520 636 9560 684
rect 9520 604 9524 636
rect 9556 604 9560 636
rect 9520 556 9560 604
rect 9520 524 9524 556
rect 9556 524 9560 556
rect 9520 476 9560 524
rect 9520 444 9524 476
rect 9556 444 9560 476
rect 9520 396 9560 444
rect 9520 364 9524 396
rect 9556 364 9560 396
rect 9520 316 9560 364
rect 9520 284 9524 316
rect 9556 284 9560 316
rect 9520 236 9560 284
rect 9520 204 9524 236
rect 9556 204 9560 236
rect 9520 156 9560 204
rect 9520 124 9524 156
rect 9556 124 9560 156
rect 9520 76 9560 124
rect 9520 44 9524 76
rect 9556 44 9560 76
rect 9520 -4 9560 44
rect 9520 -36 9524 -4
rect 9556 -36 9560 -4
rect 9520 -84 9560 -36
rect 9520 -116 9524 -84
rect 9556 -116 9560 -84
rect 9520 -120 9560 -116
rect 9600 1036 9640 1040
rect 9600 1004 9604 1036
rect 9636 1004 9640 1036
rect 9600 956 9640 1004
rect 9600 924 9604 956
rect 9636 924 9640 956
rect 9600 876 9640 924
rect 9600 844 9604 876
rect 9636 844 9640 876
rect 9600 796 9640 844
rect 9600 764 9604 796
rect 9636 764 9640 796
rect 9600 716 9640 764
rect 9600 684 9604 716
rect 9636 684 9640 716
rect 9600 636 9640 684
rect 9600 604 9604 636
rect 9636 604 9640 636
rect 9600 556 9640 604
rect 9600 524 9604 556
rect 9636 524 9640 556
rect 9600 476 9640 524
rect 9600 444 9604 476
rect 9636 444 9640 476
rect 9600 396 9640 444
rect 9600 364 9604 396
rect 9636 364 9640 396
rect 9600 316 9640 364
rect 9600 284 9604 316
rect 9636 284 9640 316
rect 9600 236 9640 284
rect 9600 204 9604 236
rect 9636 204 9640 236
rect 9600 156 9640 204
rect 9600 124 9604 156
rect 9636 124 9640 156
rect 9600 76 9640 124
rect 9600 44 9604 76
rect 9636 44 9640 76
rect 9600 -4 9640 44
rect 9600 -36 9604 -4
rect 9636 -36 9640 -4
rect 9600 -84 9640 -36
rect 9600 -116 9604 -84
rect 9636 -116 9640 -84
rect 9600 -120 9640 -116
rect 9680 1036 9720 1040
rect 9680 1004 9684 1036
rect 9716 1004 9720 1036
rect 9680 956 9720 1004
rect 9680 924 9684 956
rect 9716 924 9720 956
rect 9680 876 9720 924
rect 9680 844 9684 876
rect 9716 844 9720 876
rect 9680 796 9720 844
rect 9680 764 9684 796
rect 9716 764 9720 796
rect 9680 716 9720 764
rect 9680 684 9684 716
rect 9716 684 9720 716
rect 9680 636 9720 684
rect 9680 604 9684 636
rect 9716 604 9720 636
rect 9680 556 9720 604
rect 9680 524 9684 556
rect 9716 524 9720 556
rect 9680 476 9720 524
rect 9680 444 9684 476
rect 9716 444 9720 476
rect 9680 396 9720 444
rect 9680 364 9684 396
rect 9716 364 9720 396
rect 9680 316 9720 364
rect 9680 284 9684 316
rect 9716 284 9720 316
rect 9680 236 9720 284
rect 9680 204 9684 236
rect 9716 204 9720 236
rect 9680 156 9720 204
rect 9680 124 9684 156
rect 9716 124 9720 156
rect 9680 76 9720 124
rect 9680 44 9684 76
rect 9716 44 9720 76
rect 9680 -4 9720 44
rect 9680 -36 9684 -4
rect 9716 -36 9720 -4
rect 9680 -84 9720 -36
rect 9680 -116 9684 -84
rect 9716 -116 9720 -84
rect 9680 -120 9720 -116
rect 9760 1036 9800 1040
rect 9760 1004 9764 1036
rect 9796 1004 9800 1036
rect 9760 956 9800 1004
rect 9760 924 9764 956
rect 9796 924 9800 956
rect 9760 876 9800 924
rect 9760 844 9764 876
rect 9796 844 9800 876
rect 9760 796 9800 844
rect 9760 764 9764 796
rect 9796 764 9800 796
rect 9760 716 9800 764
rect 9760 684 9764 716
rect 9796 684 9800 716
rect 9760 636 9800 684
rect 9760 604 9764 636
rect 9796 604 9800 636
rect 9760 556 9800 604
rect 9760 524 9764 556
rect 9796 524 9800 556
rect 9760 476 9800 524
rect 9760 444 9764 476
rect 9796 444 9800 476
rect 9760 396 9800 444
rect 9760 364 9764 396
rect 9796 364 9800 396
rect 9760 316 9800 364
rect 9760 284 9764 316
rect 9796 284 9800 316
rect 9760 236 9800 284
rect 9760 204 9764 236
rect 9796 204 9800 236
rect 9760 156 9800 204
rect 9760 124 9764 156
rect 9796 124 9800 156
rect 9760 76 9800 124
rect 9760 44 9764 76
rect 9796 44 9800 76
rect 9760 -4 9800 44
rect 9760 -36 9764 -4
rect 9796 -36 9800 -4
rect 9760 -84 9800 -36
rect 9760 -116 9764 -84
rect 9796 -116 9800 -84
rect 9760 -120 9800 -116
rect 9840 1036 9880 1040
rect 9840 1004 9844 1036
rect 9876 1004 9880 1036
rect 9840 956 9880 1004
rect 9840 924 9844 956
rect 9876 924 9880 956
rect 9840 876 9880 924
rect 9840 844 9844 876
rect 9876 844 9880 876
rect 9840 796 9880 844
rect 9840 764 9844 796
rect 9876 764 9880 796
rect 9840 716 9880 764
rect 9840 684 9844 716
rect 9876 684 9880 716
rect 9840 636 9880 684
rect 9840 604 9844 636
rect 9876 604 9880 636
rect 9840 556 9880 604
rect 9840 524 9844 556
rect 9876 524 9880 556
rect 9840 476 9880 524
rect 9840 444 9844 476
rect 9876 444 9880 476
rect 9840 396 9880 444
rect 9840 364 9844 396
rect 9876 364 9880 396
rect 9840 316 9880 364
rect 9840 284 9844 316
rect 9876 284 9880 316
rect 9840 236 9880 284
rect 9840 204 9844 236
rect 9876 204 9880 236
rect 9840 156 9880 204
rect 9840 124 9844 156
rect 9876 124 9880 156
rect 9840 76 9880 124
rect 9840 44 9844 76
rect 9876 44 9880 76
rect 9840 -4 9880 44
rect 9840 -36 9844 -4
rect 9876 -36 9880 -4
rect 9840 -84 9880 -36
rect 9840 -116 9844 -84
rect 9876 -116 9880 -84
rect 9840 -120 9880 -116
rect 9920 1036 9960 1040
rect 9920 1004 9924 1036
rect 9956 1004 9960 1036
rect 9920 956 9960 1004
rect 9920 924 9924 956
rect 9956 924 9960 956
rect 9920 876 9960 924
rect 9920 844 9924 876
rect 9956 844 9960 876
rect 9920 796 9960 844
rect 9920 764 9924 796
rect 9956 764 9960 796
rect 9920 716 9960 764
rect 9920 684 9924 716
rect 9956 684 9960 716
rect 9920 636 9960 684
rect 9920 604 9924 636
rect 9956 604 9960 636
rect 9920 556 9960 604
rect 9920 524 9924 556
rect 9956 524 9960 556
rect 9920 476 9960 524
rect 9920 444 9924 476
rect 9956 444 9960 476
rect 9920 396 9960 444
rect 9920 364 9924 396
rect 9956 364 9960 396
rect 9920 316 9960 364
rect 9920 284 9924 316
rect 9956 284 9960 316
rect 9920 236 9960 284
rect 9920 204 9924 236
rect 9956 204 9960 236
rect 9920 156 9960 204
rect 9920 124 9924 156
rect 9956 124 9960 156
rect 9920 76 9960 124
rect 9920 44 9924 76
rect 9956 44 9960 76
rect 9920 -4 9960 44
rect 9920 -36 9924 -4
rect 9956 -36 9960 -4
rect 9920 -84 9960 -36
rect 9920 -116 9924 -84
rect 9956 -116 9960 -84
rect 9920 -120 9960 -116
rect 10000 1036 10040 1040
rect 10000 1004 10004 1036
rect 10036 1004 10040 1036
rect 10000 956 10040 1004
rect 10000 924 10004 956
rect 10036 924 10040 956
rect 10000 876 10040 924
rect 10000 844 10004 876
rect 10036 844 10040 876
rect 10000 796 10040 844
rect 10000 764 10004 796
rect 10036 764 10040 796
rect 10000 716 10040 764
rect 10000 684 10004 716
rect 10036 684 10040 716
rect 10000 636 10040 684
rect 10000 604 10004 636
rect 10036 604 10040 636
rect 10000 556 10040 604
rect 10000 524 10004 556
rect 10036 524 10040 556
rect 10000 476 10040 524
rect 10000 444 10004 476
rect 10036 444 10040 476
rect 10000 396 10040 444
rect 10000 364 10004 396
rect 10036 364 10040 396
rect 10000 316 10040 364
rect 10000 284 10004 316
rect 10036 284 10040 316
rect 10000 236 10040 284
rect 10000 204 10004 236
rect 10036 204 10040 236
rect 10000 156 10040 204
rect 10000 124 10004 156
rect 10036 124 10040 156
rect 10000 76 10040 124
rect 10000 44 10004 76
rect 10036 44 10040 76
rect 10000 -4 10040 44
rect 10000 -36 10004 -4
rect 10036 -36 10040 -4
rect 10000 -84 10040 -36
rect 10000 -116 10004 -84
rect 10036 -116 10040 -84
rect 10000 -120 10040 -116
rect 10080 1036 10120 1040
rect 10080 1004 10084 1036
rect 10116 1004 10120 1036
rect 10080 956 10120 1004
rect 10080 924 10084 956
rect 10116 924 10120 956
rect 10080 876 10120 924
rect 10080 844 10084 876
rect 10116 844 10120 876
rect 10080 796 10120 844
rect 10080 764 10084 796
rect 10116 764 10120 796
rect 10080 716 10120 764
rect 10080 684 10084 716
rect 10116 684 10120 716
rect 10080 636 10120 684
rect 10080 604 10084 636
rect 10116 604 10120 636
rect 10080 556 10120 604
rect 10080 524 10084 556
rect 10116 524 10120 556
rect 10080 476 10120 524
rect 10080 444 10084 476
rect 10116 444 10120 476
rect 10080 396 10120 444
rect 10080 364 10084 396
rect 10116 364 10120 396
rect 10080 316 10120 364
rect 10080 284 10084 316
rect 10116 284 10120 316
rect 10080 236 10120 284
rect 10080 204 10084 236
rect 10116 204 10120 236
rect 10080 156 10120 204
rect 10080 124 10084 156
rect 10116 124 10120 156
rect 10080 76 10120 124
rect 10080 44 10084 76
rect 10116 44 10120 76
rect 10080 -4 10120 44
rect 10080 -36 10084 -4
rect 10116 -36 10120 -4
rect 10080 -84 10120 -36
rect 10080 -116 10084 -84
rect 10116 -116 10120 -84
rect 10080 -120 10120 -116
rect 10160 1036 10200 1040
rect 10160 1004 10164 1036
rect 10196 1004 10200 1036
rect 10160 956 10200 1004
rect 10160 924 10164 956
rect 10196 924 10200 956
rect 10160 876 10200 924
rect 10160 844 10164 876
rect 10196 844 10200 876
rect 10160 796 10200 844
rect 10160 764 10164 796
rect 10196 764 10200 796
rect 10160 716 10200 764
rect 10160 684 10164 716
rect 10196 684 10200 716
rect 10160 636 10200 684
rect 10160 604 10164 636
rect 10196 604 10200 636
rect 10160 556 10200 604
rect 10160 524 10164 556
rect 10196 524 10200 556
rect 10160 476 10200 524
rect 10160 444 10164 476
rect 10196 444 10200 476
rect 10160 396 10200 444
rect 10160 364 10164 396
rect 10196 364 10200 396
rect 10160 316 10200 364
rect 10160 284 10164 316
rect 10196 284 10200 316
rect 10160 236 10200 284
rect 10160 204 10164 236
rect 10196 204 10200 236
rect 10160 156 10200 204
rect 10160 124 10164 156
rect 10196 124 10200 156
rect 10160 76 10200 124
rect 10160 44 10164 76
rect 10196 44 10200 76
rect 10160 -4 10200 44
rect 10160 -36 10164 -4
rect 10196 -36 10200 -4
rect 10160 -84 10200 -36
rect 10160 -116 10164 -84
rect 10196 -116 10200 -84
rect 10160 -120 10200 -116
rect 10240 1036 10280 1040
rect 10240 1004 10244 1036
rect 10276 1004 10280 1036
rect 10240 956 10280 1004
rect 10240 924 10244 956
rect 10276 924 10280 956
rect 10240 876 10280 924
rect 10240 844 10244 876
rect 10276 844 10280 876
rect 10240 796 10280 844
rect 10240 764 10244 796
rect 10276 764 10280 796
rect 10240 716 10280 764
rect 10240 684 10244 716
rect 10276 684 10280 716
rect 10240 636 10280 684
rect 10240 604 10244 636
rect 10276 604 10280 636
rect 10240 556 10280 604
rect 10240 524 10244 556
rect 10276 524 10280 556
rect 10240 476 10280 524
rect 10240 444 10244 476
rect 10276 444 10280 476
rect 10240 396 10280 444
rect 10240 364 10244 396
rect 10276 364 10280 396
rect 10240 316 10280 364
rect 10240 284 10244 316
rect 10276 284 10280 316
rect 10240 236 10280 284
rect 10240 204 10244 236
rect 10276 204 10280 236
rect 10240 156 10280 204
rect 10240 124 10244 156
rect 10276 124 10280 156
rect 10240 76 10280 124
rect 10240 44 10244 76
rect 10276 44 10280 76
rect 10240 -4 10280 44
rect 10240 -36 10244 -4
rect 10276 -36 10280 -4
rect 10240 -84 10280 -36
rect 10240 -116 10244 -84
rect 10276 -116 10280 -84
rect 10240 -120 10280 -116
rect 10320 1036 10360 1040
rect 10320 1004 10324 1036
rect 10356 1004 10360 1036
rect 10320 956 10360 1004
rect 10320 924 10324 956
rect 10356 924 10360 956
rect 10320 876 10360 924
rect 10320 844 10324 876
rect 10356 844 10360 876
rect 10320 796 10360 844
rect 10320 764 10324 796
rect 10356 764 10360 796
rect 10320 716 10360 764
rect 10320 684 10324 716
rect 10356 684 10360 716
rect 10320 636 10360 684
rect 10320 604 10324 636
rect 10356 604 10360 636
rect 10320 556 10360 604
rect 10320 524 10324 556
rect 10356 524 10360 556
rect 10320 476 10360 524
rect 10320 444 10324 476
rect 10356 444 10360 476
rect 10320 396 10360 444
rect 10320 364 10324 396
rect 10356 364 10360 396
rect 10320 316 10360 364
rect 10320 284 10324 316
rect 10356 284 10360 316
rect 10320 236 10360 284
rect 10320 204 10324 236
rect 10356 204 10360 236
rect 10320 156 10360 204
rect 10320 124 10324 156
rect 10356 124 10360 156
rect 10320 76 10360 124
rect 10320 44 10324 76
rect 10356 44 10360 76
rect 10320 -4 10360 44
rect 10320 -36 10324 -4
rect 10356 -36 10360 -4
rect 10320 -84 10360 -36
rect 10320 -116 10324 -84
rect 10356 -116 10360 -84
rect 10320 -120 10360 -116
rect 10400 1036 10440 1040
rect 10400 1004 10404 1036
rect 10436 1004 10440 1036
rect 10400 956 10440 1004
rect 10400 924 10404 956
rect 10436 924 10440 956
rect 10400 876 10440 924
rect 10400 844 10404 876
rect 10436 844 10440 876
rect 10400 796 10440 844
rect 10400 764 10404 796
rect 10436 764 10440 796
rect 10400 716 10440 764
rect 10400 684 10404 716
rect 10436 684 10440 716
rect 10400 636 10440 684
rect 10400 604 10404 636
rect 10436 604 10440 636
rect 10400 556 10440 604
rect 10400 524 10404 556
rect 10436 524 10440 556
rect 10400 476 10440 524
rect 10400 444 10404 476
rect 10436 444 10440 476
rect 10400 396 10440 444
rect 10400 364 10404 396
rect 10436 364 10440 396
rect 10400 316 10440 364
rect 10400 284 10404 316
rect 10436 284 10440 316
rect 10400 236 10440 284
rect 10400 204 10404 236
rect 10436 204 10440 236
rect 10400 156 10440 204
rect 10400 124 10404 156
rect 10436 124 10440 156
rect 10400 76 10440 124
rect 10400 44 10404 76
rect 10436 44 10440 76
rect 10400 -4 10440 44
rect 10400 -36 10404 -4
rect 10436 -36 10440 -4
rect 10400 -84 10440 -36
rect 10400 -116 10404 -84
rect 10436 -116 10440 -84
rect 10400 -120 10440 -116
rect 10480 1036 10520 1040
rect 10480 1004 10484 1036
rect 10516 1004 10520 1036
rect 10480 956 10520 1004
rect 10480 924 10484 956
rect 10516 924 10520 956
rect 10480 876 10520 924
rect 10480 844 10484 876
rect 10516 844 10520 876
rect 10480 796 10520 844
rect 10480 764 10484 796
rect 10516 764 10520 796
rect 10480 716 10520 764
rect 10480 684 10484 716
rect 10516 684 10520 716
rect 10480 636 10520 684
rect 10480 604 10484 636
rect 10516 604 10520 636
rect 10480 556 10520 604
rect 10480 524 10484 556
rect 10516 524 10520 556
rect 10480 476 10520 524
rect 10480 444 10484 476
rect 10516 444 10520 476
rect 10480 396 10520 444
rect 10480 364 10484 396
rect 10516 364 10520 396
rect 10480 316 10520 364
rect 10480 284 10484 316
rect 10516 284 10520 316
rect 10480 236 10520 284
rect 10480 204 10484 236
rect 10516 204 10520 236
rect 10480 156 10520 204
rect 10480 124 10484 156
rect 10516 124 10520 156
rect 10480 76 10520 124
rect 10480 44 10484 76
rect 10516 44 10520 76
rect 10480 -4 10520 44
rect 10480 -36 10484 -4
rect 10516 -36 10520 -4
rect 10480 -84 10520 -36
rect 10480 -116 10484 -84
rect 10516 -116 10520 -84
rect 10480 -120 10520 -116
rect 10560 -120 10600 1040
rect 10640 1036 10680 1040
rect 10640 1004 10644 1036
rect 10676 1004 10680 1036
rect 10640 956 10680 1004
rect 10640 924 10644 956
rect 10676 924 10680 956
rect 10640 876 10680 924
rect 10640 844 10644 876
rect 10676 844 10680 876
rect 10640 796 10680 844
rect 10640 764 10644 796
rect 10676 764 10680 796
rect 10640 716 10680 764
rect 10640 684 10644 716
rect 10676 684 10680 716
rect 10640 636 10680 684
rect 10640 604 10644 636
rect 10676 604 10680 636
rect 10640 556 10680 604
rect 10640 524 10644 556
rect 10676 524 10680 556
rect 10640 476 10680 524
rect 10640 444 10644 476
rect 10676 444 10680 476
rect 10640 396 10680 444
rect 10640 364 10644 396
rect 10676 364 10680 396
rect 10640 316 10680 364
rect 10640 284 10644 316
rect 10676 284 10680 316
rect 10640 236 10680 284
rect 10640 204 10644 236
rect 10676 204 10680 236
rect 10640 156 10680 204
rect 10640 124 10644 156
rect 10676 124 10680 156
rect 10640 76 10680 124
rect 10640 44 10644 76
rect 10676 44 10680 76
rect 10640 -4 10680 44
rect 10640 -36 10644 -4
rect 10676 -36 10680 -4
rect 10640 -84 10680 -36
rect 10640 -116 10644 -84
rect 10676 -116 10680 -84
rect 10640 -120 10680 -116
rect 10720 155 10760 1080
rect 10720 125 10725 155
rect 10755 125 10760 155
rect 10720 -120 10760 125
rect 10800 1036 10840 1040
rect 10800 1004 10804 1036
rect 10836 1004 10840 1036
rect 10800 956 10840 1004
rect 10800 924 10804 956
rect 10836 924 10840 956
rect 10800 876 10840 924
rect 10800 844 10804 876
rect 10836 844 10840 876
rect 10800 796 10840 844
rect 10800 764 10804 796
rect 10836 764 10840 796
rect 10800 716 10840 764
rect 10800 684 10804 716
rect 10836 684 10840 716
rect 10800 636 10840 684
rect 10800 604 10804 636
rect 10836 604 10840 636
rect 10800 556 10840 604
rect 10800 524 10804 556
rect 10836 524 10840 556
rect 10800 476 10840 524
rect 10800 444 10804 476
rect 10836 444 10840 476
rect 10800 396 10840 444
rect 10800 364 10804 396
rect 10836 364 10840 396
rect 10800 316 10840 364
rect 10800 284 10804 316
rect 10836 284 10840 316
rect 10800 236 10840 284
rect 10800 204 10804 236
rect 10836 204 10840 236
rect 10800 156 10840 204
rect 10800 124 10804 156
rect 10836 124 10840 156
rect 10800 76 10840 124
rect 10800 44 10804 76
rect 10836 44 10840 76
rect 10800 -4 10840 44
rect 10800 -36 10804 -4
rect 10836 -36 10840 -4
rect 10800 -84 10840 -36
rect 10800 -116 10804 -84
rect 10836 -116 10840 -84
rect 10800 -120 10840 -116
rect 10880 315 10920 1080
rect 10880 285 10885 315
rect 10915 285 10920 315
rect 10880 -120 10920 285
rect 10960 1036 11000 1080
rect 10960 1004 10964 1036
rect 10996 1004 11000 1036
rect 10960 956 11000 1004
rect 10960 924 10964 956
rect 10996 924 11000 956
rect 10960 876 11000 924
rect 10960 844 10964 876
rect 10996 844 11000 876
rect 10960 796 11000 844
rect 10960 764 10964 796
rect 10996 764 11000 796
rect 10960 716 11000 764
rect 10960 684 10964 716
rect 10996 684 11000 716
rect 10960 636 11000 684
rect 10960 604 10964 636
rect 10996 604 11000 636
rect 10960 556 11000 604
rect 10960 524 10964 556
rect 10996 524 11000 556
rect 10960 476 11000 524
rect 10960 444 10964 476
rect 10996 444 11000 476
rect 10960 396 11000 444
rect 10960 364 10964 396
rect 10996 364 11000 396
rect 10960 316 11000 364
rect 10960 284 10964 316
rect 10996 284 11000 316
rect 10960 236 11000 284
rect 10960 204 10964 236
rect 10996 204 11000 236
rect 10960 156 11000 204
rect 10960 124 10964 156
rect 10996 124 11000 156
rect 10960 76 11000 124
rect 10960 44 10964 76
rect 10996 44 11000 76
rect 10960 -4 11000 44
rect 10960 -36 10964 -4
rect 10996 -36 11000 -4
rect 10960 -84 11000 -36
rect 10960 -116 10964 -84
rect 10996 -116 11000 -84
rect 10960 -120 11000 -116
<< via3 >>
rect -716 1035 -684 1036
rect -716 1005 -715 1035
rect -715 1005 -685 1035
rect -685 1005 -684 1035
rect -716 1004 -684 1005
rect -716 955 -684 956
rect -716 925 -715 955
rect -715 925 -685 955
rect -685 925 -684 955
rect -716 924 -684 925
rect -716 875 -684 876
rect -716 845 -715 875
rect -715 845 -685 875
rect -685 845 -684 875
rect -716 844 -684 845
rect -716 764 -684 796
rect -716 684 -684 716
rect -716 635 -684 636
rect -716 605 -715 635
rect -715 605 -685 635
rect -685 605 -684 635
rect -716 604 -684 605
rect -716 555 -684 556
rect -716 525 -715 555
rect -715 525 -685 555
rect -685 525 -684 555
rect -716 524 -684 525
rect -716 475 -684 476
rect -716 445 -715 475
rect -715 445 -685 475
rect -685 445 -684 475
rect -716 444 -684 445
rect -716 395 -684 396
rect -716 365 -715 395
rect -715 365 -685 395
rect -685 365 -684 395
rect -716 364 -684 365
rect -716 315 -684 316
rect -716 285 -715 315
rect -715 285 -685 315
rect -685 285 -684 315
rect -716 284 -684 285
rect -716 235 -684 236
rect -716 205 -715 235
rect -715 205 -685 235
rect -685 205 -684 235
rect -716 204 -684 205
rect -716 155 -684 156
rect -716 125 -715 155
rect -715 125 -685 155
rect -685 125 -684 155
rect -716 124 -684 125
rect -716 75 -684 76
rect -716 45 -715 75
rect -715 45 -685 75
rect -685 45 -684 75
rect -716 44 -684 45
rect -716 -5 -684 -4
rect -716 -35 -715 -5
rect -715 -35 -685 -5
rect -685 -35 -684 -5
rect -716 -36 -684 -35
rect -716 -85 -684 -84
rect -716 -115 -715 -85
rect -715 -115 -685 -85
rect -685 -115 -684 -85
rect -716 -116 -684 -115
rect -556 1035 -524 1036
rect -556 1005 -555 1035
rect -555 1005 -525 1035
rect -525 1005 -524 1035
rect -556 1004 -524 1005
rect -556 955 -524 956
rect -556 925 -555 955
rect -555 925 -525 955
rect -525 925 -524 955
rect -556 924 -524 925
rect -556 875 -524 876
rect -556 845 -555 875
rect -555 845 -525 875
rect -525 845 -524 875
rect -556 844 -524 845
rect -556 764 -524 796
rect -556 684 -524 716
rect -556 635 -524 636
rect -556 605 -555 635
rect -555 605 -525 635
rect -525 605 -524 635
rect -556 604 -524 605
rect -556 555 -524 556
rect -556 525 -555 555
rect -555 525 -525 555
rect -525 525 -524 555
rect -556 524 -524 525
rect -556 475 -524 476
rect -556 445 -555 475
rect -555 445 -525 475
rect -525 445 -524 475
rect -556 444 -524 445
rect -556 395 -524 396
rect -556 365 -555 395
rect -555 365 -525 395
rect -525 365 -524 395
rect -556 364 -524 365
rect -556 315 -524 316
rect -556 285 -555 315
rect -555 285 -525 315
rect -525 285 -524 315
rect -556 284 -524 285
rect -556 235 -524 236
rect -556 205 -555 235
rect -555 205 -525 235
rect -525 205 -524 235
rect -556 204 -524 205
rect -556 155 -524 156
rect -556 125 -555 155
rect -555 125 -525 155
rect -525 125 -524 155
rect -556 124 -524 125
rect -556 75 -524 76
rect -556 45 -555 75
rect -555 45 -525 75
rect -525 45 -524 75
rect -556 44 -524 45
rect -556 -5 -524 -4
rect -556 -35 -555 -5
rect -555 -35 -525 -5
rect -525 -35 -524 -5
rect -556 -36 -524 -35
rect -556 -85 -524 -84
rect -556 -115 -555 -85
rect -555 -115 -525 -85
rect -525 -115 -524 -85
rect -556 -116 -524 -115
rect -396 1035 -364 1036
rect -396 1005 -395 1035
rect -395 1005 -365 1035
rect -365 1005 -364 1035
rect -396 1004 -364 1005
rect -396 955 -364 956
rect -396 925 -395 955
rect -395 925 -365 955
rect -365 925 -364 955
rect -396 924 -364 925
rect -396 875 -364 876
rect -396 845 -395 875
rect -395 845 -365 875
rect -365 845 -364 875
rect -396 844 -364 845
rect -396 764 -364 796
rect -396 684 -364 716
rect -396 635 -364 636
rect -396 605 -395 635
rect -395 605 -365 635
rect -365 605 -364 635
rect -396 604 -364 605
rect -396 555 -364 556
rect -396 525 -395 555
rect -395 525 -365 555
rect -365 525 -364 555
rect -396 524 -364 525
rect -396 444 -364 476
rect -396 395 -364 396
rect -396 365 -395 395
rect -395 365 -365 395
rect -365 365 -364 395
rect -396 364 -364 365
rect -396 315 -364 316
rect -396 285 -395 315
rect -395 285 -365 315
rect -365 285 -364 315
rect -396 284 -364 285
rect -396 235 -364 236
rect -396 205 -395 235
rect -395 205 -365 235
rect -365 205 -364 235
rect -396 204 -364 205
rect -396 155 -364 156
rect -396 125 -395 155
rect -395 125 -365 155
rect -365 125 -364 155
rect -396 124 -364 125
rect -396 75 -364 76
rect -396 45 -395 75
rect -395 45 -365 75
rect -365 45 -364 75
rect -396 44 -364 45
rect -396 -5 -364 -4
rect -396 -35 -395 -5
rect -395 -35 -365 -5
rect -365 -35 -364 -5
rect -396 -36 -364 -35
rect -396 -85 -364 -84
rect -396 -115 -395 -85
rect -395 -115 -365 -85
rect -365 -115 -364 -85
rect -396 -116 -364 -115
rect -316 1035 -284 1036
rect -316 1005 -315 1035
rect -315 1005 -285 1035
rect -285 1005 -284 1035
rect -316 1004 -284 1005
rect -316 955 -284 956
rect -316 925 -315 955
rect -315 925 -285 955
rect -285 925 -284 955
rect -316 924 -284 925
rect -316 875 -284 876
rect -316 845 -315 875
rect -315 845 -285 875
rect -285 845 -284 875
rect -316 844 -284 845
rect -316 764 -284 796
rect -316 684 -284 716
rect -316 635 -284 636
rect -316 605 -315 635
rect -315 605 -285 635
rect -285 605 -284 635
rect -316 604 -284 605
rect -316 555 -284 556
rect -316 525 -315 555
rect -315 525 -285 555
rect -285 525 -284 555
rect -316 524 -284 525
rect -316 444 -284 476
rect -316 395 -284 396
rect -316 365 -315 395
rect -315 365 -285 395
rect -285 365 -284 395
rect -316 364 -284 365
rect -316 284 -284 316
rect -316 235 -284 236
rect -316 205 -315 235
rect -315 205 -285 235
rect -285 205 -284 235
rect -316 204 -284 205
rect -316 124 -284 156
rect -316 75 -284 76
rect -316 45 -315 75
rect -315 45 -285 75
rect -285 45 -284 75
rect -316 44 -284 45
rect -316 -5 -284 -4
rect -316 -35 -315 -5
rect -315 -35 -285 -5
rect -285 -35 -284 -5
rect -316 -36 -284 -35
rect -316 -85 -284 -84
rect -316 -115 -315 -85
rect -315 -115 -285 -85
rect -285 -115 -284 -85
rect -316 -116 -284 -115
rect -236 1035 -204 1036
rect -236 1005 -235 1035
rect -235 1005 -205 1035
rect -205 1005 -204 1035
rect -236 1004 -204 1005
rect -236 955 -204 956
rect -236 925 -235 955
rect -235 925 -205 955
rect -205 925 -204 955
rect -236 924 -204 925
rect -236 875 -204 876
rect -236 845 -235 875
rect -235 845 -205 875
rect -205 845 -204 875
rect -236 844 -204 845
rect -236 764 -204 796
rect -236 684 -204 716
rect -236 635 -204 636
rect -236 605 -235 635
rect -235 605 -205 635
rect -205 605 -204 635
rect -236 604 -204 605
rect -236 555 -204 556
rect -236 525 -235 555
rect -235 525 -205 555
rect -205 525 -204 555
rect -236 524 -204 525
rect -236 444 -204 476
rect -236 395 -204 396
rect -236 365 -235 395
rect -235 365 -205 395
rect -205 365 -204 395
rect -236 364 -204 365
rect -236 284 -204 316
rect -236 235 -204 236
rect -236 205 -235 235
rect -235 205 -205 235
rect -205 205 -204 235
rect -236 204 -204 205
rect -236 124 -204 156
rect -236 75 -204 76
rect -236 45 -235 75
rect -235 45 -205 75
rect -205 45 -204 75
rect -236 44 -204 45
rect -236 -5 -204 -4
rect -236 -35 -235 -5
rect -235 -35 -205 -5
rect -205 -35 -204 -5
rect -236 -36 -204 -35
rect -236 -85 -204 -84
rect -236 -115 -235 -85
rect -235 -115 -205 -85
rect -205 -115 -204 -85
rect -236 -116 -204 -115
rect -156 1035 -124 1036
rect -156 1005 -155 1035
rect -155 1005 -125 1035
rect -125 1005 -124 1035
rect -156 1004 -124 1005
rect -156 955 -124 956
rect -156 925 -155 955
rect -155 925 -125 955
rect -125 925 -124 955
rect -156 924 -124 925
rect -156 875 -124 876
rect -156 845 -155 875
rect -155 845 -125 875
rect -125 845 -124 875
rect -156 844 -124 845
rect -156 764 -124 796
rect -156 684 -124 716
rect -156 635 -124 636
rect -156 605 -155 635
rect -155 605 -125 635
rect -125 605 -124 635
rect -156 604 -124 605
rect -156 555 -124 556
rect -156 525 -155 555
rect -155 525 -125 555
rect -125 525 -124 555
rect -156 524 -124 525
rect -156 444 -124 476
rect -156 395 -124 396
rect -156 365 -155 395
rect -155 365 -125 395
rect -125 365 -124 395
rect -156 364 -124 365
rect -156 284 -124 316
rect -156 235 -124 236
rect -156 205 -155 235
rect -155 205 -125 235
rect -125 205 -124 235
rect -156 204 -124 205
rect -156 124 -124 156
rect -156 75 -124 76
rect -156 45 -155 75
rect -155 45 -125 75
rect -125 45 -124 75
rect -156 44 -124 45
rect -156 -5 -124 -4
rect -156 -35 -155 -5
rect -155 -35 -125 -5
rect -125 -35 -124 -5
rect -156 -36 -124 -35
rect -156 -85 -124 -84
rect -156 -115 -155 -85
rect -155 -115 -125 -85
rect -125 -115 -124 -85
rect -156 -116 -124 -115
rect -76 1035 -44 1036
rect -76 1005 -75 1035
rect -75 1005 -45 1035
rect -45 1005 -44 1035
rect -76 1004 -44 1005
rect -76 955 -44 956
rect -76 925 -75 955
rect -75 925 -45 955
rect -45 925 -44 955
rect -76 924 -44 925
rect -76 875 -44 876
rect -76 845 -75 875
rect -75 845 -45 875
rect -45 845 -44 875
rect -76 844 -44 845
rect -76 764 -44 796
rect -76 684 -44 716
rect -76 635 -44 636
rect -76 605 -75 635
rect -75 605 -45 635
rect -45 605 -44 635
rect -76 604 -44 605
rect -76 555 -44 556
rect -76 525 -75 555
rect -75 525 -45 555
rect -45 525 -44 555
rect -76 524 -44 525
rect -76 444 -44 476
rect -76 395 -44 396
rect -76 365 -75 395
rect -75 365 -45 395
rect -45 365 -44 395
rect -76 364 -44 365
rect -76 284 -44 316
rect -76 235 -44 236
rect -76 205 -75 235
rect -75 205 -45 235
rect -45 205 -44 235
rect -76 204 -44 205
rect -76 124 -44 156
rect -76 75 -44 76
rect -76 45 -75 75
rect -75 45 -45 75
rect -45 45 -44 75
rect -76 44 -44 45
rect -76 -5 -44 -4
rect -76 -35 -75 -5
rect -75 -35 -45 -5
rect -45 -35 -44 -5
rect -76 -36 -44 -35
rect -76 -85 -44 -84
rect -76 -115 -75 -85
rect -75 -115 -45 -85
rect -45 -115 -44 -85
rect -76 -116 -44 -115
rect 4 1035 36 1036
rect 4 1005 5 1035
rect 5 1005 35 1035
rect 35 1005 36 1035
rect 4 1004 36 1005
rect 4 955 36 956
rect 4 925 5 955
rect 5 925 35 955
rect 35 925 36 955
rect 4 924 36 925
rect 4 875 36 876
rect 4 845 5 875
rect 5 845 35 875
rect 35 845 36 875
rect 4 844 36 845
rect 4 764 36 796
rect 4 684 36 716
rect 4 635 36 636
rect 4 605 5 635
rect 5 605 35 635
rect 35 605 36 635
rect 4 604 36 605
rect 4 555 36 556
rect 4 525 5 555
rect 5 525 35 555
rect 35 525 36 555
rect 4 524 36 525
rect 4 444 36 476
rect 4 395 36 396
rect 4 365 5 395
rect 5 365 35 395
rect 35 365 36 395
rect 4 364 36 365
rect 4 284 36 316
rect 4 235 36 236
rect 4 205 5 235
rect 5 205 35 235
rect 35 205 36 235
rect 4 204 36 205
rect 4 124 36 156
rect 4 75 36 76
rect 4 45 5 75
rect 5 45 35 75
rect 35 45 36 75
rect 4 44 36 45
rect 4 -5 36 -4
rect 4 -35 5 -5
rect 5 -35 35 -5
rect 35 -35 36 -5
rect 4 -36 36 -35
rect 4 -85 36 -84
rect 4 -115 5 -85
rect 5 -115 35 -85
rect 35 -115 36 -85
rect 4 -116 36 -115
rect 84 1035 116 1036
rect 84 1005 85 1035
rect 85 1005 115 1035
rect 115 1005 116 1035
rect 84 1004 116 1005
rect 84 955 116 956
rect 84 925 85 955
rect 85 925 115 955
rect 115 925 116 955
rect 84 924 116 925
rect 84 875 116 876
rect 84 845 85 875
rect 85 845 115 875
rect 115 845 116 875
rect 84 844 116 845
rect 84 764 116 796
rect 84 684 116 716
rect 84 635 116 636
rect 84 605 85 635
rect 85 605 115 635
rect 115 605 116 635
rect 84 604 116 605
rect 84 555 116 556
rect 84 525 85 555
rect 85 525 115 555
rect 115 525 116 555
rect 84 524 116 525
rect 84 444 116 476
rect 84 395 116 396
rect 84 365 85 395
rect 85 365 115 395
rect 115 365 116 395
rect 84 364 116 365
rect 84 284 116 316
rect 84 235 116 236
rect 84 205 85 235
rect 85 205 115 235
rect 115 205 116 235
rect 84 204 116 205
rect 84 124 116 156
rect 84 75 116 76
rect 84 45 85 75
rect 85 45 115 75
rect 115 45 116 75
rect 84 44 116 45
rect 84 -5 116 -4
rect 84 -35 85 -5
rect 85 -35 115 -5
rect 115 -35 116 -5
rect 84 -36 116 -35
rect 84 -85 116 -84
rect 84 -115 85 -85
rect 85 -115 115 -85
rect 115 -115 116 -85
rect 84 -116 116 -115
rect 164 1035 196 1036
rect 164 1005 165 1035
rect 165 1005 195 1035
rect 195 1005 196 1035
rect 164 1004 196 1005
rect 164 955 196 956
rect 164 925 165 955
rect 165 925 195 955
rect 195 925 196 955
rect 164 924 196 925
rect 164 875 196 876
rect 164 845 165 875
rect 165 845 195 875
rect 195 845 196 875
rect 164 844 196 845
rect 164 764 196 796
rect 164 684 196 716
rect 164 635 196 636
rect 164 605 165 635
rect 165 605 195 635
rect 195 605 196 635
rect 164 604 196 605
rect 164 555 196 556
rect 164 525 165 555
rect 165 525 195 555
rect 195 525 196 555
rect 164 524 196 525
rect 164 444 196 476
rect 164 395 196 396
rect 164 365 165 395
rect 165 365 195 395
rect 195 365 196 395
rect 164 364 196 365
rect 164 284 196 316
rect 164 235 196 236
rect 164 205 165 235
rect 165 205 195 235
rect 195 205 196 235
rect 164 204 196 205
rect 164 124 196 156
rect 164 75 196 76
rect 164 45 165 75
rect 165 45 195 75
rect 195 45 196 75
rect 164 44 196 45
rect 164 -5 196 -4
rect 164 -35 165 -5
rect 165 -35 195 -5
rect 195 -35 196 -5
rect 164 -36 196 -35
rect 164 -85 196 -84
rect 164 -115 165 -85
rect 165 -115 195 -85
rect 195 -115 196 -85
rect 164 -116 196 -115
rect 244 1035 276 1036
rect 244 1005 245 1035
rect 245 1005 275 1035
rect 275 1005 276 1035
rect 244 1004 276 1005
rect 244 955 276 956
rect 244 925 245 955
rect 245 925 275 955
rect 275 925 276 955
rect 244 924 276 925
rect 244 875 276 876
rect 244 845 245 875
rect 245 845 275 875
rect 275 845 276 875
rect 244 844 276 845
rect 244 764 276 796
rect 244 684 276 716
rect 244 635 276 636
rect 244 605 245 635
rect 245 605 275 635
rect 275 605 276 635
rect 244 604 276 605
rect 244 555 276 556
rect 244 525 245 555
rect 245 525 275 555
rect 275 525 276 555
rect 244 524 276 525
rect 244 444 276 476
rect 244 395 276 396
rect 244 365 245 395
rect 245 365 275 395
rect 275 365 276 395
rect 244 364 276 365
rect 244 284 276 316
rect 244 235 276 236
rect 244 205 245 235
rect 245 205 275 235
rect 275 205 276 235
rect 244 204 276 205
rect 244 124 276 156
rect 244 75 276 76
rect 244 45 245 75
rect 245 45 275 75
rect 275 45 276 75
rect 244 44 276 45
rect 244 -5 276 -4
rect 244 -35 245 -5
rect 245 -35 275 -5
rect 275 -35 276 -5
rect 244 -36 276 -35
rect 244 -85 276 -84
rect 244 -115 245 -85
rect 245 -115 275 -85
rect 275 -115 276 -85
rect 244 -116 276 -115
rect 324 1035 356 1036
rect 324 1005 325 1035
rect 325 1005 355 1035
rect 355 1005 356 1035
rect 324 1004 356 1005
rect 324 955 356 956
rect 324 925 325 955
rect 325 925 355 955
rect 355 925 356 955
rect 324 924 356 925
rect 324 875 356 876
rect 324 845 325 875
rect 325 845 355 875
rect 355 845 356 875
rect 324 844 356 845
rect 324 764 356 796
rect 324 684 356 716
rect 324 635 356 636
rect 324 605 325 635
rect 325 605 355 635
rect 355 605 356 635
rect 324 604 356 605
rect 324 555 356 556
rect 324 525 325 555
rect 325 525 355 555
rect 355 525 356 555
rect 324 524 356 525
rect 324 444 356 476
rect 324 395 356 396
rect 324 365 325 395
rect 325 365 355 395
rect 355 365 356 395
rect 324 364 356 365
rect 324 284 356 316
rect 324 235 356 236
rect 324 205 325 235
rect 325 205 355 235
rect 355 205 356 235
rect 324 204 356 205
rect 324 124 356 156
rect 324 75 356 76
rect 324 45 325 75
rect 325 45 355 75
rect 355 45 356 75
rect 324 44 356 45
rect 324 -5 356 -4
rect 324 -35 325 -5
rect 325 -35 355 -5
rect 355 -35 356 -5
rect 324 -36 356 -35
rect 324 -85 356 -84
rect 324 -115 325 -85
rect 325 -115 355 -85
rect 355 -115 356 -85
rect 324 -116 356 -115
rect 404 1035 436 1036
rect 404 1005 405 1035
rect 405 1005 435 1035
rect 435 1005 436 1035
rect 404 1004 436 1005
rect 404 955 436 956
rect 404 925 405 955
rect 405 925 435 955
rect 435 925 436 955
rect 404 924 436 925
rect 404 875 436 876
rect 404 845 405 875
rect 405 845 435 875
rect 435 845 436 875
rect 404 844 436 845
rect 404 764 436 796
rect 404 684 436 716
rect 404 635 436 636
rect 404 605 405 635
rect 405 605 435 635
rect 435 605 436 635
rect 404 604 436 605
rect 404 555 436 556
rect 404 525 405 555
rect 405 525 435 555
rect 435 525 436 555
rect 404 524 436 525
rect 404 444 436 476
rect 404 395 436 396
rect 404 365 405 395
rect 405 365 435 395
rect 435 365 436 395
rect 404 364 436 365
rect 404 284 436 316
rect 404 235 436 236
rect 404 205 405 235
rect 405 205 435 235
rect 435 205 436 235
rect 404 204 436 205
rect 404 124 436 156
rect 404 75 436 76
rect 404 45 405 75
rect 405 45 435 75
rect 435 45 436 75
rect 404 44 436 45
rect 404 -5 436 -4
rect 404 -35 405 -5
rect 405 -35 435 -5
rect 435 -35 436 -5
rect 404 -36 436 -35
rect 404 -85 436 -84
rect 404 -115 405 -85
rect 405 -115 435 -85
rect 435 -115 436 -85
rect 404 -116 436 -115
rect 484 1035 516 1036
rect 484 1005 485 1035
rect 485 1005 515 1035
rect 515 1005 516 1035
rect 484 1004 516 1005
rect 484 955 516 956
rect 484 925 485 955
rect 485 925 515 955
rect 515 925 516 955
rect 484 924 516 925
rect 484 875 516 876
rect 484 845 485 875
rect 485 845 515 875
rect 515 845 516 875
rect 484 844 516 845
rect 484 764 516 796
rect 484 684 516 716
rect 484 635 516 636
rect 484 605 485 635
rect 485 605 515 635
rect 515 605 516 635
rect 484 604 516 605
rect 484 555 516 556
rect 484 525 485 555
rect 485 525 515 555
rect 515 525 516 555
rect 484 524 516 525
rect 484 444 516 476
rect 484 395 516 396
rect 484 365 485 395
rect 485 365 515 395
rect 515 365 516 395
rect 484 364 516 365
rect 484 284 516 316
rect 484 235 516 236
rect 484 205 485 235
rect 485 205 515 235
rect 515 205 516 235
rect 484 204 516 205
rect 484 124 516 156
rect 484 75 516 76
rect 484 45 485 75
rect 485 45 515 75
rect 515 45 516 75
rect 484 44 516 45
rect 484 -5 516 -4
rect 484 -35 485 -5
rect 485 -35 515 -5
rect 515 -35 516 -5
rect 484 -36 516 -35
rect 484 -85 516 -84
rect 484 -115 485 -85
rect 485 -115 515 -85
rect 515 -115 516 -85
rect 484 -116 516 -115
rect 564 1035 596 1036
rect 564 1005 565 1035
rect 565 1005 595 1035
rect 595 1005 596 1035
rect 564 1004 596 1005
rect 564 955 596 956
rect 564 925 565 955
rect 565 925 595 955
rect 595 925 596 955
rect 564 924 596 925
rect 564 875 596 876
rect 564 845 565 875
rect 565 845 595 875
rect 595 845 596 875
rect 564 844 596 845
rect 564 764 596 796
rect 564 684 596 716
rect 564 635 596 636
rect 564 605 565 635
rect 565 605 595 635
rect 595 605 596 635
rect 564 604 596 605
rect 564 555 596 556
rect 564 525 565 555
rect 565 525 595 555
rect 595 525 596 555
rect 564 524 596 525
rect 564 444 596 476
rect 564 395 596 396
rect 564 365 565 395
rect 565 365 595 395
rect 595 365 596 395
rect 564 364 596 365
rect 564 284 596 316
rect 564 235 596 236
rect 564 205 565 235
rect 565 205 595 235
rect 595 205 596 235
rect 564 204 596 205
rect 564 124 596 156
rect 564 75 596 76
rect 564 45 565 75
rect 565 45 595 75
rect 595 45 596 75
rect 564 44 596 45
rect 564 -5 596 -4
rect 564 -35 565 -5
rect 565 -35 595 -5
rect 595 -35 596 -5
rect 564 -36 596 -35
rect 564 -85 596 -84
rect 564 -115 565 -85
rect 565 -115 595 -85
rect 595 -115 596 -85
rect 564 -116 596 -115
rect 644 1035 676 1036
rect 644 1005 645 1035
rect 645 1005 675 1035
rect 675 1005 676 1035
rect 644 1004 676 1005
rect 644 955 676 956
rect 644 925 645 955
rect 645 925 675 955
rect 675 925 676 955
rect 644 924 676 925
rect 644 875 676 876
rect 644 845 645 875
rect 645 845 675 875
rect 675 845 676 875
rect 644 844 676 845
rect 644 764 676 796
rect 644 684 676 716
rect 644 635 676 636
rect 644 605 645 635
rect 645 605 675 635
rect 675 605 676 635
rect 644 604 676 605
rect 644 555 676 556
rect 644 525 645 555
rect 645 525 675 555
rect 675 525 676 555
rect 644 524 676 525
rect 644 444 676 476
rect 644 395 676 396
rect 644 365 645 395
rect 645 365 675 395
rect 675 365 676 395
rect 644 364 676 365
rect 644 284 676 316
rect 644 235 676 236
rect 644 205 645 235
rect 645 205 675 235
rect 675 205 676 235
rect 644 204 676 205
rect 644 124 676 156
rect 644 75 676 76
rect 644 45 645 75
rect 645 45 675 75
rect 675 45 676 75
rect 644 44 676 45
rect 644 -5 676 -4
rect 644 -35 645 -5
rect 645 -35 675 -5
rect 675 -35 676 -5
rect 644 -36 676 -35
rect 644 -85 676 -84
rect 644 -115 645 -85
rect 645 -115 675 -85
rect 675 -115 676 -85
rect 644 -116 676 -115
rect 724 1035 756 1036
rect 724 1005 725 1035
rect 725 1005 755 1035
rect 755 1005 756 1035
rect 724 1004 756 1005
rect 724 955 756 956
rect 724 925 725 955
rect 725 925 755 955
rect 755 925 756 955
rect 724 924 756 925
rect 724 875 756 876
rect 724 845 725 875
rect 725 845 755 875
rect 755 845 756 875
rect 724 844 756 845
rect 724 764 756 796
rect 724 684 756 716
rect 724 635 756 636
rect 724 605 725 635
rect 725 605 755 635
rect 755 605 756 635
rect 724 604 756 605
rect 724 555 756 556
rect 724 525 725 555
rect 725 525 755 555
rect 755 525 756 555
rect 724 524 756 525
rect 724 444 756 476
rect 724 395 756 396
rect 724 365 725 395
rect 725 365 755 395
rect 755 365 756 395
rect 724 364 756 365
rect 724 284 756 316
rect 724 235 756 236
rect 724 205 725 235
rect 725 205 755 235
rect 755 205 756 235
rect 724 204 756 205
rect 724 124 756 156
rect 724 75 756 76
rect 724 45 725 75
rect 725 45 755 75
rect 755 45 756 75
rect 724 44 756 45
rect 724 -5 756 -4
rect 724 -35 725 -5
rect 725 -35 755 -5
rect 755 -35 756 -5
rect 724 -36 756 -35
rect 724 -85 756 -84
rect 724 -115 725 -85
rect 725 -115 755 -85
rect 755 -115 756 -85
rect 724 -116 756 -115
rect 804 1035 836 1036
rect 804 1005 805 1035
rect 805 1005 835 1035
rect 835 1005 836 1035
rect 804 1004 836 1005
rect 804 955 836 956
rect 804 925 805 955
rect 805 925 835 955
rect 835 925 836 955
rect 804 924 836 925
rect 804 875 836 876
rect 804 845 805 875
rect 805 845 835 875
rect 835 845 836 875
rect 804 844 836 845
rect 804 764 836 796
rect 804 684 836 716
rect 804 635 836 636
rect 804 605 805 635
rect 805 605 835 635
rect 835 605 836 635
rect 804 604 836 605
rect 804 555 836 556
rect 804 525 805 555
rect 805 525 835 555
rect 835 525 836 555
rect 804 524 836 525
rect 804 444 836 476
rect 804 395 836 396
rect 804 365 805 395
rect 805 365 835 395
rect 835 365 836 395
rect 804 364 836 365
rect 804 284 836 316
rect 804 235 836 236
rect 804 205 805 235
rect 805 205 835 235
rect 835 205 836 235
rect 804 204 836 205
rect 804 124 836 156
rect 804 75 836 76
rect 804 45 805 75
rect 805 45 835 75
rect 835 45 836 75
rect 804 44 836 45
rect 804 -5 836 -4
rect 804 -35 805 -5
rect 805 -35 835 -5
rect 835 -35 836 -5
rect 804 -36 836 -35
rect 804 -85 836 -84
rect 804 -115 805 -85
rect 805 -115 835 -85
rect 835 -115 836 -85
rect 804 -116 836 -115
rect 884 1035 916 1036
rect 884 1005 885 1035
rect 885 1005 915 1035
rect 915 1005 916 1035
rect 884 1004 916 1005
rect 884 955 916 956
rect 884 925 885 955
rect 885 925 915 955
rect 915 925 916 955
rect 884 924 916 925
rect 884 875 916 876
rect 884 845 885 875
rect 885 845 915 875
rect 915 845 916 875
rect 884 844 916 845
rect 884 764 916 796
rect 884 684 916 716
rect 884 635 916 636
rect 884 605 885 635
rect 885 605 915 635
rect 915 605 916 635
rect 884 604 916 605
rect 884 555 916 556
rect 884 525 885 555
rect 885 525 915 555
rect 915 525 916 555
rect 884 524 916 525
rect 884 444 916 476
rect 884 395 916 396
rect 884 365 885 395
rect 885 365 915 395
rect 915 365 916 395
rect 884 364 916 365
rect 884 284 916 316
rect 884 235 916 236
rect 884 205 885 235
rect 885 205 915 235
rect 915 205 916 235
rect 884 204 916 205
rect 884 124 916 156
rect 884 75 916 76
rect 884 45 885 75
rect 885 45 915 75
rect 915 45 916 75
rect 884 44 916 45
rect 884 -5 916 -4
rect 884 -35 885 -5
rect 885 -35 915 -5
rect 915 -35 916 -5
rect 884 -36 916 -35
rect 884 -85 916 -84
rect 884 -115 885 -85
rect 885 -115 915 -85
rect 915 -115 916 -85
rect 884 -116 916 -115
rect 964 1035 996 1036
rect 964 1005 965 1035
rect 965 1005 995 1035
rect 995 1005 996 1035
rect 964 1004 996 1005
rect 964 955 996 956
rect 964 925 965 955
rect 965 925 995 955
rect 995 925 996 955
rect 964 924 996 925
rect 964 875 996 876
rect 964 845 965 875
rect 965 845 995 875
rect 995 845 996 875
rect 964 844 996 845
rect 964 764 996 796
rect 964 684 996 716
rect 964 635 996 636
rect 964 605 965 635
rect 965 605 995 635
rect 995 605 996 635
rect 964 604 996 605
rect 964 555 996 556
rect 964 525 965 555
rect 965 525 995 555
rect 995 525 996 555
rect 964 524 996 525
rect 964 444 996 476
rect 964 395 996 396
rect 964 365 965 395
rect 965 365 995 395
rect 995 365 996 395
rect 964 364 996 365
rect 964 284 996 316
rect 964 235 996 236
rect 964 205 965 235
rect 965 205 995 235
rect 995 205 996 235
rect 964 204 996 205
rect 964 124 996 156
rect 964 75 996 76
rect 964 45 965 75
rect 965 45 995 75
rect 995 45 996 75
rect 964 44 996 45
rect 964 -5 996 -4
rect 964 -35 965 -5
rect 965 -35 995 -5
rect 995 -35 996 -5
rect 964 -36 996 -35
rect 964 -85 996 -84
rect 964 -115 965 -85
rect 965 -115 995 -85
rect 995 -115 996 -85
rect 964 -116 996 -115
rect 1044 1035 1076 1036
rect 1044 1005 1045 1035
rect 1045 1005 1075 1035
rect 1075 1005 1076 1035
rect 1044 1004 1076 1005
rect 1044 955 1076 956
rect 1044 925 1045 955
rect 1045 925 1075 955
rect 1075 925 1076 955
rect 1044 924 1076 925
rect 1044 875 1076 876
rect 1044 845 1045 875
rect 1045 845 1075 875
rect 1075 845 1076 875
rect 1044 844 1076 845
rect 1044 764 1076 796
rect 1044 684 1076 716
rect 1044 635 1076 636
rect 1044 605 1045 635
rect 1045 605 1075 635
rect 1075 605 1076 635
rect 1044 604 1076 605
rect 1044 555 1076 556
rect 1044 525 1045 555
rect 1045 525 1075 555
rect 1075 525 1076 555
rect 1044 524 1076 525
rect 1044 444 1076 476
rect 1044 395 1076 396
rect 1044 365 1045 395
rect 1045 365 1075 395
rect 1075 365 1076 395
rect 1044 364 1076 365
rect 1044 284 1076 316
rect 1044 235 1076 236
rect 1044 205 1045 235
rect 1045 205 1075 235
rect 1075 205 1076 235
rect 1044 204 1076 205
rect 1044 124 1076 156
rect 1044 75 1076 76
rect 1044 45 1045 75
rect 1045 45 1075 75
rect 1075 45 1076 75
rect 1044 44 1076 45
rect 1044 -5 1076 -4
rect 1044 -35 1045 -5
rect 1045 -35 1075 -5
rect 1075 -35 1076 -5
rect 1044 -36 1076 -35
rect 1044 -85 1076 -84
rect 1044 -115 1045 -85
rect 1045 -115 1075 -85
rect 1075 -115 1076 -85
rect 1044 -116 1076 -115
rect 1124 1035 1156 1036
rect 1124 1005 1125 1035
rect 1125 1005 1155 1035
rect 1155 1005 1156 1035
rect 1124 1004 1156 1005
rect 1124 955 1156 956
rect 1124 925 1125 955
rect 1125 925 1155 955
rect 1155 925 1156 955
rect 1124 924 1156 925
rect 1124 875 1156 876
rect 1124 845 1125 875
rect 1125 845 1155 875
rect 1155 845 1156 875
rect 1124 844 1156 845
rect 1124 764 1156 796
rect 1124 684 1156 716
rect 1124 635 1156 636
rect 1124 605 1125 635
rect 1125 605 1155 635
rect 1155 605 1156 635
rect 1124 604 1156 605
rect 1124 555 1156 556
rect 1124 525 1125 555
rect 1125 525 1155 555
rect 1155 525 1156 555
rect 1124 524 1156 525
rect 1124 444 1156 476
rect 1124 395 1156 396
rect 1124 365 1125 395
rect 1125 365 1155 395
rect 1155 365 1156 395
rect 1124 364 1156 365
rect 1124 284 1156 316
rect 1124 235 1156 236
rect 1124 205 1125 235
rect 1125 205 1155 235
rect 1155 205 1156 235
rect 1124 204 1156 205
rect 1124 124 1156 156
rect 1124 75 1156 76
rect 1124 45 1125 75
rect 1125 45 1155 75
rect 1155 45 1156 75
rect 1124 44 1156 45
rect 1124 -5 1156 -4
rect 1124 -35 1125 -5
rect 1125 -35 1155 -5
rect 1155 -35 1156 -5
rect 1124 -36 1156 -35
rect 1124 -85 1156 -84
rect 1124 -115 1125 -85
rect 1125 -115 1155 -85
rect 1155 -115 1156 -85
rect 1124 -116 1156 -115
rect 1204 1035 1236 1036
rect 1204 1005 1205 1035
rect 1205 1005 1235 1035
rect 1235 1005 1236 1035
rect 1204 1004 1236 1005
rect 1204 955 1236 956
rect 1204 925 1205 955
rect 1205 925 1235 955
rect 1235 925 1236 955
rect 1204 924 1236 925
rect 1204 875 1236 876
rect 1204 845 1205 875
rect 1205 845 1235 875
rect 1235 845 1236 875
rect 1204 844 1236 845
rect 1204 764 1236 796
rect 1204 684 1236 716
rect 1204 635 1236 636
rect 1204 605 1205 635
rect 1205 605 1235 635
rect 1235 605 1236 635
rect 1204 604 1236 605
rect 1204 555 1236 556
rect 1204 525 1205 555
rect 1205 525 1235 555
rect 1235 525 1236 555
rect 1204 524 1236 525
rect 1204 444 1236 476
rect 1204 395 1236 396
rect 1204 365 1205 395
rect 1205 365 1235 395
rect 1235 365 1236 395
rect 1204 364 1236 365
rect 1204 284 1236 316
rect 1204 235 1236 236
rect 1204 205 1205 235
rect 1205 205 1235 235
rect 1235 205 1236 235
rect 1204 204 1236 205
rect 1204 124 1236 156
rect 1204 75 1236 76
rect 1204 45 1205 75
rect 1205 45 1235 75
rect 1235 45 1236 75
rect 1204 44 1236 45
rect 1204 -5 1236 -4
rect 1204 -35 1205 -5
rect 1205 -35 1235 -5
rect 1235 -35 1236 -5
rect 1204 -36 1236 -35
rect 1204 -85 1236 -84
rect 1204 -115 1205 -85
rect 1205 -115 1235 -85
rect 1235 -115 1236 -85
rect 1204 -116 1236 -115
rect 1284 1035 1316 1036
rect 1284 1005 1285 1035
rect 1285 1005 1315 1035
rect 1315 1005 1316 1035
rect 1284 1004 1316 1005
rect 1284 955 1316 956
rect 1284 925 1285 955
rect 1285 925 1315 955
rect 1315 925 1316 955
rect 1284 924 1316 925
rect 1284 875 1316 876
rect 1284 845 1285 875
rect 1285 845 1315 875
rect 1315 845 1316 875
rect 1284 844 1316 845
rect 1284 764 1316 796
rect 1284 684 1316 716
rect 1284 635 1316 636
rect 1284 605 1285 635
rect 1285 605 1315 635
rect 1315 605 1316 635
rect 1284 604 1316 605
rect 1284 555 1316 556
rect 1284 525 1285 555
rect 1285 525 1315 555
rect 1315 525 1316 555
rect 1284 524 1316 525
rect 1284 444 1316 476
rect 1284 395 1316 396
rect 1284 365 1285 395
rect 1285 365 1315 395
rect 1315 365 1316 395
rect 1284 364 1316 365
rect 1284 284 1316 316
rect 1284 235 1316 236
rect 1284 205 1285 235
rect 1285 205 1315 235
rect 1315 205 1316 235
rect 1284 204 1316 205
rect 1284 124 1316 156
rect 1284 75 1316 76
rect 1284 45 1285 75
rect 1285 45 1315 75
rect 1315 45 1316 75
rect 1284 44 1316 45
rect 1284 -5 1316 -4
rect 1284 -35 1285 -5
rect 1285 -35 1315 -5
rect 1315 -35 1316 -5
rect 1284 -36 1316 -35
rect 1284 -85 1316 -84
rect 1284 -115 1285 -85
rect 1285 -115 1315 -85
rect 1315 -115 1316 -85
rect 1284 -116 1316 -115
rect 1364 1035 1396 1036
rect 1364 1005 1365 1035
rect 1365 1005 1395 1035
rect 1395 1005 1396 1035
rect 1364 1004 1396 1005
rect 1364 955 1396 956
rect 1364 925 1365 955
rect 1365 925 1395 955
rect 1395 925 1396 955
rect 1364 924 1396 925
rect 1364 875 1396 876
rect 1364 845 1365 875
rect 1365 845 1395 875
rect 1395 845 1396 875
rect 1364 844 1396 845
rect 1364 764 1396 796
rect 1364 684 1396 716
rect 1364 635 1396 636
rect 1364 605 1365 635
rect 1365 605 1395 635
rect 1395 605 1396 635
rect 1364 604 1396 605
rect 1364 555 1396 556
rect 1364 525 1365 555
rect 1365 525 1395 555
rect 1395 525 1396 555
rect 1364 524 1396 525
rect 1364 444 1396 476
rect 1364 395 1396 396
rect 1364 365 1365 395
rect 1365 365 1395 395
rect 1395 365 1396 395
rect 1364 364 1396 365
rect 1364 284 1396 316
rect 1364 235 1396 236
rect 1364 205 1365 235
rect 1365 205 1395 235
rect 1395 205 1396 235
rect 1364 204 1396 205
rect 1364 124 1396 156
rect 1364 75 1396 76
rect 1364 45 1365 75
rect 1365 45 1395 75
rect 1395 45 1396 75
rect 1364 44 1396 45
rect 1364 -5 1396 -4
rect 1364 -35 1365 -5
rect 1365 -35 1395 -5
rect 1395 -35 1396 -5
rect 1364 -36 1396 -35
rect 1364 -85 1396 -84
rect 1364 -115 1365 -85
rect 1365 -115 1395 -85
rect 1395 -115 1396 -85
rect 1364 -116 1396 -115
rect 1444 1035 1476 1036
rect 1444 1005 1445 1035
rect 1445 1005 1475 1035
rect 1475 1005 1476 1035
rect 1444 1004 1476 1005
rect 1444 955 1476 956
rect 1444 925 1445 955
rect 1445 925 1475 955
rect 1475 925 1476 955
rect 1444 924 1476 925
rect 1444 875 1476 876
rect 1444 845 1445 875
rect 1445 845 1475 875
rect 1475 845 1476 875
rect 1444 844 1476 845
rect 1444 764 1476 796
rect 1444 684 1476 716
rect 1444 635 1476 636
rect 1444 605 1445 635
rect 1445 605 1475 635
rect 1475 605 1476 635
rect 1444 604 1476 605
rect 1444 555 1476 556
rect 1444 525 1445 555
rect 1445 525 1475 555
rect 1475 525 1476 555
rect 1444 524 1476 525
rect 1444 444 1476 476
rect 1444 395 1476 396
rect 1444 365 1445 395
rect 1445 365 1475 395
rect 1475 365 1476 395
rect 1444 364 1476 365
rect 1444 284 1476 316
rect 1444 235 1476 236
rect 1444 205 1445 235
rect 1445 205 1475 235
rect 1475 205 1476 235
rect 1444 204 1476 205
rect 1444 124 1476 156
rect 1444 75 1476 76
rect 1444 45 1445 75
rect 1445 45 1475 75
rect 1475 45 1476 75
rect 1444 44 1476 45
rect 1444 -5 1476 -4
rect 1444 -35 1445 -5
rect 1445 -35 1475 -5
rect 1475 -35 1476 -5
rect 1444 -36 1476 -35
rect 1444 -85 1476 -84
rect 1444 -115 1445 -85
rect 1445 -115 1475 -85
rect 1475 -115 1476 -85
rect 1444 -116 1476 -115
rect 1524 1035 1556 1036
rect 1524 1005 1525 1035
rect 1525 1005 1555 1035
rect 1555 1005 1556 1035
rect 1524 1004 1556 1005
rect 1524 955 1556 956
rect 1524 925 1525 955
rect 1525 925 1555 955
rect 1555 925 1556 955
rect 1524 924 1556 925
rect 1524 875 1556 876
rect 1524 845 1525 875
rect 1525 845 1555 875
rect 1555 845 1556 875
rect 1524 844 1556 845
rect 1524 764 1556 796
rect 1524 684 1556 716
rect 1524 635 1556 636
rect 1524 605 1525 635
rect 1525 605 1555 635
rect 1555 605 1556 635
rect 1524 604 1556 605
rect 1524 555 1556 556
rect 1524 525 1525 555
rect 1525 525 1555 555
rect 1555 525 1556 555
rect 1524 524 1556 525
rect 1524 444 1556 476
rect 1524 395 1556 396
rect 1524 365 1525 395
rect 1525 365 1555 395
rect 1555 365 1556 395
rect 1524 364 1556 365
rect 1524 284 1556 316
rect 1524 235 1556 236
rect 1524 205 1525 235
rect 1525 205 1555 235
rect 1555 205 1556 235
rect 1524 204 1556 205
rect 1524 124 1556 156
rect 1524 75 1556 76
rect 1524 45 1525 75
rect 1525 45 1555 75
rect 1555 45 1556 75
rect 1524 44 1556 45
rect 1524 -5 1556 -4
rect 1524 -35 1525 -5
rect 1525 -35 1555 -5
rect 1555 -35 1556 -5
rect 1524 -36 1556 -35
rect 1524 -85 1556 -84
rect 1524 -115 1525 -85
rect 1525 -115 1555 -85
rect 1555 -115 1556 -85
rect 1524 -116 1556 -115
rect 1604 1035 1636 1036
rect 1604 1005 1605 1035
rect 1605 1005 1635 1035
rect 1635 1005 1636 1035
rect 1604 1004 1636 1005
rect 1604 955 1636 956
rect 1604 925 1605 955
rect 1605 925 1635 955
rect 1635 925 1636 955
rect 1604 924 1636 925
rect 1604 875 1636 876
rect 1604 845 1605 875
rect 1605 845 1635 875
rect 1635 845 1636 875
rect 1604 844 1636 845
rect 1604 764 1636 796
rect 1604 684 1636 716
rect 1604 635 1636 636
rect 1604 605 1605 635
rect 1605 605 1635 635
rect 1635 605 1636 635
rect 1604 604 1636 605
rect 1604 555 1636 556
rect 1604 525 1605 555
rect 1605 525 1635 555
rect 1635 525 1636 555
rect 1604 524 1636 525
rect 1604 444 1636 476
rect 1604 395 1636 396
rect 1604 365 1605 395
rect 1605 365 1635 395
rect 1635 365 1636 395
rect 1604 364 1636 365
rect 1604 284 1636 316
rect 1604 235 1636 236
rect 1604 205 1605 235
rect 1605 205 1635 235
rect 1635 205 1636 235
rect 1604 204 1636 205
rect 1604 124 1636 156
rect 1604 75 1636 76
rect 1604 45 1605 75
rect 1605 45 1635 75
rect 1635 45 1636 75
rect 1604 44 1636 45
rect 1604 -5 1636 -4
rect 1604 -35 1605 -5
rect 1605 -35 1635 -5
rect 1635 -35 1636 -5
rect 1604 -36 1636 -35
rect 1604 -85 1636 -84
rect 1604 -115 1605 -85
rect 1605 -115 1635 -85
rect 1635 -115 1636 -85
rect 1604 -116 1636 -115
rect 1684 1035 1716 1036
rect 1684 1005 1685 1035
rect 1685 1005 1715 1035
rect 1715 1005 1716 1035
rect 1684 1004 1716 1005
rect 1684 955 1716 956
rect 1684 925 1685 955
rect 1685 925 1715 955
rect 1715 925 1716 955
rect 1684 924 1716 925
rect 1684 875 1716 876
rect 1684 845 1685 875
rect 1685 845 1715 875
rect 1715 845 1716 875
rect 1684 844 1716 845
rect 1684 764 1716 796
rect 1684 684 1716 716
rect 1684 635 1716 636
rect 1684 605 1685 635
rect 1685 605 1715 635
rect 1715 605 1716 635
rect 1684 604 1716 605
rect 1684 555 1716 556
rect 1684 525 1685 555
rect 1685 525 1715 555
rect 1715 525 1716 555
rect 1684 524 1716 525
rect 1684 444 1716 476
rect 1684 395 1716 396
rect 1684 365 1685 395
rect 1685 365 1715 395
rect 1715 365 1716 395
rect 1684 364 1716 365
rect 1684 284 1716 316
rect 1684 235 1716 236
rect 1684 205 1685 235
rect 1685 205 1715 235
rect 1715 205 1716 235
rect 1684 204 1716 205
rect 1684 124 1716 156
rect 1684 75 1716 76
rect 1684 45 1685 75
rect 1685 45 1715 75
rect 1715 45 1716 75
rect 1684 44 1716 45
rect 1684 -5 1716 -4
rect 1684 -35 1685 -5
rect 1685 -35 1715 -5
rect 1715 -35 1716 -5
rect 1684 -36 1716 -35
rect 1684 -85 1716 -84
rect 1684 -115 1685 -85
rect 1685 -115 1715 -85
rect 1715 -115 1716 -85
rect 1684 -116 1716 -115
rect 1764 1035 1796 1036
rect 1764 1005 1765 1035
rect 1765 1005 1795 1035
rect 1795 1005 1796 1035
rect 1764 1004 1796 1005
rect 1764 955 1796 956
rect 1764 925 1765 955
rect 1765 925 1795 955
rect 1795 925 1796 955
rect 1764 924 1796 925
rect 1764 875 1796 876
rect 1764 845 1765 875
rect 1765 845 1795 875
rect 1795 845 1796 875
rect 1764 844 1796 845
rect 1764 764 1796 796
rect 1764 684 1796 716
rect 1764 635 1796 636
rect 1764 605 1765 635
rect 1765 605 1795 635
rect 1795 605 1796 635
rect 1764 604 1796 605
rect 1764 555 1796 556
rect 1764 525 1765 555
rect 1765 525 1795 555
rect 1795 525 1796 555
rect 1764 524 1796 525
rect 1764 444 1796 476
rect 1764 395 1796 396
rect 1764 365 1765 395
rect 1765 365 1795 395
rect 1795 365 1796 395
rect 1764 364 1796 365
rect 1764 284 1796 316
rect 1764 235 1796 236
rect 1764 205 1765 235
rect 1765 205 1795 235
rect 1795 205 1796 235
rect 1764 204 1796 205
rect 1764 124 1796 156
rect 1764 75 1796 76
rect 1764 45 1765 75
rect 1765 45 1795 75
rect 1795 45 1796 75
rect 1764 44 1796 45
rect 1764 -5 1796 -4
rect 1764 -35 1765 -5
rect 1765 -35 1795 -5
rect 1795 -35 1796 -5
rect 1764 -36 1796 -35
rect 1764 -85 1796 -84
rect 1764 -115 1765 -85
rect 1765 -115 1795 -85
rect 1795 -115 1796 -85
rect 1764 -116 1796 -115
rect 1844 1035 1876 1036
rect 1844 1005 1845 1035
rect 1845 1005 1875 1035
rect 1875 1005 1876 1035
rect 1844 1004 1876 1005
rect 1844 955 1876 956
rect 1844 925 1845 955
rect 1845 925 1875 955
rect 1875 925 1876 955
rect 1844 924 1876 925
rect 1844 875 1876 876
rect 1844 845 1845 875
rect 1845 845 1875 875
rect 1875 845 1876 875
rect 1844 844 1876 845
rect 1844 764 1876 796
rect 1844 684 1876 716
rect 1844 635 1876 636
rect 1844 605 1845 635
rect 1845 605 1875 635
rect 1875 605 1876 635
rect 1844 604 1876 605
rect 1844 555 1876 556
rect 1844 525 1845 555
rect 1845 525 1875 555
rect 1875 525 1876 555
rect 1844 524 1876 525
rect 1844 444 1876 476
rect 1844 395 1876 396
rect 1844 365 1845 395
rect 1845 365 1875 395
rect 1875 365 1876 395
rect 1844 364 1876 365
rect 1844 284 1876 316
rect 1844 235 1876 236
rect 1844 205 1845 235
rect 1845 205 1875 235
rect 1875 205 1876 235
rect 1844 204 1876 205
rect 1844 124 1876 156
rect 1844 75 1876 76
rect 1844 45 1845 75
rect 1845 45 1875 75
rect 1875 45 1876 75
rect 1844 44 1876 45
rect 1844 -5 1876 -4
rect 1844 -35 1845 -5
rect 1845 -35 1875 -5
rect 1875 -35 1876 -5
rect 1844 -36 1876 -35
rect 1844 -85 1876 -84
rect 1844 -115 1845 -85
rect 1845 -115 1875 -85
rect 1875 -115 1876 -85
rect 1844 -116 1876 -115
rect 1924 1035 1956 1036
rect 1924 1005 1925 1035
rect 1925 1005 1955 1035
rect 1955 1005 1956 1035
rect 1924 1004 1956 1005
rect 1924 955 1956 956
rect 1924 925 1925 955
rect 1925 925 1955 955
rect 1955 925 1956 955
rect 1924 924 1956 925
rect 1924 875 1956 876
rect 1924 845 1925 875
rect 1925 845 1955 875
rect 1955 845 1956 875
rect 1924 844 1956 845
rect 1924 764 1956 796
rect 1924 684 1956 716
rect 1924 635 1956 636
rect 1924 605 1925 635
rect 1925 605 1955 635
rect 1955 605 1956 635
rect 1924 604 1956 605
rect 1924 555 1956 556
rect 1924 525 1925 555
rect 1925 525 1955 555
rect 1955 525 1956 555
rect 1924 524 1956 525
rect 1924 444 1956 476
rect 1924 395 1956 396
rect 1924 365 1925 395
rect 1925 365 1955 395
rect 1955 365 1956 395
rect 1924 364 1956 365
rect 1924 284 1956 316
rect 1924 235 1956 236
rect 1924 205 1925 235
rect 1925 205 1955 235
rect 1955 205 1956 235
rect 1924 204 1956 205
rect 1924 124 1956 156
rect 1924 75 1956 76
rect 1924 45 1925 75
rect 1925 45 1955 75
rect 1955 45 1956 75
rect 1924 44 1956 45
rect 1924 -5 1956 -4
rect 1924 -35 1925 -5
rect 1925 -35 1955 -5
rect 1955 -35 1956 -5
rect 1924 -36 1956 -35
rect 1924 -85 1956 -84
rect 1924 -115 1925 -85
rect 1925 -115 1955 -85
rect 1955 -115 1956 -85
rect 1924 -116 1956 -115
rect 2004 1035 2036 1036
rect 2004 1005 2005 1035
rect 2005 1005 2035 1035
rect 2035 1005 2036 1035
rect 2004 1004 2036 1005
rect 2004 955 2036 956
rect 2004 925 2005 955
rect 2005 925 2035 955
rect 2035 925 2036 955
rect 2004 924 2036 925
rect 2004 875 2036 876
rect 2004 845 2005 875
rect 2005 845 2035 875
rect 2035 845 2036 875
rect 2004 844 2036 845
rect 2004 764 2036 796
rect 2004 684 2036 716
rect 2004 635 2036 636
rect 2004 605 2005 635
rect 2005 605 2035 635
rect 2035 605 2036 635
rect 2004 604 2036 605
rect 2004 555 2036 556
rect 2004 525 2005 555
rect 2005 525 2035 555
rect 2035 525 2036 555
rect 2004 524 2036 525
rect 2004 444 2036 476
rect 2004 395 2036 396
rect 2004 365 2005 395
rect 2005 365 2035 395
rect 2035 365 2036 395
rect 2004 364 2036 365
rect 2004 284 2036 316
rect 2004 235 2036 236
rect 2004 205 2005 235
rect 2005 205 2035 235
rect 2035 205 2036 235
rect 2004 204 2036 205
rect 2004 124 2036 156
rect 2004 75 2036 76
rect 2004 45 2005 75
rect 2005 45 2035 75
rect 2035 45 2036 75
rect 2004 44 2036 45
rect 2004 -5 2036 -4
rect 2004 -35 2005 -5
rect 2005 -35 2035 -5
rect 2035 -35 2036 -5
rect 2004 -36 2036 -35
rect 2004 -85 2036 -84
rect 2004 -115 2005 -85
rect 2005 -115 2035 -85
rect 2035 -115 2036 -85
rect 2004 -116 2036 -115
rect 2084 1035 2116 1036
rect 2084 1005 2085 1035
rect 2085 1005 2115 1035
rect 2115 1005 2116 1035
rect 2084 1004 2116 1005
rect 2084 955 2116 956
rect 2084 925 2085 955
rect 2085 925 2115 955
rect 2115 925 2116 955
rect 2084 924 2116 925
rect 2084 875 2116 876
rect 2084 845 2085 875
rect 2085 845 2115 875
rect 2115 845 2116 875
rect 2084 844 2116 845
rect 2084 764 2116 796
rect 2084 684 2116 716
rect 2084 635 2116 636
rect 2084 605 2085 635
rect 2085 605 2115 635
rect 2115 605 2116 635
rect 2084 604 2116 605
rect 2084 555 2116 556
rect 2084 525 2085 555
rect 2085 525 2115 555
rect 2115 525 2116 555
rect 2084 524 2116 525
rect 2084 444 2116 476
rect 2084 395 2116 396
rect 2084 365 2085 395
rect 2085 365 2115 395
rect 2115 365 2116 395
rect 2084 364 2116 365
rect 2084 284 2116 316
rect 2084 235 2116 236
rect 2084 205 2085 235
rect 2085 205 2115 235
rect 2115 205 2116 235
rect 2084 204 2116 205
rect 2084 124 2116 156
rect 2084 75 2116 76
rect 2084 45 2085 75
rect 2085 45 2115 75
rect 2115 45 2116 75
rect 2084 44 2116 45
rect 2084 -5 2116 -4
rect 2084 -35 2085 -5
rect 2085 -35 2115 -5
rect 2115 -35 2116 -5
rect 2084 -36 2116 -35
rect 2084 -85 2116 -84
rect 2084 -115 2085 -85
rect 2085 -115 2115 -85
rect 2115 -115 2116 -85
rect 2084 -116 2116 -115
rect 2164 1035 2196 1036
rect 2164 1005 2165 1035
rect 2165 1005 2195 1035
rect 2195 1005 2196 1035
rect 2164 1004 2196 1005
rect 2164 955 2196 956
rect 2164 925 2165 955
rect 2165 925 2195 955
rect 2195 925 2196 955
rect 2164 924 2196 925
rect 2164 875 2196 876
rect 2164 845 2165 875
rect 2165 845 2195 875
rect 2195 845 2196 875
rect 2164 844 2196 845
rect 2164 764 2196 796
rect 2164 684 2196 716
rect 2164 635 2196 636
rect 2164 605 2165 635
rect 2165 605 2195 635
rect 2195 605 2196 635
rect 2164 604 2196 605
rect 2164 555 2196 556
rect 2164 525 2165 555
rect 2165 525 2195 555
rect 2195 525 2196 555
rect 2164 524 2196 525
rect 2164 444 2196 476
rect 2164 395 2196 396
rect 2164 365 2165 395
rect 2165 365 2195 395
rect 2195 365 2196 395
rect 2164 364 2196 365
rect 2164 284 2196 316
rect 2164 235 2196 236
rect 2164 205 2165 235
rect 2165 205 2195 235
rect 2195 205 2196 235
rect 2164 204 2196 205
rect 2164 124 2196 156
rect 2164 75 2196 76
rect 2164 45 2165 75
rect 2165 45 2195 75
rect 2195 45 2196 75
rect 2164 44 2196 45
rect 2164 -5 2196 -4
rect 2164 -35 2165 -5
rect 2165 -35 2195 -5
rect 2195 -35 2196 -5
rect 2164 -36 2196 -35
rect 2164 -85 2196 -84
rect 2164 -115 2165 -85
rect 2165 -115 2195 -85
rect 2195 -115 2196 -85
rect 2164 -116 2196 -115
rect 2244 1035 2276 1036
rect 2244 1005 2245 1035
rect 2245 1005 2275 1035
rect 2275 1005 2276 1035
rect 2244 1004 2276 1005
rect 2244 955 2276 956
rect 2244 925 2245 955
rect 2245 925 2275 955
rect 2275 925 2276 955
rect 2244 924 2276 925
rect 2244 875 2276 876
rect 2244 845 2245 875
rect 2245 845 2275 875
rect 2275 845 2276 875
rect 2244 844 2276 845
rect 2244 764 2276 796
rect 2244 684 2276 716
rect 2244 635 2276 636
rect 2244 605 2245 635
rect 2245 605 2275 635
rect 2275 605 2276 635
rect 2244 604 2276 605
rect 2244 555 2276 556
rect 2244 525 2245 555
rect 2245 525 2275 555
rect 2275 525 2276 555
rect 2244 524 2276 525
rect 2244 444 2276 476
rect 2244 395 2276 396
rect 2244 365 2245 395
rect 2245 365 2275 395
rect 2275 365 2276 395
rect 2244 364 2276 365
rect 2244 284 2276 316
rect 2244 235 2276 236
rect 2244 205 2245 235
rect 2245 205 2275 235
rect 2275 205 2276 235
rect 2244 204 2276 205
rect 2244 124 2276 156
rect 2244 75 2276 76
rect 2244 45 2245 75
rect 2245 45 2275 75
rect 2275 45 2276 75
rect 2244 44 2276 45
rect 2244 -5 2276 -4
rect 2244 -35 2245 -5
rect 2245 -35 2275 -5
rect 2275 -35 2276 -5
rect 2244 -36 2276 -35
rect 2244 -85 2276 -84
rect 2244 -115 2245 -85
rect 2245 -115 2275 -85
rect 2275 -115 2276 -85
rect 2244 -116 2276 -115
rect 2324 1035 2356 1036
rect 2324 1005 2325 1035
rect 2325 1005 2355 1035
rect 2355 1005 2356 1035
rect 2324 1004 2356 1005
rect 2324 955 2356 956
rect 2324 925 2325 955
rect 2325 925 2355 955
rect 2355 925 2356 955
rect 2324 924 2356 925
rect 2324 875 2356 876
rect 2324 845 2325 875
rect 2325 845 2355 875
rect 2355 845 2356 875
rect 2324 844 2356 845
rect 2324 764 2356 796
rect 2324 684 2356 716
rect 2324 635 2356 636
rect 2324 605 2325 635
rect 2325 605 2355 635
rect 2355 605 2356 635
rect 2324 604 2356 605
rect 2324 555 2356 556
rect 2324 525 2325 555
rect 2325 525 2355 555
rect 2355 525 2356 555
rect 2324 524 2356 525
rect 2324 444 2356 476
rect 2324 395 2356 396
rect 2324 365 2325 395
rect 2325 365 2355 395
rect 2355 365 2356 395
rect 2324 364 2356 365
rect 2324 284 2356 316
rect 2324 235 2356 236
rect 2324 205 2325 235
rect 2325 205 2355 235
rect 2355 205 2356 235
rect 2324 204 2356 205
rect 2324 124 2356 156
rect 2324 75 2356 76
rect 2324 45 2325 75
rect 2325 45 2355 75
rect 2355 45 2356 75
rect 2324 44 2356 45
rect 2324 -5 2356 -4
rect 2324 -35 2325 -5
rect 2325 -35 2355 -5
rect 2355 -35 2356 -5
rect 2324 -36 2356 -35
rect 2324 -85 2356 -84
rect 2324 -115 2325 -85
rect 2325 -115 2355 -85
rect 2355 -115 2356 -85
rect 2324 -116 2356 -115
rect 2404 1035 2436 1036
rect 2404 1005 2405 1035
rect 2405 1005 2435 1035
rect 2435 1005 2436 1035
rect 2404 1004 2436 1005
rect 2404 955 2436 956
rect 2404 925 2405 955
rect 2405 925 2435 955
rect 2435 925 2436 955
rect 2404 924 2436 925
rect 2404 875 2436 876
rect 2404 845 2405 875
rect 2405 845 2435 875
rect 2435 845 2436 875
rect 2404 844 2436 845
rect 2404 764 2436 796
rect 2404 684 2436 716
rect 2404 635 2436 636
rect 2404 605 2405 635
rect 2405 605 2435 635
rect 2435 605 2436 635
rect 2404 604 2436 605
rect 2404 555 2436 556
rect 2404 525 2405 555
rect 2405 525 2435 555
rect 2435 525 2436 555
rect 2404 524 2436 525
rect 2404 444 2436 476
rect 2404 395 2436 396
rect 2404 365 2405 395
rect 2405 365 2435 395
rect 2435 365 2436 395
rect 2404 364 2436 365
rect 2404 284 2436 316
rect 2404 235 2436 236
rect 2404 205 2405 235
rect 2405 205 2435 235
rect 2435 205 2436 235
rect 2404 204 2436 205
rect 2404 124 2436 156
rect 2404 75 2436 76
rect 2404 45 2405 75
rect 2405 45 2435 75
rect 2435 45 2436 75
rect 2404 44 2436 45
rect 2404 -5 2436 -4
rect 2404 -35 2405 -5
rect 2405 -35 2435 -5
rect 2435 -35 2436 -5
rect 2404 -36 2436 -35
rect 2404 -85 2436 -84
rect 2404 -115 2405 -85
rect 2405 -115 2435 -85
rect 2435 -115 2436 -85
rect 2404 -116 2436 -115
rect 2484 1035 2516 1036
rect 2484 1005 2485 1035
rect 2485 1005 2515 1035
rect 2515 1005 2516 1035
rect 2484 1004 2516 1005
rect 2484 955 2516 956
rect 2484 925 2485 955
rect 2485 925 2515 955
rect 2515 925 2516 955
rect 2484 924 2516 925
rect 2484 875 2516 876
rect 2484 845 2485 875
rect 2485 845 2515 875
rect 2515 845 2516 875
rect 2484 844 2516 845
rect 2484 764 2516 796
rect 2484 684 2516 716
rect 2484 635 2516 636
rect 2484 605 2485 635
rect 2485 605 2515 635
rect 2515 605 2516 635
rect 2484 604 2516 605
rect 2484 555 2516 556
rect 2484 525 2485 555
rect 2485 525 2515 555
rect 2515 525 2516 555
rect 2484 524 2516 525
rect 2484 444 2516 476
rect 2484 395 2516 396
rect 2484 365 2485 395
rect 2485 365 2515 395
rect 2515 365 2516 395
rect 2484 364 2516 365
rect 2484 284 2516 316
rect 2484 235 2516 236
rect 2484 205 2485 235
rect 2485 205 2515 235
rect 2515 205 2516 235
rect 2484 204 2516 205
rect 2484 124 2516 156
rect 2484 75 2516 76
rect 2484 45 2485 75
rect 2485 45 2515 75
rect 2515 45 2516 75
rect 2484 44 2516 45
rect 2484 -5 2516 -4
rect 2484 -35 2485 -5
rect 2485 -35 2515 -5
rect 2515 -35 2516 -5
rect 2484 -36 2516 -35
rect 2484 -85 2516 -84
rect 2484 -115 2485 -85
rect 2485 -115 2515 -85
rect 2515 -115 2516 -85
rect 2484 -116 2516 -115
rect 2564 1035 2596 1036
rect 2564 1005 2565 1035
rect 2565 1005 2595 1035
rect 2595 1005 2596 1035
rect 2564 1004 2596 1005
rect 2564 955 2596 956
rect 2564 925 2565 955
rect 2565 925 2595 955
rect 2595 925 2596 955
rect 2564 924 2596 925
rect 2564 875 2596 876
rect 2564 845 2565 875
rect 2565 845 2595 875
rect 2595 845 2596 875
rect 2564 844 2596 845
rect 2564 764 2596 796
rect 2564 684 2596 716
rect 2564 635 2596 636
rect 2564 605 2565 635
rect 2565 605 2595 635
rect 2595 605 2596 635
rect 2564 604 2596 605
rect 2564 555 2596 556
rect 2564 525 2565 555
rect 2565 525 2595 555
rect 2595 525 2596 555
rect 2564 524 2596 525
rect 2564 444 2596 476
rect 2564 395 2596 396
rect 2564 365 2565 395
rect 2565 365 2595 395
rect 2595 365 2596 395
rect 2564 364 2596 365
rect 2564 284 2596 316
rect 2564 235 2596 236
rect 2564 205 2565 235
rect 2565 205 2595 235
rect 2595 205 2596 235
rect 2564 204 2596 205
rect 2564 124 2596 156
rect 2564 75 2596 76
rect 2564 45 2565 75
rect 2565 45 2595 75
rect 2595 45 2596 75
rect 2564 44 2596 45
rect 2564 -5 2596 -4
rect 2564 -35 2565 -5
rect 2565 -35 2595 -5
rect 2595 -35 2596 -5
rect 2564 -36 2596 -35
rect 2564 -85 2596 -84
rect 2564 -115 2565 -85
rect 2565 -115 2595 -85
rect 2595 -115 2596 -85
rect 2564 -116 2596 -115
rect 2644 1035 2676 1036
rect 2644 1005 2645 1035
rect 2645 1005 2675 1035
rect 2675 1005 2676 1035
rect 2644 1004 2676 1005
rect 2644 955 2676 956
rect 2644 925 2645 955
rect 2645 925 2675 955
rect 2675 925 2676 955
rect 2644 924 2676 925
rect 2644 875 2676 876
rect 2644 845 2645 875
rect 2645 845 2675 875
rect 2675 845 2676 875
rect 2644 844 2676 845
rect 2644 764 2676 796
rect 2644 684 2676 716
rect 2644 635 2676 636
rect 2644 605 2645 635
rect 2645 605 2675 635
rect 2675 605 2676 635
rect 2644 604 2676 605
rect 2644 555 2676 556
rect 2644 525 2645 555
rect 2645 525 2675 555
rect 2675 525 2676 555
rect 2644 524 2676 525
rect 2644 444 2676 476
rect 2644 395 2676 396
rect 2644 365 2645 395
rect 2645 365 2675 395
rect 2675 365 2676 395
rect 2644 364 2676 365
rect 2644 284 2676 316
rect 2644 235 2676 236
rect 2644 205 2645 235
rect 2645 205 2675 235
rect 2675 205 2676 235
rect 2644 204 2676 205
rect 2644 124 2676 156
rect 2644 75 2676 76
rect 2644 45 2645 75
rect 2645 45 2675 75
rect 2675 45 2676 75
rect 2644 44 2676 45
rect 2644 -5 2676 -4
rect 2644 -35 2645 -5
rect 2645 -35 2675 -5
rect 2675 -35 2676 -5
rect 2644 -36 2676 -35
rect 2644 -85 2676 -84
rect 2644 -115 2645 -85
rect 2645 -115 2675 -85
rect 2675 -115 2676 -85
rect 2644 -116 2676 -115
rect 2724 1035 2756 1036
rect 2724 1005 2725 1035
rect 2725 1005 2755 1035
rect 2755 1005 2756 1035
rect 2724 1004 2756 1005
rect 2724 955 2756 956
rect 2724 925 2725 955
rect 2725 925 2755 955
rect 2755 925 2756 955
rect 2724 924 2756 925
rect 2724 875 2756 876
rect 2724 845 2725 875
rect 2725 845 2755 875
rect 2755 845 2756 875
rect 2724 844 2756 845
rect 2724 764 2756 796
rect 2724 684 2756 716
rect 2724 635 2756 636
rect 2724 605 2725 635
rect 2725 605 2755 635
rect 2755 605 2756 635
rect 2724 604 2756 605
rect 2724 555 2756 556
rect 2724 525 2725 555
rect 2725 525 2755 555
rect 2755 525 2756 555
rect 2724 524 2756 525
rect 2724 444 2756 476
rect 2724 395 2756 396
rect 2724 365 2725 395
rect 2725 365 2755 395
rect 2755 365 2756 395
rect 2724 364 2756 365
rect 2724 284 2756 316
rect 2724 235 2756 236
rect 2724 205 2725 235
rect 2725 205 2755 235
rect 2755 205 2756 235
rect 2724 204 2756 205
rect 2724 124 2756 156
rect 2724 75 2756 76
rect 2724 45 2725 75
rect 2725 45 2755 75
rect 2755 45 2756 75
rect 2724 44 2756 45
rect 2724 -5 2756 -4
rect 2724 -35 2725 -5
rect 2725 -35 2755 -5
rect 2755 -35 2756 -5
rect 2724 -36 2756 -35
rect 2724 -85 2756 -84
rect 2724 -115 2725 -85
rect 2725 -115 2755 -85
rect 2755 -115 2756 -85
rect 2724 -116 2756 -115
rect 2804 1035 2836 1036
rect 2804 1005 2805 1035
rect 2805 1005 2835 1035
rect 2835 1005 2836 1035
rect 2804 1004 2836 1005
rect 2804 955 2836 956
rect 2804 925 2805 955
rect 2805 925 2835 955
rect 2835 925 2836 955
rect 2804 924 2836 925
rect 2804 875 2836 876
rect 2804 845 2805 875
rect 2805 845 2835 875
rect 2835 845 2836 875
rect 2804 844 2836 845
rect 2804 764 2836 796
rect 2804 684 2836 716
rect 2804 635 2836 636
rect 2804 605 2805 635
rect 2805 605 2835 635
rect 2835 605 2836 635
rect 2804 604 2836 605
rect 2804 555 2836 556
rect 2804 525 2805 555
rect 2805 525 2835 555
rect 2835 525 2836 555
rect 2804 524 2836 525
rect 2804 444 2836 476
rect 2804 395 2836 396
rect 2804 365 2805 395
rect 2805 365 2835 395
rect 2835 365 2836 395
rect 2804 364 2836 365
rect 2804 284 2836 316
rect 2804 235 2836 236
rect 2804 205 2805 235
rect 2805 205 2835 235
rect 2835 205 2836 235
rect 2804 204 2836 205
rect 2804 124 2836 156
rect 2804 75 2836 76
rect 2804 45 2805 75
rect 2805 45 2835 75
rect 2835 45 2836 75
rect 2804 44 2836 45
rect 2804 -5 2836 -4
rect 2804 -35 2805 -5
rect 2805 -35 2835 -5
rect 2835 -35 2836 -5
rect 2804 -36 2836 -35
rect 2804 -85 2836 -84
rect 2804 -115 2805 -85
rect 2805 -115 2835 -85
rect 2835 -115 2836 -85
rect 2804 -116 2836 -115
rect 2884 1035 2916 1036
rect 2884 1005 2885 1035
rect 2885 1005 2915 1035
rect 2915 1005 2916 1035
rect 2884 1004 2916 1005
rect 2884 955 2916 956
rect 2884 925 2885 955
rect 2885 925 2915 955
rect 2915 925 2916 955
rect 2884 924 2916 925
rect 2884 875 2916 876
rect 2884 845 2885 875
rect 2885 845 2915 875
rect 2915 845 2916 875
rect 2884 844 2916 845
rect 2884 764 2916 796
rect 2884 684 2916 716
rect 2884 635 2916 636
rect 2884 605 2885 635
rect 2885 605 2915 635
rect 2915 605 2916 635
rect 2884 604 2916 605
rect 2884 555 2916 556
rect 2884 525 2885 555
rect 2885 525 2915 555
rect 2915 525 2916 555
rect 2884 524 2916 525
rect 2884 444 2916 476
rect 2884 395 2916 396
rect 2884 365 2885 395
rect 2885 365 2915 395
rect 2915 365 2916 395
rect 2884 364 2916 365
rect 2884 284 2916 316
rect 2884 235 2916 236
rect 2884 205 2885 235
rect 2885 205 2915 235
rect 2915 205 2916 235
rect 2884 204 2916 205
rect 2884 124 2916 156
rect 2884 75 2916 76
rect 2884 45 2885 75
rect 2885 45 2915 75
rect 2915 45 2916 75
rect 2884 44 2916 45
rect 2884 -5 2916 -4
rect 2884 -35 2885 -5
rect 2885 -35 2915 -5
rect 2915 -35 2916 -5
rect 2884 -36 2916 -35
rect 2884 -85 2916 -84
rect 2884 -115 2885 -85
rect 2885 -115 2915 -85
rect 2915 -115 2916 -85
rect 2884 -116 2916 -115
rect 2964 1035 2996 1036
rect 2964 1005 2965 1035
rect 2965 1005 2995 1035
rect 2995 1005 2996 1035
rect 2964 1004 2996 1005
rect 2964 955 2996 956
rect 2964 925 2965 955
rect 2965 925 2995 955
rect 2995 925 2996 955
rect 2964 924 2996 925
rect 2964 875 2996 876
rect 2964 845 2965 875
rect 2965 845 2995 875
rect 2995 845 2996 875
rect 2964 844 2996 845
rect 2964 764 2996 796
rect 2964 684 2996 716
rect 2964 635 2996 636
rect 2964 605 2965 635
rect 2965 605 2995 635
rect 2995 605 2996 635
rect 2964 604 2996 605
rect 2964 555 2996 556
rect 2964 525 2965 555
rect 2965 525 2995 555
rect 2995 525 2996 555
rect 2964 524 2996 525
rect 2964 444 2996 476
rect 2964 395 2996 396
rect 2964 365 2965 395
rect 2965 365 2995 395
rect 2995 365 2996 395
rect 2964 364 2996 365
rect 2964 284 2996 316
rect 2964 235 2996 236
rect 2964 205 2965 235
rect 2965 205 2995 235
rect 2995 205 2996 235
rect 2964 204 2996 205
rect 2964 124 2996 156
rect 2964 75 2996 76
rect 2964 45 2965 75
rect 2965 45 2995 75
rect 2995 45 2996 75
rect 2964 44 2996 45
rect 2964 -5 2996 -4
rect 2964 -35 2965 -5
rect 2965 -35 2995 -5
rect 2995 -35 2996 -5
rect 2964 -36 2996 -35
rect 2964 -85 2996 -84
rect 2964 -115 2965 -85
rect 2965 -115 2995 -85
rect 2995 -115 2996 -85
rect 2964 -116 2996 -115
rect 3044 1035 3076 1036
rect 3044 1005 3045 1035
rect 3045 1005 3075 1035
rect 3075 1005 3076 1035
rect 3044 1004 3076 1005
rect 3044 955 3076 956
rect 3044 925 3045 955
rect 3045 925 3075 955
rect 3075 925 3076 955
rect 3044 924 3076 925
rect 3044 875 3076 876
rect 3044 845 3045 875
rect 3045 845 3075 875
rect 3075 845 3076 875
rect 3044 844 3076 845
rect 3044 764 3076 796
rect 3044 684 3076 716
rect 3044 635 3076 636
rect 3044 605 3045 635
rect 3045 605 3075 635
rect 3075 605 3076 635
rect 3044 604 3076 605
rect 3044 555 3076 556
rect 3044 525 3045 555
rect 3045 525 3075 555
rect 3075 525 3076 555
rect 3044 524 3076 525
rect 3044 444 3076 476
rect 3044 395 3076 396
rect 3044 365 3045 395
rect 3045 365 3075 395
rect 3075 365 3076 395
rect 3044 364 3076 365
rect 3044 284 3076 316
rect 3044 235 3076 236
rect 3044 205 3045 235
rect 3045 205 3075 235
rect 3075 205 3076 235
rect 3044 204 3076 205
rect 3044 124 3076 156
rect 3044 75 3076 76
rect 3044 45 3045 75
rect 3045 45 3075 75
rect 3075 45 3076 75
rect 3044 44 3076 45
rect 3044 -5 3076 -4
rect 3044 -35 3045 -5
rect 3045 -35 3075 -5
rect 3075 -35 3076 -5
rect 3044 -36 3076 -35
rect 3044 -85 3076 -84
rect 3044 -115 3045 -85
rect 3045 -115 3075 -85
rect 3075 -115 3076 -85
rect 3044 -116 3076 -115
rect 3124 1035 3156 1036
rect 3124 1005 3125 1035
rect 3125 1005 3155 1035
rect 3155 1005 3156 1035
rect 3124 1004 3156 1005
rect 3124 955 3156 956
rect 3124 925 3125 955
rect 3125 925 3155 955
rect 3155 925 3156 955
rect 3124 924 3156 925
rect 3124 875 3156 876
rect 3124 845 3125 875
rect 3125 845 3155 875
rect 3155 845 3156 875
rect 3124 844 3156 845
rect 3124 764 3156 796
rect 3124 684 3156 716
rect 3124 635 3156 636
rect 3124 605 3125 635
rect 3125 605 3155 635
rect 3155 605 3156 635
rect 3124 604 3156 605
rect 3124 555 3156 556
rect 3124 525 3125 555
rect 3125 525 3155 555
rect 3155 525 3156 555
rect 3124 524 3156 525
rect 3124 444 3156 476
rect 3124 395 3156 396
rect 3124 365 3125 395
rect 3125 365 3155 395
rect 3155 365 3156 395
rect 3124 364 3156 365
rect 3124 284 3156 316
rect 3124 235 3156 236
rect 3124 205 3125 235
rect 3125 205 3155 235
rect 3155 205 3156 235
rect 3124 204 3156 205
rect 3124 124 3156 156
rect 3124 75 3156 76
rect 3124 45 3125 75
rect 3125 45 3155 75
rect 3155 45 3156 75
rect 3124 44 3156 45
rect 3124 -5 3156 -4
rect 3124 -35 3125 -5
rect 3125 -35 3155 -5
rect 3155 -35 3156 -5
rect 3124 -36 3156 -35
rect 3124 -85 3156 -84
rect 3124 -115 3125 -85
rect 3125 -115 3155 -85
rect 3155 -115 3156 -85
rect 3124 -116 3156 -115
rect 3204 1035 3236 1036
rect 3204 1005 3205 1035
rect 3205 1005 3235 1035
rect 3235 1005 3236 1035
rect 3204 1004 3236 1005
rect 3204 955 3236 956
rect 3204 925 3205 955
rect 3205 925 3235 955
rect 3235 925 3236 955
rect 3204 924 3236 925
rect 3204 875 3236 876
rect 3204 845 3205 875
rect 3205 845 3235 875
rect 3235 845 3236 875
rect 3204 844 3236 845
rect 3204 764 3236 796
rect 3204 684 3236 716
rect 3204 635 3236 636
rect 3204 605 3205 635
rect 3205 605 3235 635
rect 3235 605 3236 635
rect 3204 604 3236 605
rect 3204 555 3236 556
rect 3204 525 3205 555
rect 3205 525 3235 555
rect 3235 525 3236 555
rect 3204 524 3236 525
rect 3204 444 3236 476
rect 3204 395 3236 396
rect 3204 365 3205 395
rect 3205 365 3235 395
rect 3235 365 3236 395
rect 3204 364 3236 365
rect 3204 284 3236 316
rect 3204 235 3236 236
rect 3204 205 3205 235
rect 3205 205 3235 235
rect 3235 205 3236 235
rect 3204 204 3236 205
rect 3204 124 3236 156
rect 3204 75 3236 76
rect 3204 45 3205 75
rect 3205 45 3235 75
rect 3235 45 3236 75
rect 3204 44 3236 45
rect 3204 -5 3236 -4
rect 3204 -35 3205 -5
rect 3205 -35 3235 -5
rect 3235 -35 3236 -5
rect 3204 -36 3236 -35
rect 3204 -85 3236 -84
rect 3204 -115 3205 -85
rect 3205 -115 3235 -85
rect 3235 -115 3236 -85
rect 3204 -116 3236 -115
rect 3284 1035 3316 1036
rect 3284 1005 3285 1035
rect 3285 1005 3315 1035
rect 3315 1005 3316 1035
rect 3284 1004 3316 1005
rect 3284 955 3316 956
rect 3284 925 3285 955
rect 3285 925 3315 955
rect 3315 925 3316 955
rect 3284 924 3316 925
rect 3284 875 3316 876
rect 3284 845 3285 875
rect 3285 845 3315 875
rect 3315 845 3316 875
rect 3284 844 3316 845
rect 3284 764 3316 796
rect 3284 684 3316 716
rect 3284 635 3316 636
rect 3284 605 3285 635
rect 3285 605 3315 635
rect 3315 605 3316 635
rect 3284 604 3316 605
rect 3284 555 3316 556
rect 3284 525 3285 555
rect 3285 525 3315 555
rect 3315 525 3316 555
rect 3284 524 3316 525
rect 3284 444 3316 476
rect 3284 395 3316 396
rect 3284 365 3285 395
rect 3285 365 3315 395
rect 3315 365 3316 395
rect 3284 364 3316 365
rect 3284 284 3316 316
rect 3284 235 3316 236
rect 3284 205 3285 235
rect 3285 205 3315 235
rect 3315 205 3316 235
rect 3284 204 3316 205
rect 3284 124 3316 156
rect 3284 75 3316 76
rect 3284 45 3285 75
rect 3285 45 3315 75
rect 3315 45 3316 75
rect 3284 44 3316 45
rect 3284 -5 3316 -4
rect 3284 -35 3285 -5
rect 3285 -35 3315 -5
rect 3315 -35 3316 -5
rect 3284 -36 3316 -35
rect 3284 -85 3316 -84
rect 3284 -115 3285 -85
rect 3285 -115 3315 -85
rect 3315 -115 3316 -85
rect 3284 -116 3316 -115
rect 3364 1035 3396 1036
rect 3364 1005 3365 1035
rect 3365 1005 3395 1035
rect 3395 1005 3396 1035
rect 3364 1004 3396 1005
rect 3364 955 3396 956
rect 3364 925 3365 955
rect 3365 925 3395 955
rect 3395 925 3396 955
rect 3364 924 3396 925
rect 3364 875 3396 876
rect 3364 845 3365 875
rect 3365 845 3395 875
rect 3395 845 3396 875
rect 3364 844 3396 845
rect 3364 764 3396 796
rect 3364 684 3396 716
rect 3364 635 3396 636
rect 3364 605 3365 635
rect 3365 605 3395 635
rect 3395 605 3396 635
rect 3364 604 3396 605
rect 3364 555 3396 556
rect 3364 525 3365 555
rect 3365 525 3395 555
rect 3395 525 3396 555
rect 3364 524 3396 525
rect 3364 444 3396 476
rect 3364 395 3396 396
rect 3364 365 3365 395
rect 3365 365 3395 395
rect 3395 365 3396 395
rect 3364 364 3396 365
rect 3364 284 3396 316
rect 3364 235 3396 236
rect 3364 205 3365 235
rect 3365 205 3395 235
rect 3395 205 3396 235
rect 3364 204 3396 205
rect 3364 124 3396 156
rect 3364 75 3396 76
rect 3364 45 3365 75
rect 3365 45 3395 75
rect 3395 45 3396 75
rect 3364 44 3396 45
rect 3364 -5 3396 -4
rect 3364 -35 3365 -5
rect 3365 -35 3395 -5
rect 3395 -35 3396 -5
rect 3364 -36 3396 -35
rect 3364 -85 3396 -84
rect 3364 -115 3365 -85
rect 3365 -115 3395 -85
rect 3395 -115 3396 -85
rect 3364 -116 3396 -115
rect 3444 1035 3476 1036
rect 3444 1005 3445 1035
rect 3445 1005 3475 1035
rect 3475 1005 3476 1035
rect 3444 1004 3476 1005
rect 3444 955 3476 956
rect 3444 925 3445 955
rect 3445 925 3475 955
rect 3475 925 3476 955
rect 3444 924 3476 925
rect 3444 875 3476 876
rect 3444 845 3445 875
rect 3445 845 3475 875
rect 3475 845 3476 875
rect 3444 844 3476 845
rect 3444 764 3476 796
rect 3444 684 3476 716
rect 3444 635 3476 636
rect 3444 605 3445 635
rect 3445 605 3475 635
rect 3475 605 3476 635
rect 3444 604 3476 605
rect 3444 555 3476 556
rect 3444 525 3445 555
rect 3445 525 3475 555
rect 3475 525 3476 555
rect 3444 524 3476 525
rect 3444 444 3476 476
rect 3444 395 3476 396
rect 3444 365 3445 395
rect 3445 365 3475 395
rect 3475 365 3476 395
rect 3444 364 3476 365
rect 3444 284 3476 316
rect 3444 235 3476 236
rect 3444 205 3445 235
rect 3445 205 3475 235
rect 3475 205 3476 235
rect 3444 204 3476 205
rect 3444 124 3476 156
rect 3444 75 3476 76
rect 3444 45 3445 75
rect 3445 45 3475 75
rect 3475 45 3476 75
rect 3444 44 3476 45
rect 3444 -5 3476 -4
rect 3444 -35 3445 -5
rect 3445 -35 3475 -5
rect 3475 -35 3476 -5
rect 3444 -36 3476 -35
rect 3444 -85 3476 -84
rect 3444 -115 3445 -85
rect 3445 -115 3475 -85
rect 3475 -115 3476 -85
rect 3444 -116 3476 -115
rect 3524 1035 3556 1036
rect 3524 1005 3525 1035
rect 3525 1005 3555 1035
rect 3555 1005 3556 1035
rect 3524 1004 3556 1005
rect 3524 955 3556 956
rect 3524 925 3525 955
rect 3525 925 3555 955
rect 3555 925 3556 955
rect 3524 924 3556 925
rect 3524 875 3556 876
rect 3524 845 3525 875
rect 3525 845 3555 875
rect 3555 845 3556 875
rect 3524 844 3556 845
rect 3524 764 3556 796
rect 3524 684 3556 716
rect 3524 635 3556 636
rect 3524 605 3525 635
rect 3525 605 3555 635
rect 3555 605 3556 635
rect 3524 604 3556 605
rect 3524 555 3556 556
rect 3524 525 3525 555
rect 3525 525 3555 555
rect 3555 525 3556 555
rect 3524 524 3556 525
rect 3524 444 3556 476
rect 3524 395 3556 396
rect 3524 365 3525 395
rect 3525 365 3555 395
rect 3555 365 3556 395
rect 3524 364 3556 365
rect 3524 284 3556 316
rect 3524 235 3556 236
rect 3524 205 3525 235
rect 3525 205 3555 235
rect 3555 205 3556 235
rect 3524 204 3556 205
rect 3524 124 3556 156
rect 3524 75 3556 76
rect 3524 45 3525 75
rect 3525 45 3555 75
rect 3555 45 3556 75
rect 3524 44 3556 45
rect 3524 -5 3556 -4
rect 3524 -35 3525 -5
rect 3525 -35 3555 -5
rect 3555 -35 3556 -5
rect 3524 -36 3556 -35
rect 3524 -85 3556 -84
rect 3524 -115 3525 -85
rect 3525 -115 3555 -85
rect 3555 -115 3556 -85
rect 3524 -116 3556 -115
rect 3604 1035 3636 1036
rect 3604 1005 3605 1035
rect 3605 1005 3635 1035
rect 3635 1005 3636 1035
rect 3604 1004 3636 1005
rect 3604 955 3636 956
rect 3604 925 3605 955
rect 3605 925 3635 955
rect 3635 925 3636 955
rect 3604 924 3636 925
rect 3604 875 3636 876
rect 3604 845 3605 875
rect 3605 845 3635 875
rect 3635 845 3636 875
rect 3604 844 3636 845
rect 3604 764 3636 796
rect 3604 684 3636 716
rect 3604 635 3636 636
rect 3604 605 3605 635
rect 3605 605 3635 635
rect 3635 605 3636 635
rect 3604 604 3636 605
rect 3604 555 3636 556
rect 3604 525 3605 555
rect 3605 525 3635 555
rect 3635 525 3636 555
rect 3604 524 3636 525
rect 3604 444 3636 476
rect 3604 395 3636 396
rect 3604 365 3605 395
rect 3605 365 3635 395
rect 3635 365 3636 395
rect 3604 364 3636 365
rect 3604 284 3636 316
rect 3604 235 3636 236
rect 3604 205 3605 235
rect 3605 205 3635 235
rect 3635 205 3636 235
rect 3604 204 3636 205
rect 3604 124 3636 156
rect 3604 75 3636 76
rect 3604 45 3605 75
rect 3605 45 3635 75
rect 3635 45 3636 75
rect 3604 44 3636 45
rect 3604 -5 3636 -4
rect 3604 -35 3605 -5
rect 3605 -35 3635 -5
rect 3635 -35 3636 -5
rect 3604 -36 3636 -35
rect 3604 -85 3636 -84
rect 3604 -115 3605 -85
rect 3605 -115 3635 -85
rect 3635 -115 3636 -85
rect 3604 -116 3636 -115
rect 3684 1035 3716 1036
rect 3684 1005 3685 1035
rect 3685 1005 3715 1035
rect 3715 1005 3716 1035
rect 3684 1004 3716 1005
rect 3684 955 3716 956
rect 3684 925 3685 955
rect 3685 925 3715 955
rect 3715 925 3716 955
rect 3684 924 3716 925
rect 3684 875 3716 876
rect 3684 845 3685 875
rect 3685 845 3715 875
rect 3715 845 3716 875
rect 3684 844 3716 845
rect 3684 764 3716 796
rect 3684 684 3716 716
rect 3684 635 3716 636
rect 3684 605 3685 635
rect 3685 605 3715 635
rect 3715 605 3716 635
rect 3684 604 3716 605
rect 3684 555 3716 556
rect 3684 525 3685 555
rect 3685 525 3715 555
rect 3715 525 3716 555
rect 3684 524 3716 525
rect 3684 444 3716 476
rect 3684 395 3716 396
rect 3684 365 3685 395
rect 3685 365 3715 395
rect 3715 365 3716 395
rect 3684 364 3716 365
rect 3684 284 3716 316
rect 3684 235 3716 236
rect 3684 205 3685 235
rect 3685 205 3715 235
rect 3715 205 3716 235
rect 3684 204 3716 205
rect 3684 124 3716 156
rect 3684 75 3716 76
rect 3684 45 3685 75
rect 3685 45 3715 75
rect 3715 45 3716 75
rect 3684 44 3716 45
rect 3684 -5 3716 -4
rect 3684 -35 3685 -5
rect 3685 -35 3715 -5
rect 3715 -35 3716 -5
rect 3684 -36 3716 -35
rect 3684 -85 3716 -84
rect 3684 -115 3685 -85
rect 3685 -115 3715 -85
rect 3715 -115 3716 -85
rect 3684 -116 3716 -115
rect 3764 1035 3796 1036
rect 3764 1005 3765 1035
rect 3765 1005 3795 1035
rect 3795 1005 3796 1035
rect 3764 1004 3796 1005
rect 3764 955 3796 956
rect 3764 925 3765 955
rect 3765 925 3795 955
rect 3795 925 3796 955
rect 3764 924 3796 925
rect 3764 875 3796 876
rect 3764 845 3765 875
rect 3765 845 3795 875
rect 3795 845 3796 875
rect 3764 844 3796 845
rect 3764 764 3796 796
rect 3764 684 3796 716
rect 3764 635 3796 636
rect 3764 605 3765 635
rect 3765 605 3795 635
rect 3795 605 3796 635
rect 3764 604 3796 605
rect 3764 555 3796 556
rect 3764 525 3765 555
rect 3765 525 3795 555
rect 3795 525 3796 555
rect 3764 524 3796 525
rect 3764 444 3796 476
rect 3764 395 3796 396
rect 3764 365 3765 395
rect 3765 365 3795 395
rect 3795 365 3796 395
rect 3764 364 3796 365
rect 3764 284 3796 316
rect 3764 235 3796 236
rect 3764 205 3765 235
rect 3765 205 3795 235
rect 3795 205 3796 235
rect 3764 204 3796 205
rect 3764 124 3796 156
rect 3764 75 3796 76
rect 3764 45 3765 75
rect 3765 45 3795 75
rect 3795 45 3796 75
rect 3764 44 3796 45
rect 3764 -5 3796 -4
rect 3764 -35 3765 -5
rect 3765 -35 3795 -5
rect 3795 -35 3796 -5
rect 3764 -36 3796 -35
rect 3764 -85 3796 -84
rect 3764 -115 3765 -85
rect 3765 -115 3795 -85
rect 3795 -115 3796 -85
rect 3764 -116 3796 -115
rect 3844 1035 3876 1036
rect 3844 1005 3845 1035
rect 3845 1005 3875 1035
rect 3875 1005 3876 1035
rect 3844 1004 3876 1005
rect 3844 955 3876 956
rect 3844 925 3845 955
rect 3845 925 3875 955
rect 3875 925 3876 955
rect 3844 924 3876 925
rect 3844 875 3876 876
rect 3844 845 3845 875
rect 3845 845 3875 875
rect 3875 845 3876 875
rect 3844 844 3876 845
rect 3844 764 3876 796
rect 3844 684 3876 716
rect 3844 635 3876 636
rect 3844 605 3845 635
rect 3845 605 3875 635
rect 3875 605 3876 635
rect 3844 604 3876 605
rect 3844 555 3876 556
rect 3844 525 3845 555
rect 3845 525 3875 555
rect 3875 525 3876 555
rect 3844 524 3876 525
rect 3844 444 3876 476
rect 3844 395 3876 396
rect 3844 365 3845 395
rect 3845 365 3875 395
rect 3875 365 3876 395
rect 3844 364 3876 365
rect 3844 284 3876 316
rect 3844 235 3876 236
rect 3844 205 3845 235
rect 3845 205 3875 235
rect 3875 205 3876 235
rect 3844 204 3876 205
rect 3844 124 3876 156
rect 3844 75 3876 76
rect 3844 45 3845 75
rect 3845 45 3875 75
rect 3875 45 3876 75
rect 3844 44 3876 45
rect 3844 -5 3876 -4
rect 3844 -35 3845 -5
rect 3845 -35 3875 -5
rect 3875 -35 3876 -5
rect 3844 -36 3876 -35
rect 3844 -85 3876 -84
rect 3844 -115 3845 -85
rect 3845 -115 3875 -85
rect 3875 -115 3876 -85
rect 3844 -116 3876 -115
rect 3924 1035 3956 1036
rect 3924 1005 3925 1035
rect 3925 1005 3955 1035
rect 3955 1005 3956 1035
rect 3924 1004 3956 1005
rect 3924 955 3956 956
rect 3924 925 3925 955
rect 3925 925 3955 955
rect 3955 925 3956 955
rect 3924 924 3956 925
rect 3924 875 3956 876
rect 3924 845 3925 875
rect 3925 845 3955 875
rect 3955 845 3956 875
rect 3924 844 3956 845
rect 3924 764 3956 796
rect 3924 684 3956 716
rect 3924 635 3956 636
rect 3924 605 3925 635
rect 3925 605 3955 635
rect 3955 605 3956 635
rect 3924 604 3956 605
rect 3924 555 3956 556
rect 3924 525 3925 555
rect 3925 525 3955 555
rect 3955 525 3956 555
rect 3924 524 3956 525
rect 3924 444 3956 476
rect 3924 395 3956 396
rect 3924 365 3925 395
rect 3925 365 3955 395
rect 3955 365 3956 395
rect 3924 364 3956 365
rect 3924 284 3956 316
rect 3924 235 3956 236
rect 3924 205 3925 235
rect 3925 205 3955 235
rect 3955 205 3956 235
rect 3924 204 3956 205
rect 3924 124 3956 156
rect 3924 75 3956 76
rect 3924 45 3925 75
rect 3925 45 3955 75
rect 3955 45 3956 75
rect 3924 44 3956 45
rect 3924 -5 3956 -4
rect 3924 -35 3925 -5
rect 3925 -35 3955 -5
rect 3955 -35 3956 -5
rect 3924 -36 3956 -35
rect 3924 -85 3956 -84
rect 3924 -115 3925 -85
rect 3925 -115 3955 -85
rect 3955 -115 3956 -85
rect 3924 -116 3956 -115
rect 4004 1035 4036 1036
rect 4004 1005 4005 1035
rect 4005 1005 4035 1035
rect 4035 1005 4036 1035
rect 4004 1004 4036 1005
rect 4004 955 4036 956
rect 4004 925 4005 955
rect 4005 925 4035 955
rect 4035 925 4036 955
rect 4004 924 4036 925
rect 4004 875 4036 876
rect 4004 845 4005 875
rect 4005 845 4035 875
rect 4035 845 4036 875
rect 4004 844 4036 845
rect 4004 764 4036 796
rect 4004 684 4036 716
rect 4004 635 4036 636
rect 4004 605 4005 635
rect 4005 605 4035 635
rect 4035 605 4036 635
rect 4004 604 4036 605
rect 4004 555 4036 556
rect 4004 525 4005 555
rect 4005 525 4035 555
rect 4035 525 4036 555
rect 4004 524 4036 525
rect 4004 444 4036 476
rect 4004 395 4036 396
rect 4004 365 4005 395
rect 4005 365 4035 395
rect 4035 365 4036 395
rect 4004 364 4036 365
rect 4004 284 4036 316
rect 4004 235 4036 236
rect 4004 205 4005 235
rect 4005 205 4035 235
rect 4035 205 4036 235
rect 4004 204 4036 205
rect 4004 124 4036 156
rect 4004 75 4036 76
rect 4004 45 4005 75
rect 4005 45 4035 75
rect 4035 45 4036 75
rect 4004 44 4036 45
rect 4004 -5 4036 -4
rect 4004 -35 4005 -5
rect 4005 -35 4035 -5
rect 4035 -35 4036 -5
rect 4004 -36 4036 -35
rect 4004 -85 4036 -84
rect 4004 -115 4005 -85
rect 4005 -115 4035 -85
rect 4035 -115 4036 -85
rect 4004 -116 4036 -115
rect 4084 1035 4116 1036
rect 4084 1005 4085 1035
rect 4085 1005 4115 1035
rect 4115 1005 4116 1035
rect 4084 1004 4116 1005
rect 4084 955 4116 956
rect 4084 925 4085 955
rect 4085 925 4115 955
rect 4115 925 4116 955
rect 4084 924 4116 925
rect 4084 875 4116 876
rect 4084 845 4085 875
rect 4085 845 4115 875
rect 4115 845 4116 875
rect 4084 844 4116 845
rect 4084 764 4116 796
rect 4084 684 4116 716
rect 4084 635 4116 636
rect 4084 605 4085 635
rect 4085 605 4115 635
rect 4115 605 4116 635
rect 4084 604 4116 605
rect 4084 555 4116 556
rect 4084 525 4085 555
rect 4085 525 4115 555
rect 4115 525 4116 555
rect 4084 524 4116 525
rect 4084 444 4116 476
rect 4084 395 4116 396
rect 4084 365 4085 395
rect 4085 365 4115 395
rect 4115 365 4116 395
rect 4084 364 4116 365
rect 4084 284 4116 316
rect 4084 235 4116 236
rect 4084 205 4085 235
rect 4085 205 4115 235
rect 4115 205 4116 235
rect 4084 204 4116 205
rect 4084 124 4116 156
rect 4084 75 4116 76
rect 4084 45 4085 75
rect 4085 45 4115 75
rect 4115 45 4116 75
rect 4084 44 4116 45
rect 4084 -5 4116 -4
rect 4084 -35 4085 -5
rect 4085 -35 4115 -5
rect 4115 -35 4116 -5
rect 4084 -36 4116 -35
rect 4084 -85 4116 -84
rect 4084 -115 4085 -85
rect 4085 -115 4115 -85
rect 4115 -115 4116 -85
rect 4084 -116 4116 -115
rect 4164 1035 4196 1036
rect 4164 1005 4165 1035
rect 4165 1005 4195 1035
rect 4195 1005 4196 1035
rect 4164 1004 4196 1005
rect 4164 955 4196 956
rect 4164 925 4165 955
rect 4165 925 4195 955
rect 4195 925 4196 955
rect 4164 924 4196 925
rect 4164 875 4196 876
rect 4164 845 4165 875
rect 4165 845 4195 875
rect 4195 845 4196 875
rect 4164 844 4196 845
rect 4164 764 4196 796
rect 4164 684 4196 716
rect 4164 635 4196 636
rect 4164 605 4165 635
rect 4165 605 4195 635
rect 4195 605 4196 635
rect 4164 604 4196 605
rect 4164 555 4196 556
rect 4164 525 4165 555
rect 4165 525 4195 555
rect 4195 525 4196 555
rect 4164 524 4196 525
rect 4164 444 4196 476
rect 4164 395 4196 396
rect 4164 365 4165 395
rect 4165 365 4195 395
rect 4195 365 4196 395
rect 4164 364 4196 365
rect 4164 284 4196 316
rect 4164 235 4196 236
rect 4164 205 4165 235
rect 4165 205 4195 235
rect 4195 205 4196 235
rect 4164 204 4196 205
rect 4164 124 4196 156
rect 4164 75 4196 76
rect 4164 45 4165 75
rect 4165 45 4195 75
rect 4195 45 4196 75
rect 4164 44 4196 45
rect 4164 -5 4196 -4
rect 4164 -35 4165 -5
rect 4165 -35 4195 -5
rect 4195 -35 4196 -5
rect 4164 -36 4196 -35
rect 4164 -85 4196 -84
rect 4164 -115 4165 -85
rect 4165 -115 4195 -85
rect 4195 -115 4196 -85
rect 4164 -116 4196 -115
rect 4244 1035 4276 1036
rect 4244 1005 4245 1035
rect 4245 1005 4275 1035
rect 4275 1005 4276 1035
rect 4244 1004 4276 1005
rect 4244 955 4276 956
rect 4244 925 4245 955
rect 4245 925 4275 955
rect 4275 925 4276 955
rect 4244 924 4276 925
rect 4244 875 4276 876
rect 4244 845 4245 875
rect 4245 845 4275 875
rect 4275 845 4276 875
rect 4244 844 4276 845
rect 4244 764 4276 796
rect 4244 684 4276 716
rect 4244 635 4276 636
rect 4244 605 4245 635
rect 4245 605 4275 635
rect 4275 605 4276 635
rect 4244 604 4276 605
rect 4244 555 4276 556
rect 4244 525 4245 555
rect 4245 525 4275 555
rect 4275 525 4276 555
rect 4244 524 4276 525
rect 4244 444 4276 476
rect 4244 395 4276 396
rect 4244 365 4245 395
rect 4245 365 4275 395
rect 4275 365 4276 395
rect 4244 364 4276 365
rect 4244 284 4276 316
rect 4244 235 4276 236
rect 4244 205 4245 235
rect 4245 205 4275 235
rect 4275 205 4276 235
rect 4244 204 4276 205
rect 4244 124 4276 156
rect 4244 75 4276 76
rect 4244 45 4245 75
rect 4245 45 4275 75
rect 4275 45 4276 75
rect 4244 44 4276 45
rect 4244 -5 4276 -4
rect 4244 -35 4245 -5
rect 4245 -35 4275 -5
rect 4275 -35 4276 -5
rect 4244 -36 4276 -35
rect 4244 -85 4276 -84
rect 4244 -115 4245 -85
rect 4245 -115 4275 -85
rect 4275 -115 4276 -85
rect 4244 -116 4276 -115
rect 4324 1035 4356 1036
rect 4324 1005 4325 1035
rect 4325 1005 4355 1035
rect 4355 1005 4356 1035
rect 4324 1004 4356 1005
rect 4324 955 4356 956
rect 4324 925 4325 955
rect 4325 925 4355 955
rect 4355 925 4356 955
rect 4324 924 4356 925
rect 4324 875 4356 876
rect 4324 845 4325 875
rect 4325 845 4355 875
rect 4355 845 4356 875
rect 4324 844 4356 845
rect 4324 764 4356 796
rect 4324 684 4356 716
rect 4324 635 4356 636
rect 4324 605 4325 635
rect 4325 605 4355 635
rect 4355 605 4356 635
rect 4324 604 4356 605
rect 4324 555 4356 556
rect 4324 525 4325 555
rect 4325 525 4355 555
rect 4355 525 4356 555
rect 4324 524 4356 525
rect 4324 444 4356 476
rect 4324 395 4356 396
rect 4324 365 4325 395
rect 4325 365 4355 395
rect 4355 365 4356 395
rect 4324 364 4356 365
rect 4324 284 4356 316
rect 4324 235 4356 236
rect 4324 205 4325 235
rect 4325 205 4355 235
rect 4355 205 4356 235
rect 4324 204 4356 205
rect 4324 124 4356 156
rect 4324 75 4356 76
rect 4324 45 4325 75
rect 4325 45 4355 75
rect 4355 45 4356 75
rect 4324 44 4356 45
rect 4324 -5 4356 -4
rect 4324 -35 4325 -5
rect 4325 -35 4355 -5
rect 4355 -35 4356 -5
rect 4324 -36 4356 -35
rect 4324 -85 4356 -84
rect 4324 -115 4325 -85
rect 4325 -115 4355 -85
rect 4355 -115 4356 -85
rect 4324 -116 4356 -115
rect 4404 1035 4436 1036
rect 4404 1005 4405 1035
rect 4405 1005 4435 1035
rect 4435 1005 4436 1035
rect 4404 1004 4436 1005
rect 4404 955 4436 956
rect 4404 925 4405 955
rect 4405 925 4435 955
rect 4435 925 4436 955
rect 4404 924 4436 925
rect 4404 875 4436 876
rect 4404 845 4405 875
rect 4405 845 4435 875
rect 4435 845 4436 875
rect 4404 844 4436 845
rect 4404 764 4436 796
rect 4404 684 4436 716
rect 4404 635 4436 636
rect 4404 605 4405 635
rect 4405 605 4435 635
rect 4435 605 4436 635
rect 4404 604 4436 605
rect 4404 555 4436 556
rect 4404 525 4405 555
rect 4405 525 4435 555
rect 4435 525 4436 555
rect 4404 524 4436 525
rect 4404 444 4436 476
rect 4404 395 4436 396
rect 4404 365 4405 395
rect 4405 365 4435 395
rect 4435 365 4436 395
rect 4404 364 4436 365
rect 4404 284 4436 316
rect 4404 235 4436 236
rect 4404 205 4405 235
rect 4405 205 4435 235
rect 4435 205 4436 235
rect 4404 204 4436 205
rect 4404 124 4436 156
rect 4404 75 4436 76
rect 4404 45 4405 75
rect 4405 45 4435 75
rect 4435 45 4436 75
rect 4404 44 4436 45
rect 4404 -5 4436 -4
rect 4404 -35 4405 -5
rect 4405 -35 4435 -5
rect 4435 -35 4436 -5
rect 4404 -36 4436 -35
rect 4404 -85 4436 -84
rect 4404 -115 4405 -85
rect 4405 -115 4435 -85
rect 4435 -115 4436 -85
rect 4404 -116 4436 -115
rect 4484 1035 4516 1036
rect 4484 1005 4485 1035
rect 4485 1005 4515 1035
rect 4515 1005 4516 1035
rect 4484 1004 4516 1005
rect 4484 955 4516 956
rect 4484 925 4485 955
rect 4485 925 4515 955
rect 4515 925 4516 955
rect 4484 924 4516 925
rect 4484 875 4516 876
rect 4484 845 4485 875
rect 4485 845 4515 875
rect 4515 845 4516 875
rect 4484 844 4516 845
rect 4484 764 4516 796
rect 4484 684 4516 716
rect 4484 635 4516 636
rect 4484 605 4485 635
rect 4485 605 4515 635
rect 4515 605 4516 635
rect 4484 604 4516 605
rect 4484 555 4516 556
rect 4484 525 4485 555
rect 4485 525 4515 555
rect 4515 525 4516 555
rect 4484 524 4516 525
rect 4484 444 4516 476
rect 4484 395 4516 396
rect 4484 365 4485 395
rect 4485 365 4515 395
rect 4515 365 4516 395
rect 4484 364 4516 365
rect 4484 284 4516 316
rect 4484 235 4516 236
rect 4484 205 4485 235
rect 4485 205 4515 235
rect 4515 205 4516 235
rect 4484 204 4516 205
rect 4484 124 4516 156
rect 4484 75 4516 76
rect 4484 45 4485 75
rect 4485 45 4515 75
rect 4515 45 4516 75
rect 4484 44 4516 45
rect 4484 -5 4516 -4
rect 4484 -35 4485 -5
rect 4485 -35 4515 -5
rect 4515 -35 4516 -5
rect 4484 -36 4516 -35
rect 4484 -85 4516 -84
rect 4484 -115 4485 -85
rect 4485 -115 4515 -85
rect 4515 -115 4516 -85
rect 4484 -116 4516 -115
rect 4564 1035 4596 1036
rect 4564 1005 4565 1035
rect 4565 1005 4595 1035
rect 4595 1005 4596 1035
rect 4564 1004 4596 1005
rect 4564 955 4596 956
rect 4564 925 4565 955
rect 4565 925 4595 955
rect 4595 925 4596 955
rect 4564 924 4596 925
rect 4564 875 4596 876
rect 4564 845 4565 875
rect 4565 845 4595 875
rect 4595 845 4596 875
rect 4564 844 4596 845
rect 4564 764 4596 796
rect 4564 684 4596 716
rect 4564 635 4596 636
rect 4564 605 4565 635
rect 4565 605 4595 635
rect 4595 605 4596 635
rect 4564 604 4596 605
rect 4564 555 4596 556
rect 4564 525 4565 555
rect 4565 525 4595 555
rect 4595 525 4596 555
rect 4564 524 4596 525
rect 4564 444 4596 476
rect 4564 395 4596 396
rect 4564 365 4565 395
rect 4565 365 4595 395
rect 4595 365 4596 395
rect 4564 364 4596 365
rect 4564 284 4596 316
rect 4564 235 4596 236
rect 4564 205 4565 235
rect 4565 205 4595 235
rect 4595 205 4596 235
rect 4564 204 4596 205
rect 4564 124 4596 156
rect 4564 75 4596 76
rect 4564 45 4565 75
rect 4565 45 4595 75
rect 4595 45 4596 75
rect 4564 44 4596 45
rect 4564 -5 4596 -4
rect 4564 -35 4565 -5
rect 4565 -35 4595 -5
rect 4595 -35 4596 -5
rect 4564 -36 4596 -35
rect 4564 -85 4596 -84
rect 4564 -115 4565 -85
rect 4565 -115 4595 -85
rect 4595 -115 4596 -85
rect 4564 -116 4596 -115
rect 4644 1035 4676 1036
rect 4644 1005 4645 1035
rect 4645 1005 4675 1035
rect 4675 1005 4676 1035
rect 4644 1004 4676 1005
rect 4644 955 4676 956
rect 4644 925 4645 955
rect 4645 925 4675 955
rect 4675 925 4676 955
rect 4644 924 4676 925
rect 4644 875 4676 876
rect 4644 845 4645 875
rect 4645 845 4675 875
rect 4675 845 4676 875
rect 4644 844 4676 845
rect 4644 764 4676 796
rect 4644 684 4676 716
rect 4644 635 4676 636
rect 4644 605 4645 635
rect 4645 605 4675 635
rect 4675 605 4676 635
rect 4644 604 4676 605
rect 4644 555 4676 556
rect 4644 525 4645 555
rect 4645 525 4675 555
rect 4675 525 4676 555
rect 4644 524 4676 525
rect 4644 444 4676 476
rect 4644 395 4676 396
rect 4644 365 4645 395
rect 4645 365 4675 395
rect 4675 365 4676 395
rect 4644 364 4676 365
rect 4644 284 4676 316
rect 4644 235 4676 236
rect 4644 205 4645 235
rect 4645 205 4675 235
rect 4675 205 4676 235
rect 4644 204 4676 205
rect 4644 124 4676 156
rect 4644 75 4676 76
rect 4644 45 4645 75
rect 4645 45 4675 75
rect 4675 45 4676 75
rect 4644 44 4676 45
rect 4644 -5 4676 -4
rect 4644 -35 4645 -5
rect 4645 -35 4675 -5
rect 4675 -35 4676 -5
rect 4644 -36 4676 -35
rect 4644 -85 4676 -84
rect 4644 -115 4645 -85
rect 4645 -115 4675 -85
rect 4675 -115 4676 -85
rect 4644 -116 4676 -115
rect 4724 1035 4756 1036
rect 4724 1005 4725 1035
rect 4725 1005 4755 1035
rect 4755 1005 4756 1035
rect 4724 1004 4756 1005
rect 4724 955 4756 956
rect 4724 925 4725 955
rect 4725 925 4755 955
rect 4755 925 4756 955
rect 4724 924 4756 925
rect 4724 875 4756 876
rect 4724 845 4725 875
rect 4725 845 4755 875
rect 4755 845 4756 875
rect 4724 844 4756 845
rect 4724 764 4756 796
rect 4724 684 4756 716
rect 4724 635 4756 636
rect 4724 605 4725 635
rect 4725 605 4755 635
rect 4755 605 4756 635
rect 4724 604 4756 605
rect 4724 555 4756 556
rect 4724 525 4725 555
rect 4725 525 4755 555
rect 4755 525 4756 555
rect 4724 524 4756 525
rect 4724 444 4756 476
rect 4724 395 4756 396
rect 4724 365 4725 395
rect 4725 365 4755 395
rect 4755 365 4756 395
rect 4724 364 4756 365
rect 4724 284 4756 316
rect 4724 235 4756 236
rect 4724 205 4725 235
rect 4725 205 4755 235
rect 4755 205 4756 235
rect 4724 204 4756 205
rect 4724 124 4756 156
rect 4724 75 4756 76
rect 4724 45 4725 75
rect 4725 45 4755 75
rect 4755 45 4756 75
rect 4724 44 4756 45
rect 4724 -5 4756 -4
rect 4724 -35 4725 -5
rect 4725 -35 4755 -5
rect 4755 -35 4756 -5
rect 4724 -36 4756 -35
rect 4724 -85 4756 -84
rect 4724 -115 4725 -85
rect 4725 -115 4755 -85
rect 4755 -115 4756 -85
rect 4724 -116 4756 -115
rect 4804 1035 4836 1036
rect 4804 1005 4805 1035
rect 4805 1005 4835 1035
rect 4835 1005 4836 1035
rect 4804 1004 4836 1005
rect 4804 955 4836 956
rect 4804 925 4805 955
rect 4805 925 4835 955
rect 4835 925 4836 955
rect 4804 924 4836 925
rect 4804 875 4836 876
rect 4804 845 4805 875
rect 4805 845 4835 875
rect 4835 845 4836 875
rect 4804 844 4836 845
rect 4804 764 4836 796
rect 4804 684 4836 716
rect 4804 635 4836 636
rect 4804 605 4805 635
rect 4805 605 4835 635
rect 4835 605 4836 635
rect 4804 604 4836 605
rect 4804 555 4836 556
rect 4804 525 4805 555
rect 4805 525 4835 555
rect 4835 525 4836 555
rect 4804 524 4836 525
rect 4804 444 4836 476
rect 4804 395 4836 396
rect 4804 365 4805 395
rect 4805 365 4835 395
rect 4835 365 4836 395
rect 4804 364 4836 365
rect 4804 284 4836 316
rect 4804 235 4836 236
rect 4804 205 4805 235
rect 4805 205 4835 235
rect 4835 205 4836 235
rect 4804 204 4836 205
rect 4804 124 4836 156
rect 4804 75 4836 76
rect 4804 45 4805 75
rect 4805 45 4835 75
rect 4835 45 4836 75
rect 4804 44 4836 45
rect 4804 -5 4836 -4
rect 4804 -35 4805 -5
rect 4805 -35 4835 -5
rect 4835 -35 4836 -5
rect 4804 -36 4836 -35
rect 4804 -85 4836 -84
rect 4804 -115 4805 -85
rect 4805 -115 4835 -85
rect 4835 -115 4836 -85
rect 4804 -116 4836 -115
rect 4884 1035 4916 1036
rect 4884 1005 4885 1035
rect 4885 1005 4915 1035
rect 4915 1005 4916 1035
rect 4884 1004 4916 1005
rect 4884 955 4916 956
rect 4884 925 4885 955
rect 4885 925 4915 955
rect 4915 925 4916 955
rect 4884 924 4916 925
rect 4884 875 4916 876
rect 4884 845 4885 875
rect 4885 845 4915 875
rect 4915 845 4916 875
rect 4884 844 4916 845
rect 4884 764 4916 796
rect 4884 684 4916 716
rect 4884 635 4916 636
rect 4884 605 4885 635
rect 4885 605 4915 635
rect 4915 605 4916 635
rect 4884 604 4916 605
rect 4884 555 4916 556
rect 4884 525 4885 555
rect 4885 525 4915 555
rect 4915 525 4916 555
rect 4884 524 4916 525
rect 4884 444 4916 476
rect 4884 395 4916 396
rect 4884 365 4885 395
rect 4885 365 4915 395
rect 4915 365 4916 395
rect 4884 364 4916 365
rect 4884 284 4916 316
rect 4884 235 4916 236
rect 4884 205 4885 235
rect 4885 205 4915 235
rect 4915 205 4916 235
rect 4884 204 4916 205
rect 4884 124 4916 156
rect 4884 75 4916 76
rect 4884 45 4885 75
rect 4885 45 4915 75
rect 4915 45 4916 75
rect 4884 44 4916 45
rect 4884 -5 4916 -4
rect 4884 -35 4885 -5
rect 4885 -35 4915 -5
rect 4915 -35 4916 -5
rect 4884 -36 4916 -35
rect 4884 -85 4916 -84
rect 4884 -115 4885 -85
rect 4885 -115 4915 -85
rect 4915 -115 4916 -85
rect 4884 -116 4916 -115
rect 4964 1035 4996 1036
rect 4964 1005 4965 1035
rect 4965 1005 4995 1035
rect 4995 1005 4996 1035
rect 4964 1004 4996 1005
rect 4964 955 4996 956
rect 4964 925 4965 955
rect 4965 925 4995 955
rect 4995 925 4996 955
rect 4964 924 4996 925
rect 4964 875 4996 876
rect 4964 845 4965 875
rect 4965 845 4995 875
rect 4995 845 4996 875
rect 4964 844 4996 845
rect 4964 764 4996 796
rect 4964 684 4996 716
rect 4964 635 4996 636
rect 4964 605 4965 635
rect 4965 605 4995 635
rect 4995 605 4996 635
rect 4964 604 4996 605
rect 4964 555 4996 556
rect 4964 525 4965 555
rect 4965 525 4995 555
rect 4995 525 4996 555
rect 4964 524 4996 525
rect 4964 444 4996 476
rect 4964 395 4996 396
rect 4964 365 4965 395
rect 4965 365 4995 395
rect 4995 365 4996 395
rect 4964 364 4996 365
rect 4964 284 4996 316
rect 4964 235 4996 236
rect 4964 205 4965 235
rect 4965 205 4995 235
rect 4995 205 4996 235
rect 4964 204 4996 205
rect 4964 124 4996 156
rect 4964 75 4996 76
rect 4964 45 4965 75
rect 4965 45 4995 75
rect 4995 45 4996 75
rect 4964 44 4996 45
rect 4964 -5 4996 -4
rect 4964 -35 4965 -5
rect 4965 -35 4995 -5
rect 4995 -35 4996 -5
rect 4964 -36 4996 -35
rect 4964 -85 4996 -84
rect 4964 -115 4965 -85
rect 4965 -115 4995 -85
rect 4995 -115 4996 -85
rect 4964 -116 4996 -115
rect 5044 1035 5076 1036
rect 5044 1005 5045 1035
rect 5045 1005 5075 1035
rect 5075 1005 5076 1035
rect 5044 1004 5076 1005
rect 5044 955 5076 956
rect 5044 925 5045 955
rect 5045 925 5075 955
rect 5075 925 5076 955
rect 5044 924 5076 925
rect 5044 875 5076 876
rect 5044 845 5045 875
rect 5045 845 5075 875
rect 5075 845 5076 875
rect 5044 844 5076 845
rect 5044 764 5076 796
rect 5044 684 5076 716
rect 5044 635 5076 636
rect 5044 605 5045 635
rect 5045 605 5075 635
rect 5075 605 5076 635
rect 5044 604 5076 605
rect 5044 555 5076 556
rect 5044 525 5045 555
rect 5045 525 5075 555
rect 5075 525 5076 555
rect 5044 524 5076 525
rect 5044 444 5076 476
rect 5044 395 5076 396
rect 5044 365 5045 395
rect 5045 365 5075 395
rect 5075 365 5076 395
rect 5044 364 5076 365
rect 5044 284 5076 316
rect 5044 235 5076 236
rect 5044 205 5045 235
rect 5045 205 5075 235
rect 5075 205 5076 235
rect 5044 204 5076 205
rect 5044 124 5076 156
rect 5044 75 5076 76
rect 5044 45 5045 75
rect 5045 45 5075 75
rect 5075 45 5076 75
rect 5044 44 5076 45
rect 5044 -5 5076 -4
rect 5044 -35 5045 -5
rect 5045 -35 5075 -5
rect 5075 -35 5076 -5
rect 5044 -36 5076 -35
rect 5044 -85 5076 -84
rect 5044 -115 5045 -85
rect 5045 -115 5075 -85
rect 5075 -115 5076 -85
rect 5044 -116 5076 -115
rect 5124 1035 5156 1036
rect 5124 1005 5125 1035
rect 5125 1005 5155 1035
rect 5155 1005 5156 1035
rect 5124 1004 5156 1005
rect 5124 955 5156 956
rect 5124 925 5125 955
rect 5125 925 5155 955
rect 5155 925 5156 955
rect 5124 924 5156 925
rect 5124 875 5156 876
rect 5124 845 5125 875
rect 5125 845 5155 875
rect 5155 845 5156 875
rect 5124 844 5156 845
rect 5124 764 5156 796
rect 5124 684 5156 716
rect 5124 635 5156 636
rect 5124 605 5125 635
rect 5125 605 5155 635
rect 5155 605 5156 635
rect 5124 604 5156 605
rect 5124 555 5156 556
rect 5124 525 5125 555
rect 5125 525 5155 555
rect 5155 525 5156 555
rect 5124 524 5156 525
rect 5124 444 5156 476
rect 5124 395 5156 396
rect 5124 365 5125 395
rect 5125 365 5155 395
rect 5155 365 5156 395
rect 5124 364 5156 365
rect 5124 284 5156 316
rect 5124 235 5156 236
rect 5124 205 5125 235
rect 5125 205 5155 235
rect 5155 205 5156 235
rect 5124 204 5156 205
rect 5124 124 5156 156
rect 5124 75 5156 76
rect 5124 45 5125 75
rect 5125 45 5155 75
rect 5155 45 5156 75
rect 5124 44 5156 45
rect 5124 -5 5156 -4
rect 5124 -35 5125 -5
rect 5125 -35 5155 -5
rect 5155 -35 5156 -5
rect 5124 -36 5156 -35
rect 5124 -85 5156 -84
rect 5124 -115 5125 -85
rect 5125 -115 5155 -85
rect 5155 -115 5156 -85
rect 5124 -116 5156 -115
rect 5204 1035 5236 1036
rect 5204 1005 5205 1035
rect 5205 1005 5235 1035
rect 5235 1005 5236 1035
rect 5204 1004 5236 1005
rect 5204 955 5236 956
rect 5204 925 5205 955
rect 5205 925 5235 955
rect 5235 925 5236 955
rect 5204 924 5236 925
rect 5204 875 5236 876
rect 5204 845 5205 875
rect 5205 845 5235 875
rect 5235 845 5236 875
rect 5204 844 5236 845
rect 5204 764 5236 796
rect 5204 684 5236 716
rect 5204 635 5236 636
rect 5204 605 5205 635
rect 5205 605 5235 635
rect 5235 605 5236 635
rect 5204 604 5236 605
rect 5204 555 5236 556
rect 5204 525 5205 555
rect 5205 525 5235 555
rect 5235 525 5236 555
rect 5204 524 5236 525
rect 5204 444 5236 476
rect 5204 395 5236 396
rect 5204 365 5205 395
rect 5205 365 5235 395
rect 5235 365 5236 395
rect 5204 364 5236 365
rect 5204 284 5236 316
rect 5204 235 5236 236
rect 5204 205 5205 235
rect 5205 205 5235 235
rect 5235 205 5236 235
rect 5204 204 5236 205
rect 5204 124 5236 156
rect 5204 75 5236 76
rect 5204 45 5205 75
rect 5205 45 5235 75
rect 5235 45 5236 75
rect 5204 44 5236 45
rect 5204 -5 5236 -4
rect 5204 -35 5205 -5
rect 5205 -35 5235 -5
rect 5235 -35 5236 -5
rect 5204 -36 5236 -35
rect 5204 -85 5236 -84
rect 5204 -115 5205 -85
rect 5205 -115 5235 -85
rect 5235 -115 5236 -85
rect 5204 -116 5236 -115
rect 5284 1035 5316 1036
rect 5284 1005 5285 1035
rect 5285 1005 5315 1035
rect 5315 1005 5316 1035
rect 5284 1004 5316 1005
rect 5284 955 5316 956
rect 5284 925 5285 955
rect 5285 925 5315 955
rect 5315 925 5316 955
rect 5284 924 5316 925
rect 5284 875 5316 876
rect 5284 845 5285 875
rect 5285 845 5315 875
rect 5315 845 5316 875
rect 5284 844 5316 845
rect 5284 764 5316 796
rect 5284 684 5316 716
rect 5284 635 5316 636
rect 5284 605 5285 635
rect 5285 605 5315 635
rect 5315 605 5316 635
rect 5284 604 5316 605
rect 5284 555 5316 556
rect 5284 525 5285 555
rect 5285 525 5315 555
rect 5315 525 5316 555
rect 5284 524 5316 525
rect 5284 444 5316 476
rect 5284 395 5316 396
rect 5284 365 5285 395
rect 5285 365 5315 395
rect 5315 365 5316 395
rect 5284 364 5316 365
rect 5284 284 5316 316
rect 5284 235 5316 236
rect 5284 205 5285 235
rect 5285 205 5315 235
rect 5315 205 5316 235
rect 5284 204 5316 205
rect 5284 124 5316 156
rect 5284 75 5316 76
rect 5284 45 5285 75
rect 5285 45 5315 75
rect 5315 45 5316 75
rect 5284 44 5316 45
rect 5284 -5 5316 -4
rect 5284 -35 5285 -5
rect 5285 -35 5315 -5
rect 5315 -35 5316 -5
rect 5284 -36 5316 -35
rect 5284 -85 5316 -84
rect 5284 -115 5285 -85
rect 5285 -115 5315 -85
rect 5315 -115 5316 -85
rect 5284 -116 5316 -115
rect 5364 1035 5396 1036
rect 5364 1005 5365 1035
rect 5365 1005 5395 1035
rect 5395 1005 5396 1035
rect 5364 1004 5396 1005
rect 5364 955 5396 956
rect 5364 925 5365 955
rect 5365 925 5395 955
rect 5395 925 5396 955
rect 5364 924 5396 925
rect 5364 875 5396 876
rect 5364 845 5365 875
rect 5365 845 5395 875
rect 5395 845 5396 875
rect 5364 844 5396 845
rect 5364 764 5396 796
rect 5364 684 5396 716
rect 5364 635 5396 636
rect 5364 605 5365 635
rect 5365 605 5395 635
rect 5395 605 5396 635
rect 5364 604 5396 605
rect 5364 555 5396 556
rect 5364 525 5365 555
rect 5365 525 5395 555
rect 5395 525 5396 555
rect 5364 524 5396 525
rect 5364 444 5396 476
rect 5364 395 5396 396
rect 5364 365 5365 395
rect 5365 365 5395 395
rect 5395 365 5396 395
rect 5364 364 5396 365
rect 5364 284 5396 316
rect 5364 235 5396 236
rect 5364 205 5365 235
rect 5365 205 5395 235
rect 5395 205 5396 235
rect 5364 204 5396 205
rect 5364 124 5396 156
rect 5364 75 5396 76
rect 5364 45 5365 75
rect 5365 45 5395 75
rect 5395 45 5396 75
rect 5364 44 5396 45
rect 5364 -5 5396 -4
rect 5364 -35 5365 -5
rect 5365 -35 5395 -5
rect 5395 -35 5396 -5
rect 5364 -36 5396 -35
rect 5364 -85 5396 -84
rect 5364 -115 5365 -85
rect 5365 -115 5395 -85
rect 5395 -115 5396 -85
rect 5364 -116 5396 -115
rect 5444 1035 5476 1036
rect 5444 1005 5445 1035
rect 5445 1005 5475 1035
rect 5475 1005 5476 1035
rect 5444 1004 5476 1005
rect 5444 955 5476 956
rect 5444 925 5445 955
rect 5445 925 5475 955
rect 5475 925 5476 955
rect 5444 924 5476 925
rect 5444 875 5476 876
rect 5444 845 5445 875
rect 5445 845 5475 875
rect 5475 845 5476 875
rect 5444 844 5476 845
rect 5444 764 5476 796
rect 5444 684 5476 716
rect 5444 635 5476 636
rect 5444 605 5445 635
rect 5445 605 5475 635
rect 5475 605 5476 635
rect 5444 604 5476 605
rect 5444 555 5476 556
rect 5444 525 5445 555
rect 5445 525 5475 555
rect 5475 525 5476 555
rect 5444 524 5476 525
rect 5444 444 5476 476
rect 5444 395 5476 396
rect 5444 365 5445 395
rect 5445 365 5475 395
rect 5475 365 5476 395
rect 5444 364 5476 365
rect 5444 284 5476 316
rect 5444 235 5476 236
rect 5444 205 5445 235
rect 5445 205 5475 235
rect 5475 205 5476 235
rect 5444 204 5476 205
rect 5444 124 5476 156
rect 5444 75 5476 76
rect 5444 45 5445 75
rect 5445 45 5475 75
rect 5475 45 5476 75
rect 5444 44 5476 45
rect 5444 -5 5476 -4
rect 5444 -35 5445 -5
rect 5445 -35 5475 -5
rect 5475 -35 5476 -5
rect 5444 -36 5476 -35
rect 5444 -85 5476 -84
rect 5444 -115 5445 -85
rect 5445 -115 5475 -85
rect 5475 -115 5476 -85
rect 5444 -116 5476 -115
rect 5524 1035 5556 1036
rect 5524 1005 5525 1035
rect 5525 1005 5555 1035
rect 5555 1005 5556 1035
rect 5524 1004 5556 1005
rect 5524 955 5556 956
rect 5524 925 5525 955
rect 5525 925 5555 955
rect 5555 925 5556 955
rect 5524 924 5556 925
rect 5524 875 5556 876
rect 5524 845 5525 875
rect 5525 845 5555 875
rect 5555 845 5556 875
rect 5524 844 5556 845
rect 5524 764 5556 796
rect 5524 684 5556 716
rect 5524 635 5556 636
rect 5524 605 5525 635
rect 5525 605 5555 635
rect 5555 605 5556 635
rect 5524 604 5556 605
rect 5524 555 5556 556
rect 5524 525 5525 555
rect 5525 525 5555 555
rect 5555 525 5556 555
rect 5524 524 5556 525
rect 5524 444 5556 476
rect 5524 395 5556 396
rect 5524 365 5525 395
rect 5525 365 5555 395
rect 5555 365 5556 395
rect 5524 364 5556 365
rect 5524 284 5556 316
rect 5524 235 5556 236
rect 5524 205 5525 235
rect 5525 205 5555 235
rect 5555 205 5556 235
rect 5524 204 5556 205
rect 5524 124 5556 156
rect 5524 75 5556 76
rect 5524 45 5525 75
rect 5525 45 5555 75
rect 5555 45 5556 75
rect 5524 44 5556 45
rect 5524 -5 5556 -4
rect 5524 -35 5525 -5
rect 5525 -35 5555 -5
rect 5555 -35 5556 -5
rect 5524 -36 5556 -35
rect 5524 -85 5556 -84
rect 5524 -115 5525 -85
rect 5525 -115 5555 -85
rect 5555 -115 5556 -85
rect 5524 -116 5556 -115
rect 5604 1035 5636 1036
rect 5604 1005 5605 1035
rect 5605 1005 5635 1035
rect 5635 1005 5636 1035
rect 5604 1004 5636 1005
rect 5604 955 5636 956
rect 5604 925 5605 955
rect 5605 925 5635 955
rect 5635 925 5636 955
rect 5604 924 5636 925
rect 5604 875 5636 876
rect 5604 845 5605 875
rect 5605 845 5635 875
rect 5635 845 5636 875
rect 5604 844 5636 845
rect 5604 764 5636 796
rect 5604 684 5636 716
rect 5604 635 5636 636
rect 5604 605 5605 635
rect 5605 605 5635 635
rect 5635 605 5636 635
rect 5604 604 5636 605
rect 5604 555 5636 556
rect 5604 525 5605 555
rect 5605 525 5635 555
rect 5635 525 5636 555
rect 5604 524 5636 525
rect 5604 444 5636 476
rect 5604 395 5636 396
rect 5604 365 5605 395
rect 5605 365 5635 395
rect 5635 365 5636 395
rect 5604 364 5636 365
rect 5604 284 5636 316
rect 5604 235 5636 236
rect 5604 205 5605 235
rect 5605 205 5635 235
rect 5635 205 5636 235
rect 5604 204 5636 205
rect 5604 124 5636 156
rect 5604 75 5636 76
rect 5604 45 5605 75
rect 5605 45 5635 75
rect 5635 45 5636 75
rect 5604 44 5636 45
rect 5604 -5 5636 -4
rect 5604 -35 5605 -5
rect 5605 -35 5635 -5
rect 5635 -35 5636 -5
rect 5604 -36 5636 -35
rect 5604 -85 5636 -84
rect 5604 -115 5605 -85
rect 5605 -115 5635 -85
rect 5635 -115 5636 -85
rect 5604 -116 5636 -115
rect 5684 1035 5716 1036
rect 5684 1005 5685 1035
rect 5685 1005 5715 1035
rect 5715 1005 5716 1035
rect 5684 1004 5716 1005
rect 5684 955 5716 956
rect 5684 925 5685 955
rect 5685 925 5715 955
rect 5715 925 5716 955
rect 5684 924 5716 925
rect 5684 875 5716 876
rect 5684 845 5685 875
rect 5685 845 5715 875
rect 5715 845 5716 875
rect 5684 844 5716 845
rect 5684 764 5716 796
rect 5684 684 5716 716
rect 5684 635 5716 636
rect 5684 605 5685 635
rect 5685 605 5715 635
rect 5715 605 5716 635
rect 5684 604 5716 605
rect 5684 555 5716 556
rect 5684 525 5685 555
rect 5685 525 5715 555
rect 5715 525 5716 555
rect 5684 524 5716 525
rect 5684 444 5716 476
rect 5684 395 5716 396
rect 5684 365 5685 395
rect 5685 365 5715 395
rect 5715 365 5716 395
rect 5684 364 5716 365
rect 5684 284 5716 316
rect 5684 235 5716 236
rect 5684 205 5685 235
rect 5685 205 5715 235
rect 5715 205 5716 235
rect 5684 204 5716 205
rect 5684 124 5716 156
rect 5684 75 5716 76
rect 5684 45 5685 75
rect 5685 45 5715 75
rect 5715 45 5716 75
rect 5684 44 5716 45
rect 5684 -5 5716 -4
rect 5684 -35 5685 -5
rect 5685 -35 5715 -5
rect 5715 -35 5716 -5
rect 5684 -36 5716 -35
rect 5684 -85 5716 -84
rect 5684 -115 5685 -85
rect 5685 -115 5715 -85
rect 5715 -115 5716 -85
rect 5684 -116 5716 -115
rect 5764 1035 5796 1036
rect 5764 1005 5765 1035
rect 5765 1005 5795 1035
rect 5795 1005 5796 1035
rect 5764 1004 5796 1005
rect 5764 955 5796 956
rect 5764 925 5765 955
rect 5765 925 5795 955
rect 5795 925 5796 955
rect 5764 924 5796 925
rect 5764 875 5796 876
rect 5764 845 5765 875
rect 5765 845 5795 875
rect 5795 845 5796 875
rect 5764 844 5796 845
rect 5764 764 5796 796
rect 5764 684 5796 716
rect 5764 635 5796 636
rect 5764 605 5765 635
rect 5765 605 5795 635
rect 5795 605 5796 635
rect 5764 604 5796 605
rect 5764 555 5796 556
rect 5764 525 5765 555
rect 5765 525 5795 555
rect 5795 525 5796 555
rect 5764 524 5796 525
rect 5764 444 5796 476
rect 5764 395 5796 396
rect 5764 365 5765 395
rect 5765 365 5795 395
rect 5795 365 5796 395
rect 5764 364 5796 365
rect 5764 284 5796 316
rect 5764 235 5796 236
rect 5764 205 5765 235
rect 5765 205 5795 235
rect 5795 205 5796 235
rect 5764 204 5796 205
rect 5764 124 5796 156
rect 5764 75 5796 76
rect 5764 45 5765 75
rect 5765 45 5795 75
rect 5795 45 5796 75
rect 5764 44 5796 45
rect 5764 -5 5796 -4
rect 5764 -35 5765 -5
rect 5765 -35 5795 -5
rect 5795 -35 5796 -5
rect 5764 -36 5796 -35
rect 5764 -85 5796 -84
rect 5764 -115 5765 -85
rect 5765 -115 5795 -85
rect 5795 -115 5796 -85
rect 5764 -116 5796 -115
rect 5844 1035 5876 1036
rect 5844 1005 5845 1035
rect 5845 1005 5875 1035
rect 5875 1005 5876 1035
rect 5844 1004 5876 1005
rect 5844 955 5876 956
rect 5844 925 5845 955
rect 5845 925 5875 955
rect 5875 925 5876 955
rect 5844 924 5876 925
rect 5844 875 5876 876
rect 5844 845 5845 875
rect 5845 845 5875 875
rect 5875 845 5876 875
rect 5844 844 5876 845
rect 5844 764 5876 796
rect 5844 684 5876 716
rect 5844 635 5876 636
rect 5844 605 5845 635
rect 5845 605 5875 635
rect 5875 605 5876 635
rect 5844 604 5876 605
rect 5844 555 5876 556
rect 5844 525 5845 555
rect 5845 525 5875 555
rect 5875 525 5876 555
rect 5844 524 5876 525
rect 5844 444 5876 476
rect 5844 395 5876 396
rect 5844 365 5845 395
rect 5845 365 5875 395
rect 5875 365 5876 395
rect 5844 364 5876 365
rect 5844 284 5876 316
rect 5844 235 5876 236
rect 5844 205 5845 235
rect 5845 205 5875 235
rect 5875 205 5876 235
rect 5844 204 5876 205
rect 5844 124 5876 156
rect 5844 75 5876 76
rect 5844 45 5845 75
rect 5845 45 5875 75
rect 5875 45 5876 75
rect 5844 44 5876 45
rect 5844 -5 5876 -4
rect 5844 -35 5845 -5
rect 5845 -35 5875 -5
rect 5875 -35 5876 -5
rect 5844 -36 5876 -35
rect 5844 -85 5876 -84
rect 5844 -115 5845 -85
rect 5845 -115 5875 -85
rect 5875 -115 5876 -85
rect 5844 -116 5876 -115
rect 5924 1035 5956 1036
rect 5924 1005 5925 1035
rect 5925 1005 5955 1035
rect 5955 1005 5956 1035
rect 5924 1004 5956 1005
rect 5924 955 5956 956
rect 5924 925 5925 955
rect 5925 925 5955 955
rect 5955 925 5956 955
rect 5924 924 5956 925
rect 5924 875 5956 876
rect 5924 845 5925 875
rect 5925 845 5955 875
rect 5955 845 5956 875
rect 5924 844 5956 845
rect 5924 764 5956 796
rect 5924 684 5956 716
rect 5924 635 5956 636
rect 5924 605 5925 635
rect 5925 605 5955 635
rect 5955 605 5956 635
rect 5924 604 5956 605
rect 5924 555 5956 556
rect 5924 525 5925 555
rect 5925 525 5955 555
rect 5955 525 5956 555
rect 5924 524 5956 525
rect 5924 444 5956 476
rect 5924 395 5956 396
rect 5924 365 5925 395
rect 5925 365 5955 395
rect 5955 365 5956 395
rect 5924 364 5956 365
rect 5924 284 5956 316
rect 5924 235 5956 236
rect 5924 205 5925 235
rect 5925 205 5955 235
rect 5955 205 5956 235
rect 5924 204 5956 205
rect 5924 124 5956 156
rect 5924 75 5956 76
rect 5924 45 5925 75
rect 5925 45 5955 75
rect 5955 45 5956 75
rect 5924 44 5956 45
rect 5924 -5 5956 -4
rect 5924 -35 5925 -5
rect 5925 -35 5955 -5
rect 5955 -35 5956 -5
rect 5924 -36 5956 -35
rect 5924 -85 5956 -84
rect 5924 -115 5925 -85
rect 5925 -115 5955 -85
rect 5955 -115 5956 -85
rect 5924 -116 5956 -115
rect 6004 1035 6036 1036
rect 6004 1005 6005 1035
rect 6005 1005 6035 1035
rect 6035 1005 6036 1035
rect 6004 1004 6036 1005
rect 6004 955 6036 956
rect 6004 925 6005 955
rect 6005 925 6035 955
rect 6035 925 6036 955
rect 6004 924 6036 925
rect 6004 875 6036 876
rect 6004 845 6005 875
rect 6005 845 6035 875
rect 6035 845 6036 875
rect 6004 844 6036 845
rect 6004 764 6036 796
rect 6004 684 6036 716
rect 6004 635 6036 636
rect 6004 605 6005 635
rect 6005 605 6035 635
rect 6035 605 6036 635
rect 6004 604 6036 605
rect 6004 555 6036 556
rect 6004 525 6005 555
rect 6005 525 6035 555
rect 6035 525 6036 555
rect 6004 524 6036 525
rect 6004 444 6036 476
rect 6004 395 6036 396
rect 6004 365 6005 395
rect 6005 365 6035 395
rect 6035 365 6036 395
rect 6004 364 6036 365
rect 6004 284 6036 316
rect 6004 235 6036 236
rect 6004 205 6005 235
rect 6005 205 6035 235
rect 6035 205 6036 235
rect 6004 204 6036 205
rect 6004 124 6036 156
rect 6004 75 6036 76
rect 6004 45 6005 75
rect 6005 45 6035 75
rect 6035 45 6036 75
rect 6004 44 6036 45
rect 6004 -5 6036 -4
rect 6004 -35 6005 -5
rect 6005 -35 6035 -5
rect 6035 -35 6036 -5
rect 6004 -36 6036 -35
rect 6004 -85 6036 -84
rect 6004 -115 6005 -85
rect 6005 -115 6035 -85
rect 6035 -115 6036 -85
rect 6004 -116 6036 -115
rect 6084 1035 6116 1036
rect 6084 1005 6085 1035
rect 6085 1005 6115 1035
rect 6115 1005 6116 1035
rect 6084 1004 6116 1005
rect 6084 955 6116 956
rect 6084 925 6085 955
rect 6085 925 6115 955
rect 6115 925 6116 955
rect 6084 924 6116 925
rect 6084 875 6116 876
rect 6084 845 6085 875
rect 6085 845 6115 875
rect 6115 845 6116 875
rect 6084 844 6116 845
rect 6084 764 6116 796
rect 6084 684 6116 716
rect 6084 635 6116 636
rect 6084 605 6085 635
rect 6085 605 6115 635
rect 6115 605 6116 635
rect 6084 604 6116 605
rect 6084 555 6116 556
rect 6084 525 6085 555
rect 6085 525 6115 555
rect 6115 525 6116 555
rect 6084 524 6116 525
rect 6084 444 6116 476
rect 6084 395 6116 396
rect 6084 365 6085 395
rect 6085 365 6115 395
rect 6115 365 6116 395
rect 6084 364 6116 365
rect 6084 284 6116 316
rect 6084 235 6116 236
rect 6084 205 6085 235
rect 6085 205 6115 235
rect 6115 205 6116 235
rect 6084 204 6116 205
rect 6084 124 6116 156
rect 6084 75 6116 76
rect 6084 45 6085 75
rect 6085 45 6115 75
rect 6115 45 6116 75
rect 6084 44 6116 45
rect 6084 -5 6116 -4
rect 6084 -35 6085 -5
rect 6085 -35 6115 -5
rect 6115 -35 6116 -5
rect 6084 -36 6116 -35
rect 6084 -85 6116 -84
rect 6084 -115 6085 -85
rect 6085 -115 6115 -85
rect 6115 -115 6116 -85
rect 6084 -116 6116 -115
rect 6164 1035 6196 1036
rect 6164 1005 6165 1035
rect 6165 1005 6195 1035
rect 6195 1005 6196 1035
rect 6164 1004 6196 1005
rect 6164 955 6196 956
rect 6164 925 6165 955
rect 6165 925 6195 955
rect 6195 925 6196 955
rect 6164 924 6196 925
rect 6164 875 6196 876
rect 6164 845 6165 875
rect 6165 845 6195 875
rect 6195 845 6196 875
rect 6164 844 6196 845
rect 6164 764 6196 796
rect 6164 684 6196 716
rect 6164 635 6196 636
rect 6164 605 6165 635
rect 6165 605 6195 635
rect 6195 605 6196 635
rect 6164 604 6196 605
rect 6164 555 6196 556
rect 6164 525 6165 555
rect 6165 525 6195 555
rect 6195 525 6196 555
rect 6164 524 6196 525
rect 6164 444 6196 476
rect 6164 395 6196 396
rect 6164 365 6165 395
rect 6165 365 6195 395
rect 6195 365 6196 395
rect 6164 364 6196 365
rect 6164 284 6196 316
rect 6164 235 6196 236
rect 6164 205 6165 235
rect 6165 205 6195 235
rect 6195 205 6196 235
rect 6164 204 6196 205
rect 6164 124 6196 156
rect 6164 75 6196 76
rect 6164 45 6165 75
rect 6165 45 6195 75
rect 6195 45 6196 75
rect 6164 44 6196 45
rect 6164 -5 6196 -4
rect 6164 -35 6165 -5
rect 6165 -35 6195 -5
rect 6195 -35 6196 -5
rect 6164 -36 6196 -35
rect 6164 -85 6196 -84
rect 6164 -115 6165 -85
rect 6165 -115 6195 -85
rect 6195 -115 6196 -85
rect 6164 -116 6196 -115
rect 6244 1035 6276 1036
rect 6244 1005 6245 1035
rect 6245 1005 6275 1035
rect 6275 1005 6276 1035
rect 6244 1004 6276 1005
rect 6244 955 6276 956
rect 6244 925 6245 955
rect 6245 925 6275 955
rect 6275 925 6276 955
rect 6244 924 6276 925
rect 6244 875 6276 876
rect 6244 845 6245 875
rect 6245 845 6275 875
rect 6275 845 6276 875
rect 6244 844 6276 845
rect 6244 764 6276 796
rect 6244 684 6276 716
rect 6244 635 6276 636
rect 6244 605 6245 635
rect 6245 605 6275 635
rect 6275 605 6276 635
rect 6244 604 6276 605
rect 6244 555 6276 556
rect 6244 525 6245 555
rect 6245 525 6275 555
rect 6275 525 6276 555
rect 6244 524 6276 525
rect 6244 444 6276 476
rect 6244 395 6276 396
rect 6244 365 6245 395
rect 6245 365 6275 395
rect 6275 365 6276 395
rect 6244 364 6276 365
rect 6244 284 6276 316
rect 6244 235 6276 236
rect 6244 205 6245 235
rect 6245 205 6275 235
rect 6275 205 6276 235
rect 6244 204 6276 205
rect 6244 124 6276 156
rect 6244 75 6276 76
rect 6244 45 6245 75
rect 6245 45 6275 75
rect 6275 45 6276 75
rect 6244 44 6276 45
rect 6244 -5 6276 -4
rect 6244 -35 6245 -5
rect 6245 -35 6275 -5
rect 6275 -35 6276 -5
rect 6244 -36 6276 -35
rect 6244 -85 6276 -84
rect 6244 -115 6245 -85
rect 6245 -115 6275 -85
rect 6275 -115 6276 -85
rect 6244 -116 6276 -115
rect 6324 1035 6356 1036
rect 6324 1005 6325 1035
rect 6325 1005 6355 1035
rect 6355 1005 6356 1035
rect 6324 1004 6356 1005
rect 6324 955 6356 956
rect 6324 925 6325 955
rect 6325 925 6355 955
rect 6355 925 6356 955
rect 6324 924 6356 925
rect 6324 875 6356 876
rect 6324 845 6325 875
rect 6325 845 6355 875
rect 6355 845 6356 875
rect 6324 844 6356 845
rect 6324 764 6356 796
rect 6324 684 6356 716
rect 6324 635 6356 636
rect 6324 605 6325 635
rect 6325 605 6355 635
rect 6355 605 6356 635
rect 6324 604 6356 605
rect 6324 555 6356 556
rect 6324 525 6325 555
rect 6325 525 6355 555
rect 6355 525 6356 555
rect 6324 524 6356 525
rect 6324 444 6356 476
rect 6324 395 6356 396
rect 6324 365 6325 395
rect 6325 365 6355 395
rect 6355 365 6356 395
rect 6324 364 6356 365
rect 6324 284 6356 316
rect 6324 235 6356 236
rect 6324 205 6325 235
rect 6325 205 6355 235
rect 6355 205 6356 235
rect 6324 204 6356 205
rect 6324 124 6356 156
rect 6324 75 6356 76
rect 6324 45 6325 75
rect 6325 45 6355 75
rect 6355 45 6356 75
rect 6324 44 6356 45
rect 6324 -5 6356 -4
rect 6324 -35 6325 -5
rect 6325 -35 6355 -5
rect 6355 -35 6356 -5
rect 6324 -36 6356 -35
rect 6324 -85 6356 -84
rect 6324 -115 6325 -85
rect 6325 -115 6355 -85
rect 6355 -115 6356 -85
rect 6324 -116 6356 -115
rect 6404 1035 6436 1036
rect 6404 1005 6405 1035
rect 6405 1005 6435 1035
rect 6435 1005 6436 1035
rect 6404 1004 6436 1005
rect 6404 955 6436 956
rect 6404 925 6405 955
rect 6405 925 6435 955
rect 6435 925 6436 955
rect 6404 924 6436 925
rect 6404 875 6436 876
rect 6404 845 6405 875
rect 6405 845 6435 875
rect 6435 845 6436 875
rect 6404 844 6436 845
rect 6404 764 6436 796
rect 6404 684 6436 716
rect 6404 635 6436 636
rect 6404 605 6405 635
rect 6405 605 6435 635
rect 6435 605 6436 635
rect 6404 604 6436 605
rect 6404 555 6436 556
rect 6404 525 6405 555
rect 6405 525 6435 555
rect 6435 525 6436 555
rect 6404 524 6436 525
rect 6404 444 6436 476
rect 6404 395 6436 396
rect 6404 365 6405 395
rect 6405 365 6435 395
rect 6435 365 6436 395
rect 6404 364 6436 365
rect 6404 284 6436 316
rect 6404 235 6436 236
rect 6404 205 6405 235
rect 6405 205 6435 235
rect 6435 205 6436 235
rect 6404 204 6436 205
rect 6404 124 6436 156
rect 6404 75 6436 76
rect 6404 45 6405 75
rect 6405 45 6435 75
rect 6435 45 6436 75
rect 6404 44 6436 45
rect 6404 -5 6436 -4
rect 6404 -35 6405 -5
rect 6405 -35 6435 -5
rect 6435 -35 6436 -5
rect 6404 -36 6436 -35
rect 6404 -85 6436 -84
rect 6404 -115 6405 -85
rect 6405 -115 6435 -85
rect 6435 -115 6436 -85
rect 6404 -116 6436 -115
rect 6484 1035 6516 1036
rect 6484 1005 6485 1035
rect 6485 1005 6515 1035
rect 6515 1005 6516 1035
rect 6484 1004 6516 1005
rect 6484 955 6516 956
rect 6484 925 6485 955
rect 6485 925 6515 955
rect 6515 925 6516 955
rect 6484 924 6516 925
rect 6484 875 6516 876
rect 6484 845 6485 875
rect 6485 845 6515 875
rect 6515 845 6516 875
rect 6484 844 6516 845
rect 6484 764 6516 796
rect 6484 684 6516 716
rect 6484 635 6516 636
rect 6484 605 6485 635
rect 6485 605 6515 635
rect 6515 605 6516 635
rect 6484 604 6516 605
rect 6484 555 6516 556
rect 6484 525 6485 555
rect 6485 525 6515 555
rect 6515 525 6516 555
rect 6484 524 6516 525
rect 6484 444 6516 476
rect 6484 395 6516 396
rect 6484 365 6485 395
rect 6485 365 6515 395
rect 6515 365 6516 395
rect 6484 364 6516 365
rect 6484 284 6516 316
rect 6484 235 6516 236
rect 6484 205 6485 235
rect 6485 205 6515 235
rect 6515 205 6516 235
rect 6484 204 6516 205
rect 6484 124 6516 156
rect 6484 75 6516 76
rect 6484 45 6485 75
rect 6485 45 6515 75
rect 6515 45 6516 75
rect 6484 44 6516 45
rect 6484 -5 6516 -4
rect 6484 -35 6485 -5
rect 6485 -35 6515 -5
rect 6515 -35 6516 -5
rect 6484 -36 6516 -35
rect 6484 -85 6516 -84
rect 6484 -115 6485 -85
rect 6485 -115 6515 -85
rect 6515 -115 6516 -85
rect 6484 -116 6516 -115
rect 6564 1035 6596 1036
rect 6564 1005 6565 1035
rect 6565 1005 6595 1035
rect 6595 1005 6596 1035
rect 6564 1004 6596 1005
rect 6564 955 6596 956
rect 6564 925 6565 955
rect 6565 925 6595 955
rect 6595 925 6596 955
rect 6564 924 6596 925
rect 6564 875 6596 876
rect 6564 845 6565 875
rect 6565 845 6595 875
rect 6595 845 6596 875
rect 6564 844 6596 845
rect 6564 764 6596 796
rect 6564 684 6596 716
rect 6564 635 6596 636
rect 6564 605 6565 635
rect 6565 605 6595 635
rect 6595 605 6596 635
rect 6564 604 6596 605
rect 6564 555 6596 556
rect 6564 525 6565 555
rect 6565 525 6595 555
rect 6595 525 6596 555
rect 6564 524 6596 525
rect 6564 444 6596 476
rect 6564 395 6596 396
rect 6564 365 6565 395
rect 6565 365 6595 395
rect 6595 365 6596 395
rect 6564 364 6596 365
rect 6564 284 6596 316
rect 6564 235 6596 236
rect 6564 205 6565 235
rect 6565 205 6595 235
rect 6595 205 6596 235
rect 6564 204 6596 205
rect 6564 124 6596 156
rect 6564 75 6596 76
rect 6564 45 6565 75
rect 6565 45 6595 75
rect 6595 45 6596 75
rect 6564 44 6596 45
rect 6564 -5 6596 -4
rect 6564 -35 6565 -5
rect 6565 -35 6595 -5
rect 6595 -35 6596 -5
rect 6564 -36 6596 -35
rect 6564 -85 6596 -84
rect 6564 -115 6565 -85
rect 6565 -115 6595 -85
rect 6595 -115 6596 -85
rect 6564 -116 6596 -115
rect 6644 1035 6676 1036
rect 6644 1005 6645 1035
rect 6645 1005 6675 1035
rect 6675 1005 6676 1035
rect 6644 1004 6676 1005
rect 6644 955 6676 956
rect 6644 925 6645 955
rect 6645 925 6675 955
rect 6675 925 6676 955
rect 6644 924 6676 925
rect 6644 875 6676 876
rect 6644 845 6645 875
rect 6645 845 6675 875
rect 6675 845 6676 875
rect 6644 844 6676 845
rect 6644 764 6676 796
rect 6644 684 6676 716
rect 6644 635 6676 636
rect 6644 605 6645 635
rect 6645 605 6675 635
rect 6675 605 6676 635
rect 6644 604 6676 605
rect 6644 555 6676 556
rect 6644 525 6645 555
rect 6645 525 6675 555
rect 6675 525 6676 555
rect 6644 524 6676 525
rect 6644 444 6676 476
rect 6644 395 6676 396
rect 6644 365 6645 395
rect 6645 365 6675 395
rect 6675 365 6676 395
rect 6644 364 6676 365
rect 6644 284 6676 316
rect 6644 235 6676 236
rect 6644 205 6645 235
rect 6645 205 6675 235
rect 6675 205 6676 235
rect 6644 204 6676 205
rect 6644 124 6676 156
rect 6644 75 6676 76
rect 6644 45 6645 75
rect 6645 45 6675 75
rect 6675 45 6676 75
rect 6644 44 6676 45
rect 6644 -5 6676 -4
rect 6644 -35 6645 -5
rect 6645 -35 6675 -5
rect 6675 -35 6676 -5
rect 6644 -36 6676 -35
rect 6644 -85 6676 -84
rect 6644 -115 6645 -85
rect 6645 -115 6675 -85
rect 6675 -115 6676 -85
rect 6644 -116 6676 -115
rect 6724 1035 6756 1036
rect 6724 1005 6725 1035
rect 6725 1005 6755 1035
rect 6755 1005 6756 1035
rect 6724 1004 6756 1005
rect 6724 955 6756 956
rect 6724 925 6725 955
rect 6725 925 6755 955
rect 6755 925 6756 955
rect 6724 924 6756 925
rect 6724 875 6756 876
rect 6724 845 6725 875
rect 6725 845 6755 875
rect 6755 845 6756 875
rect 6724 844 6756 845
rect 6724 764 6756 796
rect 6724 684 6756 716
rect 6724 635 6756 636
rect 6724 605 6725 635
rect 6725 605 6755 635
rect 6755 605 6756 635
rect 6724 604 6756 605
rect 6724 555 6756 556
rect 6724 525 6725 555
rect 6725 525 6755 555
rect 6755 525 6756 555
rect 6724 524 6756 525
rect 6724 444 6756 476
rect 6724 395 6756 396
rect 6724 365 6725 395
rect 6725 365 6755 395
rect 6755 365 6756 395
rect 6724 364 6756 365
rect 6724 284 6756 316
rect 6724 235 6756 236
rect 6724 205 6725 235
rect 6725 205 6755 235
rect 6755 205 6756 235
rect 6724 204 6756 205
rect 6724 124 6756 156
rect 6724 75 6756 76
rect 6724 45 6725 75
rect 6725 45 6755 75
rect 6755 45 6756 75
rect 6724 44 6756 45
rect 6724 -5 6756 -4
rect 6724 -35 6725 -5
rect 6725 -35 6755 -5
rect 6755 -35 6756 -5
rect 6724 -36 6756 -35
rect 6724 -85 6756 -84
rect 6724 -115 6725 -85
rect 6725 -115 6755 -85
rect 6755 -115 6756 -85
rect 6724 -116 6756 -115
rect 6804 1035 6836 1036
rect 6804 1005 6805 1035
rect 6805 1005 6835 1035
rect 6835 1005 6836 1035
rect 6804 1004 6836 1005
rect 6804 955 6836 956
rect 6804 925 6805 955
rect 6805 925 6835 955
rect 6835 925 6836 955
rect 6804 924 6836 925
rect 6804 875 6836 876
rect 6804 845 6805 875
rect 6805 845 6835 875
rect 6835 845 6836 875
rect 6804 844 6836 845
rect 6804 764 6836 796
rect 6804 684 6836 716
rect 6804 635 6836 636
rect 6804 605 6805 635
rect 6805 605 6835 635
rect 6835 605 6836 635
rect 6804 604 6836 605
rect 6804 555 6836 556
rect 6804 525 6805 555
rect 6805 525 6835 555
rect 6835 525 6836 555
rect 6804 524 6836 525
rect 6804 444 6836 476
rect 6804 395 6836 396
rect 6804 365 6805 395
rect 6805 365 6835 395
rect 6835 365 6836 395
rect 6804 364 6836 365
rect 6804 284 6836 316
rect 6804 235 6836 236
rect 6804 205 6805 235
rect 6805 205 6835 235
rect 6835 205 6836 235
rect 6804 204 6836 205
rect 6804 124 6836 156
rect 6804 75 6836 76
rect 6804 45 6805 75
rect 6805 45 6835 75
rect 6835 45 6836 75
rect 6804 44 6836 45
rect 6804 -5 6836 -4
rect 6804 -35 6805 -5
rect 6805 -35 6835 -5
rect 6835 -35 6836 -5
rect 6804 -36 6836 -35
rect 6804 -85 6836 -84
rect 6804 -115 6805 -85
rect 6805 -115 6835 -85
rect 6835 -115 6836 -85
rect 6804 -116 6836 -115
rect 6884 1035 6916 1036
rect 6884 1005 6885 1035
rect 6885 1005 6915 1035
rect 6915 1005 6916 1035
rect 6884 1004 6916 1005
rect 6884 955 6916 956
rect 6884 925 6885 955
rect 6885 925 6915 955
rect 6915 925 6916 955
rect 6884 924 6916 925
rect 6884 875 6916 876
rect 6884 845 6885 875
rect 6885 845 6915 875
rect 6915 845 6916 875
rect 6884 844 6916 845
rect 6884 764 6916 796
rect 6884 684 6916 716
rect 6884 635 6916 636
rect 6884 605 6885 635
rect 6885 605 6915 635
rect 6915 605 6916 635
rect 6884 604 6916 605
rect 6884 555 6916 556
rect 6884 525 6885 555
rect 6885 525 6915 555
rect 6915 525 6916 555
rect 6884 524 6916 525
rect 6884 444 6916 476
rect 6884 395 6916 396
rect 6884 365 6885 395
rect 6885 365 6915 395
rect 6915 365 6916 395
rect 6884 364 6916 365
rect 6884 284 6916 316
rect 6884 235 6916 236
rect 6884 205 6885 235
rect 6885 205 6915 235
rect 6915 205 6916 235
rect 6884 204 6916 205
rect 6884 124 6916 156
rect 6884 75 6916 76
rect 6884 45 6885 75
rect 6885 45 6915 75
rect 6915 45 6916 75
rect 6884 44 6916 45
rect 6884 -5 6916 -4
rect 6884 -35 6885 -5
rect 6885 -35 6915 -5
rect 6915 -35 6916 -5
rect 6884 -36 6916 -35
rect 6884 -85 6916 -84
rect 6884 -115 6885 -85
rect 6885 -115 6915 -85
rect 6915 -115 6916 -85
rect 6884 -116 6916 -115
rect 6964 1035 6996 1036
rect 6964 1005 6965 1035
rect 6965 1005 6995 1035
rect 6995 1005 6996 1035
rect 6964 1004 6996 1005
rect 6964 955 6996 956
rect 6964 925 6965 955
rect 6965 925 6995 955
rect 6995 925 6996 955
rect 6964 924 6996 925
rect 6964 875 6996 876
rect 6964 845 6965 875
rect 6965 845 6995 875
rect 6995 845 6996 875
rect 6964 844 6996 845
rect 6964 764 6996 796
rect 6964 684 6996 716
rect 6964 635 6996 636
rect 6964 605 6965 635
rect 6965 605 6995 635
rect 6995 605 6996 635
rect 6964 604 6996 605
rect 6964 555 6996 556
rect 6964 525 6965 555
rect 6965 525 6995 555
rect 6995 525 6996 555
rect 6964 524 6996 525
rect 6964 444 6996 476
rect 6964 395 6996 396
rect 6964 365 6965 395
rect 6965 365 6995 395
rect 6995 365 6996 395
rect 6964 364 6996 365
rect 6964 284 6996 316
rect 6964 235 6996 236
rect 6964 205 6965 235
rect 6965 205 6995 235
rect 6995 205 6996 235
rect 6964 204 6996 205
rect 6964 124 6996 156
rect 6964 75 6996 76
rect 6964 45 6965 75
rect 6965 45 6995 75
rect 6995 45 6996 75
rect 6964 44 6996 45
rect 6964 -5 6996 -4
rect 6964 -35 6965 -5
rect 6965 -35 6995 -5
rect 6995 -35 6996 -5
rect 6964 -36 6996 -35
rect 6964 -85 6996 -84
rect 6964 -115 6965 -85
rect 6965 -115 6995 -85
rect 6995 -115 6996 -85
rect 6964 -116 6996 -115
rect 7044 1035 7076 1036
rect 7044 1005 7045 1035
rect 7045 1005 7075 1035
rect 7075 1005 7076 1035
rect 7044 1004 7076 1005
rect 7044 955 7076 956
rect 7044 925 7045 955
rect 7045 925 7075 955
rect 7075 925 7076 955
rect 7044 924 7076 925
rect 7044 875 7076 876
rect 7044 845 7045 875
rect 7045 845 7075 875
rect 7075 845 7076 875
rect 7044 844 7076 845
rect 7044 764 7076 796
rect 7044 684 7076 716
rect 7044 635 7076 636
rect 7044 605 7045 635
rect 7045 605 7075 635
rect 7075 605 7076 635
rect 7044 604 7076 605
rect 7044 555 7076 556
rect 7044 525 7045 555
rect 7045 525 7075 555
rect 7075 525 7076 555
rect 7044 524 7076 525
rect 7044 444 7076 476
rect 7044 395 7076 396
rect 7044 365 7045 395
rect 7045 365 7075 395
rect 7075 365 7076 395
rect 7044 364 7076 365
rect 7044 284 7076 316
rect 7044 235 7076 236
rect 7044 205 7045 235
rect 7045 205 7075 235
rect 7075 205 7076 235
rect 7044 204 7076 205
rect 7044 124 7076 156
rect 7044 75 7076 76
rect 7044 45 7045 75
rect 7045 45 7075 75
rect 7075 45 7076 75
rect 7044 44 7076 45
rect 7044 -5 7076 -4
rect 7044 -35 7045 -5
rect 7045 -35 7075 -5
rect 7075 -35 7076 -5
rect 7044 -36 7076 -35
rect 7044 -85 7076 -84
rect 7044 -115 7045 -85
rect 7045 -115 7075 -85
rect 7075 -115 7076 -85
rect 7044 -116 7076 -115
rect 7124 1035 7156 1036
rect 7124 1005 7125 1035
rect 7125 1005 7155 1035
rect 7155 1005 7156 1035
rect 7124 1004 7156 1005
rect 7124 955 7156 956
rect 7124 925 7125 955
rect 7125 925 7155 955
rect 7155 925 7156 955
rect 7124 924 7156 925
rect 7124 875 7156 876
rect 7124 845 7125 875
rect 7125 845 7155 875
rect 7155 845 7156 875
rect 7124 844 7156 845
rect 7124 764 7156 796
rect 7124 684 7156 716
rect 7124 635 7156 636
rect 7124 605 7125 635
rect 7125 605 7155 635
rect 7155 605 7156 635
rect 7124 604 7156 605
rect 7124 555 7156 556
rect 7124 525 7125 555
rect 7125 525 7155 555
rect 7155 525 7156 555
rect 7124 524 7156 525
rect 7124 444 7156 476
rect 7124 395 7156 396
rect 7124 365 7125 395
rect 7125 365 7155 395
rect 7155 365 7156 395
rect 7124 364 7156 365
rect 7124 284 7156 316
rect 7124 235 7156 236
rect 7124 205 7125 235
rect 7125 205 7155 235
rect 7155 205 7156 235
rect 7124 204 7156 205
rect 7124 124 7156 156
rect 7124 75 7156 76
rect 7124 45 7125 75
rect 7125 45 7155 75
rect 7155 45 7156 75
rect 7124 44 7156 45
rect 7124 -5 7156 -4
rect 7124 -35 7125 -5
rect 7125 -35 7155 -5
rect 7155 -35 7156 -5
rect 7124 -36 7156 -35
rect 7124 -85 7156 -84
rect 7124 -115 7125 -85
rect 7125 -115 7155 -85
rect 7155 -115 7156 -85
rect 7124 -116 7156 -115
rect 7204 1035 7236 1036
rect 7204 1005 7205 1035
rect 7205 1005 7235 1035
rect 7235 1005 7236 1035
rect 7204 1004 7236 1005
rect 7204 955 7236 956
rect 7204 925 7205 955
rect 7205 925 7235 955
rect 7235 925 7236 955
rect 7204 924 7236 925
rect 7204 875 7236 876
rect 7204 845 7205 875
rect 7205 845 7235 875
rect 7235 845 7236 875
rect 7204 844 7236 845
rect 7204 764 7236 796
rect 7204 684 7236 716
rect 7204 635 7236 636
rect 7204 605 7205 635
rect 7205 605 7235 635
rect 7235 605 7236 635
rect 7204 604 7236 605
rect 7204 555 7236 556
rect 7204 525 7205 555
rect 7205 525 7235 555
rect 7235 525 7236 555
rect 7204 524 7236 525
rect 7204 444 7236 476
rect 7204 395 7236 396
rect 7204 365 7205 395
rect 7205 365 7235 395
rect 7235 365 7236 395
rect 7204 364 7236 365
rect 7204 284 7236 316
rect 7204 235 7236 236
rect 7204 205 7205 235
rect 7205 205 7235 235
rect 7235 205 7236 235
rect 7204 204 7236 205
rect 7204 124 7236 156
rect 7204 75 7236 76
rect 7204 45 7205 75
rect 7205 45 7235 75
rect 7235 45 7236 75
rect 7204 44 7236 45
rect 7204 -5 7236 -4
rect 7204 -35 7205 -5
rect 7205 -35 7235 -5
rect 7235 -35 7236 -5
rect 7204 -36 7236 -35
rect 7204 -85 7236 -84
rect 7204 -115 7205 -85
rect 7205 -115 7235 -85
rect 7235 -115 7236 -85
rect 7204 -116 7236 -115
rect 7284 1035 7316 1036
rect 7284 1005 7285 1035
rect 7285 1005 7315 1035
rect 7315 1005 7316 1035
rect 7284 1004 7316 1005
rect 7284 955 7316 956
rect 7284 925 7285 955
rect 7285 925 7315 955
rect 7315 925 7316 955
rect 7284 924 7316 925
rect 7284 875 7316 876
rect 7284 845 7285 875
rect 7285 845 7315 875
rect 7315 845 7316 875
rect 7284 844 7316 845
rect 7284 764 7316 796
rect 7284 684 7316 716
rect 7284 635 7316 636
rect 7284 605 7285 635
rect 7285 605 7315 635
rect 7315 605 7316 635
rect 7284 604 7316 605
rect 7284 555 7316 556
rect 7284 525 7285 555
rect 7285 525 7315 555
rect 7315 525 7316 555
rect 7284 524 7316 525
rect 7284 444 7316 476
rect 7284 395 7316 396
rect 7284 365 7285 395
rect 7285 365 7315 395
rect 7315 365 7316 395
rect 7284 364 7316 365
rect 7284 284 7316 316
rect 7284 235 7316 236
rect 7284 205 7285 235
rect 7285 205 7315 235
rect 7315 205 7316 235
rect 7284 204 7316 205
rect 7284 124 7316 156
rect 7284 75 7316 76
rect 7284 45 7285 75
rect 7285 45 7315 75
rect 7315 45 7316 75
rect 7284 44 7316 45
rect 7284 -5 7316 -4
rect 7284 -35 7285 -5
rect 7285 -35 7315 -5
rect 7315 -35 7316 -5
rect 7284 -36 7316 -35
rect 7284 -85 7316 -84
rect 7284 -115 7285 -85
rect 7285 -115 7315 -85
rect 7315 -115 7316 -85
rect 7284 -116 7316 -115
rect 7364 1035 7396 1036
rect 7364 1005 7365 1035
rect 7365 1005 7395 1035
rect 7395 1005 7396 1035
rect 7364 1004 7396 1005
rect 7364 955 7396 956
rect 7364 925 7365 955
rect 7365 925 7395 955
rect 7395 925 7396 955
rect 7364 924 7396 925
rect 7364 875 7396 876
rect 7364 845 7365 875
rect 7365 845 7395 875
rect 7395 845 7396 875
rect 7364 844 7396 845
rect 7364 764 7396 796
rect 7364 684 7396 716
rect 7364 635 7396 636
rect 7364 605 7365 635
rect 7365 605 7395 635
rect 7395 605 7396 635
rect 7364 604 7396 605
rect 7364 555 7396 556
rect 7364 525 7365 555
rect 7365 525 7395 555
rect 7395 525 7396 555
rect 7364 524 7396 525
rect 7364 444 7396 476
rect 7364 395 7396 396
rect 7364 365 7365 395
rect 7365 365 7395 395
rect 7395 365 7396 395
rect 7364 364 7396 365
rect 7364 284 7396 316
rect 7364 235 7396 236
rect 7364 205 7365 235
rect 7365 205 7395 235
rect 7395 205 7396 235
rect 7364 204 7396 205
rect 7364 124 7396 156
rect 7364 75 7396 76
rect 7364 45 7365 75
rect 7365 45 7395 75
rect 7395 45 7396 75
rect 7364 44 7396 45
rect 7364 -5 7396 -4
rect 7364 -35 7365 -5
rect 7365 -35 7395 -5
rect 7395 -35 7396 -5
rect 7364 -36 7396 -35
rect 7364 -85 7396 -84
rect 7364 -115 7365 -85
rect 7365 -115 7395 -85
rect 7395 -115 7396 -85
rect 7364 -116 7396 -115
rect 7444 1035 7476 1036
rect 7444 1005 7445 1035
rect 7445 1005 7475 1035
rect 7475 1005 7476 1035
rect 7444 1004 7476 1005
rect 7444 955 7476 956
rect 7444 925 7445 955
rect 7445 925 7475 955
rect 7475 925 7476 955
rect 7444 924 7476 925
rect 7444 875 7476 876
rect 7444 845 7445 875
rect 7445 845 7475 875
rect 7475 845 7476 875
rect 7444 844 7476 845
rect 7444 764 7476 796
rect 7444 684 7476 716
rect 7444 635 7476 636
rect 7444 605 7445 635
rect 7445 605 7475 635
rect 7475 605 7476 635
rect 7444 604 7476 605
rect 7444 555 7476 556
rect 7444 525 7445 555
rect 7445 525 7475 555
rect 7475 525 7476 555
rect 7444 524 7476 525
rect 7444 444 7476 476
rect 7444 395 7476 396
rect 7444 365 7445 395
rect 7445 365 7475 395
rect 7475 365 7476 395
rect 7444 364 7476 365
rect 7444 284 7476 316
rect 7444 235 7476 236
rect 7444 205 7445 235
rect 7445 205 7475 235
rect 7475 205 7476 235
rect 7444 204 7476 205
rect 7444 124 7476 156
rect 7444 75 7476 76
rect 7444 45 7445 75
rect 7445 45 7475 75
rect 7475 45 7476 75
rect 7444 44 7476 45
rect 7444 -5 7476 -4
rect 7444 -35 7445 -5
rect 7445 -35 7475 -5
rect 7475 -35 7476 -5
rect 7444 -36 7476 -35
rect 7444 -85 7476 -84
rect 7444 -115 7445 -85
rect 7445 -115 7475 -85
rect 7475 -115 7476 -85
rect 7444 -116 7476 -115
rect 7524 1035 7556 1036
rect 7524 1005 7525 1035
rect 7525 1005 7555 1035
rect 7555 1005 7556 1035
rect 7524 1004 7556 1005
rect 7524 955 7556 956
rect 7524 925 7525 955
rect 7525 925 7555 955
rect 7555 925 7556 955
rect 7524 924 7556 925
rect 7524 875 7556 876
rect 7524 845 7525 875
rect 7525 845 7555 875
rect 7555 845 7556 875
rect 7524 844 7556 845
rect 7524 764 7556 796
rect 7524 684 7556 716
rect 7524 635 7556 636
rect 7524 605 7525 635
rect 7525 605 7555 635
rect 7555 605 7556 635
rect 7524 604 7556 605
rect 7524 555 7556 556
rect 7524 525 7525 555
rect 7525 525 7555 555
rect 7555 525 7556 555
rect 7524 524 7556 525
rect 7524 444 7556 476
rect 7524 395 7556 396
rect 7524 365 7525 395
rect 7525 365 7555 395
rect 7555 365 7556 395
rect 7524 364 7556 365
rect 7524 284 7556 316
rect 7524 235 7556 236
rect 7524 205 7525 235
rect 7525 205 7555 235
rect 7555 205 7556 235
rect 7524 204 7556 205
rect 7524 124 7556 156
rect 7524 75 7556 76
rect 7524 45 7525 75
rect 7525 45 7555 75
rect 7555 45 7556 75
rect 7524 44 7556 45
rect 7524 -5 7556 -4
rect 7524 -35 7525 -5
rect 7525 -35 7555 -5
rect 7555 -35 7556 -5
rect 7524 -36 7556 -35
rect 7524 -85 7556 -84
rect 7524 -115 7525 -85
rect 7525 -115 7555 -85
rect 7555 -115 7556 -85
rect 7524 -116 7556 -115
rect 7604 1035 7636 1036
rect 7604 1005 7605 1035
rect 7605 1005 7635 1035
rect 7635 1005 7636 1035
rect 7604 1004 7636 1005
rect 7604 955 7636 956
rect 7604 925 7605 955
rect 7605 925 7635 955
rect 7635 925 7636 955
rect 7604 924 7636 925
rect 7604 875 7636 876
rect 7604 845 7605 875
rect 7605 845 7635 875
rect 7635 845 7636 875
rect 7604 844 7636 845
rect 7604 764 7636 796
rect 7604 684 7636 716
rect 7604 635 7636 636
rect 7604 605 7605 635
rect 7605 605 7635 635
rect 7635 605 7636 635
rect 7604 604 7636 605
rect 7604 555 7636 556
rect 7604 525 7605 555
rect 7605 525 7635 555
rect 7635 525 7636 555
rect 7604 524 7636 525
rect 7604 444 7636 476
rect 7604 395 7636 396
rect 7604 365 7605 395
rect 7605 365 7635 395
rect 7635 365 7636 395
rect 7604 364 7636 365
rect 7604 284 7636 316
rect 7604 235 7636 236
rect 7604 205 7605 235
rect 7605 205 7635 235
rect 7635 205 7636 235
rect 7604 204 7636 205
rect 7604 124 7636 156
rect 7604 75 7636 76
rect 7604 45 7605 75
rect 7605 45 7635 75
rect 7635 45 7636 75
rect 7604 44 7636 45
rect 7604 -5 7636 -4
rect 7604 -35 7605 -5
rect 7605 -35 7635 -5
rect 7635 -35 7636 -5
rect 7604 -36 7636 -35
rect 7604 -85 7636 -84
rect 7604 -115 7605 -85
rect 7605 -115 7635 -85
rect 7635 -115 7636 -85
rect 7604 -116 7636 -115
rect 7684 1035 7716 1036
rect 7684 1005 7685 1035
rect 7685 1005 7715 1035
rect 7715 1005 7716 1035
rect 7684 1004 7716 1005
rect 7684 955 7716 956
rect 7684 925 7685 955
rect 7685 925 7715 955
rect 7715 925 7716 955
rect 7684 924 7716 925
rect 7684 875 7716 876
rect 7684 845 7685 875
rect 7685 845 7715 875
rect 7715 845 7716 875
rect 7684 844 7716 845
rect 7684 764 7716 796
rect 7684 684 7716 716
rect 7684 635 7716 636
rect 7684 605 7685 635
rect 7685 605 7715 635
rect 7715 605 7716 635
rect 7684 604 7716 605
rect 7684 555 7716 556
rect 7684 525 7685 555
rect 7685 525 7715 555
rect 7715 525 7716 555
rect 7684 524 7716 525
rect 7684 444 7716 476
rect 7684 395 7716 396
rect 7684 365 7685 395
rect 7685 365 7715 395
rect 7715 365 7716 395
rect 7684 364 7716 365
rect 7684 284 7716 316
rect 7684 235 7716 236
rect 7684 205 7685 235
rect 7685 205 7715 235
rect 7715 205 7716 235
rect 7684 204 7716 205
rect 7684 124 7716 156
rect 7684 75 7716 76
rect 7684 45 7685 75
rect 7685 45 7715 75
rect 7715 45 7716 75
rect 7684 44 7716 45
rect 7684 -5 7716 -4
rect 7684 -35 7685 -5
rect 7685 -35 7715 -5
rect 7715 -35 7716 -5
rect 7684 -36 7716 -35
rect 7684 -85 7716 -84
rect 7684 -115 7685 -85
rect 7685 -115 7715 -85
rect 7715 -115 7716 -85
rect 7684 -116 7716 -115
rect 7764 1035 7796 1036
rect 7764 1005 7765 1035
rect 7765 1005 7795 1035
rect 7795 1005 7796 1035
rect 7764 1004 7796 1005
rect 7764 955 7796 956
rect 7764 925 7765 955
rect 7765 925 7795 955
rect 7795 925 7796 955
rect 7764 924 7796 925
rect 7764 875 7796 876
rect 7764 845 7765 875
rect 7765 845 7795 875
rect 7795 845 7796 875
rect 7764 844 7796 845
rect 7764 764 7796 796
rect 7764 684 7796 716
rect 7764 635 7796 636
rect 7764 605 7765 635
rect 7765 605 7795 635
rect 7795 605 7796 635
rect 7764 604 7796 605
rect 7764 555 7796 556
rect 7764 525 7765 555
rect 7765 525 7795 555
rect 7795 525 7796 555
rect 7764 524 7796 525
rect 7764 444 7796 476
rect 7764 395 7796 396
rect 7764 365 7765 395
rect 7765 365 7795 395
rect 7795 365 7796 395
rect 7764 364 7796 365
rect 7764 284 7796 316
rect 7764 235 7796 236
rect 7764 205 7765 235
rect 7765 205 7795 235
rect 7795 205 7796 235
rect 7764 204 7796 205
rect 7764 124 7796 156
rect 7764 75 7796 76
rect 7764 45 7765 75
rect 7765 45 7795 75
rect 7795 45 7796 75
rect 7764 44 7796 45
rect 7764 -5 7796 -4
rect 7764 -35 7765 -5
rect 7765 -35 7795 -5
rect 7795 -35 7796 -5
rect 7764 -36 7796 -35
rect 7764 -85 7796 -84
rect 7764 -115 7765 -85
rect 7765 -115 7795 -85
rect 7795 -115 7796 -85
rect 7764 -116 7796 -115
rect 7844 1035 7876 1036
rect 7844 1005 7845 1035
rect 7845 1005 7875 1035
rect 7875 1005 7876 1035
rect 7844 1004 7876 1005
rect 7844 955 7876 956
rect 7844 925 7845 955
rect 7845 925 7875 955
rect 7875 925 7876 955
rect 7844 924 7876 925
rect 7844 875 7876 876
rect 7844 845 7845 875
rect 7845 845 7875 875
rect 7875 845 7876 875
rect 7844 844 7876 845
rect 7844 764 7876 796
rect 7844 684 7876 716
rect 7844 635 7876 636
rect 7844 605 7845 635
rect 7845 605 7875 635
rect 7875 605 7876 635
rect 7844 604 7876 605
rect 7844 555 7876 556
rect 7844 525 7845 555
rect 7845 525 7875 555
rect 7875 525 7876 555
rect 7844 524 7876 525
rect 7844 444 7876 476
rect 7844 395 7876 396
rect 7844 365 7845 395
rect 7845 365 7875 395
rect 7875 365 7876 395
rect 7844 364 7876 365
rect 7844 284 7876 316
rect 7844 235 7876 236
rect 7844 205 7845 235
rect 7845 205 7875 235
rect 7875 205 7876 235
rect 7844 204 7876 205
rect 7844 124 7876 156
rect 7844 75 7876 76
rect 7844 45 7845 75
rect 7845 45 7875 75
rect 7875 45 7876 75
rect 7844 44 7876 45
rect 7844 -5 7876 -4
rect 7844 -35 7845 -5
rect 7845 -35 7875 -5
rect 7875 -35 7876 -5
rect 7844 -36 7876 -35
rect 7844 -85 7876 -84
rect 7844 -115 7845 -85
rect 7845 -115 7875 -85
rect 7875 -115 7876 -85
rect 7844 -116 7876 -115
rect 7924 1035 7956 1036
rect 7924 1005 7925 1035
rect 7925 1005 7955 1035
rect 7955 1005 7956 1035
rect 7924 1004 7956 1005
rect 7924 955 7956 956
rect 7924 925 7925 955
rect 7925 925 7955 955
rect 7955 925 7956 955
rect 7924 924 7956 925
rect 7924 875 7956 876
rect 7924 845 7925 875
rect 7925 845 7955 875
rect 7955 845 7956 875
rect 7924 844 7956 845
rect 7924 764 7956 796
rect 7924 684 7956 716
rect 7924 635 7956 636
rect 7924 605 7925 635
rect 7925 605 7955 635
rect 7955 605 7956 635
rect 7924 604 7956 605
rect 7924 555 7956 556
rect 7924 525 7925 555
rect 7925 525 7955 555
rect 7955 525 7956 555
rect 7924 524 7956 525
rect 7924 444 7956 476
rect 7924 395 7956 396
rect 7924 365 7925 395
rect 7925 365 7955 395
rect 7955 365 7956 395
rect 7924 364 7956 365
rect 7924 284 7956 316
rect 7924 235 7956 236
rect 7924 205 7925 235
rect 7925 205 7955 235
rect 7955 205 7956 235
rect 7924 204 7956 205
rect 7924 124 7956 156
rect 7924 75 7956 76
rect 7924 45 7925 75
rect 7925 45 7955 75
rect 7955 45 7956 75
rect 7924 44 7956 45
rect 7924 -5 7956 -4
rect 7924 -35 7925 -5
rect 7925 -35 7955 -5
rect 7955 -35 7956 -5
rect 7924 -36 7956 -35
rect 7924 -85 7956 -84
rect 7924 -115 7925 -85
rect 7925 -115 7955 -85
rect 7955 -115 7956 -85
rect 7924 -116 7956 -115
rect 8004 1035 8036 1036
rect 8004 1005 8005 1035
rect 8005 1005 8035 1035
rect 8035 1005 8036 1035
rect 8004 1004 8036 1005
rect 8004 955 8036 956
rect 8004 925 8005 955
rect 8005 925 8035 955
rect 8035 925 8036 955
rect 8004 924 8036 925
rect 8004 875 8036 876
rect 8004 845 8005 875
rect 8005 845 8035 875
rect 8035 845 8036 875
rect 8004 844 8036 845
rect 8004 764 8036 796
rect 8004 684 8036 716
rect 8004 635 8036 636
rect 8004 605 8005 635
rect 8005 605 8035 635
rect 8035 605 8036 635
rect 8004 604 8036 605
rect 8004 555 8036 556
rect 8004 525 8005 555
rect 8005 525 8035 555
rect 8035 525 8036 555
rect 8004 524 8036 525
rect 8004 444 8036 476
rect 8004 395 8036 396
rect 8004 365 8005 395
rect 8005 365 8035 395
rect 8035 365 8036 395
rect 8004 364 8036 365
rect 8004 284 8036 316
rect 8004 235 8036 236
rect 8004 205 8005 235
rect 8005 205 8035 235
rect 8035 205 8036 235
rect 8004 204 8036 205
rect 8004 124 8036 156
rect 8004 75 8036 76
rect 8004 45 8005 75
rect 8005 45 8035 75
rect 8035 45 8036 75
rect 8004 44 8036 45
rect 8004 -5 8036 -4
rect 8004 -35 8005 -5
rect 8005 -35 8035 -5
rect 8035 -35 8036 -5
rect 8004 -36 8036 -35
rect 8004 -85 8036 -84
rect 8004 -115 8005 -85
rect 8005 -115 8035 -85
rect 8035 -115 8036 -85
rect 8004 -116 8036 -115
rect 8084 1035 8116 1036
rect 8084 1005 8085 1035
rect 8085 1005 8115 1035
rect 8115 1005 8116 1035
rect 8084 1004 8116 1005
rect 8084 955 8116 956
rect 8084 925 8085 955
rect 8085 925 8115 955
rect 8115 925 8116 955
rect 8084 924 8116 925
rect 8084 875 8116 876
rect 8084 845 8085 875
rect 8085 845 8115 875
rect 8115 845 8116 875
rect 8084 844 8116 845
rect 8084 764 8116 796
rect 8084 684 8116 716
rect 8084 635 8116 636
rect 8084 605 8085 635
rect 8085 605 8115 635
rect 8115 605 8116 635
rect 8084 604 8116 605
rect 8084 555 8116 556
rect 8084 525 8085 555
rect 8085 525 8115 555
rect 8115 525 8116 555
rect 8084 524 8116 525
rect 8084 444 8116 476
rect 8084 395 8116 396
rect 8084 365 8085 395
rect 8085 365 8115 395
rect 8115 365 8116 395
rect 8084 364 8116 365
rect 8084 284 8116 316
rect 8084 235 8116 236
rect 8084 205 8085 235
rect 8085 205 8115 235
rect 8115 205 8116 235
rect 8084 204 8116 205
rect 8084 124 8116 156
rect 8084 75 8116 76
rect 8084 45 8085 75
rect 8085 45 8115 75
rect 8115 45 8116 75
rect 8084 44 8116 45
rect 8084 -5 8116 -4
rect 8084 -35 8085 -5
rect 8085 -35 8115 -5
rect 8115 -35 8116 -5
rect 8084 -36 8116 -35
rect 8084 -85 8116 -84
rect 8084 -115 8085 -85
rect 8085 -115 8115 -85
rect 8115 -115 8116 -85
rect 8084 -116 8116 -115
rect 8164 1035 8196 1036
rect 8164 1005 8165 1035
rect 8165 1005 8195 1035
rect 8195 1005 8196 1035
rect 8164 1004 8196 1005
rect 8164 955 8196 956
rect 8164 925 8165 955
rect 8165 925 8195 955
rect 8195 925 8196 955
rect 8164 924 8196 925
rect 8164 875 8196 876
rect 8164 845 8165 875
rect 8165 845 8195 875
rect 8195 845 8196 875
rect 8164 844 8196 845
rect 8164 764 8196 796
rect 8164 684 8196 716
rect 8164 635 8196 636
rect 8164 605 8165 635
rect 8165 605 8195 635
rect 8195 605 8196 635
rect 8164 604 8196 605
rect 8164 555 8196 556
rect 8164 525 8165 555
rect 8165 525 8195 555
rect 8195 525 8196 555
rect 8164 524 8196 525
rect 8164 444 8196 476
rect 8164 395 8196 396
rect 8164 365 8165 395
rect 8165 365 8195 395
rect 8195 365 8196 395
rect 8164 364 8196 365
rect 8164 284 8196 316
rect 8164 235 8196 236
rect 8164 205 8165 235
rect 8165 205 8195 235
rect 8195 205 8196 235
rect 8164 204 8196 205
rect 8164 124 8196 156
rect 8164 75 8196 76
rect 8164 45 8165 75
rect 8165 45 8195 75
rect 8195 45 8196 75
rect 8164 44 8196 45
rect 8164 -5 8196 -4
rect 8164 -35 8165 -5
rect 8165 -35 8195 -5
rect 8195 -35 8196 -5
rect 8164 -36 8196 -35
rect 8164 -85 8196 -84
rect 8164 -115 8165 -85
rect 8165 -115 8195 -85
rect 8195 -115 8196 -85
rect 8164 -116 8196 -115
rect 8244 1035 8276 1036
rect 8244 1005 8245 1035
rect 8245 1005 8275 1035
rect 8275 1005 8276 1035
rect 8244 1004 8276 1005
rect 8244 955 8276 956
rect 8244 925 8245 955
rect 8245 925 8275 955
rect 8275 925 8276 955
rect 8244 924 8276 925
rect 8244 875 8276 876
rect 8244 845 8245 875
rect 8245 845 8275 875
rect 8275 845 8276 875
rect 8244 844 8276 845
rect 8244 764 8276 796
rect 8244 684 8276 716
rect 8244 635 8276 636
rect 8244 605 8245 635
rect 8245 605 8275 635
rect 8275 605 8276 635
rect 8244 604 8276 605
rect 8244 555 8276 556
rect 8244 525 8245 555
rect 8245 525 8275 555
rect 8275 525 8276 555
rect 8244 524 8276 525
rect 8244 444 8276 476
rect 8244 395 8276 396
rect 8244 365 8245 395
rect 8245 365 8275 395
rect 8275 365 8276 395
rect 8244 364 8276 365
rect 8244 284 8276 316
rect 8244 235 8276 236
rect 8244 205 8245 235
rect 8245 205 8275 235
rect 8275 205 8276 235
rect 8244 204 8276 205
rect 8244 124 8276 156
rect 8244 75 8276 76
rect 8244 45 8245 75
rect 8245 45 8275 75
rect 8275 45 8276 75
rect 8244 44 8276 45
rect 8244 -5 8276 -4
rect 8244 -35 8245 -5
rect 8245 -35 8275 -5
rect 8275 -35 8276 -5
rect 8244 -36 8276 -35
rect 8244 -85 8276 -84
rect 8244 -115 8245 -85
rect 8245 -115 8275 -85
rect 8275 -115 8276 -85
rect 8244 -116 8276 -115
rect 8324 1035 8356 1036
rect 8324 1005 8325 1035
rect 8325 1005 8355 1035
rect 8355 1005 8356 1035
rect 8324 1004 8356 1005
rect 8324 955 8356 956
rect 8324 925 8325 955
rect 8325 925 8355 955
rect 8355 925 8356 955
rect 8324 924 8356 925
rect 8324 875 8356 876
rect 8324 845 8325 875
rect 8325 845 8355 875
rect 8355 845 8356 875
rect 8324 844 8356 845
rect 8324 764 8356 796
rect 8324 684 8356 716
rect 8324 635 8356 636
rect 8324 605 8325 635
rect 8325 605 8355 635
rect 8355 605 8356 635
rect 8324 604 8356 605
rect 8324 555 8356 556
rect 8324 525 8325 555
rect 8325 525 8355 555
rect 8355 525 8356 555
rect 8324 524 8356 525
rect 8324 444 8356 476
rect 8324 395 8356 396
rect 8324 365 8325 395
rect 8325 365 8355 395
rect 8355 365 8356 395
rect 8324 364 8356 365
rect 8324 284 8356 316
rect 8324 235 8356 236
rect 8324 205 8325 235
rect 8325 205 8355 235
rect 8355 205 8356 235
rect 8324 204 8356 205
rect 8324 124 8356 156
rect 8324 75 8356 76
rect 8324 45 8325 75
rect 8325 45 8355 75
rect 8355 45 8356 75
rect 8324 44 8356 45
rect 8324 -5 8356 -4
rect 8324 -35 8325 -5
rect 8325 -35 8355 -5
rect 8355 -35 8356 -5
rect 8324 -36 8356 -35
rect 8324 -85 8356 -84
rect 8324 -115 8325 -85
rect 8325 -115 8355 -85
rect 8355 -115 8356 -85
rect 8324 -116 8356 -115
rect 8404 1035 8436 1036
rect 8404 1005 8405 1035
rect 8405 1005 8435 1035
rect 8435 1005 8436 1035
rect 8404 1004 8436 1005
rect 8404 955 8436 956
rect 8404 925 8405 955
rect 8405 925 8435 955
rect 8435 925 8436 955
rect 8404 924 8436 925
rect 8404 875 8436 876
rect 8404 845 8405 875
rect 8405 845 8435 875
rect 8435 845 8436 875
rect 8404 844 8436 845
rect 8404 764 8436 796
rect 8404 684 8436 716
rect 8404 635 8436 636
rect 8404 605 8405 635
rect 8405 605 8435 635
rect 8435 605 8436 635
rect 8404 604 8436 605
rect 8404 555 8436 556
rect 8404 525 8405 555
rect 8405 525 8435 555
rect 8435 525 8436 555
rect 8404 524 8436 525
rect 8404 444 8436 476
rect 8404 395 8436 396
rect 8404 365 8405 395
rect 8405 365 8435 395
rect 8435 365 8436 395
rect 8404 364 8436 365
rect 8404 284 8436 316
rect 8404 235 8436 236
rect 8404 205 8405 235
rect 8405 205 8435 235
rect 8435 205 8436 235
rect 8404 204 8436 205
rect 8404 124 8436 156
rect 8404 75 8436 76
rect 8404 45 8405 75
rect 8405 45 8435 75
rect 8435 45 8436 75
rect 8404 44 8436 45
rect 8404 -5 8436 -4
rect 8404 -35 8405 -5
rect 8405 -35 8435 -5
rect 8435 -35 8436 -5
rect 8404 -36 8436 -35
rect 8404 -85 8436 -84
rect 8404 -115 8405 -85
rect 8405 -115 8435 -85
rect 8435 -115 8436 -85
rect 8404 -116 8436 -115
rect 8484 1035 8516 1036
rect 8484 1005 8485 1035
rect 8485 1005 8515 1035
rect 8515 1005 8516 1035
rect 8484 1004 8516 1005
rect 8484 955 8516 956
rect 8484 925 8485 955
rect 8485 925 8515 955
rect 8515 925 8516 955
rect 8484 924 8516 925
rect 8484 875 8516 876
rect 8484 845 8485 875
rect 8485 845 8515 875
rect 8515 845 8516 875
rect 8484 844 8516 845
rect 8484 764 8516 796
rect 8484 684 8516 716
rect 8484 635 8516 636
rect 8484 605 8485 635
rect 8485 605 8515 635
rect 8515 605 8516 635
rect 8484 604 8516 605
rect 8484 555 8516 556
rect 8484 525 8485 555
rect 8485 525 8515 555
rect 8515 525 8516 555
rect 8484 524 8516 525
rect 8484 444 8516 476
rect 8484 395 8516 396
rect 8484 365 8485 395
rect 8485 365 8515 395
rect 8515 365 8516 395
rect 8484 364 8516 365
rect 8484 284 8516 316
rect 8484 235 8516 236
rect 8484 205 8485 235
rect 8485 205 8515 235
rect 8515 205 8516 235
rect 8484 204 8516 205
rect 8484 124 8516 156
rect 8484 75 8516 76
rect 8484 45 8485 75
rect 8485 45 8515 75
rect 8515 45 8516 75
rect 8484 44 8516 45
rect 8484 -5 8516 -4
rect 8484 -35 8485 -5
rect 8485 -35 8515 -5
rect 8515 -35 8516 -5
rect 8484 -36 8516 -35
rect 8484 -85 8516 -84
rect 8484 -115 8485 -85
rect 8485 -115 8515 -85
rect 8515 -115 8516 -85
rect 8484 -116 8516 -115
rect 8564 1035 8596 1036
rect 8564 1005 8565 1035
rect 8565 1005 8595 1035
rect 8595 1005 8596 1035
rect 8564 1004 8596 1005
rect 8564 955 8596 956
rect 8564 925 8565 955
rect 8565 925 8595 955
rect 8595 925 8596 955
rect 8564 924 8596 925
rect 8564 875 8596 876
rect 8564 845 8565 875
rect 8565 845 8595 875
rect 8595 845 8596 875
rect 8564 844 8596 845
rect 8564 764 8596 796
rect 8564 684 8596 716
rect 8564 635 8596 636
rect 8564 605 8565 635
rect 8565 605 8595 635
rect 8595 605 8596 635
rect 8564 604 8596 605
rect 8564 555 8596 556
rect 8564 525 8565 555
rect 8565 525 8595 555
rect 8595 525 8596 555
rect 8564 524 8596 525
rect 8564 444 8596 476
rect 8564 395 8596 396
rect 8564 365 8565 395
rect 8565 365 8595 395
rect 8595 365 8596 395
rect 8564 364 8596 365
rect 8564 284 8596 316
rect 8564 235 8596 236
rect 8564 205 8565 235
rect 8565 205 8595 235
rect 8595 205 8596 235
rect 8564 204 8596 205
rect 8564 124 8596 156
rect 8564 75 8596 76
rect 8564 45 8565 75
rect 8565 45 8595 75
rect 8595 45 8596 75
rect 8564 44 8596 45
rect 8564 -5 8596 -4
rect 8564 -35 8565 -5
rect 8565 -35 8595 -5
rect 8595 -35 8596 -5
rect 8564 -36 8596 -35
rect 8564 -85 8596 -84
rect 8564 -115 8565 -85
rect 8565 -115 8595 -85
rect 8595 -115 8596 -85
rect 8564 -116 8596 -115
rect 8644 1035 8676 1036
rect 8644 1005 8645 1035
rect 8645 1005 8675 1035
rect 8675 1005 8676 1035
rect 8644 1004 8676 1005
rect 8644 955 8676 956
rect 8644 925 8645 955
rect 8645 925 8675 955
rect 8675 925 8676 955
rect 8644 924 8676 925
rect 8644 875 8676 876
rect 8644 845 8645 875
rect 8645 845 8675 875
rect 8675 845 8676 875
rect 8644 844 8676 845
rect 8644 764 8676 796
rect 8644 684 8676 716
rect 8644 635 8676 636
rect 8644 605 8645 635
rect 8645 605 8675 635
rect 8675 605 8676 635
rect 8644 604 8676 605
rect 8644 555 8676 556
rect 8644 525 8645 555
rect 8645 525 8675 555
rect 8675 525 8676 555
rect 8644 524 8676 525
rect 8644 444 8676 476
rect 8644 395 8676 396
rect 8644 365 8645 395
rect 8645 365 8675 395
rect 8675 365 8676 395
rect 8644 364 8676 365
rect 8644 284 8676 316
rect 8644 235 8676 236
rect 8644 205 8645 235
rect 8645 205 8675 235
rect 8675 205 8676 235
rect 8644 204 8676 205
rect 8644 124 8676 156
rect 8644 75 8676 76
rect 8644 45 8645 75
rect 8645 45 8675 75
rect 8675 45 8676 75
rect 8644 44 8676 45
rect 8644 -5 8676 -4
rect 8644 -35 8645 -5
rect 8645 -35 8675 -5
rect 8675 -35 8676 -5
rect 8644 -36 8676 -35
rect 8644 -85 8676 -84
rect 8644 -115 8645 -85
rect 8645 -115 8675 -85
rect 8675 -115 8676 -85
rect 8644 -116 8676 -115
rect 8724 1035 8756 1036
rect 8724 1005 8725 1035
rect 8725 1005 8755 1035
rect 8755 1005 8756 1035
rect 8724 1004 8756 1005
rect 8724 955 8756 956
rect 8724 925 8725 955
rect 8725 925 8755 955
rect 8755 925 8756 955
rect 8724 924 8756 925
rect 8724 875 8756 876
rect 8724 845 8725 875
rect 8725 845 8755 875
rect 8755 845 8756 875
rect 8724 844 8756 845
rect 8724 764 8756 796
rect 8724 684 8756 716
rect 8724 635 8756 636
rect 8724 605 8725 635
rect 8725 605 8755 635
rect 8755 605 8756 635
rect 8724 604 8756 605
rect 8724 555 8756 556
rect 8724 525 8725 555
rect 8725 525 8755 555
rect 8755 525 8756 555
rect 8724 524 8756 525
rect 8724 444 8756 476
rect 8724 395 8756 396
rect 8724 365 8725 395
rect 8725 365 8755 395
rect 8755 365 8756 395
rect 8724 364 8756 365
rect 8724 284 8756 316
rect 8724 235 8756 236
rect 8724 205 8725 235
rect 8725 205 8755 235
rect 8755 205 8756 235
rect 8724 204 8756 205
rect 8724 124 8756 156
rect 8724 75 8756 76
rect 8724 45 8725 75
rect 8725 45 8755 75
rect 8755 45 8756 75
rect 8724 44 8756 45
rect 8724 -5 8756 -4
rect 8724 -35 8725 -5
rect 8725 -35 8755 -5
rect 8755 -35 8756 -5
rect 8724 -36 8756 -35
rect 8724 -85 8756 -84
rect 8724 -115 8725 -85
rect 8725 -115 8755 -85
rect 8755 -115 8756 -85
rect 8724 -116 8756 -115
rect 8804 1035 8836 1036
rect 8804 1005 8805 1035
rect 8805 1005 8835 1035
rect 8835 1005 8836 1035
rect 8804 1004 8836 1005
rect 8804 955 8836 956
rect 8804 925 8805 955
rect 8805 925 8835 955
rect 8835 925 8836 955
rect 8804 924 8836 925
rect 8804 875 8836 876
rect 8804 845 8805 875
rect 8805 845 8835 875
rect 8835 845 8836 875
rect 8804 844 8836 845
rect 8804 764 8836 796
rect 8804 684 8836 716
rect 8804 635 8836 636
rect 8804 605 8805 635
rect 8805 605 8835 635
rect 8835 605 8836 635
rect 8804 604 8836 605
rect 8804 555 8836 556
rect 8804 525 8805 555
rect 8805 525 8835 555
rect 8835 525 8836 555
rect 8804 524 8836 525
rect 8804 444 8836 476
rect 8804 395 8836 396
rect 8804 365 8805 395
rect 8805 365 8835 395
rect 8835 365 8836 395
rect 8804 364 8836 365
rect 8804 284 8836 316
rect 8804 235 8836 236
rect 8804 205 8805 235
rect 8805 205 8835 235
rect 8835 205 8836 235
rect 8804 204 8836 205
rect 8804 124 8836 156
rect 8804 75 8836 76
rect 8804 45 8805 75
rect 8805 45 8835 75
rect 8835 45 8836 75
rect 8804 44 8836 45
rect 8804 -5 8836 -4
rect 8804 -35 8805 -5
rect 8805 -35 8835 -5
rect 8835 -35 8836 -5
rect 8804 -36 8836 -35
rect 8804 -85 8836 -84
rect 8804 -115 8805 -85
rect 8805 -115 8835 -85
rect 8835 -115 8836 -85
rect 8804 -116 8836 -115
rect 8884 1035 8916 1036
rect 8884 1005 8885 1035
rect 8885 1005 8915 1035
rect 8915 1005 8916 1035
rect 8884 1004 8916 1005
rect 8884 955 8916 956
rect 8884 925 8885 955
rect 8885 925 8915 955
rect 8915 925 8916 955
rect 8884 924 8916 925
rect 8884 875 8916 876
rect 8884 845 8885 875
rect 8885 845 8915 875
rect 8915 845 8916 875
rect 8884 844 8916 845
rect 8884 764 8916 796
rect 8884 684 8916 716
rect 8884 635 8916 636
rect 8884 605 8885 635
rect 8885 605 8915 635
rect 8915 605 8916 635
rect 8884 604 8916 605
rect 8884 555 8916 556
rect 8884 525 8885 555
rect 8885 525 8915 555
rect 8915 525 8916 555
rect 8884 524 8916 525
rect 8884 444 8916 476
rect 8884 395 8916 396
rect 8884 365 8885 395
rect 8885 365 8915 395
rect 8915 365 8916 395
rect 8884 364 8916 365
rect 8884 284 8916 316
rect 8884 235 8916 236
rect 8884 205 8885 235
rect 8885 205 8915 235
rect 8915 205 8916 235
rect 8884 204 8916 205
rect 8884 124 8916 156
rect 8884 75 8916 76
rect 8884 45 8885 75
rect 8885 45 8915 75
rect 8915 45 8916 75
rect 8884 44 8916 45
rect 8884 -5 8916 -4
rect 8884 -35 8885 -5
rect 8885 -35 8915 -5
rect 8915 -35 8916 -5
rect 8884 -36 8916 -35
rect 8884 -85 8916 -84
rect 8884 -115 8885 -85
rect 8885 -115 8915 -85
rect 8915 -115 8916 -85
rect 8884 -116 8916 -115
rect 8964 1035 8996 1036
rect 8964 1005 8965 1035
rect 8965 1005 8995 1035
rect 8995 1005 8996 1035
rect 8964 1004 8996 1005
rect 8964 955 8996 956
rect 8964 925 8965 955
rect 8965 925 8995 955
rect 8995 925 8996 955
rect 8964 924 8996 925
rect 8964 875 8996 876
rect 8964 845 8965 875
rect 8965 845 8995 875
rect 8995 845 8996 875
rect 8964 844 8996 845
rect 8964 764 8996 796
rect 8964 684 8996 716
rect 8964 635 8996 636
rect 8964 605 8965 635
rect 8965 605 8995 635
rect 8995 605 8996 635
rect 8964 604 8996 605
rect 8964 555 8996 556
rect 8964 525 8965 555
rect 8965 525 8995 555
rect 8995 525 8996 555
rect 8964 524 8996 525
rect 8964 444 8996 476
rect 8964 395 8996 396
rect 8964 365 8965 395
rect 8965 365 8995 395
rect 8995 365 8996 395
rect 8964 364 8996 365
rect 8964 284 8996 316
rect 8964 235 8996 236
rect 8964 205 8965 235
rect 8965 205 8995 235
rect 8995 205 8996 235
rect 8964 204 8996 205
rect 8964 124 8996 156
rect 8964 75 8996 76
rect 8964 45 8965 75
rect 8965 45 8995 75
rect 8995 45 8996 75
rect 8964 44 8996 45
rect 8964 -5 8996 -4
rect 8964 -35 8965 -5
rect 8965 -35 8995 -5
rect 8995 -35 8996 -5
rect 8964 -36 8996 -35
rect 8964 -85 8996 -84
rect 8964 -115 8965 -85
rect 8965 -115 8995 -85
rect 8995 -115 8996 -85
rect 8964 -116 8996 -115
rect 9044 1035 9076 1036
rect 9044 1005 9045 1035
rect 9045 1005 9075 1035
rect 9075 1005 9076 1035
rect 9044 1004 9076 1005
rect 9044 955 9076 956
rect 9044 925 9045 955
rect 9045 925 9075 955
rect 9075 925 9076 955
rect 9044 924 9076 925
rect 9044 875 9076 876
rect 9044 845 9045 875
rect 9045 845 9075 875
rect 9075 845 9076 875
rect 9044 844 9076 845
rect 9044 764 9076 796
rect 9044 684 9076 716
rect 9044 635 9076 636
rect 9044 605 9045 635
rect 9045 605 9075 635
rect 9075 605 9076 635
rect 9044 604 9076 605
rect 9044 555 9076 556
rect 9044 525 9045 555
rect 9045 525 9075 555
rect 9075 525 9076 555
rect 9044 524 9076 525
rect 9044 444 9076 476
rect 9044 395 9076 396
rect 9044 365 9045 395
rect 9045 365 9075 395
rect 9075 365 9076 395
rect 9044 364 9076 365
rect 9044 284 9076 316
rect 9044 235 9076 236
rect 9044 205 9045 235
rect 9045 205 9075 235
rect 9075 205 9076 235
rect 9044 204 9076 205
rect 9044 124 9076 156
rect 9044 75 9076 76
rect 9044 45 9045 75
rect 9045 45 9075 75
rect 9075 45 9076 75
rect 9044 44 9076 45
rect 9044 -5 9076 -4
rect 9044 -35 9045 -5
rect 9045 -35 9075 -5
rect 9075 -35 9076 -5
rect 9044 -36 9076 -35
rect 9044 -85 9076 -84
rect 9044 -115 9045 -85
rect 9045 -115 9075 -85
rect 9075 -115 9076 -85
rect 9044 -116 9076 -115
rect 9124 1035 9156 1036
rect 9124 1005 9125 1035
rect 9125 1005 9155 1035
rect 9155 1005 9156 1035
rect 9124 1004 9156 1005
rect 9124 955 9156 956
rect 9124 925 9125 955
rect 9125 925 9155 955
rect 9155 925 9156 955
rect 9124 924 9156 925
rect 9124 875 9156 876
rect 9124 845 9125 875
rect 9125 845 9155 875
rect 9155 845 9156 875
rect 9124 844 9156 845
rect 9124 764 9156 796
rect 9124 684 9156 716
rect 9124 635 9156 636
rect 9124 605 9125 635
rect 9125 605 9155 635
rect 9155 605 9156 635
rect 9124 604 9156 605
rect 9124 555 9156 556
rect 9124 525 9125 555
rect 9125 525 9155 555
rect 9155 525 9156 555
rect 9124 524 9156 525
rect 9124 444 9156 476
rect 9124 395 9156 396
rect 9124 365 9125 395
rect 9125 365 9155 395
rect 9155 365 9156 395
rect 9124 364 9156 365
rect 9124 284 9156 316
rect 9124 235 9156 236
rect 9124 205 9125 235
rect 9125 205 9155 235
rect 9155 205 9156 235
rect 9124 204 9156 205
rect 9124 124 9156 156
rect 9124 75 9156 76
rect 9124 45 9125 75
rect 9125 45 9155 75
rect 9155 45 9156 75
rect 9124 44 9156 45
rect 9124 -5 9156 -4
rect 9124 -35 9125 -5
rect 9125 -35 9155 -5
rect 9155 -35 9156 -5
rect 9124 -36 9156 -35
rect 9124 -85 9156 -84
rect 9124 -115 9125 -85
rect 9125 -115 9155 -85
rect 9155 -115 9156 -85
rect 9124 -116 9156 -115
rect 9204 1035 9236 1036
rect 9204 1005 9205 1035
rect 9205 1005 9235 1035
rect 9235 1005 9236 1035
rect 9204 1004 9236 1005
rect 9204 955 9236 956
rect 9204 925 9205 955
rect 9205 925 9235 955
rect 9235 925 9236 955
rect 9204 924 9236 925
rect 9204 875 9236 876
rect 9204 845 9205 875
rect 9205 845 9235 875
rect 9235 845 9236 875
rect 9204 844 9236 845
rect 9204 764 9236 796
rect 9204 684 9236 716
rect 9204 635 9236 636
rect 9204 605 9205 635
rect 9205 605 9235 635
rect 9235 605 9236 635
rect 9204 604 9236 605
rect 9204 555 9236 556
rect 9204 525 9205 555
rect 9205 525 9235 555
rect 9235 525 9236 555
rect 9204 524 9236 525
rect 9204 444 9236 476
rect 9204 395 9236 396
rect 9204 365 9205 395
rect 9205 365 9235 395
rect 9235 365 9236 395
rect 9204 364 9236 365
rect 9204 284 9236 316
rect 9204 235 9236 236
rect 9204 205 9205 235
rect 9205 205 9235 235
rect 9235 205 9236 235
rect 9204 204 9236 205
rect 9204 124 9236 156
rect 9204 75 9236 76
rect 9204 45 9205 75
rect 9205 45 9235 75
rect 9235 45 9236 75
rect 9204 44 9236 45
rect 9204 -5 9236 -4
rect 9204 -35 9205 -5
rect 9205 -35 9235 -5
rect 9235 -35 9236 -5
rect 9204 -36 9236 -35
rect 9204 -85 9236 -84
rect 9204 -115 9205 -85
rect 9205 -115 9235 -85
rect 9235 -115 9236 -85
rect 9204 -116 9236 -115
rect 9284 1035 9316 1036
rect 9284 1005 9285 1035
rect 9285 1005 9315 1035
rect 9315 1005 9316 1035
rect 9284 1004 9316 1005
rect 9284 955 9316 956
rect 9284 925 9285 955
rect 9285 925 9315 955
rect 9315 925 9316 955
rect 9284 924 9316 925
rect 9284 875 9316 876
rect 9284 845 9285 875
rect 9285 845 9315 875
rect 9315 845 9316 875
rect 9284 844 9316 845
rect 9284 764 9316 796
rect 9284 684 9316 716
rect 9284 635 9316 636
rect 9284 605 9285 635
rect 9285 605 9315 635
rect 9315 605 9316 635
rect 9284 604 9316 605
rect 9284 555 9316 556
rect 9284 525 9285 555
rect 9285 525 9315 555
rect 9315 525 9316 555
rect 9284 524 9316 525
rect 9284 444 9316 476
rect 9284 395 9316 396
rect 9284 365 9285 395
rect 9285 365 9315 395
rect 9315 365 9316 395
rect 9284 364 9316 365
rect 9284 284 9316 316
rect 9284 235 9316 236
rect 9284 205 9285 235
rect 9285 205 9315 235
rect 9315 205 9316 235
rect 9284 204 9316 205
rect 9284 124 9316 156
rect 9284 75 9316 76
rect 9284 45 9285 75
rect 9285 45 9315 75
rect 9315 45 9316 75
rect 9284 44 9316 45
rect 9284 -5 9316 -4
rect 9284 -35 9285 -5
rect 9285 -35 9315 -5
rect 9315 -35 9316 -5
rect 9284 -36 9316 -35
rect 9284 -85 9316 -84
rect 9284 -115 9285 -85
rect 9285 -115 9315 -85
rect 9315 -115 9316 -85
rect 9284 -116 9316 -115
rect 9364 1035 9396 1036
rect 9364 1005 9365 1035
rect 9365 1005 9395 1035
rect 9395 1005 9396 1035
rect 9364 1004 9396 1005
rect 9364 955 9396 956
rect 9364 925 9365 955
rect 9365 925 9395 955
rect 9395 925 9396 955
rect 9364 924 9396 925
rect 9364 875 9396 876
rect 9364 845 9365 875
rect 9365 845 9395 875
rect 9395 845 9396 875
rect 9364 844 9396 845
rect 9364 764 9396 796
rect 9364 684 9396 716
rect 9364 635 9396 636
rect 9364 605 9365 635
rect 9365 605 9395 635
rect 9395 605 9396 635
rect 9364 604 9396 605
rect 9364 555 9396 556
rect 9364 525 9365 555
rect 9365 525 9395 555
rect 9395 525 9396 555
rect 9364 524 9396 525
rect 9364 444 9396 476
rect 9364 395 9396 396
rect 9364 365 9365 395
rect 9365 365 9395 395
rect 9395 365 9396 395
rect 9364 364 9396 365
rect 9364 284 9396 316
rect 9364 235 9396 236
rect 9364 205 9365 235
rect 9365 205 9395 235
rect 9395 205 9396 235
rect 9364 204 9396 205
rect 9364 124 9396 156
rect 9364 75 9396 76
rect 9364 45 9365 75
rect 9365 45 9395 75
rect 9395 45 9396 75
rect 9364 44 9396 45
rect 9364 -5 9396 -4
rect 9364 -35 9365 -5
rect 9365 -35 9395 -5
rect 9395 -35 9396 -5
rect 9364 -36 9396 -35
rect 9364 -85 9396 -84
rect 9364 -115 9365 -85
rect 9365 -115 9395 -85
rect 9395 -115 9396 -85
rect 9364 -116 9396 -115
rect 9444 1035 9476 1036
rect 9444 1005 9445 1035
rect 9445 1005 9475 1035
rect 9475 1005 9476 1035
rect 9444 1004 9476 1005
rect 9444 955 9476 956
rect 9444 925 9445 955
rect 9445 925 9475 955
rect 9475 925 9476 955
rect 9444 924 9476 925
rect 9444 875 9476 876
rect 9444 845 9445 875
rect 9445 845 9475 875
rect 9475 845 9476 875
rect 9444 844 9476 845
rect 9444 764 9476 796
rect 9444 684 9476 716
rect 9444 635 9476 636
rect 9444 605 9445 635
rect 9445 605 9475 635
rect 9475 605 9476 635
rect 9444 604 9476 605
rect 9444 555 9476 556
rect 9444 525 9445 555
rect 9445 525 9475 555
rect 9475 525 9476 555
rect 9444 524 9476 525
rect 9444 444 9476 476
rect 9444 395 9476 396
rect 9444 365 9445 395
rect 9445 365 9475 395
rect 9475 365 9476 395
rect 9444 364 9476 365
rect 9444 284 9476 316
rect 9444 235 9476 236
rect 9444 205 9445 235
rect 9445 205 9475 235
rect 9475 205 9476 235
rect 9444 204 9476 205
rect 9444 124 9476 156
rect 9444 75 9476 76
rect 9444 45 9445 75
rect 9445 45 9475 75
rect 9475 45 9476 75
rect 9444 44 9476 45
rect 9444 -5 9476 -4
rect 9444 -35 9445 -5
rect 9445 -35 9475 -5
rect 9475 -35 9476 -5
rect 9444 -36 9476 -35
rect 9444 -85 9476 -84
rect 9444 -115 9445 -85
rect 9445 -115 9475 -85
rect 9475 -115 9476 -85
rect 9444 -116 9476 -115
rect 9524 1035 9556 1036
rect 9524 1005 9525 1035
rect 9525 1005 9555 1035
rect 9555 1005 9556 1035
rect 9524 1004 9556 1005
rect 9524 955 9556 956
rect 9524 925 9525 955
rect 9525 925 9555 955
rect 9555 925 9556 955
rect 9524 924 9556 925
rect 9524 875 9556 876
rect 9524 845 9525 875
rect 9525 845 9555 875
rect 9555 845 9556 875
rect 9524 844 9556 845
rect 9524 764 9556 796
rect 9524 684 9556 716
rect 9524 635 9556 636
rect 9524 605 9525 635
rect 9525 605 9555 635
rect 9555 605 9556 635
rect 9524 604 9556 605
rect 9524 555 9556 556
rect 9524 525 9525 555
rect 9525 525 9555 555
rect 9555 525 9556 555
rect 9524 524 9556 525
rect 9524 444 9556 476
rect 9524 395 9556 396
rect 9524 365 9525 395
rect 9525 365 9555 395
rect 9555 365 9556 395
rect 9524 364 9556 365
rect 9524 284 9556 316
rect 9524 235 9556 236
rect 9524 205 9525 235
rect 9525 205 9555 235
rect 9555 205 9556 235
rect 9524 204 9556 205
rect 9524 124 9556 156
rect 9524 75 9556 76
rect 9524 45 9525 75
rect 9525 45 9555 75
rect 9555 45 9556 75
rect 9524 44 9556 45
rect 9524 -5 9556 -4
rect 9524 -35 9525 -5
rect 9525 -35 9555 -5
rect 9555 -35 9556 -5
rect 9524 -36 9556 -35
rect 9524 -85 9556 -84
rect 9524 -115 9525 -85
rect 9525 -115 9555 -85
rect 9555 -115 9556 -85
rect 9524 -116 9556 -115
rect 9604 1035 9636 1036
rect 9604 1005 9605 1035
rect 9605 1005 9635 1035
rect 9635 1005 9636 1035
rect 9604 1004 9636 1005
rect 9604 955 9636 956
rect 9604 925 9605 955
rect 9605 925 9635 955
rect 9635 925 9636 955
rect 9604 924 9636 925
rect 9604 875 9636 876
rect 9604 845 9605 875
rect 9605 845 9635 875
rect 9635 845 9636 875
rect 9604 844 9636 845
rect 9604 764 9636 796
rect 9604 684 9636 716
rect 9604 635 9636 636
rect 9604 605 9605 635
rect 9605 605 9635 635
rect 9635 605 9636 635
rect 9604 604 9636 605
rect 9604 555 9636 556
rect 9604 525 9605 555
rect 9605 525 9635 555
rect 9635 525 9636 555
rect 9604 524 9636 525
rect 9604 444 9636 476
rect 9604 395 9636 396
rect 9604 365 9605 395
rect 9605 365 9635 395
rect 9635 365 9636 395
rect 9604 364 9636 365
rect 9604 284 9636 316
rect 9604 235 9636 236
rect 9604 205 9605 235
rect 9605 205 9635 235
rect 9635 205 9636 235
rect 9604 204 9636 205
rect 9604 124 9636 156
rect 9604 75 9636 76
rect 9604 45 9605 75
rect 9605 45 9635 75
rect 9635 45 9636 75
rect 9604 44 9636 45
rect 9604 -5 9636 -4
rect 9604 -35 9605 -5
rect 9605 -35 9635 -5
rect 9635 -35 9636 -5
rect 9604 -36 9636 -35
rect 9604 -85 9636 -84
rect 9604 -115 9605 -85
rect 9605 -115 9635 -85
rect 9635 -115 9636 -85
rect 9604 -116 9636 -115
rect 9684 1035 9716 1036
rect 9684 1005 9685 1035
rect 9685 1005 9715 1035
rect 9715 1005 9716 1035
rect 9684 1004 9716 1005
rect 9684 955 9716 956
rect 9684 925 9685 955
rect 9685 925 9715 955
rect 9715 925 9716 955
rect 9684 924 9716 925
rect 9684 875 9716 876
rect 9684 845 9685 875
rect 9685 845 9715 875
rect 9715 845 9716 875
rect 9684 844 9716 845
rect 9684 764 9716 796
rect 9684 684 9716 716
rect 9684 635 9716 636
rect 9684 605 9685 635
rect 9685 605 9715 635
rect 9715 605 9716 635
rect 9684 604 9716 605
rect 9684 555 9716 556
rect 9684 525 9685 555
rect 9685 525 9715 555
rect 9715 525 9716 555
rect 9684 524 9716 525
rect 9684 444 9716 476
rect 9684 395 9716 396
rect 9684 365 9685 395
rect 9685 365 9715 395
rect 9715 365 9716 395
rect 9684 364 9716 365
rect 9684 284 9716 316
rect 9684 235 9716 236
rect 9684 205 9685 235
rect 9685 205 9715 235
rect 9715 205 9716 235
rect 9684 204 9716 205
rect 9684 124 9716 156
rect 9684 75 9716 76
rect 9684 45 9685 75
rect 9685 45 9715 75
rect 9715 45 9716 75
rect 9684 44 9716 45
rect 9684 -5 9716 -4
rect 9684 -35 9685 -5
rect 9685 -35 9715 -5
rect 9715 -35 9716 -5
rect 9684 -36 9716 -35
rect 9684 -85 9716 -84
rect 9684 -115 9685 -85
rect 9685 -115 9715 -85
rect 9715 -115 9716 -85
rect 9684 -116 9716 -115
rect 9764 1035 9796 1036
rect 9764 1005 9765 1035
rect 9765 1005 9795 1035
rect 9795 1005 9796 1035
rect 9764 1004 9796 1005
rect 9764 955 9796 956
rect 9764 925 9765 955
rect 9765 925 9795 955
rect 9795 925 9796 955
rect 9764 924 9796 925
rect 9764 875 9796 876
rect 9764 845 9765 875
rect 9765 845 9795 875
rect 9795 845 9796 875
rect 9764 844 9796 845
rect 9764 764 9796 796
rect 9764 684 9796 716
rect 9764 635 9796 636
rect 9764 605 9765 635
rect 9765 605 9795 635
rect 9795 605 9796 635
rect 9764 604 9796 605
rect 9764 555 9796 556
rect 9764 525 9765 555
rect 9765 525 9795 555
rect 9795 525 9796 555
rect 9764 524 9796 525
rect 9764 444 9796 476
rect 9764 395 9796 396
rect 9764 365 9765 395
rect 9765 365 9795 395
rect 9795 365 9796 395
rect 9764 364 9796 365
rect 9764 284 9796 316
rect 9764 235 9796 236
rect 9764 205 9765 235
rect 9765 205 9795 235
rect 9795 205 9796 235
rect 9764 204 9796 205
rect 9764 124 9796 156
rect 9764 75 9796 76
rect 9764 45 9765 75
rect 9765 45 9795 75
rect 9795 45 9796 75
rect 9764 44 9796 45
rect 9764 -5 9796 -4
rect 9764 -35 9765 -5
rect 9765 -35 9795 -5
rect 9795 -35 9796 -5
rect 9764 -36 9796 -35
rect 9764 -85 9796 -84
rect 9764 -115 9765 -85
rect 9765 -115 9795 -85
rect 9795 -115 9796 -85
rect 9764 -116 9796 -115
rect 9844 1035 9876 1036
rect 9844 1005 9845 1035
rect 9845 1005 9875 1035
rect 9875 1005 9876 1035
rect 9844 1004 9876 1005
rect 9844 955 9876 956
rect 9844 925 9845 955
rect 9845 925 9875 955
rect 9875 925 9876 955
rect 9844 924 9876 925
rect 9844 875 9876 876
rect 9844 845 9845 875
rect 9845 845 9875 875
rect 9875 845 9876 875
rect 9844 844 9876 845
rect 9844 764 9876 796
rect 9844 684 9876 716
rect 9844 635 9876 636
rect 9844 605 9845 635
rect 9845 605 9875 635
rect 9875 605 9876 635
rect 9844 604 9876 605
rect 9844 555 9876 556
rect 9844 525 9845 555
rect 9845 525 9875 555
rect 9875 525 9876 555
rect 9844 524 9876 525
rect 9844 444 9876 476
rect 9844 395 9876 396
rect 9844 365 9845 395
rect 9845 365 9875 395
rect 9875 365 9876 395
rect 9844 364 9876 365
rect 9844 284 9876 316
rect 9844 235 9876 236
rect 9844 205 9845 235
rect 9845 205 9875 235
rect 9875 205 9876 235
rect 9844 204 9876 205
rect 9844 124 9876 156
rect 9844 75 9876 76
rect 9844 45 9845 75
rect 9845 45 9875 75
rect 9875 45 9876 75
rect 9844 44 9876 45
rect 9844 -5 9876 -4
rect 9844 -35 9845 -5
rect 9845 -35 9875 -5
rect 9875 -35 9876 -5
rect 9844 -36 9876 -35
rect 9844 -85 9876 -84
rect 9844 -115 9845 -85
rect 9845 -115 9875 -85
rect 9875 -115 9876 -85
rect 9844 -116 9876 -115
rect 9924 1035 9956 1036
rect 9924 1005 9925 1035
rect 9925 1005 9955 1035
rect 9955 1005 9956 1035
rect 9924 1004 9956 1005
rect 9924 955 9956 956
rect 9924 925 9925 955
rect 9925 925 9955 955
rect 9955 925 9956 955
rect 9924 924 9956 925
rect 9924 875 9956 876
rect 9924 845 9925 875
rect 9925 845 9955 875
rect 9955 845 9956 875
rect 9924 844 9956 845
rect 9924 764 9956 796
rect 9924 684 9956 716
rect 9924 635 9956 636
rect 9924 605 9925 635
rect 9925 605 9955 635
rect 9955 605 9956 635
rect 9924 604 9956 605
rect 9924 555 9956 556
rect 9924 525 9925 555
rect 9925 525 9955 555
rect 9955 525 9956 555
rect 9924 524 9956 525
rect 9924 444 9956 476
rect 9924 395 9956 396
rect 9924 365 9925 395
rect 9925 365 9955 395
rect 9955 365 9956 395
rect 9924 364 9956 365
rect 9924 284 9956 316
rect 9924 235 9956 236
rect 9924 205 9925 235
rect 9925 205 9955 235
rect 9955 205 9956 235
rect 9924 204 9956 205
rect 9924 124 9956 156
rect 9924 75 9956 76
rect 9924 45 9925 75
rect 9925 45 9955 75
rect 9955 45 9956 75
rect 9924 44 9956 45
rect 9924 -5 9956 -4
rect 9924 -35 9925 -5
rect 9925 -35 9955 -5
rect 9955 -35 9956 -5
rect 9924 -36 9956 -35
rect 9924 -85 9956 -84
rect 9924 -115 9925 -85
rect 9925 -115 9955 -85
rect 9955 -115 9956 -85
rect 9924 -116 9956 -115
rect 10004 1035 10036 1036
rect 10004 1005 10005 1035
rect 10005 1005 10035 1035
rect 10035 1005 10036 1035
rect 10004 1004 10036 1005
rect 10004 955 10036 956
rect 10004 925 10005 955
rect 10005 925 10035 955
rect 10035 925 10036 955
rect 10004 924 10036 925
rect 10004 875 10036 876
rect 10004 845 10005 875
rect 10005 845 10035 875
rect 10035 845 10036 875
rect 10004 844 10036 845
rect 10004 764 10036 796
rect 10004 684 10036 716
rect 10004 635 10036 636
rect 10004 605 10005 635
rect 10005 605 10035 635
rect 10035 605 10036 635
rect 10004 604 10036 605
rect 10004 555 10036 556
rect 10004 525 10005 555
rect 10005 525 10035 555
rect 10035 525 10036 555
rect 10004 524 10036 525
rect 10004 444 10036 476
rect 10004 395 10036 396
rect 10004 365 10005 395
rect 10005 365 10035 395
rect 10035 365 10036 395
rect 10004 364 10036 365
rect 10004 284 10036 316
rect 10004 235 10036 236
rect 10004 205 10005 235
rect 10005 205 10035 235
rect 10035 205 10036 235
rect 10004 204 10036 205
rect 10004 124 10036 156
rect 10004 75 10036 76
rect 10004 45 10005 75
rect 10005 45 10035 75
rect 10035 45 10036 75
rect 10004 44 10036 45
rect 10004 -5 10036 -4
rect 10004 -35 10005 -5
rect 10005 -35 10035 -5
rect 10035 -35 10036 -5
rect 10004 -36 10036 -35
rect 10004 -85 10036 -84
rect 10004 -115 10005 -85
rect 10005 -115 10035 -85
rect 10035 -115 10036 -85
rect 10004 -116 10036 -115
rect 10084 1035 10116 1036
rect 10084 1005 10085 1035
rect 10085 1005 10115 1035
rect 10115 1005 10116 1035
rect 10084 1004 10116 1005
rect 10084 955 10116 956
rect 10084 925 10085 955
rect 10085 925 10115 955
rect 10115 925 10116 955
rect 10084 924 10116 925
rect 10084 875 10116 876
rect 10084 845 10085 875
rect 10085 845 10115 875
rect 10115 845 10116 875
rect 10084 844 10116 845
rect 10084 764 10116 796
rect 10084 684 10116 716
rect 10084 635 10116 636
rect 10084 605 10085 635
rect 10085 605 10115 635
rect 10115 605 10116 635
rect 10084 604 10116 605
rect 10084 555 10116 556
rect 10084 525 10085 555
rect 10085 525 10115 555
rect 10115 525 10116 555
rect 10084 524 10116 525
rect 10084 444 10116 476
rect 10084 395 10116 396
rect 10084 365 10085 395
rect 10085 365 10115 395
rect 10115 365 10116 395
rect 10084 364 10116 365
rect 10084 284 10116 316
rect 10084 235 10116 236
rect 10084 205 10085 235
rect 10085 205 10115 235
rect 10115 205 10116 235
rect 10084 204 10116 205
rect 10084 124 10116 156
rect 10084 75 10116 76
rect 10084 45 10085 75
rect 10085 45 10115 75
rect 10115 45 10116 75
rect 10084 44 10116 45
rect 10084 -5 10116 -4
rect 10084 -35 10085 -5
rect 10085 -35 10115 -5
rect 10115 -35 10116 -5
rect 10084 -36 10116 -35
rect 10084 -85 10116 -84
rect 10084 -115 10085 -85
rect 10085 -115 10115 -85
rect 10115 -115 10116 -85
rect 10084 -116 10116 -115
rect 10164 1035 10196 1036
rect 10164 1005 10165 1035
rect 10165 1005 10195 1035
rect 10195 1005 10196 1035
rect 10164 1004 10196 1005
rect 10164 955 10196 956
rect 10164 925 10165 955
rect 10165 925 10195 955
rect 10195 925 10196 955
rect 10164 924 10196 925
rect 10164 875 10196 876
rect 10164 845 10165 875
rect 10165 845 10195 875
rect 10195 845 10196 875
rect 10164 844 10196 845
rect 10164 764 10196 796
rect 10164 684 10196 716
rect 10164 635 10196 636
rect 10164 605 10165 635
rect 10165 605 10195 635
rect 10195 605 10196 635
rect 10164 604 10196 605
rect 10164 555 10196 556
rect 10164 525 10165 555
rect 10165 525 10195 555
rect 10195 525 10196 555
rect 10164 524 10196 525
rect 10164 444 10196 476
rect 10164 395 10196 396
rect 10164 365 10165 395
rect 10165 365 10195 395
rect 10195 365 10196 395
rect 10164 364 10196 365
rect 10164 284 10196 316
rect 10164 235 10196 236
rect 10164 205 10165 235
rect 10165 205 10195 235
rect 10195 205 10196 235
rect 10164 204 10196 205
rect 10164 124 10196 156
rect 10164 75 10196 76
rect 10164 45 10165 75
rect 10165 45 10195 75
rect 10195 45 10196 75
rect 10164 44 10196 45
rect 10164 -5 10196 -4
rect 10164 -35 10165 -5
rect 10165 -35 10195 -5
rect 10195 -35 10196 -5
rect 10164 -36 10196 -35
rect 10164 -85 10196 -84
rect 10164 -115 10165 -85
rect 10165 -115 10195 -85
rect 10195 -115 10196 -85
rect 10164 -116 10196 -115
rect 10244 1035 10276 1036
rect 10244 1005 10245 1035
rect 10245 1005 10275 1035
rect 10275 1005 10276 1035
rect 10244 1004 10276 1005
rect 10244 955 10276 956
rect 10244 925 10245 955
rect 10245 925 10275 955
rect 10275 925 10276 955
rect 10244 924 10276 925
rect 10244 875 10276 876
rect 10244 845 10245 875
rect 10245 845 10275 875
rect 10275 845 10276 875
rect 10244 844 10276 845
rect 10244 764 10276 796
rect 10244 684 10276 716
rect 10244 635 10276 636
rect 10244 605 10245 635
rect 10245 605 10275 635
rect 10275 605 10276 635
rect 10244 604 10276 605
rect 10244 555 10276 556
rect 10244 525 10245 555
rect 10245 525 10275 555
rect 10275 525 10276 555
rect 10244 524 10276 525
rect 10244 444 10276 476
rect 10244 395 10276 396
rect 10244 365 10245 395
rect 10245 365 10275 395
rect 10275 365 10276 395
rect 10244 364 10276 365
rect 10244 284 10276 316
rect 10244 235 10276 236
rect 10244 205 10245 235
rect 10245 205 10275 235
rect 10275 205 10276 235
rect 10244 204 10276 205
rect 10244 124 10276 156
rect 10244 75 10276 76
rect 10244 45 10245 75
rect 10245 45 10275 75
rect 10275 45 10276 75
rect 10244 44 10276 45
rect 10244 -5 10276 -4
rect 10244 -35 10245 -5
rect 10245 -35 10275 -5
rect 10275 -35 10276 -5
rect 10244 -36 10276 -35
rect 10244 -85 10276 -84
rect 10244 -115 10245 -85
rect 10245 -115 10275 -85
rect 10275 -115 10276 -85
rect 10244 -116 10276 -115
rect 10324 1035 10356 1036
rect 10324 1005 10325 1035
rect 10325 1005 10355 1035
rect 10355 1005 10356 1035
rect 10324 1004 10356 1005
rect 10324 955 10356 956
rect 10324 925 10325 955
rect 10325 925 10355 955
rect 10355 925 10356 955
rect 10324 924 10356 925
rect 10324 875 10356 876
rect 10324 845 10325 875
rect 10325 845 10355 875
rect 10355 845 10356 875
rect 10324 844 10356 845
rect 10324 764 10356 796
rect 10324 684 10356 716
rect 10324 635 10356 636
rect 10324 605 10325 635
rect 10325 605 10355 635
rect 10355 605 10356 635
rect 10324 604 10356 605
rect 10324 555 10356 556
rect 10324 525 10325 555
rect 10325 525 10355 555
rect 10355 525 10356 555
rect 10324 524 10356 525
rect 10324 444 10356 476
rect 10324 395 10356 396
rect 10324 365 10325 395
rect 10325 365 10355 395
rect 10355 365 10356 395
rect 10324 364 10356 365
rect 10324 284 10356 316
rect 10324 235 10356 236
rect 10324 205 10325 235
rect 10325 205 10355 235
rect 10355 205 10356 235
rect 10324 204 10356 205
rect 10324 124 10356 156
rect 10324 75 10356 76
rect 10324 45 10325 75
rect 10325 45 10355 75
rect 10355 45 10356 75
rect 10324 44 10356 45
rect 10324 -5 10356 -4
rect 10324 -35 10325 -5
rect 10325 -35 10355 -5
rect 10355 -35 10356 -5
rect 10324 -36 10356 -35
rect 10324 -85 10356 -84
rect 10324 -115 10325 -85
rect 10325 -115 10355 -85
rect 10355 -115 10356 -85
rect 10324 -116 10356 -115
rect 10404 1035 10436 1036
rect 10404 1005 10405 1035
rect 10405 1005 10435 1035
rect 10435 1005 10436 1035
rect 10404 1004 10436 1005
rect 10404 955 10436 956
rect 10404 925 10405 955
rect 10405 925 10435 955
rect 10435 925 10436 955
rect 10404 924 10436 925
rect 10404 875 10436 876
rect 10404 845 10405 875
rect 10405 845 10435 875
rect 10435 845 10436 875
rect 10404 844 10436 845
rect 10404 764 10436 796
rect 10404 684 10436 716
rect 10404 635 10436 636
rect 10404 605 10405 635
rect 10405 605 10435 635
rect 10435 605 10436 635
rect 10404 604 10436 605
rect 10404 555 10436 556
rect 10404 525 10405 555
rect 10405 525 10435 555
rect 10435 525 10436 555
rect 10404 524 10436 525
rect 10404 444 10436 476
rect 10404 395 10436 396
rect 10404 365 10405 395
rect 10405 365 10435 395
rect 10435 365 10436 395
rect 10404 364 10436 365
rect 10404 284 10436 316
rect 10404 235 10436 236
rect 10404 205 10405 235
rect 10405 205 10435 235
rect 10435 205 10436 235
rect 10404 204 10436 205
rect 10404 124 10436 156
rect 10404 75 10436 76
rect 10404 45 10405 75
rect 10405 45 10435 75
rect 10435 45 10436 75
rect 10404 44 10436 45
rect 10404 -5 10436 -4
rect 10404 -35 10405 -5
rect 10405 -35 10435 -5
rect 10435 -35 10436 -5
rect 10404 -36 10436 -35
rect 10404 -85 10436 -84
rect 10404 -115 10405 -85
rect 10405 -115 10435 -85
rect 10435 -115 10436 -85
rect 10404 -116 10436 -115
rect 10484 1035 10516 1036
rect 10484 1005 10485 1035
rect 10485 1005 10515 1035
rect 10515 1005 10516 1035
rect 10484 1004 10516 1005
rect 10484 955 10516 956
rect 10484 925 10485 955
rect 10485 925 10515 955
rect 10515 925 10516 955
rect 10484 924 10516 925
rect 10484 875 10516 876
rect 10484 845 10485 875
rect 10485 845 10515 875
rect 10515 845 10516 875
rect 10484 844 10516 845
rect 10484 764 10516 796
rect 10484 684 10516 716
rect 10484 635 10516 636
rect 10484 605 10485 635
rect 10485 605 10515 635
rect 10515 605 10516 635
rect 10484 604 10516 605
rect 10484 555 10516 556
rect 10484 525 10485 555
rect 10485 525 10515 555
rect 10515 525 10516 555
rect 10484 524 10516 525
rect 10484 444 10516 476
rect 10484 395 10516 396
rect 10484 365 10485 395
rect 10485 365 10515 395
rect 10515 365 10516 395
rect 10484 364 10516 365
rect 10484 284 10516 316
rect 10484 235 10516 236
rect 10484 205 10485 235
rect 10485 205 10515 235
rect 10515 205 10516 235
rect 10484 204 10516 205
rect 10484 124 10516 156
rect 10484 75 10516 76
rect 10484 45 10485 75
rect 10485 45 10515 75
rect 10515 45 10516 75
rect 10484 44 10516 45
rect 10484 -5 10516 -4
rect 10484 -35 10485 -5
rect 10485 -35 10515 -5
rect 10515 -35 10516 -5
rect 10484 -36 10516 -35
rect 10484 -85 10516 -84
rect 10484 -115 10485 -85
rect 10485 -115 10515 -85
rect 10515 -115 10516 -85
rect 10484 -116 10516 -115
rect 10644 1035 10676 1036
rect 10644 1005 10645 1035
rect 10645 1005 10675 1035
rect 10675 1005 10676 1035
rect 10644 1004 10676 1005
rect 10644 955 10676 956
rect 10644 925 10645 955
rect 10645 925 10675 955
rect 10675 925 10676 955
rect 10644 924 10676 925
rect 10644 875 10676 876
rect 10644 845 10645 875
rect 10645 845 10675 875
rect 10675 845 10676 875
rect 10644 844 10676 845
rect 10644 795 10676 796
rect 10644 765 10645 795
rect 10645 765 10675 795
rect 10675 765 10676 795
rect 10644 764 10676 765
rect 10644 715 10676 716
rect 10644 685 10645 715
rect 10645 685 10675 715
rect 10675 685 10676 715
rect 10644 684 10676 685
rect 10644 635 10676 636
rect 10644 605 10645 635
rect 10645 605 10675 635
rect 10675 605 10676 635
rect 10644 604 10676 605
rect 10644 555 10676 556
rect 10644 525 10645 555
rect 10645 525 10675 555
rect 10675 525 10676 555
rect 10644 524 10676 525
rect 10644 475 10676 476
rect 10644 445 10645 475
rect 10645 445 10675 475
rect 10675 445 10676 475
rect 10644 444 10676 445
rect 10644 395 10676 396
rect 10644 365 10645 395
rect 10645 365 10675 395
rect 10675 365 10676 395
rect 10644 364 10676 365
rect 10644 284 10676 316
rect 10644 235 10676 236
rect 10644 205 10645 235
rect 10645 205 10675 235
rect 10675 205 10676 235
rect 10644 204 10676 205
rect 10644 124 10676 156
rect 10644 75 10676 76
rect 10644 45 10645 75
rect 10645 45 10675 75
rect 10675 45 10676 75
rect 10644 44 10676 45
rect 10644 -5 10676 -4
rect 10644 -35 10645 -5
rect 10645 -35 10675 -5
rect 10675 -35 10676 -5
rect 10644 -36 10676 -35
rect 10644 -85 10676 -84
rect 10644 -115 10645 -85
rect 10645 -115 10675 -85
rect 10675 -115 10676 -85
rect 10644 -116 10676 -115
rect 10804 1035 10836 1036
rect 10804 1005 10805 1035
rect 10805 1005 10835 1035
rect 10835 1005 10836 1035
rect 10804 1004 10836 1005
rect 10804 955 10836 956
rect 10804 925 10805 955
rect 10805 925 10835 955
rect 10835 925 10836 955
rect 10804 924 10836 925
rect 10804 875 10836 876
rect 10804 845 10805 875
rect 10805 845 10835 875
rect 10835 845 10836 875
rect 10804 844 10836 845
rect 10804 795 10836 796
rect 10804 765 10805 795
rect 10805 765 10835 795
rect 10835 765 10836 795
rect 10804 764 10836 765
rect 10804 715 10836 716
rect 10804 685 10805 715
rect 10805 685 10835 715
rect 10835 685 10836 715
rect 10804 684 10836 685
rect 10804 635 10836 636
rect 10804 605 10805 635
rect 10805 605 10835 635
rect 10835 605 10836 635
rect 10804 604 10836 605
rect 10804 555 10836 556
rect 10804 525 10805 555
rect 10805 525 10835 555
rect 10835 525 10836 555
rect 10804 524 10836 525
rect 10804 475 10836 476
rect 10804 445 10805 475
rect 10805 445 10835 475
rect 10835 445 10836 475
rect 10804 444 10836 445
rect 10804 395 10836 396
rect 10804 365 10805 395
rect 10805 365 10835 395
rect 10835 365 10836 395
rect 10804 364 10836 365
rect 10804 284 10836 316
rect 10804 235 10836 236
rect 10804 205 10805 235
rect 10805 205 10835 235
rect 10835 205 10836 235
rect 10804 204 10836 205
rect 10804 155 10836 156
rect 10804 125 10805 155
rect 10805 125 10835 155
rect 10835 125 10836 155
rect 10804 124 10836 125
rect 10804 75 10836 76
rect 10804 45 10805 75
rect 10805 45 10835 75
rect 10835 45 10836 75
rect 10804 44 10836 45
rect 10804 -5 10836 -4
rect 10804 -35 10805 -5
rect 10805 -35 10835 -5
rect 10835 -35 10836 -5
rect 10804 -36 10836 -35
rect 10804 -85 10836 -84
rect 10804 -115 10805 -85
rect 10805 -115 10835 -85
rect 10835 -115 10836 -85
rect 10804 -116 10836 -115
rect 10964 1035 10996 1036
rect 10964 1005 10965 1035
rect 10965 1005 10995 1035
rect 10995 1005 10996 1035
rect 10964 1004 10996 1005
rect 10964 955 10996 956
rect 10964 925 10965 955
rect 10965 925 10995 955
rect 10995 925 10996 955
rect 10964 924 10996 925
rect 10964 875 10996 876
rect 10964 845 10965 875
rect 10965 845 10995 875
rect 10995 845 10996 875
rect 10964 844 10996 845
rect 10964 795 10996 796
rect 10964 765 10965 795
rect 10965 765 10995 795
rect 10995 765 10996 795
rect 10964 764 10996 765
rect 10964 715 10996 716
rect 10964 685 10965 715
rect 10965 685 10995 715
rect 10995 685 10996 715
rect 10964 684 10996 685
rect 10964 635 10996 636
rect 10964 605 10965 635
rect 10965 605 10995 635
rect 10995 605 10996 635
rect 10964 604 10996 605
rect 10964 555 10996 556
rect 10964 525 10965 555
rect 10965 525 10995 555
rect 10995 525 10996 555
rect 10964 524 10996 525
rect 10964 475 10996 476
rect 10964 445 10965 475
rect 10965 445 10995 475
rect 10995 445 10996 475
rect 10964 444 10996 445
rect 10964 395 10996 396
rect 10964 365 10965 395
rect 10965 365 10995 395
rect 10995 365 10996 395
rect 10964 364 10996 365
rect 10964 284 10996 316
rect 10964 235 10996 236
rect 10964 205 10965 235
rect 10965 205 10995 235
rect 10995 205 10996 235
rect 10964 204 10996 205
rect 10964 155 10996 156
rect 10964 125 10965 155
rect 10965 125 10995 155
rect 10995 125 10996 155
rect 10964 124 10996 125
rect 10964 75 10996 76
rect 10964 45 10965 75
rect 10965 45 10995 75
rect 10995 45 10996 75
rect 10964 44 10996 45
rect 10964 -5 10996 -4
rect 10964 -35 10965 -5
rect 10965 -35 10995 -5
rect 10995 -35 10996 -5
rect 10964 -36 10996 -35
rect 10964 -85 10996 -84
rect 10964 -115 10965 -85
rect 10965 -115 10995 -85
rect 10995 -115 10996 -85
rect 10964 -116 10996 -115
<< metal4 >>
rect -720 1036 11000 1040
rect -720 1004 -716 1036
rect -684 1004 -556 1036
rect -524 1004 -396 1036
rect -364 1004 -316 1036
rect -284 1004 -236 1036
rect -204 1004 -156 1036
rect -124 1004 -76 1036
rect -44 1004 4 1036
rect 36 1004 84 1036
rect 116 1004 164 1036
rect 196 1004 244 1036
rect 276 1004 324 1036
rect 356 1004 404 1036
rect 436 1004 484 1036
rect 516 1004 564 1036
rect 596 1004 644 1036
rect 676 1004 724 1036
rect 756 1004 804 1036
rect 836 1004 884 1036
rect 916 1004 964 1036
rect 996 1004 1044 1036
rect 1076 1004 1124 1036
rect 1156 1004 1204 1036
rect 1236 1004 1284 1036
rect 1316 1004 1364 1036
rect 1396 1004 1444 1036
rect 1476 1004 1524 1036
rect 1556 1004 1604 1036
rect 1636 1004 1684 1036
rect 1716 1004 1764 1036
rect 1796 1004 1844 1036
rect 1876 1004 1924 1036
rect 1956 1004 2004 1036
rect 2036 1004 2084 1036
rect 2116 1004 2164 1036
rect 2196 1004 2244 1036
rect 2276 1004 2324 1036
rect 2356 1004 2404 1036
rect 2436 1004 2484 1036
rect 2516 1004 2564 1036
rect 2596 1004 2644 1036
rect 2676 1004 2724 1036
rect 2756 1004 2804 1036
rect 2836 1004 2884 1036
rect 2916 1004 2964 1036
rect 2996 1004 3044 1036
rect 3076 1004 3124 1036
rect 3156 1004 3204 1036
rect 3236 1004 3284 1036
rect 3316 1004 3364 1036
rect 3396 1004 3444 1036
rect 3476 1004 3524 1036
rect 3556 1004 3604 1036
rect 3636 1004 3684 1036
rect 3716 1004 3764 1036
rect 3796 1004 3844 1036
rect 3876 1004 3924 1036
rect 3956 1004 4004 1036
rect 4036 1004 4084 1036
rect 4116 1004 4164 1036
rect 4196 1004 4244 1036
rect 4276 1004 4324 1036
rect 4356 1004 4404 1036
rect 4436 1004 4484 1036
rect 4516 1004 4564 1036
rect 4596 1004 4644 1036
rect 4676 1004 4724 1036
rect 4756 1004 4804 1036
rect 4836 1004 4884 1036
rect 4916 1004 4964 1036
rect 4996 1004 5044 1036
rect 5076 1004 5124 1036
rect 5156 1004 5204 1036
rect 5236 1004 5284 1036
rect 5316 1004 5364 1036
rect 5396 1004 5444 1036
rect 5476 1004 5524 1036
rect 5556 1004 5604 1036
rect 5636 1004 5684 1036
rect 5716 1004 5764 1036
rect 5796 1004 5844 1036
rect 5876 1004 5924 1036
rect 5956 1004 6004 1036
rect 6036 1004 6084 1036
rect 6116 1004 6164 1036
rect 6196 1004 6244 1036
rect 6276 1004 6324 1036
rect 6356 1004 6404 1036
rect 6436 1004 6484 1036
rect 6516 1004 6564 1036
rect 6596 1004 6644 1036
rect 6676 1004 6724 1036
rect 6756 1004 6804 1036
rect 6836 1004 6884 1036
rect 6916 1004 6964 1036
rect 6996 1004 7044 1036
rect 7076 1004 7124 1036
rect 7156 1004 7204 1036
rect 7236 1004 7284 1036
rect 7316 1004 7364 1036
rect 7396 1004 7444 1036
rect 7476 1004 7524 1036
rect 7556 1004 7604 1036
rect 7636 1004 7684 1036
rect 7716 1004 7764 1036
rect 7796 1004 7844 1036
rect 7876 1004 7924 1036
rect 7956 1004 8004 1036
rect 8036 1004 8084 1036
rect 8116 1004 8164 1036
rect 8196 1004 8244 1036
rect 8276 1004 8324 1036
rect 8356 1004 8404 1036
rect 8436 1004 8484 1036
rect 8516 1004 8564 1036
rect 8596 1004 8644 1036
rect 8676 1004 8724 1036
rect 8756 1004 8804 1036
rect 8836 1004 8884 1036
rect 8916 1004 8964 1036
rect 8996 1004 9044 1036
rect 9076 1004 9124 1036
rect 9156 1004 9204 1036
rect 9236 1004 9284 1036
rect 9316 1004 9364 1036
rect 9396 1004 9444 1036
rect 9476 1004 9524 1036
rect 9556 1004 9604 1036
rect 9636 1004 9684 1036
rect 9716 1004 9764 1036
rect 9796 1004 9844 1036
rect 9876 1004 9924 1036
rect 9956 1004 10004 1036
rect 10036 1004 10084 1036
rect 10116 1004 10164 1036
rect 10196 1004 10244 1036
rect 10276 1004 10324 1036
rect 10356 1004 10404 1036
rect 10436 1004 10484 1036
rect 10516 1004 10644 1036
rect 10676 1004 10804 1036
rect 10836 1004 10964 1036
rect 10996 1004 11000 1036
rect -720 1000 11000 1004
rect -720 956 11000 960
rect -720 924 -716 956
rect -684 924 -556 956
rect -524 924 -396 956
rect -364 924 -316 956
rect -284 924 -236 956
rect -204 924 -156 956
rect -124 924 -76 956
rect -44 924 4 956
rect 36 924 84 956
rect 116 924 164 956
rect 196 924 244 956
rect 276 924 324 956
rect 356 924 404 956
rect 436 924 484 956
rect 516 924 564 956
rect 596 924 644 956
rect 676 924 724 956
rect 756 924 804 956
rect 836 924 884 956
rect 916 924 964 956
rect 996 924 1044 956
rect 1076 924 1124 956
rect 1156 924 1204 956
rect 1236 924 1284 956
rect 1316 924 1364 956
rect 1396 924 1444 956
rect 1476 924 1524 956
rect 1556 924 1604 956
rect 1636 924 1684 956
rect 1716 924 1764 956
rect 1796 924 1844 956
rect 1876 924 1924 956
rect 1956 924 2004 956
rect 2036 924 2084 956
rect 2116 924 2164 956
rect 2196 924 2244 956
rect 2276 924 2324 956
rect 2356 924 2404 956
rect 2436 924 2484 956
rect 2516 924 2564 956
rect 2596 924 2644 956
rect 2676 924 2724 956
rect 2756 924 2804 956
rect 2836 924 2884 956
rect 2916 924 2964 956
rect 2996 924 3044 956
rect 3076 924 3124 956
rect 3156 924 3204 956
rect 3236 924 3284 956
rect 3316 924 3364 956
rect 3396 924 3444 956
rect 3476 924 3524 956
rect 3556 924 3604 956
rect 3636 924 3684 956
rect 3716 924 3764 956
rect 3796 924 3844 956
rect 3876 924 3924 956
rect 3956 924 4004 956
rect 4036 924 4084 956
rect 4116 924 4164 956
rect 4196 924 4244 956
rect 4276 924 4324 956
rect 4356 924 4404 956
rect 4436 924 4484 956
rect 4516 924 4564 956
rect 4596 924 4644 956
rect 4676 924 4724 956
rect 4756 924 4804 956
rect 4836 924 4884 956
rect 4916 924 4964 956
rect 4996 924 5044 956
rect 5076 924 5124 956
rect 5156 924 5204 956
rect 5236 924 5284 956
rect 5316 924 5364 956
rect 5396 924 5444 956
rect 5476 924 5524 956
rect 5556 924 5604 956
rect 5636 924 5684 956
rect 5716 924 5764 956
rect 5796 924 5844 956
rect 5876 924 5924 956
rect 5956 924 6004 956
rect 6036 924 6084 956
rect 6116 924 6164 956
rect 6196 924 6244 956
rect 6276 924 6324 956
rect 6356 924 6404 956
rect 6436 924 6484 956
rect 6516 924 6564 956
rect 6596 924 6644 956
rect 6676 924 6724 956
rect 6756 924 6804 956
rect 6836 924 6884 956
rect 6916 924 6964 956
rect 6996 924 7044 956
rect 7076 924 7124 956
rect 7156 924 7204 956
rect 7236 924 7284 956
rect 7316 924 7364 956
rect 7396 924 7444 956
rect 7476 924 7524 956
rect 7556 924 7604 956
rect 7636 924 7684 956
rect 7716 924 7764 956
rect 7796 924 7844 956
rect 7876 924 7924 956
rect 7956 924 8004 956
rect 8036 924 8084 956
rect 8116 924 8164 956
rect 8196 924 8244 956
rect 8276 924 8324 956
rect 8356 924 8404 956
rect 8436 924 8484 956
rect 8516 924 8564 956
rect 8596 924 8644 956
rect 8676 924 8724 956
rect 8756 924 8804 956
rect 8836 924 8884 956
rect 8916 924 8964 956
rect 8996 924 9044 956
rect 9076 924 9124 956
rect 9156 924 9204 956
rect 9236 924 9284 956
rect 9316 924 9364 956
rect 9396 924 9444 956
rect 9476 924 9524 956
rect 9556 924 9604 956
rect 9636 924 9684 956
rect 9716 924 9764 956
rect 9796 924 9844 956
rect 9876 924 9924 956
rect 9956 924 10004 956
rect 10036 924 10084 956
rect 10116 924 10164 956
rect 10196 924 10244 956
rect 10276 924 10324 956
rect 10356 924 10404 956
rect 10436 924 10484 956
rect 10516 924 10644 956
rect 10676 924 10804 956
rect 10836 924 10964 956
rect 10996 924 11000 956
rect -720 920 11000 924
rect -720 876 11000 880
rect -720 844 -716 876
rect -684 844 -556 876
rect -524 844 -396 876
rect -364 844 -316 876
rect -284 844 -236 876
rect -204 844 -156 876
rect -124 844 -76 876
rect -44 844 4 876
rect 36 844 84 876
rect 116 844 164 876
rect 196 844 244 876
rect 276 844 324 876
rect 356 844 404 876
rect 436 844 484 876
rect 516 844 564 876
rect 596 844 644 876
rect 676 844 724 876
rect 756 844 804 876
rect 836 844 884 876
rect 916 844 964 876
rect 996 844 1044 876
rect 1076 844 1124 876
rect 1156 844 1204 876
rect 1236 844 1284 876
rect 1316 844 1364 876
rect 1396 844 1444 876
rect 1476 844 1524 876
rect 1556 844 1604 876
rect 1636 844 1684 876
rect 1716 844 1764 876
rect 1796 844 1844 876
rect 1876 844 1924 876
rect 1956 844 2004 876
rect 2036 844 2084 876
rect 2116 844 2164 876
rect 2196 844 2244 876
rect 2276 844 2324 876
rect 2356 844 2404 876
rect 2436 844 2484 876
rect 2516 844 2564 876
rect 2596 844 2644 876
rect 2676 844 2724 876
rect 2756 844 2804 876
rect 2836 844 2884 876
rect 2916 844 2964 876
rect 2996 844 3044 876
rect 3076 844 3124 876
rect 3156 844 3204 876
rect 3236 844 3284 876
rect 3316 844 3364 876
rect 3396 844 3444 876
rect 3476 844 3524 876
rect 3556 844 3604 876
rect 3636 844 3684 876
rect 3716 844 3764 876
rect 3796 844 3844 876
rect 3876 844 3924 876
rect 3956 844 4004 876
rect 4036 844 4084 876
rect 4116 844 4164 876
rect 4196 844 4244 876
rect 4276 844 4324 876
rect 4356 844 4404 876
rect 4436 844 4484 876
rect 4516 844 4564 876
rect 4596 844 4644 876
rect 4676 844 4724 876
rect 4756 844 4804 876
rect 4836 844 4884 876
rect 4916 844 4964 876
rect 4996 844 5044 876
rect 5076 844 5124 876
rect 5156 844 5204 876
rect 5236 844 5284 876
rect 5316 844 5364 876
rect 5396 844 5444 876
rect 5476 844 5524 876
rect 5556 844 5604 876
rect 5636 844 5684 876
rect 5716 844 5764 876
rect 5796 844 5844 876
rect 5876 844 5924 876
rect 5956 844 6004 876
rect 6036 844 6084 876
rect 6116 844 6164 876
rect 6196 844 6244 876
rect 6276 844 6324 876
rect 6356 844 6404 876
rect 6436 844 6484 876
rect 6516 844 6564 876
rect 6596 844 6644 876
rect 6676 844 6724 876
rect 6756 844 6804 876
rect 6836 844 6884 876
rect 6916 844 6964 876
rect 6996 844 7044 876
rect 7076 844 7124 876
rect 7156 844 7204 876
rect 7236 844 7284 876
rect 7316 844 7364 876
rect 7396 844 7444 876
rect 7476 844 7524 876
rect 7556 844 7604 876
rect 7636 844 7684 876
rect 7716 844 7764 876
rect 7796 844 7844 876
rect 7876 844 7924 876
rect 7956 844 8004 876
rect 8036 844 8084 876
rect 8116 844 8164 876
rect 8196 844 8244 876
rect 8276 844 8324 876
rect 8356 844 8404 876
rect 8436 844 8484 876
rect 8516 844 8564 876
rect 8596 844 8644 876
rect 8676 844 8724 876
rect 8756 844 8804 876
rect 8836 844 8884 876
rect 8916 844 8964 876
rect 8996 844 9044 876
rect 9076 844 9124 876
rect 9156 844 9204 876
rect 9236 844 9284 876
rect 9316 844 9364 876
rect 9396 844 9444 876
rect 9476 844 9524 876
rect 9556 844 9604 876
rect 9636 844 9684 876
rect 9716 844 9764 876
rect 9796 844 9844 876
rect 9876 844 9924 876
rect 9956 844 10004 876
rect 10036 844 10084 876
rect 10116 844 10164 876
rect 10196 844 10244 876
rect 10276 844 10324 876
rect 10356 844 10404 876
rect 10436 844 10484 876
rect 10516 844 10644 876
rect 10676 844 10804 876
rect 10836 844 10964 876
rect 10996 844 11000 876
rect -720 840 11000 844
rect -720 796 10600 800
rect -720 764 -716 796
rect -684 764 -556 796
rect -524 764 -396 796
rect -364 764 -316 796
rect -284 764 -236 796
rect -204 764 -156 796
rect -124 764 -76 796
rect -44 764 4 796
rect 36 764 84 796
rect 116 764 164 796
rect 196 764 244 796
rect 276 764 324 796
rect 356 764 404 796
rect 436 764 484 796
rect 516 764 564 796
rect 596 764 644 796
rect 676 764 724 796
rect 756 764 804 796
rect 836 764 884 796
rect 916 764 964 796
rect 996 764 1044 796
rect 1076 764 1124 796
rect 1156 764 1204 796
rect 1236 764 1284 796
rect 1316 764 1364 796
rect 1396 764 1444 796
rect 1476 764 1524 796
rect 1556 764 1604 796
rect 1636 764 1684 796
rect 1716 764 1764 796
rect 1796 764 1844 796
rect 1876 764 1924 796
rect 1956 764 2004 796
rect 2036 764 2084 796
rect 2116 764 2164 796
rect 2196 764 2244 796
rect 2276 764 2324 796
rect 2356 764 2404 796
rect 2436 764 2484 796
rect 2516 764 2564 796
rect 2596 764 2644 796
rect 2676 764 2724 796
rect 2756 764 2804 796
rect 2836 764 2884 796
rect 2916 764 2964 796
rect 2996 764 3044 796
rect 3076 764 3124 796
rect 3156 764 3204 796
rect 3236 764 3284 796
rect 3316 764 3364 796
rect 3396 764 3444 796
rect 3476 764 3524 796
rect 3556 764 3604 796
rect 3636 764 3684 796
rect 3716 764 3764 796
rect 3796 764 3844 796
rect 3876 764 3924 796
rect 3956 764 4004 796
rect 4036 764 4084 796
rect 4116 764 4164 796
rect 4196 764 4244 796
rect 4276 764 4324 796
rect 4356 764 4404 796
rect 4436 764 4484 796
rect 4516 764 4564 796
rect 4596 764 4644 796
rect 4676 764 4724 796
rect 4756 764 4804 796
rect 4836 764 4884 796
rect 4916 764 4964 796
rect 4996 764 5044 796
rect 5076 764 5124 796
rect 5156 764 5204 796
rect 5236 764 5284 796
rect 5316 764 5364 796
rect 5396 764 5444 796
rect 5476 764 5524 796
rect 5556 764 5604 796
rect 5636 764 5684 796
rect 5716 764 5764 796
rect 5796 764 5844 796
rect 5876 764 5924 796
rect 5956 764 6004 796
rect 6036 764 6084 796
rect 6116 764 6164 796
rect 6196 764 6244 796
rect 6276 764 6324 796
rect 6356 764 6404 796
rect 6436 764 6484 796
rect 6516 764 6564 796
rect 6596 764 6644 796
rect 6676 764 6724 796
rect 6756 764 6804 796
rect 6836 764 6884 796
rect 6916 764 6964 796
rect 6996 764 7044 796
rect 7076 764 7124 796
rect 7156 764 7204 796
rect 7236 764 7284 796
rect 7316 764 7364 796
rect 7396 764 7444 796
rect 7476 764 7524 796
rect 7556 764 7604 796
rect 7636 764 7684 796
rect 7716 764 7764 796
rect 7796 764 7844 796
rect 7876 764 7924 796
rect 7956 764 8004 796
rect 8036 764 8084 796
rect 8116 764 8164 796
rect 8196 764 8244 796
rect 8276 764 8324 796
rect 8356 764 8404 796
rect 8436 764 8484 796
rect 8516 764 8564 796
rect 8596 764 8644 796
rect 8676 764 8724 796
rect 8756 764 8804 796
rect 8836 764 8884 796
rect 8916 764 8964 796
rect 8996 764 9044 796
rect 9076 764 9124 796
rect 9156 764 9204 796
rect 9236 764 9284 796
rect 9316 764 9364 796
rect 9396 764 9444 796
rect 9476 764 9524 796
rect 9556 764 9604 796
rect 9636 764 9684 796
rect 9716 764 9764 796
rect 9796 764 9844 796
rect 9876 764 9924 796
rect 9956 764 10004 796
rect 10036 764 10084 796
rect 10116 764 10164 796
rect 10196 764 10244 796
rect 10276 764 10324 796
rect 10356 764 10404 796
rect 10436 764 10484 796
rect 10516 764 10600 796
rect -720 760 10600 764
rect 10640 796 11000 800
rect 10640 764 10644 796
rect 10676 764 10804 796
rect 10836 764 10964 796
rect 10996 764 11000 796
rect 10640 760 11000 764
rect -720 716 10600 720
rect -720 684 -716 716
rect -684 684 -556 716
rect -524 684 -396 716
rect -364 684 -316 716
rect -284 684 -236 716
rect -204 684 -156 716
rect -124 684 -76 716
rect -44 684 4 716
rect 36 684 84 716
rect 116 684 164 716
rect 196 684 244 716
rect 276 684 324 716
rect 356 684 404 716
rect 436 684 484 716
rect 516 684 564 716
rect 596 684 644 716
rect 676 684 724 716
rect 756 684 804 716
rect 836 684 884 716
rect 916 684 964 716
rect 996 684 1044 716
rect 1076 684 1124 716
rect 1156 684 1204 716
rect 1236 684 1284 716
rect 1316 684 1364 716
rect 1396 684 1444 716
rect 1476 684 1524 716
rect 1556 684 1604 716
rect 1636 684 1684 716
rect 1716 684 1764 716
rect 1796 684 1844 716
rect 1876 684 1924 716
rect 1956 684 2004 716
rect 2036 684 2084 716
rect 2116 684 2164 716
rect 2196 684 2244 716
rect 2276 684 2324 716
rect 2356 684 2404 716
rect 2436 684 2484 716
rect 2516 684 2564 716
rect 2596 684 2644 716
rect 2676 684 2724 716
rect 2756 684 2804 716
rect 2836 684 2884 716
rect 2916 684 2964 716
rect 2996 684 3044 716
rect 3076 684 3124 716
rect 3156 684 3204 716
rect 3236 684 3284 716
rect 3316 684 3364 716
rect 3396 684 3444 716
rect 3476 684 3524 716
rect 3556 684 3604 716
rect 3636 684 3684 716
rect 3716 684 3764 716
rect 3796 684 3844 716
rect 3876 684 3924 716
rect 3956 684 4004 716
rect 4036 684 4084 716
rect 4116 684 4164 716
rect 4196 684 4244 716
rect 4276 684 4324 716
rect 4356 684 4404 716
rect 4436 684 4484 716
rect 4516 684 4564 716
rect 4596 684 4644 716
rect 4676 684 4724 716
rect 4756 684 4804 716
rect 4836 684 4884 716
rect 4916 684 4964 716
rect 4996 684 5044 716
rect 5076 684 5124 716
rect 5156 684 5204 716
rect 5236 684 5284 716
rect 5316 684 5364 716
rect 5396 684 5444 716
rect 5476 684 5524 716
rect 5556 684 5604 716
rect 5636 684 5684 716
rect 5716 684 5764 716
rect 5796 684 5844 716
rect 5876 684 5924 716
rect 5956 684 6004 716
rect 6036 684 6084 716
rect 6116 684 6164 716
rect 6196 684 6244 716
rect 6276 684 6324 716
rect 6356 684 6404 716
rect 6436 684 6484 716
rect 6516 684 6564 716
rect 6596 684 6644 716
rect 6676 684 6724 716
rect 6756 684 6804 716
rect 6836 684 6884 716
rect 6916 684 6964 716
rect 6996 684 7044 716
rect 7076 684 7124 716
rect 7156 684 7204 716
rect 7236 684 7284 716
rect 7316 684 7364 716
rect 7396 684 7444 716
rect 7476 684 7524 716
rect 7556 684 7604 716
rect 7636 684 7684 716
rect 7716 684 7764 716
rect 7796 684 7844 716
rect 7876 684 7924 716
rect 7956 684 8004 716
rect 8036 684 8084 716
rect 8116 684 8164 716
rect 8196 684 8244 716
rect 8276 684 8324 716
rect 8356 684 8404 716
rect 8436 684 8484 716
rect 8516 684 8564 716
rect 8596 684 8644 716
rect 8676 684 8724 716
rect 8756 684 8804 716
rect 8836 684 8884 716
rect 8916 684 8964 716
rect 8996 684 9044 716
rect 9076 684 9124 716
rect 9156 684 9204 716
rect 9236 684 9284 716
rect 9316 684 9364 716
rect 9396 684 9444 716
rect 9476 684 9524 716
rect 9556 684 9604 716
rect 9636 684 9684 716
rect 9716 684 9764 716
rect 9796 684 9844 716
rect 9876 684 9924 716
rect 9956 684 10004 716
rect 10036 684 10084 716
rect 10116 684 10164 716
rect 10196 684 10244 716
rect 10276 684 10324 716
rect 10356 684 10404 716
rect 10436 684 10484 716
rect 10516 684 10600 716
rect -720 680 10600 684
rect 10640 716 11000 720
rect 10640 684 10644 716
rect 10676 684 10804 716
rect 10836 684 10964 716
rect 10996 684 11000 716
rect 10640 680 11000 684
rect -720 636 11000 640
rect -720 604 -716 636
rect -684 604 -556 636
rect -524 604 -396 636
rect -364 604 -316 636
rect -284 604 -236 636
rect -204 604 -156 636
rect -124 604 -76 636
rect -44 604 4 636
rect 36 604 84 636
rect 116 604 164 636
rect 196 604 244 636
rect 276 604 324 636
rect 356 604 404 636
rect 436 604 484 636
rect 516 604 564 636
rect 596 604 644 636
rect 676 604 724 636
rect 756 604 804 636
rect 836 604 884 636
rect 916 604 964 636
rect 996 604 1044 636
rect 1076 604 1124 636
rect 1156 604 1204 636
rect 1236 604 1284 636
rect 1316 604 1364 636
rect 1396 604 1444 636
rect 1476 604 1524 636
rect 1556 604 1604 636
rect 1636 604 1684 636
rect 1716 604 1764 636
rect 1796 604 1844 636
rect 1876 604 1924 636
rect 1956 604 2004 636
rect 2036 604 2084 636
rect 2116 604 2164 636
rect 2196 604 2244 636
rect 2276 604 2324 636
rect 2356 604 2404 636
rect 2436 604 2484 636
rect 2516 604 2564 636
rect 2596 604 2644 636
rect 2676 604 2724 636
rect 2756 604 2804 636
rect 2836 604 2884 636
rect 2916 604 2964 636
rect 2996 604 3044 636
rect 3076 604 3124 636
rect 3156 604 3204 636
rect 3236 604 3284 636
rect 3316 604 3364 636
rect 3396 604 3444 636
rect 3476 604 3524 636
rect 3556 604 3604 636
rect 3636 604 3684 636
rect 3716 604 3764 636
rect 3796 604 3844 636
rect 3876 604 3924 636
rect 3956 604 4004 636
rect 4036 604 4084 636
rect 4116 604 4164 636
rect 4196 604 4244 636
rect 4276 604 4324 636
rect 4356 604 4404 636
rect 4436 604 4484 636
rect 4516 604 4564 636
rect 4596 604 4644 636
rect 4676 604 4724 636
rect 4756 604 4804 636
rect 4836 604 4884 636
rect 4916 604 4964 636
rect 4996 604 5044 636
rect 5076 604 5124 636
rect 5156 604 5204 636
rect 5236 604 5284 636
rect 5316 604 5364 636
rect 5396 604 5444 636
rect 5476 604 5524 636
rect 5556 604 5604 636
rect 5636 604 5684 636
rect 5716 604 5764 636
rect 5796 604 5844 636
rect 5876 604 5924 636
rect 5956 604 6004 636
rect 6036 604 6084 636
rect 6116 604 6164 636
rect 6196 604 6244 636
rect 6276 604 6324 636
rect 6356 604 6404 636
rect 6436 604 6484 636
rect 6516 604 6564 636
rect 6596 604 6644 636
rect 6676 604 6724 636
rect 6756 604 6804 636
rect 6836 604 6884 636
rect 6916 604 6964 636
rect 6996 604 7044 636
rect 7076 604 7124 636
rect 7156 604 7204 636
rect 7236 604 7284 636
rect 7316 604 7364 636
rect 7396 604 7444 636
rect 7476 604 7524 636
rect 7556 604 7604 636
rect 7636 604 7684 636
rect 7716 604 7764 636
rect 7796 604 7844 636
rect 7876 604 7924 636
rect 7956 604 8004 636
rect 8036 604 8084 636
rect 8116 604 8164 636
rect 8196 604 8244 636
rect 8276 604 8324 636
rect 8356 604 8404 636
rect 8436 604 8484 636
rect 8516 604 8564 636
rect 8596 604 8644 636
rect 8676 604 8724 636
rect 8756 604 8804 636
rect 8836 604 8884 636
rect 8916 604 8964 636
rect 8996 604 9044 636
rect 9076 604 9124 636
rect 9156 604 9204 636
rect 9236 604 9284 636
rect 9316 604 9364 636
rect 9396 604 9444 636
rect 9476 604 9524 636
rect 9556 604 9604 636
rect 9636 604 9684 636
rect 9716 604 9764 636
rect 9796 604 9844 636
rect 9876 604 9924 636
rect 9956 604 10004 636
rect 10036 604 10084 636
rect 10116 604 10164 636
rect 10196 604 10244 636
rect 10276 604 10324 636
rect 10356 604 10404 636
rect 10436 604 10484 636
rect 10516 604 10644 636
rect 10676 604 10804 636
rect 10836 604 10964 636
rect 10996 604 11000 636
rect -720 600 11000 604
rect -720 556 11000 560
rect -720 524 -716 556
rect -684 524 -556 556
rect -524 524 -396 556
rect -364 524 -316 556
rect -284 524 -236 556
rect -204 524 -156 556
rect -124 524 -76 556
rect -44 524 4 556
rect 36 524 84 556
rect 116 524 164 556
rect 196 524 244 556
rect 276 524 324 556
rect 356 524 404 556
rect 436 524 484 556
rect 516 524 564 556
rect 596 524 644 556
rect 676 524 724 556
rect 756 524 804 556
rect 836 524 884 556
rect 916 524 964 556
rect 996 524 1044 556
rect 1076 524 1124 556
rect 1156 524 1204 556
rect 1236 524 1284 556
rect 1316 524 1364 556
rect 1396 524 1444 556
rect 1476 524 1524 556
rect 1556 524 1604 556
rect 1636 524 1684 556
rect 1716 524 1764 556
rect 1796 524 1844 556
rect 1876 524 1924 556
rect 1956 524 2004 556
rect 2036 524 2084 556
rect 2116 524 2164 556
rect 2196 524 2244 556
rect 2276 524 2324 556
rect 2356 524 2404 556
rect 2436 524 2484 556
rect 2516 524 2564 556
rect 2596 524 2644 556
rect 2676 524 2724 556
rect 2756 524 2804 556
rect 2836 524 2884 556
rect 2916 524 2964 556
rect 2996 524 3044 556
rect 3076 524 3124 556
rect 3156 524 3204 556
rect 3236 524 3284 556
rect 3316 524 3364 556
rect 3396 524 3444 556
rect 3476 524 3524 556
rect 3556 524 3604 556
rect 3636 524 3684 556
rect 3716 524 3764 556
rect 3796 524 3844 556
rect 3876 524 3924 556
rect 3956 524 4004 556
rect 4036 524 4084 556
rect 4116 524 4164 556
rect 4196 524 4244 556
rect 4276 524 4324 556
rect 4356 524 4404 556
rect 4436 524 4484 556
rect 4516 524 4564 556
rect 4596 524 4644 556
rect 4676 524 4724 556
rect 4756 524 4804 556
rect 4836 524 4884 556
rect 4916 524 4964 556
rect 4996 524 5044 556
rect 5076 524 5124 556
rect 5156 524 5204 556
rect 5236 524 5284 556
rect 5316 524 5364 556
rect 5396 524 5444 556
rect 5476 524 5524 556
rect 5556 524 5604 556
rect 5636 524 5684 556
rect 5716 524 5764 556
rect 5796 524 5844 556
rect 5876 524 5924 556
rect 5956 524 6004 556
rect 6036 524 6084 556
rect 6116 524 6164 556
rect 6196 524 6244 556
rect 6276 524 6324 556
rect 6356 524 6404 556
rect 6436 524 6484 556
rect 6516 524 6564 556
rect 6596 524 6644 556
rect 6676 524 6724 556
rect 6756 524 6804 556
rect 6836 524 6884 556
rect 6916 524 6964 556
rect 6996 524 7044 556
rect 7076 524 7124 556
rect 7156 524 7204 556
rect 7236 524 7284 556
rect 7316 524 7364 556
rect 7396 524 7444 556
rect 7476 524 7524 556
rect 7556 524 7604 556
rect 7636 524 7684 556
rect 7716 524 7764 556
rect 7796 524 7844 556
rect 7876 524 7924 556
rect 7956 524 8004 556
rect 8036 524 8084 556
rect 8116 524 8164 556
rect 8196 524 8244 556
rect 8276 524 8324 556
rect 8356 524 8404 556
rect 8436 524 8484 556
rect 8516 524 8564 556
rect 8596 524 8644 556
rect 8676 524 8724 556
rect 8756 524 8804 556
rect 8836 524 8884 556
rect 8916 524 8964 556
rect 8996 524 9044 556
rect 9076 524 9124 556
rect 9156 524 9204 556
rect 9236 524 9284 556
rect 9316 524 9364 556
rect 9396 524 9444 556
rect 9476 524 9524 556
rect 9556 524 9604 556
rect 9636 524 9684 556
rect 9716 524 9764 556
rect 9796 524 9844 556
rect 9876 524 9924 556
rect 9956 524 10004 556
rect 10036 524 10084 556
rect 10116 524 10164 556
rect 10196 524 10244 556
rect 10276 524 10324 556
rect 10356 524 10404 556
rect 10436 524 10484 556
rect 10516 524 10644 556
rect 10676 524 10804 556
rect 10836 524 10964 556
rect 10996 524 11000 556
rect -720 520 11000 524
rect -720 476 10600 480
rect -720 444 -716 476
rect -684 444 -556 476
rect -524 444 -396 476
rect -364 444 -316 476
rect -284 444 -236 476
rect -204 444 -156 476
rect -124 444 -76 476
rect -44 444 4 476
rect 36 444 84 476
rect 116 444 164 476
rect 196 444 244 476
rect 276 444 324 476
rect 356 444 404 476
rect 436 444 484 476
rect 516 444 564 476
rect 596 444 644 476
rect 676 444 724 476
rect 756 444 804 476
rect 836 444 884 476
rect 916 444 964 476
rect 996 444 1044 476
rect 1076 444 1124 476
rect 1156 444 1204 476
rect 1236 444 1284 476
rect 1316 444 1364 476
rect 1396 444 1444 476
rect 1476 444 1524 476
rect 1556 444 1604 476
rect 1636 444 1684 476
rect 1716 444 1764 476
rect 1796 444 1844 476
rect 1876 444 1924 476
rect 1956 444 2004 476
rect 2036 444 2084 476
rect 2116 444 2164 476
rect 2196 444 2244 476
rect 2276 444 2324 476
rect 2356 444 2404 476
rect 2436 444 2484 476
rect 2516 444 2564 476
rect 2596 444 2644 476
rect 2676 444 2724 476
rect 2756 444 2804 476
rect 2836 444 2884 476
rect 2916 444 2964 476
rect 2996 444 3044 476
rect 3076 444 3124 476
rect 3156 444 3204 476
rect 3236 444 3284 476
rect 3316 444 3364 476
rect 3396 444 3444 476
rect 3476 444 3524 476
rect 3556 444 3604 476
rect 3636 444 3684 476
rect 3716 444 3764 476
rect 3796 444 3844 476
rect 3876 444 3924 476
rect 3956 444 4004 476
rect 4036 444 4084 476
rect 4116 444 4164 476
rect 4196 444 4244 476
rect 4276 444 4324 476
rect 4356 444 4404 476
rect 4436 444 4484 476
rect 4516 444 4564 476
rect 4596 444 4644 476
rect 4676 444 4724 476
rect 4756 444 4804 476
rect 4836 444 4884 476
rect 4916 444 4964 476
rect 4996 444 5044 476
rect 5076 444 5124 476
rect 5156 444 5204 476
rect 5236 444 5284 476
rect 5316 444 5364 476
rect 5396 444 5444 476
rect 5476 444 5524 476
rect 5556 444 5604 476
rect 5636 444 5684 476
rect 5716 444 5764 476
rect 5796 444 5844 476
rect 5876 444 5924 476
rect 5956 444 6004 476
rect 6036 444 6084 476
rect 6116 444 6164 476
rect 6196 444 6244 476
rect 6276 444 6324 476
rect 6356 444 6404 476
rect 6436 444 6484 476
rect 6516 444 6564 476
rect 6596 444 6644 476
rect 6676 444 6724 476
rect 6756 444 6804 476
rect 6836 444 6884 476
rect 6916 444 6964 476
rect 6996 444 7044 476
rect 7076 444 7124 476
rect 7156 444 7204 476
rect 7236 444 7284 476
rect 7316 444 7364 476
rect 7396 444 7444 476
rect 7476 444 7524 476
rect 7556 444 7604 476
rect 7636 444 7684 476
rect 7716 444 7764 476
rect 7796 444 7844 476
rect 7876 444 7924 476
rect 7956 444 8004 476
rect 8036 444 8084 476
rect 8116 444 8164 476
rect 8196 444 8244 476
rect 8276 444 8324 476
rect 8356 444 8404 476
rect 8436 444 8484 476
rect 8516 444 8564 476
rect 8596 444 8644 476
rect 8676 444 8724 476
rect 8756 444 8804 476
rect 8836 444 8884 476
rect 8916 444 8964 476
rect 8996 444 9044 476
rect 9076 444 9124 476
rect 9156 444 9204 476
rect 9236 444 9284 476
rect 9316 444 9364 476
rect 9396 444 9444 476
rect 9476 444 9524 476
rect 9556 444 9604 476
rect 9636 444 9684 476
rect 9716 444 9764 476
rect 9796 444 9844 476
rect 9876 444 9924 476
rect 9956 444 10004 476
rect 10036 444 10084 476
rect 10116 444 10164 476
rect 10196 444 10244 476
rect 10276 444 10324 476
rect 10356 444 10404 476
rect 10436 444 10484 476
rect 10516 444 10600 476
rect -720 440 10600 444
rect 10640 476 11000 480
rect 10640 444 10644 476
rect 10676 444 10804 476
rect 10836 444 10964 476
rect 10996 444 11000 476
rect 10640 440 11000 444
rect -720 396 11000 400
rect -720 364 -716 396
rect -684 364 -556 396
rect -524 364 -396 396
rect -364 364 -316 396
rect -284 364 -236 396
rect -204 364 -156 396
rect -124 364 -76 396
rect -44 364 4 396
rect 36 364 84 396
rect 116 364 164 396
rect 196 364 244 396
rect 276 364 324 396
rect 356 364 404 396
rect 436 364 484 396
rect 516 364 564 396
rect 596 364 644 396
rect 676 364 724 396
rect 756 364 804 396
rect 836 364 884 396
rect 916 364 964 396
rect 996 364 1044 396
rect 1076 364 1124 396
rect 1156 364 1204 396
rect 1236 364 1284 396
rect 1316 364 1364 396
rect 1396 364 1444 396
rect 1476 364 1524 396
rect 1556 364 1604 396
rect 1636 364 1684 396
rect 1716 364 1764 396
rect 1796 364 1844 396
rect 1876 364 1924 396
rect 1956 364 2004 396
rect 2036 364 2084 396
rect 2116 364 2164 396
rect 2196 364 2244 396
rect 2276 364 2324 396
rect 2356 364 2404 396
rect 2436 364 2484 396
rect 2516 364 2564 396
rect 2596 364 2644 396
rect 2676 364 2724 396
rect 2756 364 2804 396
rect 2836 364 2884 396
rect 2916 364 2964 396
rect 2996 364 3044 396
rect 3076 364 3124 396
rect 3156 364 3204 396
rect 3236 364 3284 396
rect 3316 364 3364 396
rect 3396 364 3444 396
rect 3476 364 3524 396
rect 3556 364 3604 396
rect 3636 364 3684 396
rect 3716 364 3764 396
rect 3796 364 3844 396
rect 3876 364 3924 396
rect 3956 364 4004 396
rect 4036 364 4084 396
rect 4116 364 4164 396
rect 4196 364 4244 396
rect 4276 364 4324 396
rect 4356 364 4404 396
rect 4436 364 4484 396
rect 4516 364 4564 396
rect 4596 364 4644 396
rect 4676 364 4724 396
rect 4756 364 4804 396
rect 4836 364 4884 396
rect 4916 364 4964 396
rect 4996 364 5044 396
rect 5076 364 5124 396
rect 5156 364 5204 396
rect 5236 364 5284 396
rect 5316 364 5364 396
rect 5396 364 5444 396
rect 5476 364 5524 396
rect 5556 364 5604 396
rect 5636 364 5684 396
rect 5716 364 5764 396
rect 5796 364 5844 396
rect 5876 364 5924 396
rect 5956 364 6004 396
rect 6036 364 6084 396
rect 6116 364 6164 396
rect 6196 364 6244 396
rect 6276 364 6324 396
rect 6356 364 6404 396
rect 6436 364 6484 396
rect 6516 364 6564 396
rect 6596 364 6644 396
rect 6676 364 6724 396
rect 6756 364 6804 396
rect 6836 364 6884 396
rect 6916 364 6964 396
rect 6996 364 7044 396
rect 7076 364 7124 396
rect 7156 364 7204 396
rect 7236 364 7284 396
rect 7316 364 7364 396
rect 7396 364 7444 396
rect 7476 364 7524 396
rect 7556 364 7604 396
rect 7636 364 7684 396
rect 7716 364 7764 396
rect 7796 364 7844 396
rect 7876 364 7924 396
rect 7956 364 8004 396
rect 8036 364 8084 396
rect 8116 364 8164 396
rect 8196 364 8244 396
rect 8276 364 8324 396
rect 8356 364 8404 396
rect 8436 364 8484 396
rect 8516 364 8564 396
rect 8596 364 8644 396
rect 8676 364 8724 396
rect 8756 364 8804 396
rect 8836 364 8884 396
rect 8916 364 8964 396
rect 8996 364 9044 396
rect 9076 364 9124 396
rect 9156 364 9204 396
rect 9236 364 9284 396
rect 9316 364 9364 396
rect 9396 364 9444 396
rect 9476 364 9524 396
rect 9556 364 9604 396
rect 9636 364 9684 396
rect 9716 364 9764 396
rect 9796 364 9844 396
rect 9876 364 9924 396
rect 9956 364 10004 396
rect 10036 364 10084 396
rect 10116 364 10164 396
rect 10196 364 10244 396
rect 10276 364 10324 396
rect 10356 364 10404 396
rect 10436 364 10484 396
rect 10516 364 10644 396
rect 10676 364 10804 396
rect 10836 364 10964 396
rect 10996 364 11000 396
rect -720 360 11000 364
rect -720 316 -360 320
rect -720 284 -716 316
rect -684 284 -556 316
rect -524 284 -396 316
rect -364 284 -360 316
rect -720 280 -360 284
rect -320 316 11000 320
rect -320 284 -316 316
rect -284 284 -236 316
rect -204 284 -156 316
rect -124 284 -76 316
rect -44 284 4 316
rect 36 284 84 316
rect 116 284 164 316
rect 196 284 244 316
rect 276 284 324 316
rect 356 284 404 316
rect 436 284 484 316
rect 516 284 564 316
rect 596 284 644 316
rect 676 284 724 316
rect 756 284 804 316
rect 836 284 884 316
rect 916 284 964 316
rect 996 284 1044 316
rect 1076 284 1124 316
rect 1156 284 1204 316
rect 1236 284 1284 316
rect 1316 284 1364 316
rect 1396 284 1444 316
rect 1476 284 1524 316
rect 1556 284 1604 316
rect 1636 284 1684 316
rect 1716 284 1764 316
rect 1796 284 1844 316
rect 1876 284 1924 316
rect 1956 284 2004 316
rect 2036 284 2084 316
rect 2116 284 2164 316
rect 2196 284 2244 316
rect 2276 284 2324 316
rect 2356 284 2404 316
rect 2436 284 2484 316
rect 2516 284 2564 316
rect 2596 284 2644 316
rect 2676 284 2724 316
rect 2756 284 2804 316
rect 2836 284 2884 316
rect 2916 284 2964 316
rect 2996 284 3044 316
rect 3076 284 3124 316
rect 3156 284 3204 316
rect 3236 284 3284 316
rect 3316 284 3364 316
rect 3396 284 3444 316
rect 3476 284 3524 316
rect 3556 284 3604 316
rect 3636 284 3684 316
rect 3716 284 3764 316
rect 3796 284 3844 316
rect 3876 284 3924 316
rect 3956 284 4004 316
rect 4036 284 4084 316
rect 4116 284 4164 316
rect 4196 284 4244 316
rect 4276 284 4324 316
rect 4356 284 4404 316
rect 4436 284 4484 316
rect 4516 284 4564 316
rect 4596 284 4644 316
rect 4676 284 4724 316
rect 4756 284 4804 316
rect 4836 284 4884 316
rect 4916 284 4964 316
rect 4996 284 5044 316
rect 5076 284 5124 316
rect 5156 284 5204 316
rect 5236 284 5284 316
rect 5316 284 5364 316
rect 5396 284 5444 316
rect 5476 284 5524 316
rect 5556 284 5604 316
rect 5636 284 5684 316
rect 5716 284 5764 316
rect 5796 284 5844 316
rect 5876 284 5924 316
rect 5956 284 6004 316
rect 6036 284 6084 316
rect 6116 284 6164 316
rect 6196 284 6244 316
rect 6276 284 6324 316
rect 6356 284 6404 316
rect 6436 284 6484 316
rect 6516 284 6564 316
rect 6596 284 6644 316
rect 6676 284 6724 316
rect 6756 284 6804 316
rect 6836 284 6884 316
rect 6916 284 6964 316
rect 6996 284 7044 316
rect 7076 284 7124 316
rect 7156 284 7204 316
rect 7236 284 7284 316
rect 7316 284 7364 316
rect 7396 284 7444 316
rect 7476 284 7524 316
rect 7556 284 7604 316
rect 7636 284 7684 316
rect 7716 284 7764 316
rect 7796 284 7844 316
rect 7876 284 7924 316
rect 7956 284 8004 316
rect 8036 284 8084 316
rect 8116 284 8164 316
rect 8196 284 8244 316
rect 8276 284 8324 316
rect 8356 284 8404 316
rect 8436 284 8484 316
rect 8516 284 8564 316
rect 8596 284 8644 316
rect 8676 284 8724 316
rect 8756 284 8804 316
rect 8836 284 8884 316
rect 8916 284 8964 316
rect 8996 284 9044 316
rect 9076 284 9124 316
rect 9156 284 9204 316
rect 9236 284 9284 316
rect 9316 284 9364 316
rect 9396 284 9444 316
rect 9476 284 9524 316
rect 9556 284 9604 316
rect 9636 284 9684 316
rect 9716 284 9764 316
rect 9796 284 9844 316
rect 9876 284 9924 316
rect 9956 284 10004 316
rect 10036 284 10084 316
rect 10116 284 10164 316
rect 10196 284 10244 316
rect 10276 284 10324 316
rect 10356 284 10404 316
rect 10436 284 10484 316
rect 10516 284 10644 316
rect 10676 284 10804 316
rect 10836 284 10964 316
rect 10996 284 11000 316
rect -320 280 11000 284
rect -720 236 11000 240
rect -720 204 -716 236
rect -684 204 -556 236
rect -524 204 -396 236
rect -364 204 -316 236
rect -284 204 -236 236
rect -204 204 -156 236
rect -124 204 -76 236
rect -44 204 4 236
rect 36 204 84 236
rect 116 204 164 236
rect 196 204 244 236
rect 276 204 324 236
rect 356 204 404 236
rect 436 204 484 236
rect 516 204 564 236
rect 596 204 644 236
rect 676 204 724 236
rect 756 204 804 236
rect 836 204 884 236
rect 916 204 964 236
rect 996 204 1044 236
rect 1076 204 1124 236
rect 1156 204 1204 236
rect 1236 204 1284 236
rect 1316 204 1364 236
rect 1396 204 1444 236
rect 1476 204 1524 236
rect 1556 204 1604 236
rect 1636 204 1684 236
rect 1716 204 1764 236
rect 1796 204 1844 236
rect 1876 204 1924 236
rect 1956 204 2004 236
rect 2036 204 2084 236
rect 2116 204 2164 236
rect 2196 204 2244 236
rect 2276 204 2324 236
rect 2356 204 2404 236
rect 2436 204 2484 236
rect 2516 204 2564 236
rect 2596 204 2644 236
rect 2676 204 2724 236
rect 2756 204 2804 236
rect 2836 204 2884 236
rect 2916 204 2964 236
rect 2996 204 3044 236
rect 3076 204 3124 236
rect 3156 204 3204 236
rect 3236 204 3284 236
rect 3316 204 3364 236
rect 3396 204 3444 236
rect 3476 204 3524 236
rect 3556 204 3604 236
rect 3636 204 3684 236
rect 3716 204 3764 236
rect 3796 204 3844 236
rect 3876 204 3924 236
rect 3956 204 4004 236
rect 4036 204 4084 236
rect 4116 204 4164 236
rect 4196 204 4244 236
rect 4276 204 4324 236
rect 4356 204 4404 236
rect 4436 204 4484 236
rect 4516 204 4564 236
rect 4596 204 4644 236
rect 4676 204 4724 236
rect 4756 204 4804 236
rect 4836 204 4884 236
rect 4916 204 4964 236
rect 4996 204 5044 236
rect 5076 204 5124 236
rect 5156 204 5204 236
rect 5236 204 5284 236
rect 5316 204 5364 236
rect 5396 204 5444 236
rect 5476 204 5524 236
rect 5556 204 5604 236
rect 5636 204 5684 236
rect 5716 204 5764 236
rect 5796 204 5844 236
rect 5876 204 5924 236
rect 5956 204 6004 236
rect 6036 204 6084 236
rect 6116 204 6164 236
rect 6196 204 6244 236
rect 6276 204 6324 236
rect 6356 204 6404 236
rect 6436 204 6484 236
rect 6516 204 6564 236
rect 6596 204 6644 236
rect 6676 204 6724 236
rect 6756 204 6804 236
rect 6836 204 6884 236
rect 6916 204 6964 236
rect 6996 204 7044 236
rect 7076 204 7124 236
rect 7156 204 7204 236
rect 7236 204 7284 236
rect 7316 204 7364 236
rect 7396 204 7444 236
rect 7476 204 7524 236
rect 7556 204 7604 236
rect 7636 204 7684 236
rect 7716 204 7764 236
rect 7796 204 7844 236
rect 7876 204 7924 236
rect 7956 204 8004 236
rect 8036 204 8084 236
rect 8116 204 8164 236
rect 8196 204 8244 236
rect 8276 204 8324 236
rect 8356 204 8404 236
rect 8436 204 8484 236
rect 8516 204 8564 236
rect 8596 204 8644 236
rect 8676 204 8724 236
rect 8756 204 8804 236
rect 8836 204 8884 236
rect 8916 204 8964 236
rect 8996 204 9044 236
rect 9076 204 9124 236
rect 9156 204 9204 236
rect 9236 204 9284 236
rect 9316 204 9364 236
rect 9396 204 9444 236
rect 9476 204 9524 236
rect 9556 204 9604 236
rect 9636 204 9684 236
rect 9716 204 9764 236
rect 9796 204 9844 236
rect 9876 204 9924 236
rect 9956 204 10004 236
rect 10036 204 10084 236
rect 10116 204 10164 236
rect 10196 204 10244 236
rect 10276 204 10324 236
rect 10356 204 10404 236
rect 10436 204 10484 236
rect 10516 204 10644 236
rect 10676 204 10804 236
rect 10836 204 10964 236
rect 10996 204 11000 236
rect -720 200 11000 204
rect -720 156 -360 160
rect -720 124 -716 156
rect -684 124 -556 156
rect -524 124 -396 156
rect -364 124 -360 156
rect -720 120 -360 124
rect -320 156 11000 160
rect -320 124 -316 156
rect -284 124 -236 156
rect -204 124 -156 156
rect -124 124 -76 156
rect -44 124 4 156
rect 36 124 84 156
rect 116 124 164 156
rect 196 124 244 156
rect 276 124 324 156
rect 356 124 404 156
rect 436 124 484 156
rect 516 124 564 156
rect 596 124 644 156
rect 676 124 724 156
rect 756 124 804 156
rect 836 124 884 156
rect 916 124 964 156
rect 996 124 1044 156
rect 1076 124 1124 156
rect 1156 124 1204 156
rect 1236 124 1284 156
rect 1316 124 1364 156
rect 1396 124 1444 156
rect 1476 124 1524 156
rect 1556 124 1604 156
rect 1636 124 1684 156
rect 1716 124 1764 156
rect 1796 124 1844 156
rect 1876 124 1924 156
rect 1956 124 2004 156
rect 2036 124 2084 156
rect 2116 124 2164 156
rect 2196 124 2244 156
rect 2276 124 2324 156
rect 2356 124 2404 156
rect 2436 124 2484 156
rect 2516 124 2564 156
rect 2596 124 2644 156
rect 2676 124 2724 156
rect 2756 124 2804 156
rect 2836 124 2884 156
rect 2916 124 2964 156
rect 2996 124 3044 156
rect 3076 124 3124 156
rect 3156 124 3204 156
rect 3236 124 3284 156
rect 3316 124 3364 156
rect 3396 124 3444 156
rect 3476 124 3524 156
rect 3556 124 3604 156
rect 3636 124 3684 156
rect 3716 124 3764 156
rect 3796 124 3844 156
rect 3876 124 3924 156
rect 3956 124 4004 156
rect 4036 124 4084 156
rect 4116 124 4164 156
rect 4196 124 4244 156
rect 4276 124 4324 156
rect 4356 124 4404 156
rect 4436 124 4484 156
rect 4516 124 4564 156
rect 4596 124 4644 156
rect 4676 124 4724 156
rect 4756 124 4804 156
rect 4836 124 4884 156
rect 4916 124 4964 156
rect 4996 124 5044 156
rect 5076 124 5124 156
rect 5156 124 5204 156
rect 5236 124 5284 156
rect 5316 124 5364 156
rect 5396 124 5444 156
rect 5476 124 5524 156
rect 5556 124 5604 156
rect 5636 124 5684 156
rect 5716 124 5764 156
rect 5796 124 5844 156
rect 5876 124 5924 156
rect 5956 124 6004 156
rect 6036 124 6084 156
rect 6116 124 6164 156
rect 6196 124 6244 156
rect 6276 124 6324 156
rect 6356 124 6404 156
rect 6436 124 6484 156
rect 6516 124 6564 156
rect 6596 124 6644 156
rect 6676 124 6724 156
rect 6756 124 6804 156
rect 6836 124 6884 156
rect 6916 124 6964 156
rect 6996 124 7044 156
rect 7076 124 7124 156
rect 7156 124 7204 156
rect 7236 124 7284 156
rect 7316 124 7364 156
rect 7396 124 7444 156
rect 7476 124 7524 156
rect 7556 124 7604 156
rect 7636 124 7684 156
rect 7716 124 7764 156
rect 7796 124 7844 156
rect 7876 124 7924 156
rect 7956 124 8004 156
rect 8036 124 8084 156
rect 8116 124 8164 156
rect 8196 124 8244 156
rect 8276 124 8324 156
rect 8356 124 8404 156
rect 8436 124 8484 156
rect 8516 124 8564 156
rect 8596 124 8644 156
rect 8676 124 8724 156
rect 8756 124 8804 156
rect 8836 124 8884 156
rect 8916 124 8964 156
rect 8996 124 9044 156
rect 9076 124 9124 156
rect 9156 124 9204 156
rect 9236 124 9284 156
rect 9316 124 9364 156
rect 9396 124 9444 156
rect 9476 124 9524 156
rect 9556 124 9604 156
rect 9636 124 9684 156
rect 9716 124 9764 156
rect 9796 124 9844 156
rect 9876 124 9924 156
rect 9956 124 10004 156
rect 10036 124 10084 156
rect 10116 124 10164 156
rect 10196 124 10244 156
rect 10276 124 10324 156
rect 10356 124 10404 156
rect 10436 124 10484 156
rect 10516 124 10644 156
rect 10676 124 10804 156
rect 10836 124 10964 156
rect 10996 124 11000 156
rect -320 120 11000 124
rect -720 76 11000 80
rect -720 44 -716 76
rect -684 44 -556 76
rect -524 44 -396 76
rect -364 44 -316 76
rect -284 44 -236 76
rect -204 44 -156 76
rect -124 44 -76 76
rect -44 44 4 76
rect 36 44 84 76
rect 116 44 164 76
rect 196 44 244 76
rect 276 44 324 76
rect 356 44 404 76
rect 436 44 484 76
rect 516 44 564 76
rect 596 44 644 76
rect 676 44 724 76
rect 756 44 804 76
rect 836 44 884 76
rect 916 44 964 76
rect 996 44 1044 76
rect 1076 44 1124 76
rect 1156 44 1204 76
rect 1236 44 1284 76
rect 1316 44 1364 76
rect 1396 44 1444 76
rect 1476 44 1524 76
rect 1556 44 1604 76
rect 1636 44 1684 76
rect 1716 44 1764 76
rect 1796 44 1844 76
rect 1876 44 1924 76
rect 1956 44 2004 76
rect 2036 44 2084 76
rect 2116 44 2164 76
rect 2196 44 2244 76
rect 2276 44 2324 76
rect 2356 44 2404 76
rect 2436 44 2484 76
rect 2516 44 2564 76
rect 2596 44 2644 76
rect 2676 44 2724 76
rect 2756 44 2804 76
rect 2836 44 2884 76
rect 2916 44 2964 76
rect 2996 44 3044 76
rect 3076 44 3124 76
rect 3156 44 3204 76
rect 3236 44 3284 76
rect 3316 44 3364 76
rect 3396 44 3444 76
rect 3476 44 3524 76
rect 3556 44 3604 76
rect 3636 44 3684 76
rect 3716 44 3764 76
rect 3796 44 3844 76
rect 3876 44 3924 76
rect 3956 44 4004 76
rect 4036 44 4084 76
rect 4116 44 4164 76
rect 4196 44 4244 76
rect 4276 44 4324 76
rect 4356 44 4404 76
rect 4436 44 4484 76
rect 4516 44 4564 76
rect 4596 44 4644 76
rect 4676 44 4724 76
rect 4756 44 4804 76
rect 4836 44 4884 76
rect 4916 44 4964 76
rect 4996 44 5044 76
rect 5076 44 5124 76
rect 5156 44 5204 76
rect 5236 44 5284 76
rect 5316 44 5364 76
rect 5396 44 5444 76
rect 5476 44 5524 76
rect 5556 44 5604 76
rect 5636 44 5684 76
rect 5716 44 5764 76
rect 5796 44 5844 76
rect 5876 44 5924 76
rect 5956 44 6004 76
rect 6036 44 6084 76
rect 6116 44 6164 76
rect 6196 44 6244 76
rect 6276 44 6324 76
rect 6356 44 6404 76
rect 6436 44 6484 76
rect 6516 44 6564 76
rect 6596 44 6644 76
rect 6676 44 6724 76
rect 6756 44 6804 76
rect 6836 44 6884 76
rect 6916 44 6964 76
rect 6996 44 7044 76
rect 7076 44 7124 76
rect 7156 44 7204 76
rect 7236 44 7284 76
rect 7316 44 7364 76
rect 7396 44 7444 76
rect 7476 44 7524 76
rect 7556 44 7604 76
rect 7636 44 7684 76
rect 7716 44 7764 76
rect 7796 44 7844 76
rect 7876 44 7924 76
rect 7956 44 8004 76
rect 8036 44 8084 76
rect 8116 44 8164 76
rect 8196 44 8244 76
rect 8276 44 8324 76
rect 8356 44 8404 76
rect 8436 44 8484 76
rect 8516 44 8564 76
rect 8596 44 8644 76
rect 8676 44 8724 76
rect 8756 44 8804 76
rect 8836 44 8884 76
rect 8916 44 8964 76
rect 8996 44 9044 76
rect 9076 44 9124 76
rect 9156 44 9204 76
rect 9236 44 9284 76
rect 9316 44 9364 76
rect 9396 44 9444 76
rect 9476 44 9524 76
rect 9556 44 9604 76
rect 9636 44 9684 76
rect 9716 44 9764 76
rect 9796 44 9844 76
rect 9876 44 9924 76
rect 9956 44 10004 76
rect 10036 44 10084 76
rect 10116 44 10164 76
rect 10196 44 10244 76
rect 10276 44 10324 76
rect 10356 44 10404 76
rect 10436 44 10484 76
rect 10516 44 10644 76
rect 10676 44 10804 76
rect 10836 44 10964 76
rect 10996 44 11000 76
rect -720 40 11000 44
rect -720 -4 11000 0
rect -720 -36 -716 -4
rect -684 -36 -556 -4
rect -524 -36 -396 -4
rect -364 -36 -316 -4
rect -284 -36 -236 -4
rect -204 -36 -156 -4
rect -124 -36 -76 -4
rect -44 -36 4 -4
rect 36 -36 84 -4
rect 116 -36 164 -4
rect 196 -36 244 -4
rect 276 -36 324 -4
rect 356 -36 404 -4
rect 436 -36 484 -4
rect 516 -36 564 -4
rect 596 -36 644 -4
rect 676 -36 724 -4
rect 756 -36 804 -4
rect 836 -36 884 -4
rect 916 -36 964 -4
rect 996 -36 1044 -4
rect 1076 -36 1124 -4
rect 1156 -36 1204 -4
rect 1236 -36 1284 -4
rect 1316 -36 1364 -4
rect 1396 -36 1444 -4
rect 1476 -36 1524 -4
rect 1556 -36 1604 -4
rect 1636 -36 1684 -4
rect 1716 -36 1764 -4
rect 1796 -36 1844 -4
rect 1876 -36 1924 -4
rect 1956 -36 2004 -4
rect 2036 -36 2084 -4
rect 2116 -36 2164 -4
rect 2196 -36 2244 -4
rect 2276 -36 2324 -4
rect 2356 -36 2404 -4
rect 2436 -36 2484 -4
rect 2516 -36 2564 -4
rect 2596 -36 2644 -4
rect 2676 -36 2724 -4
rect 2756 -36 2804 -4
rect 2836 -36 2884 -4
rect 2916 -36 2964 -4
rect 2996 -36 3044 -4
rect 3076 -36 3124 -4
rect 3156 -36 3204 -4
rect 3236 -36 3284 -4
rect 3316 -36 3364 -4
rect 3396 -36 3444 -4
rect 3476 -36 3524 -4
rect 3556 -36 3604 -4
rect 3636 -36 3684 -4
rect 3716 -36 3764 -4
rect 3796 -36 3844 -4
rect 3876 -36 3924 -4
rect 3956 -36 4004 -4
rect 4036 -36 4084 -4
rect 4116 -36 4164 -4
rect 4196 -36 4244 -4
rect 4276 -36 4324 -4
rect 4356 -36 4404 -4
rect 4436 -36 4484 -4
rect 4516 -36 4564 -4
rect 4596 -36 4644 -4
rect 4676 -36 4724 -4
rect 4756 -36 4804 -4
rect 4836 -36 4884 -4
rect 4916 -36 4964 -4
rect 4996 -36 5044 -4
rect 5076 -36 5124 -4
rect 5156 -36 5204 -4
rect 5236 -36 5284 -4
rect 5316 -36 5364 -4
rect 5396 -36 5444 -4
rect 5476 -36 5524 -4
rect 5556 -36 5604 -4
rect 5636 -36 5684 -4
rect 5716 -36 5764 -4
rect 5796 -36 5844 -4
rect 5876 -36 5924 -4
rect 5956 -36 6004 -4
rect 6036 -36 6084 -4
rect 6116 -36 6164 -4
rect 6196 -36 6244 -4
rect 6276 -36 6324 -4
rect 6356 -36 6404 -4
rect 6436 -36 6484 -4
rect 6516 -36 6564 -4
rect 6596 -36 6644 -4
rect 6676 -36 6724 -4
rect 6756 -36 6804 -4
rect 6836 -36 6884 -4
rect 6916 -36 6964 -4
rect 6996 -36 7044 -4
rect 7076 -36 7124 -4
rect 7156 -36 7204 -4
rect 7236 -36 7284 -4
rect 7316 -36 7364 -4
rect 7396 -36 7444 -4
rect 7476 -36 7524 -4
rect 7556 -36 7604 -4
rect 7636 -36 7684 -4
rect 7716 -36 7764 -4
rect 7796 -36 7844 -4
rect 7876 -36 7924 -4
rect 7956 -36 8004 -4
rect 8036 -36 8084 -4
rect 8116 -36 8164 -4
rect 8196 -36 8244 -4
rect 8276 -36 8324 -4
rect 8356 -36 8404 -4
rect 8436 -36 8484 -4
rect 8516 -36 8564 -4
rect 8596 -36 8644 -4
rect 8676 -36 8724 -4
rect 8756 -36 8804 -4
rect 8836 -36 8884 -4
rect 8916 -36 8964 -4
rect 8996 -36 9044 -4
rect 9076 -36 9124 -4
rect 9156 -36 9204 -4
rect 9236 -36 9284 -4
rect 9316 -36 9364 -4
rect 9396 -36 9444 -4
rect 9476 -36 9524 -4
rect 9556 -36 9604 -4
rect 9636 -36 9684 -4
rect 9716 -36 9764 -4
rect 9796 -36 9844 -4
rect 9876 -36 9924 -4
rect 9956 -36 10004 -4
rect 10036 -36 10084 -4
rect 10116 -36 10164 -4
rect 10196 -36 10244 -4
rect 10276 -36 10324 -4
rect 10356 -36 10404 -4
rect 10436 -36 10484 -4
rect 10516 -36 10644 -4
rect 10676 -36 10804 -4
rect 10836 -36 10964 -4
rect 10996 -36 11000 -4
rect -720 -40 11000 -36
rect -720 -84 11000 -80
rect -720 -116 -716 -84
rect -684 -116 -556 -84
rect -524 -116 -396 -84
rect -364 -116 -316 -84
rect -284 -116 -236 -84
rect -204 -116 -156 -84
rect -124 -116 -76 -84
rect -44 -116 4 -84
rect 36 -116 84 -84
rect 116 -116 164 -84
rect 196 -116 244 -84
rect 276 -116 324 -84
rect 356 -116 404 -84
rect 436 -116 484 -84
rect 516 -116 564 -84
rect 596 -116 644 -84
rect 676 -116 724 -84
rect 756 -116 804 -84
rect 836 -116 884 -84
rect 916 -116 964 -84
rect 996 -116 1044 -84
rect 1076 -116 1124 -84
rect 1156 -116 1204 -84
rect 1236 -116 1284 -84
rect 1316 -116 1364 -84
rect 1396 -116 1444 -84
rect 1476 -116 1524 -84
rect 1556 -116 1604 -84
rect 1636 -116 1684 -84
rect 1716 -116 1764 -84
rect 1796 -116 1844 -84
rect 1876 -116 1924 -84
rect 1956 -116 2004 -84
rect 2036 -116 2084 -84
rect 2116 -116 2164 -84
rect 2196 -116 2244 -84
rect 2276 -116 2324 -84
rect 2356 -116 2404 -84
rect 2436 -116 2484 -84
rect 2516 -116 2564 -84
rect 2596 -116 2644 -84
rect 2676 -116 2724 -84
rect 2756 -116 2804 -84
rect 2836 -116 2884 -84
rect 2916 -116 2964 -84
rect 2996 -116 3044 -84
rect 3076 -116 3124 -84
rect 3156 -116 3204 -84
rect 3236 -116 3284 -84
rect 3316 -116 3364 -84
rect 3396 -116 3444 -84
rect 3476 -116 3524 -84
rect 3556 -116 3604 -84
rect 3636 -116 3684 -84
rect 3716 -116 3764 -84
rect 3796 -116 3844 -84
rect 3876 -116 3924 -84
rect 3956 -116 4004 -84
rect 4036 -116 4084 -84
rect 4116 -116 4164 -84
rect 4196 -116 4244 -84
rect 4276 -116 4324 -84
rect 4356 -116 4404 -84
rect 4436 -116 4484 -84
rect 4516 -116 4564 -84
rect 4596 -116 4644 -84
rect 4676 -116 4724 -84
rect 4756 -116 4804 -84
rect 4836 -116 4884 -84
rect 4916 -116 4964 -84
rect 4996 -116 5044 -84
rect 5076 -116 5124 -84
rect 5156 -116 5204 -84
rect 5236 -116 5284 -84
rect 5316 -116 5364 -84
rect 5396 -116 5444 -84
rect 5476 -116 5524 -84
rect 5556 -116 5604 -84
rect 5636 -116 5684 -84
rect 5716 -116 5764 -84
rect 5796 -116 5844 -84
rect 5876 -116 5924 -84
rect 5956 -116 6004 -84
rect 6036 -116 6084 -84
rect 6116 -116 6164 -84
rect 6196 -116 6244 -84
rect 6276 -116 6324 -84
rect 6356 -116 6404 -84
rect 6436 -116 6484 -84
rect 6516 -116 6564 -84
rect 6596 -116 6644 -84
rect 6676 -116 6724 -84
rect 6756 -116 6804 -84
rect 6836 -116 6884 -84
rect 6916 -116 6964 -84
rect 6996 -116 7044 -84
rect 7076 -116 7124 -84
rect 7156 -116 7204 -84
rect 7236 -116 7284 -84
rect 7316 -116 7364 -84
rect 7396 -116 7444 -84
rect 7476 -116 7524 -84
rect 7556 -116 7604 -84
rect 7636 -116 7684 -84
rect 7716 -116 7764 -84
rect 7796 -116 7844 -84
rect 7876 -116 7924 -84
rect 7956 -116 8004 -84
rect 8036 -116 8084 -84
rect 8116 -116 8164 -84
rect 8196 -116 8244 -84
rect 8276 -116 8324 -84
rect 8356 -116 8404 -84
rect 8436 -116 8484 -84
rect 8516 -116 8564 -84
rect 8596 -116 8644 -84
rect 8676 -116 8724 -84
rect 8756 -116 8804 -84
rect 8836 -116 8884 -84
rect 8916 -116 8964 -84
rect 8996 -116 9044 -84
rect 9076 -116 9124 -84
rect 9156 -116 9204 -84
rect 9236 -116 9284 -84
rect 9316 -116 9364 -84
rect 9396 -116 9444 -84
rect 9476 -116 9524 -84
rect 9556 -116 9604 -84
rect 9636 -116 9684 -84
rect 9716 -116 9764 -84
rect 9796 -116 9844 -84
rect 9876 -116 9924 -84
rect 9956 -116 10004 -84
rect 10036 -116 10084 -84
rect 10116 -116 10164 -84
rect 10196 -116 10244 -84
rect 10276 -116 10324 -84
rect 10356 -116 10404 -84
rect 10436 -116 10484 -84
rect 10516 -116 10644 -84
rect 10676 -116 10804 -84
rect 10836 -116 10964 -84
rect 10996 -116 11000 -84
rect -720 -120 11000 -116
<< labels >>
rlabel metal3 -640 1040 -600 1080 0 ii
port 1 nsew
rlabel metal3 -480 1040 -440 1080 0 vi
port 2 nsew
rlabel metal3 10720 1040 10760 1080 0 n
rlabel metal3 10880 1040 10920 1080 0 vo
port 3 nsew
rlabel metal3 10960 1040 11000 1080 0 vssa
port 4 nsew
<< end >>
